magic
tech sky130A
magscale 1 2
timestamp 1605062100
<< locali >>
rect 5127 180249 5161 187967
rect 82223 180181 82257 187559
rect 4023 173653 4057 174163
rect 4023 164541 4057 164711
rect 4023 155361 4057 155667
rect 4023 141557 4057 146827
rect 4115 141625 4149 146759
rect 4023 123469 4057 128807
rect 4115 123537 4149 128603
rect 4023 105449 4057 110651
rect 4115 105517 4149 110583
rect 4023 97833 4057 99091
rect 4023 97765 4057 97799
rect 4023 97731 4149 97765
rect 3287 96201 3321 96303
rect 4023 96133 4057 96303
rect 4115 94705 4149 97731
rect 5805 97527 5897 97561
rect 5771 96881 5805 97323
rect 5863 97085 5897 97527
rect 81303 97085 81337 97391
rect 5863 97051 5955 97085
rect 14971 96745 15005 96983
rect 81395 96949 81429 97255
rect 83051 97017 83085 97595
rect 19571 96813 19605 96847
rect 19513 96779 19605 96813
rect 72747 96677 72781 96779
rect 26011 95589 26045 95827
rect 28311 95385 28345 95759
rect 57843 95453 57877 95555
rect 4057 94671 4149 94705
rect 4023 94229 4057 94671
rect 46619 94637 46653 94943
rect 51771 94637 51805 95079
rect 55727 94297 55761 94671
rect 55819 94433 55853 95011
rect 58947 94637 58981 94875
rect 59717 94671 59959 94705
rect 64651 93957 64685 94399
rect 69251 93481 69285 94807
rect 73667 94229 73701 96779
rect 74771 96473 74805 96847
rect 81487 96813 81521 96915
rect 80015 96473 80049 96711
rect 80107 96473 80141 96575
rect 80015 96439 80141 96473
rect 82499 96201 82533 96507
rect 77991 94637 78025 94739
rect 78175 94297 78209 94671
rect 59959 92801 59993 92903
rect 81303 92189 81337 93039
rect 81395 92393 81429 92563
rect 4023 80969 4057 89911
rect 5403 83417 5437 89911
rect 4023 56285 4057 61555
rect 83143 56421 83177 56523
rect 3563 44521 3597 44827
rect 4023 38333 4057 44759
rect 4023 16573 4057 22931
rect 4115 15281 4149 24155
rect 4023 3313 4057 13615
rect 4023 2701 4057 3279
rect 4667 2905 4701 3211
rect 5035 2633 5069 2803
rect 5771 2769 5805 3415
rect 61649 2871 61891 2905
rect 5587 2429 5621 2735
rect 57475 2565 57509 2803
rect 61833 2735 61891 2769
rect 81303 2701 81337 3347
rect 69803 2157 69837 2463
rect 78727 2157 78761 2531
rect 81395 1409 81429 3687
rect 82591 593 82625 8787
rect 82775 3517 82809 4027
rect 84063 3313 84097 3483
<< viali >>
rect 5127 187967 5161 188001
rect 3563 182731 3597 182765
rect 3563 181643 3597 181677
rect 5127 180215 5161 180249
rect 82223 187559 82257 187593
rect 3563 180147 3597 180181
rect 82223 180147 82257 180181
rect 3563 178855 3597 178889
rect 3563 176679 3597 176713
rect 3471 175591 3505 175625
rect 4023 174163 4057 174197
rect 3563 173959 3597 173993
rect 4023 173619 4057 173653
rect 4023 164711 4057 164745
rect 4023 164507 4057 164541
rect 4023 155667 4057 155701
rect 4023 155327 4057 155361
rect 4023 146827 4057 146861
rect 4115 146759 4149 146793
rect 4115 141591 4149 141625
rect 4023 141523 4057 141557
rect 4023 128807 4057 128841
rect 4115 128603 4149 128637
rect 4115 123503 4149 123537
rect 4023 123435 4057 123469
rect 3563 116431 3597 116465
rect 3471 114731 3505 114765
rect 4023 110651 4057 110685
rect 4115 110583 4149 110617
rect 4115 105483 4149 105517
rect 4023 105415 4057 105449
rect 4023 99091 4057 99125
rect 3103 98343 3137 98377
rect 3563 98343 3597 98377
rect 3563 98139 3597 98173
rect 83879 98139 83913 98173
rect 2367 97799 2401 97833
rect 2827 97799 2861 97833
rect 4023 97799 4057 97833
rect 2827 97595 2861 97629
rect 3195 97595 3229 97629
rect 1723 97459 1757 97493
rect 2091 97255 2125 97289
rect 2459 97255 2493 97289
rect 3471 97255 3505 97289
rect 987 97051 1021 97085
rect 1355 96983 1389 97017
rect 2091 96983 2125 97017
rect 2827 96847 2861 96881
rect 1723 96711 1757 96745
rect 2459 96711 2493 96745
rect 3563 96711 3597 96745
rect 3195 96303 3229 96337
rect 3287 96303 3321 96337
rect 4023 96303 4057 96337
rect 2091 96167 2125 96201
rect 2459 96167 2493 96201
rect 2827 96167 2861 96201
rect 3287 96167 3321 96201
rect 3563 96167 3597 96201
rect 4023 96099 4057 96133
rect 2827 95963 2861 95997
rect 3563 95963 3597 95997
rect 2459 95691 2493 95725
rect 3195 95419 3229 95453
rect 3563 95351 3597 95385
rect 83051 97595 83085 97629
rect 84247 97595 84281 97629
rect 5771 97527 5805 97561
rect 5771 97323 5805 97357
rect 81303 97391 81337 97425
rect 5955 97051 5989 97085
rect 81303 97051 81337 97085
rect 81395 97255 81429 97289
rect 5771 96847 5805 96881
rect 14971 96983 15005 97017
rect 83787 97527 83821 97561
rect 84155 97051 84189 97085
rect 83051 96983 83085 97017
rect 81395 96915 81429 96949
rect 81487 96915 81521 96949
rect 19571 96847 19605 96881
rect 74771 96847 74805 96881
rect 19479 96779 19513 96813
rect 72747 96779 72781 96813
rect 14971 96711 15005 96745
rect 72747 96643 72781 96677
rect 73667 96779 73701 96813
rect 26011 95827 26045 95861
rect 26011 95555 26045 95589
rect 28311 95759 28345 95793
rect 57843 95555 57877 95589
rect 57843 95419 57877 95453
rect 28311 95351 28345 95385
rect 51771 95079 51805 95113
rect 4023 94671 4057 94705
rect 46619 94943 46653 94977
rect 46619 94603 46653 94637
rect 55819 95011 55853 95045
rect 51771 94603 51805 94637
rect 55727 94671 55761 94705
rect 58947 94875 58981 94909
rect 69251 94807 69285 94841
rect 59683 94671 59717 94705
rect 59959 94671 59993 94705
rect 58947 94603 58981 94637
rect 55819 94399 55853 94433
rect 64651 94399 64685 94433
rect 55727 94263 55761 94297
rect 4023 94195 4057 94229
rect 64651 93923 64685 93957
rect 83787 96847 83821 96881
rect 81487 96779 81521 96813
rect 84615 96779 84649 96813
rect 74771 96439 74805 96473
rect 80015 96711 80049 96745
rect 84983 96711 85017 96745
rect 80107 96575 80141 96609
rect 82499 96507 82533 96541
rect 83787 96303 83821 96337
rect 84247 96303 84281 96337
rect 82499 96167 82533 96201
rect 83879 95963 83913 95997
rect 77991 94739 78025 94773
rect 77991 94603 78025 94637
rect 78175 94671 78209 94705
rect 78175 94263 78209 94297
rect 73667 94195 73701 94229
rect 69251 93447 69285 93481
rect 83787 93447 83821 93481
rect 81303 93039 81337 93073
rect 59959 92903 59993 92937
rect 59959 92767 59993 92801
rect 83787 92903 83821 92937
rect 81395 92563 81429 92597
rect 81395 92359 81429 92393
rect 81303 92155 81337 92189
rect 83879 91815 83913 91849
rect 4023 89911 4057 89945
rect 3563 88551 3597 88585
rect 3563 87803 3597 87837
rect 3563 85831 3597 85865
rect 3563 84811 3597 84845
rect 3563 83111 3597 83145
rect 3471 82159 3505 82193
rect 5403 89911 5437 89945
rect 5403 83383 5437 83417
rect 4023 80935 4057 80969
rect 3563 79847 3597 79881
rect 4023 61555 4057 61589
rect 83143 56523 83177 56557
rect 83143 56387 83177 56421
rect 4023 56251 4057 56285
rect 3563 44827 3597 44861
rect 3563 44487 3597 44521
rect 4023 44759 4057 44793
rect 4023 38299 4057 38333
rect 83879 31431 83913 31465
rect 83879 29867 83913 29901
rect 83879 28711 83913 28745
rect 83879 27079 83913 27113
rect 83787 25991 83821 26025
rect 4115 24155 4149 24189
rect 4023 22931 4057 22965
rect 3563 22523 3597 22557
rect 3563 20551 3597 20585
rect 4023 16539 4057 16573
rect 83879 23815 83913 23849
rect 83879 22931 83913 22965
rect 4115 15247 4149 15281
rect 4023 13615 4057 13649
rect 3563 5115 3597 5149
rect 3563 4571 3597 4605
rect 2827 4231 2861 4265
rect 1999 4027 2033 4061
rect 2459 4027 2493 4061
rect 2827 4027 2861 4061
rect 3563 3959 3597 3993
rect 3195 3891 3229 3925
rect 2827 3483 2861 3517
rect 82591 8787 82625 8821
rect 81395 3687 81429 3721
rect 2091 3279 2125 3313
rect 4023 3279 4057 3313
rect 1723 3211 1757 3245
rect 1355 3143 1389 3177
rect 2459 3143 2493 3177
rect 3563 3143 3597 3177
rect 1355 2939 1389 2973
rect 2827 2939 2861 2973
rect 1723 2871 1757 2905
rect 2459 2871 2493 2905
rect 3195 2871 3229 2905
rect 3563 2803 3597 2837
rect 5771 3415 5805 3449
rect 4667 3211 4701 3245
rect 4667 2871 4701 2905
rect 619 2667 653 2701
rect 2091 2667 2125 2701
rect 4023 2667 4057 2701
rect 5035 2803 5069 2837
rect 81303 3347 81337 3381
rect 61615 2871 61649 2905
rect 61891 2871 61925 2905
rect 987 2599 1021 2633
rect 5035 2599 5069 2633
rect 5587 2735 5621 2769
rect 5771 2735 5805 2769
rect 57475 2803 57509 2837
rect 61799 2735 61833 2769
rect 61891 2735 61925 2769
rect 81303 2667 81337 2701
rect 57475 2531 57509 2565
rect 78727 2531 78761 2565
rect 5587 2395 5621 2429
rect 69803 2463 69837 2497
rect 2827 2259 2861 2293
rect 2459 2123 2493 2157
rect 69803 2123 69837 2157
rect 78727 2123 78761 2157
rect 1723 2055 1757 2089
rect 2091 2055 2125 2089
rect 3563 2055 3597 2089
rect 81395 1375 81429 1409
rect 82775 4027 82809 4061
rect 83787 4027 83821 4061
rect 82775 3483 82809 3517
rect 84063 3483 84097 3517
rect 84615 3483 84649 3517
rect 84063 3279 84097 3313
rect 84155 3211 84189 3245
rect 83787 3143 83821 3177
rect 83787 2939 83821 2973
rect 84247 2939 84281 2973
rect 84983 2871 85017 2905
rect 84615 2735 84649 2769
rect 83879 2191 83913 2225
rect 84155 2123 84189 2157
rect 82591 559 82625 593
<< metal1 >>
rect 5848 188502 5854 188554
rect 5906 188542 5912 188554
rect 82484 188542 82490 188554
rect 5906 188514 82490 188542
rect 5906 188502 5912 188514
rect 82484 188502 82490 188514
rect 82542 188502 82548 188554
rect 5204 188434 5210 188486
rect 5262 188474 5268 188486
rect 84324 188474 84330 188486
rect 5262 188446 84330 188474
rect 5262 188434 5268 188446
rect 84324 188434 84330 188446
rect 84382 188434 84388 188486
rect 5296 188366 5302 188418
rect 5354 188406 5360 188418
rect 85152 188406 85158 188418
rect 5354 188378 85158 188406
rect 5354 188366 5360 188378
rect 85152 188366 85158 188378
rect 85210 188366 85216 188418
rect 2628 188298 2634 188350
rect 2686 188338 2692 188350
rect 82116 188338 82122 188350
rect 2686 188310 82122 188338
rect 2686 188298 2692 188310
rect 82116 188298 82122 188310
rect 82174 188298 82180 188350
rect 2352 188230 2358 188282
rect 2410 188270 2416 188282
rect 81840 188270 81846 188282
rect 2410 188242 81846 188270
rect 2410 188230 2416 188242
rect 81840 188230 81846 188242
rect 81898 188230 81904 188282
rect 2812 188162 2818 188214
rect 2870 188202 2876 188214
rect 82392 188202 82398 188214
rect 2870 188174 82398 188202
rect 2870 188162 2876 188174
rect 82392 188162 82398 188174
rect 82450 188162 82456 188214
rect 2076 188094 2082 188146
rect 2134 188134 2140 188146
rect 81932 188134 81938 188146
rect 2134 188106 81938 188134
rect 2134 188094 2140 188106
rect 81932 188094 81938 188106
rect 81990 188094 81996 188146
rect 2720 188026 2726 188078
rect 2778 188066 2784 188078
rect 82576 188066 82582 188078
rect 2778 188038 82582 188066
rect 2778 188026 2784 188038
rect 82576 188026 82582 188038
rect 82634 188026 82640 188078
rect 5115 188001 5173 188007
rect 5115 187967 5127 188001
rect 5161 187998 5173 188001
rect 82208 187998 82214 188010
rect 5161 187970 82214 187998
rect 5161 187967 5173 187970
rect 5115 187961 5173 187967
rect 82208 187958 82214 187970
rect 82266 187958 82272 188010
rect 2444 187890 2450 187942
rect 2502 187930 2508 187942
rect 83220 187930 83226 187942
rect 2502 187902 83226 187930
rect 2502 187890 2508 187902
rect 83220 187890 83226 187902
rect 83278 187890 83284 187942
rect 1340 187822 1346 187874
rect 1398 187862 1404 187874
rect 82300 187862 82306 187874
rect 1398 187834 82306 187862
rect 1398 187822 1404 187834
rect 82300 187822 82306 187834
rect 82358 187822 82364 187874
rect 4744 187550 4750 187602
rect 4802 187590 4808 187602
rect 82211 187593 82269 187599
rect 82211 187590 82223 187593
rect 4802 187562 82223 187590
rect 4802 187550 4808 187562
rect 82211 187559 82223 187562
rect 82257 187559 82269 187593
rect 82211 187553 82269 187559
rect 38 187500 3902 187522
rect 38 187448 2916 187500
rect 2968 187448 2980 187500
rect 3032 187448 3044 187500
rect 3096 187448 3108 187500
rect 3160 187448 3902 187500
rect 38 187426 3902 187448
rect 83298 187500 87806 187522
rect 83298 187448 86916 187500
rect 86968 187448 86980 187500
rect 87032 187448 87044 187500
rect 87096 187448 87108 187500
rect 87160 187448 87806 187500
rect 83298 187426 87806 187448
rect 5112 187346 5118 187398
rect 5170 187386 5176 187398
rect 84784 187386 84790 187398
rect 5170 187358 84790 187386
rect 5170 187346 5176 187358
rect 84784 187346 84790 187358
rect 84842 187346 84848 187398
rect 4560 187278 4566 187330
rect 4618 187318 4624 187330
rect 82024 187318 82030 187330
rect 4618 187290 82030 187318
rect 4618 187278 4624 187290
rect 82024 187278 82030 187290
rect 82082 187278 82088 187330
rect 5756 187210 5762 187262
rect 5814 187250 5820 187262
rect 84048 187250 84054 187262
rect 5814 187222 84054 187250
rect 5814 187210 5820 187222
rect 84048 187210 84054 187222
rect 84106 187210 84112 187262
rect 4468 187142 4474 187194
rect 4526 187182 4532 187194
rect 83312 187182 83318 187194
rect 4526 187154 83318 187182
rect 4526 187142 4532 187154
rect 83312 187142 83318 187154
rect 83370 187142 83376 187194
rect 4928 187074 4934 187126
rect 4986 187114 4992 187126
rect 84416 187114 84422 187126
rect 4986 187086 84422 187114
rect 4986 187074 4992 187086
rect 84416 187074 84422 187086
rect 84474 187074 84480 187126
rect 4192 187006 4198 187058
rect 4250 187046 4256 187058
rect 84324 187046 84330 187058
rect 4250 187018 84330 187046
rect 4250 187006 4256 187018
rect 84324 187006 84330 187018
rect 84382 187006 84388 187058
rect 38 186956 3902 186978
rect 38 186904 916 186956
rect 968 186904 980 186956
rect 1032 186904 1044 186956
rect 1096 186904 1108 186956
rect 1160 186904 3902 186956
rect 38 186882 3902 186904
rect 83298 186956 87806 186978
rect 83298 186904 84916 186956
rect 84968 186904 84980 186956
rect 85032 186904 85044 186956
rect 85096 186904 85108 186956
rect 85160 186904 87806 186956
rect 83298 186882 87806 186904
rect 4652 186802 4658 186854
rect 4710 186842 4716 186854
rect 84692 186842 84698 186854
rect 4710 186814 84698 186842
rect 4710 186802 4716 186814
rect 84692 186802 84698 186814
rect 84750 186802 84756 186854
rect 4100 186734 4106 186786
rect 4158 186774 4164 186786
rect 84140 186774 84146 186786
rect 4158 186746 84146 186774
rect 4158 186734 4164 186746
rect 84140 186734 84146 186746
rect 84198 186734 84204 186786
rect 4836 186666 4842 186718
rect 4894 186706 4900 186718
rect 85152 186706 85158 186718
rect 4894 186678 85158 186706
rect 4894 186666 4900 186678
rect 85152 186666 85158 186678
rect 85210 186666 85216 186718
rect 3364 186598 3370 186650
rect 3422 186638 3428 186650
rect 84508 186638 84514 186650
rect 3422 186610 84514 186638
rect 3422 186598 3428 186610
rect 84508 186598 84514 186610
rect 84566 186598 84572 186650
rect 1984 186530 1990 186582
rect 2042 186570 2048 186582
rect 83956 186570 83962 186582
rect 2042 186542 83962 186570
rect 2042 186530 2048 186542
rect 83956 186530 83962 186542
rect 84014 186530 84020 186582
rect 38 186412 3902 186434
rect 38 186360 2916 186412
rect 2968 186360 2980 186412
rect 3032 186360 3044 186412
rect 3096 186360 3108 186412
rect 3160 186360 3902 186412
rect 38 186338 3902 186360
rect 83298 186412 87806 186434
rect 83298 186360 86916 186412
rect 86968 186360 86980 186412
rect 87032 186360 87044 186412
rect 87096 186360 87108 186412
rect 87160 186360 87806 186412
rect 83298 186338 87806 186360
rect 38 185868 3902 185890
rect 38 185816 916 185868
rect 968 185816 980 185868
rect 1032 185816 1044 185868
rect 1096 185816 1108 185868
rect 1160 185816 3902 185868
rect 38 185794 3902 185816
rect 83298 185868 87806 185890
rect 83298 185816 84916 185868
rect 84968 185816 84980 185868
rect 85032 185816 85044 185868
rect 85096 185816 85108 185868
rect 85160 185816 87806 185868
rect 83298 185794 87806 185816
rect 84324 185374 84330 185426
rect 84382 185414 84388 185426
rect 84784 185414 84790 185426
rect 84382 185386 84790 185414
rect 84382 185374 84388 185386
rect 84784 185374 84790 185386
rect 84842 185374 84848 185426
rect 38 185324 3902 185346
rect 38 185272 2916 185324
rect 2968 185272 2980 185324
rect 3032 185272 3044 185324
rect 3096 185272 3108 185324
rect 3160 185272 3902 185324
rect 38 185250 3902 185272
rect 83298 185324 87806 185346
rect 83298 185272 86916 185324
rect 86968 185272 86980 185324
rect 87032 185272 87044 185324
rect 87096 185272 87108 185324
rect 87160 185272 87806 185324
rect 83298 185250 87806 185272
rect 38 184780 3902 184802
rect 38 184728 916 184780
rect 968 184728 980 184780
rect 1032 184728 1044 184780
rect 1096 184728 1108 184780
rect 1160 184728 3902 184780
rect 38 184706 3902 184728
rect 83298 184780 87806 184802
rect 83298 184728 84916 184780
rect 84968 184728 84980 184780
rect 85032 184728 85044 184780
rect 85096 184728 85108 184780
rect 85160 184728 87806 184780
rect 83298 184706 87806 184728
rect 38 184236 3902 184258
rect 38 184184 2916 184236
rect 2968 184184 2980 184236
rect 3032 184184 3044 184236
rect 3096 184184 3108 184236
rect 3160 184184 3902 184236
rect 38 184162 3902 184184
rect 83298 184236 87806 184258
rect 83298 184184 86916 184236
rect 86968 184184 86980 184236
rect 87032 184184 87044 184236
rect 87096 184184 87108 184236
rect 87160 184184 87806 184236
rect 83298 184162 87806 184184
rect 38 183692 3902 183714
rect 38 183640 916 183692
rect 968 183640 980 183692
rect 1032 183640 1044 183692
rect 1096 183640 1108 183692
rect 1160 183640 3902 183692
rect 38 183618 3902 183640
rect 83298 183692 87806 183714
rect 83298 183640 84916 183692
rect 84968 183640 84980 183692
rect 85032 183640 85044 183692
rect 85096 183640 85108 183692
rect 85160 183640 87806 183692
rect 83298 183618 87806 183640
rect 38 183148 3902 183170
rect 38 183096 2916 183148
rect 2968 183096 2980 183148
rect 3032 183096 3044 183148
rect 3096 183096 3108 183148
rect 3160 183096 3902 183148
rect 38 183074 3902 183096
rect 83298 183148 87806 183170
rect 83298 183096 86916 183148
rect 86968 183096 86980 183148
rect 87032 183096 87044 183148
rect 87096 183096 87108 183148
rect 87160 183096 87806 183148
rect 83298 183074 87806 183096
rect 3551 182765 3609 182771
rect 3551 182731 3563 182765
rect 3597 182762 3609 182765
rect 3916 182762 3922 182774
rect 3597 182734 3922 182762
rect 3597 182731 3609 182734
rect 3551 182725 3609 182731
rect 3916 182722 3922 182734
rect 3974 182722 3980 182774
rect 38 182604 3902 182626
rect 38 182552 916 182604
rect 968 182552 980 182604
rect 1032 182552 1044 182604
rect 1096 182552 1108 182604
rect 1160 182552 3902 182604
rect 38 182530 3902 182552
rect 83298 182604 87806 182626
rect 83298 182552 84916 182604
rect 84968 182552 84980 182604
rect 85032 182552 85044 182604
rect 85096 182552 85108 182604
rect 85160 182552 87806 182604
rect 83298 182530 87806 182552
rect 84232 182246 84238 182298
rect 84290 182286 84296 182298
rect 84416 182286 84422 182298
rect 84290 182258 84422 182286
rect 84290 182246 84296 182258
rect 84416 182246 84422 182258
rect 84474 182246 84480 182298
rect 84416 182110 84422 182162
rect 84474 182150 84480 182162
rect 84600 182150 84606 182162
rect 84474 182122 84606 182150
rect 84474 182110 84480 182122
rect 84600 182110 84606 182122
rect 84658 182110 84664 182162
rect 38 182060 3902 182082
rect 38 182008 2916 182060
rect 2968 182008 2980 182060
rect 3032 182008 3044 182060
rect 3096 182008 3108 182060
rect 3160 182008 3902 182060
rect 38 181986 3902 182008
rect 83298 182060 87806 182082
rect 83298 182008 86916 182060
rect 86968 182008 86980 182060
rect 87032 182008 87044 182060
rect 87096 182008 87108 182060
rect 87160 182008 87806 182060
rect 83298 181986 87806 182008
rect 3548 181674 3554 181686
rect 3509 181646 3554 181674
rect 3548 181634 3554 181646
rect 3606 181634 3612 181686
rect 38 181516 3902 181538
rect 38 181464 916 181516
rect 968 181464 980 181516
rect 1032 181464 1044 181516
rect 1096 181464 1108 181516
rect 1160 181464 3902 181516
rect 38 181442 3902 181464
rect 83298 181516 87806 181538
rect 83298 181464 84916 181516
rect 84968 181464 84980 181516
rect 85032 181464 85044 181516
rect 85096 181464 85108 181516
rect 85160 181464 87806 181516
rect 83298 181442 87806 181464
rect 38 180972 3902 180994
rect 38 180920 2916 180972
rect 2968 180920 2980 180972
rect 3032 180920 3044 180972
rect 3096 180920 3108 180972
rect 3160 180920 3902 180972
rect 38 180898 3902 180920
rect 83298 180972 87806 180994
rect 83298 180920 86916 180972
rect 86968 180920 86980 180972
rect 87032 180920 87044 180972
rect 87096 180920 87108 180972
rect 87160 180920 87806 180972
rect 83298 180898 87806 180920
rect 38 180428 3902 180450
rect 38 180376 916 180428
rect 968 180376 980 180428
rect 1032 180376 1044 180428
rect 1096 180376 1108 180428
rect 1160 180376 3902 180428
rect 38 180354 3902 180376
rect 83298 180428 87806 180450
rect 83298 180376 84916 180428
rect 84968 180376 84980 180428
rect 85032 180376 85044 180428
rect 85096 180376 85108 180428
rect 85160 180376 87806 180428
rect 83298 180354 87806 180376
rect 5115 180249 5173 180255
rect 5115 180246 5127 180249
rect 2186 180218 5127 180246
rect 2186 180190 2214 180218
rect 5115 180215 5127 180218
rect 5161 180215 5173 180249
rect 5115 180209 5173 180215
rect 2168 180138 2174 180190
rect 2226 180138 2232 180190
rect 3548 180178 3554 180190
rect 3509 180150 3554 180178
rect 3548 180138 3554 180150
rect 3606 180138 3612 180190
rect 82211 180181 82269 180187
rect 82211 180147 82223 180181
rect 82257 180178 82269 180181
rect 84324 180178 84330 180190
rect 82257 180150 84330 180178
rect 82257 180147 82269 180150
rect 82211 180141 82269 180147
rect 84324 180138 84330 180150
rect 84382 180138 84388 180190
rect 38 179884 3902 179906
rect 38 179832 2916 179884
rect 2968 179832 2980 179884
rect 3032 179832 3044 179884
rect 3096 179832 3108 179884
rect 3160 179832 3902 179884
rect 38 179810 3902 179832
rect 83298 179884 87806 179906
rect 83298 179832 86916 179884
rect 86968 179832 86980 179884
rect 87032 179832 87044 179884
rect 87096 179832 87108 179884
rect 87160 179832 87806 179884
rect 83298 179810 87806 179832
rect 38 179340 3902 179362
rect 38 179288 916 179340
rect 968 179288 980 179340
rect 1032 179288 1044 179340
rect 1096 179288 1108 179340
rect 1160 179288 3902 179340
rect 38 179266 3902 179288
rect 83298 179340 87806 179362
rect 83298 179288 84916 179340
rect 84968 179288 84980 179340
rect 85032 179288 85044 179340
rect 85096 179288 85108 179340
rect 85160 179288 87806 179340
rect 83298 179266 87806 179288
rect 3551 178889 3609 178895
rect 3551 178855 3563 178889
rect 3597 178886 3609 178889
rect 4008 178886 4014 178898
rect 3597 178858 4014 178886
rect 3597 178855 3609 178858
rect 3551 178849 3609 178855
rect 4008 178846 4014 178858
rect 4066 178846 4072 178898
rect 38 178796 3902 178818
rect 38 178744 2916 178796
rect 2968 178744 2980 178796
rect 3032 178744 3044 178796
rect 3096 178744 3108 178796
rect 3160 178744 3902 178796
rect 38 178722 3902 178744
rect 83298 178796 87806 178818
rect 83298 178744 86916 178796
rect 86968 178744 86980 178796
rect 87032 178744 87044 178796
rect 87096 178744 87108 178796
rect 87160 178744 87806 178796
rect 83298 178722 87806 178744
rect 84692 178506 84698 178558
rect 84750 178506 84756 178558
rect 84710 178354 84738 178506
rect 84692 178302 84698 178354
rect 84750 178302 84756 178354
rect 38 178252 3902 178274
rect 38 178200 916 178252
rect 968 178200 980 178252
rect 1032 178200 1044 178252
rect 1096 178200 1108 178252
rect 1160 178200 3902 178252
rect 38 178178 3902 178200
rect 83298 178252 87806 178274
rect 83298 178200 84916 178252
rect 84968 178200 84980 178252
rect 85032 178200 85044 178252
rect 85096 178200 85108 178252
rect 85160 178200 87806 178252
rect 83298 178178 87806 178200
rect 38 177708 3902 177730
rect 38 177656 2916 177708
rect 2968 177656 2980 177708
rect 3032 177656 3044 177708
rect 3096 177656 3108 177708
rect 3160 177656 3902 177708
rect 38 177634 3902 177656
rect 83298 177708 87806 177730
rect 83298 177656 86916 177708
rect 86968 177656 86980 177708
rect 87032 177656 87044 177708
rect 87096 177656 87108 177708
rect 87160 177656 87806 177708
rect 83298 177634 87806 177656
rect 38 177164 3902 177186
rect 38 177112 916 177164
rect 968 177112 980 177164
rect 1032 177112 1044 177164
rect 1096 177112 1108 177164
rect 1160 177112 3902 177164
rect 38 177090 3902 177112
rect 83298 177164 87806 177186
rect 83298 177112 84916 177164
rect 84968 177112 84980 177164
rect 85032 177112 85044 177164
rect 85096 177112 85108 177164
rect 85160 177112 87806 177164
rect 83298 177090 87806 177112
rect 3551 176713 3609 176719
rect 3551 176679 3563 176713
rect 3597 176710 3609 176713
rect 3640 176710 3646 176722
rect 3597 176682 3646 176710
rect 3597 176679 3609 176682
rect 3551 176673 3609 176679
rect 3640 176670 3646 176682
rect 3698 176670 3704 176722
rect 38 176620 3902 176642
rect 38 176568 2916 176620
rect 2968 176568 2980 176620
rect 3032 176568 3044 176620
rect 3096 176568 3108 176620
rect 3160 176568 3902 176620
rect 38 176546 3902 176568
rect 83298 176620 87806 176642
rect 83298 176568 86916 176620
rect 86968 176568 86980 176620
rect 87032 176568 87044 176620
rect 87096 176568 87108 176620
rect 87160 176568 87806 176620
rect 83298 176546 87806 176568
rect 38 176076 3902 176098
rect 38 176024 916 176076
rect 968 176024 980 176076
rect 1032 176024 1044 176076
rect 1096 176024 1108 176076
rect 1160 176024 3902 176076
rect 38 176002 3902 176024
rect 83298 176076 87806 176098
rect 83298 176024 84916 176076
rect 84968 176024 84980 176076
rect 85032 176024 85044 176076
rect 85096 176024 85108 176076
rect 85160 176024 87806 176076
rect 83298 176002 87806 176024
rect 3272 175582 3278 175634
rect 3330 175622 3336 175634
rect 3459 175625 3517 175631
rect 3459 175622 3471 175625
rect 3330 175594 3471 175622
rect 3330 175582 3336 175594
rect 3459 175591 3471 175594
rect 3505 175591 3517 175625
rect 3459 175585 3517 175591
rect 84600 175582 84606 175634
rect 84658 175622 84664 175634
rect 84784 175622 84790 175634
rect 84658 175594 84790 175622
rect 84658 175582 84664 175594
rect 84784 175582 84790 175594
rect 84842 175582 84848 175634
rect 38 175532 3902 175554
rect 38 175480 2916 175532
rect 2968 175480 2980 175532
rect 3032 175480 3044 175532
rect 3096 175480 3108 175532
rect 3160 175480 3902 175532
rect 38 175458 3902 175480
rect 83298 175532 87806 175554
rect 83298 175480 86916 175532
rect 86968 175480 86980 175532
rect 87032 175480 87044 175532
rect 87096 175480 87108 175532
rect 87160 175480 87806 175532
rect 83298 175458 87806 175480
rect 38 174988 3902 175010
rect 38 174936 916 174988
rect 968 174936 980 174988
rect 1032 174936 1044 174988
rect 1096 174936 1108 174988
rect 1160 174936 3902 174988
rect 38 174914 3902 174936
rect 83298 174988 87806 175010
rect 83298 174936 84916 174988
rect 84968 174936 84980 174988
rect 85032 174936 85044 174988
rect 85096 174936 85108 174988
rect 85160 174936 87806 174988
rect 83298 174914 87806 174936
rect 38 174444 3902 174466
rect 38 174392 2916 174444
rect 2968 174392 2980 174444
rect 3032 174392 3044 174444
rect 3096 174392 3108 174444
rect 3160 174392 3902 174444
rect 38 174370 3902 174392
rect 83298 174444 87806 174466
rect 83298 174392 86916 174444
rect 86968 174392 86980 174444
rect 87032 174392 87044 174444
rect 87096 174392 87108 174444
rect 87160 174392 87806 174444
rect 83298 174370 87806 174392
rect 3640 174154 3646 174206
rect 3698 174194 3704 174206
rect 4011 174197 4069 174203
rect 4011 174194 4023 174197
rect 3698 174166 4023 174194
rect 3698 174154 3704 174166
rect 4011 174163 4023 174166
rect 4057 174163 4069 174197
rect 4011 174157 4069 174163
rect 3551 173993 3609 173999
rect 3551 173959 3563 173993
rect 3597 173990 3609 173993
rect 3640 173990 3646 174002
rect 3597 173962 3646 173990
rect 3597 173959 3609 173962
rect 3551 173953 3609 173959
rect 3640 173950 3646 173962
rect 3698 173950 3704 174002
rect 38 173900 3902 173922
rect 38 173848 916 173900
rect 968 173848 980 173900
rect 1032 173848 1044 173900
rect 1096 173848 1108 173900
rect 1160 173848 3902 173900
rect 38 173826 3902 173848
rect 83298 173900 87806 173922
rect 83298 173848 84916 173900
rect 84968 173848 84980 173900
rect 85032 173848 85044 173900
rect 85096 173848 85108 173900
rect 85160 173848 87806 173900
rect 83298 173826 87806 173848
rect 2168 173610 2174 173662
rect 2226 173610 2232 173662
rect 3456 173610 3462 173662
rect 3514 173650 3520 173662
rect 4011 173653 4069 173659
rect 4011 173650 4023 173653
rect 3514 173622 4023 173650
rect 3514 173610 3520 173622
rect 4011 173619 4023 173622
rect 4057 173619 4069 173653
rect 4011 173613 4069 173619
rect 84324 173610 84330 173662
rect 84382 173650 84388 173662
rect 84784 173650 84790 173662
rect 84382 173622 84790 173650
rect 84382 173610 84388 173622
rect 84784 173610 84790 173622
rect 84842 173610 84848 173662
rect 2186 173582 2214 173610
rect 2260 173582 2266 173594
rect 2186 173554 2266 173582
rect 2260 173542 2266 173554
rect 2318 173542 2324 173594
rect 38 173356 3902 173378
rect 38 173304 2916 173356
rect 2968 173304 2980 173356
rect 3032 173304 3044 173356
rect 3096 173304 3108 173356
rect 3160 173304 3902 173356
rect 38 173282 3902 173304
rect 83298 173356 87806 173378
rect 83298 173304 86916 173356
rect 86968 173304 86980 173356
rect 87032 173304 87044 173356
rect 87096 173304 87108 173356
rect 87160 173304 87806 173356
rect 83298 173282 87806 173304
rect 38 172812 3902 172834
rect 38 172760 916 172812
rect 968 172760 980 172812
rect 1032 172760 1044 172812
rect 1096 172760 1108 172812
rect 1160 172760 3902 172812
rect 38 172738 3902 172760
rect 83298 172812 87806 172834
rect 83298 172760 84916 172812
rect 84968 172760 84980 172812
rect 85032 172760 85044 172812
rect 85096 172760 85108 172812
rect 85160 172760 87806 172812
rect 83298 172738 87806 172760
rect 38 172268 3902 172290
rect 38 172216 2916 172268
rect 2968 172216 2980 172268
rect 3032 172216 3044 172268
rect 3096 172216 3108 172268
rect 3160 172216 3902 172268
rect 38 172194 3902 172216
rect 83298 172268 87806 172290
rect 83298 172216 86916 172268
rect 86968 172216 86980 172268
rect 87032 172216 87044 172268
rect 87096 172216 87108 172268
rect 87160 172216 87806 172268
rect 83298 172194 87806 172216
rect 38 171724 3902 171746
rect 38 171672 916 171724
rect 968 171672 980 171724
rect 1032 171672 1044 171724
rect 1096 171672 1108 171724
rect 1160 171672 3902 171724
rect 38 171650 3902 171672
rect 83298 171724 87806 171746
rect 83298 171672 84916 171724
rect 84968 171672 84980 171724
rect 85032 171672 85044 171724
rect 85096 171672 85108 171724
rect 85160 171672 87806 171724
rect 83298 171650 87806 171672
rect 38 171180 3902 171202
rect 38 171128 2916 171180
rect 2968 171128 2980 171180
rect 3032 171128 3044 171180
rect 3096 171128 3108 171180
rect 3160 171128 3902 171180
rect 38 171106 3902 171128
rect 83298 171180 87806 171202
rect 83298 171128 86916 171180
rect 86968 171128 86980 171180
rect 87032 171128 87044 171180
rect 87096 171128 87108 171180
rect 87160 171128 87806 171180
rect 83298 171106 87806 171128
rect 84324 171026 84330 171078
rect 84382 171066 84388 171078
rect 84784 171066 84790 171078
rect 84382 171038 84790 171066
rect 84382 171026 84388 171038
rect 84784 171026 84790 171038
rect 84842 171026 84848 171078
rect 38 170636 3902 170658
rect 38 170584 916 170636
rect 968 170584 980 170636
rect 1032 170584 1044 170636
rect 1096 170584 1108 170636
rect 1160 170584 3902 170636
rect 38 170562 3902 170584
rect 83298 170636 87806 170658
rect 83298 170584 84916 170636
rect 84968 170584 84980 170636
rect 85032 170584 85044 170636
rect 85096 170584 85108 170636
rect 85160 170584 87806 170636
rect 83298 170562 87806 170584
rect 38 170092 3902 170114
rect 38 170040 2916 170092
rect 2968 170040 2980 170092
rect 3032 170040 3044 170092
rect 3096 170040 3108 170092
rect 3160 170040 3902 170092
rect 38 170018 3902 170040
rect 83298 170092 87806 170114
rect 83298 170040 86916 170092
rect 86968 170040 86980 170092
rect 87032 170040 87044 170092
rect 87096 170040 87108 170092
rect 87160 170040 87806 170092
rect 83298 170018 87806 170040
rect 38 169548 3902 169570
rect 38 169496 916 169548
rect 968 169496 980 169548
rect 1032 169496 1044 169548
rect 1096 169496 1108 169548
rect 1160 169496 3902 169548
rect 38 169474 3902 169496
rect 83298 169548 87806 169570
rect 83298 169496 84916 169548
rect 84968 169496 84980 169548
rect 85032 169496 85044 169548
rect 85096 169496 85108 169548
rect 85160 169496 87806 169548
rect 83298 169474 87806 169496
rect 38 169004 3902 169026
rect 38 168952 2916 169004
rect 2968 168952 2980 169004
rect 3032 168952 3044 169004
rect 3096 168952 3108 169004
rect 3160 168952 3902 169004
rect 38 168930 3902 168952
rect 83298 169004 87806 169026
rect 83298 168952 86916 169004
rect 86968 168952 86980 169004
rect 87032 168952 87044 169004
rect 87096 168952 87108 169004
rect 87160 168952 87806 169004
rect 83298 168930 87806 168952
rect 38 168460 3902 168482
rect 38 168408 916 168460
rect 968 168408 980 168460
rect 1032 168408 1044 168460
rect 1096 168408 1108 168460
rect 1160 168408 3902 168460
rect 38 168386 3902 168408
rect 83298 168460 87806 168482
rect 83298 168408 84916 168460
rect 84968 168408 84980 168460
rect 85032 168408 85044 168460
rect 85096 168408 85108 168460
rect 85160 168408 87806 168460
rect 83298 168386 87806 168408
rect 38 167916 3902 167938
rect 38 167864 2916 167916
rect 2968 167864 2980 167916
rect 3032 167864 3044 167916
rect 3096 167864 3108 167916
rect 3160 167864 3902 167916
rect 38 167842 3902 167864
rect 83298 167916 87806 167938
rect 83298 167864 86916 167916
rect 86968 167864 86980 167916
rect 87032 167864 87044 167916
rect 87096 167864 87108 167916
rect 87160 167864 87806 167916
rect 83298 167842 87806 167864
rect 38 167372 3902 167394
rect 38 167320 916 167372
rect 968 167320 980 167372
rect 1032 167320 1044 167372
rect 1096 167320 1108 167372
rect 1160 167320 3902 167372
rect 38 167298 3902 167320
rect 83298 167372 87806 167394
rect 83298 167320 84916 167372
rect 84968 167320 84980 167372
rect 85032 167320 85044 167372
rect 85096 167320 85108 167372
rect 85160 167320 87806 167372
rect 83298 167298 87806 167320
rect 38 166828 3902 166850
rect 38 166776 2916 166828
rect 2968 166776 2980 166828
rect 3032 166776 3044 166828
rect 3096 166776 3108 166828
rect 3160 166776 3902 166828
rect 38 166754 3902 166776
rect 83298 166828 87806 166850
rect 83298 166776 86916 166828
rect 86968 166776 86980 166828
rect 87032 166776 87044 166828
rect 87096 166776 87108 166828
rect 87160 166776 87806 166828
rect 83298 166754 87806 166776
rect 38 166284 3902 166306
rect 38 166232 916 166284
rect 968 166232 980 166284
rect 1032 166232 1044 166284
rect 1096 166232 1108 166284
rect 1160 166232 3902 166284
rect 38 166210 3902 166232
rect 83298 166284 87806 166306
rect 83298 166232 84916 166284
rect 84968 166232 84980 166284
rect 85032 166232 85044 166284
rect 85096 166232 85108 166284
rect 85160 166232 87806 166284
rect 83298 166210 87806 166232
rect 38 165740 3902 165762
rect 38 165688 2916 165740
rect 2968 165688 2980 165740
rect 3032 165688 3044 165740
rect 3096 165688 3108 165740
rect 3160 165688 3902 165740
rect 38 165666 3902 165688
rect 83298 165740 87806 165762
rect 83298 165688 86916 165740
rect 86968 165688 86980 165740
rect 87032 165688 87044 165740
rect 87096 165688 87108 165740
rect 87160 165688 87806 165740
rect 83298 165666 87806 165688
rect 38 165196 3902 165218
rect 38 165144 916 165196
rect 968 165144 980 165196
rect 1032 165144 1044 165196
rect 1096 165144 1108 165196
rect 1160 165144 3902 165196
rect 38 165122 3902 165144
rect 83298 165196 87806 165218
rect 83298 165144 84916 165196
rect 84968 165144 84980 165196
rect 85032 165144 85044 165196
rect 85096 165144 85108 165196
rect 85160 165144 87806 165196
rect 83298 165122 87806 165144
rect 83956 164838 83962 164890
rect 84014 164878 84020 164890
rect 84416 164878 84422 164890
rect 84014 164850 84422 164878
rect 84014 164838 84020 164850
rect 84416 164838 84422 164850
rect 84474 164838 84480 164890
rect 84232 164770 84238 164822
rect 84290 164770 84296 164822
rect 3732 164702 3738 164754
rect 3790 164742 3796 164754
rect 4011 164745 4069 164751
rect 4011 164742 4023 164745
rect 3790 164714 4023 164742
rect 3790 164702 3796 164714
rect 4011 164711 4023 164714
rect 4057 164711 4069 164745
rect 84250 164742 84278 164770
rect 84600 164742 84606 164754
rect 84250 164714 84606 164742
rect 4011 164705 4069 164711
rect 84600 164702 84606 164714
rect 84658 164702 84664 164754
rect 38 164652 3902 164674
rect 38 164600 2916 164652
rect 2968 164600 2980 164652
rect 3032 164600 3044 164652
rect 3096 164600 3108 164652
rect 3160 164600 3902 164652
rect 38 164578 3902 164600
rect 83298 164652 87806 164674
rect 83298 164600 86916 164652
rect 86968 164600 86980 164652
rect 87032 164600 87044 164652
rect 87096 164600 87108 164652
rect 87160 164600 87806 164652
rect 83298 164578 87806 164600
rect 3732 164498 3738 164550
rect 3790 164538 3796 164550
rect 4011 164541 4069 164547
rect 4011 164538 4023 164541
rect 3790 164510 4023 164538
rect 3790 164498 3796 164510
rect 4011 164507 4023 164510
rect 4057 164507 4069 164541
rect 4011 164501 4069 164507
rect 83956 164498 83962 164550
rect 84014 164538 84020 164550
rect 84232 164538 84238 164550
rect 84014 164510 84238 164538
rect 84014 164498 84020 164510
rect 84232 164498 84238 164510
rect 84290 164498 84296 164550
rect 84324 164498 84330 164550
rect 84382 164538 84388 164550
rect 85152 164538 85158 164550
rect 84382 164510 85158 164538
rect 84382 164498 84388 164510
rect 85152 164498 85158 164510
rect 85210 164498 85216 164550
rect 38 164108 3902 164130
rect 38 164056 916 164108
rect 968 164056 980 164108
rect 1032 164056 1044 164108
rect 1096 164056 1108 164108
rect 1160 164056 3902 164108
rect 38 164034 3902 164056
rect 83298 164108 87806 164130
rect 83298 164056 84916 164108
rect 84968 164056 84980 164108
rect 85032 164056 85044 164108
rect 85096 164056 85108 164108
rect 85160 164056 87806 164108
rect 83298 164034 87806 164056
rect 81748 163886 81754 163938
rect 81806 163926 81812 163938
rect 85152 163926 85158 163938
rect 81806 163898 85158 163926
rect 81806 163886 81812 163898
rect 85152 163886 85158 163898
rect 85210 163886 85216 163938
rect 38 163564 3902 163586
rect 38 163512 2916 163564
rect 2968 163512 2980 163564
rect 3032 163512 3044 163564
rect 3096 163512 3108 163564
rect 3160 163512 3902 163564
rect 38 163490 3902 163512
rect 83298 163564 87806 163586
rect 83298 163512 86916 163564
rect 86968 163512 86980 163564
rect 87032 163512 87044 163564
rect 87096 163512 87108 163564
rect 87160 163512 87806 163564
rect 83298 163490 87806 163512
rect 38 163020 3902 163042
rect 38 162968 916 163020
rect 968 162968 980 163020
rect 1032 162968 1044 163020
rect 1096 162968 1108 163020
rect 1160 162968 3902 163020
rect 38 162946 3902 162968
rect 83298 163020 87806 163042
rect 83298 162968 84916 163020
rect 84968 162968 84980 163020
rect 85032 162968 85044 163020
rect 85096 162968 85108 163020
rect 85160 162968 87806 163020
rect 83298 162946 87806 162968
rect 81840 162798 81846 162850
rect 81898 162838 81904 162850
rect 84324 162838 84330 162850
rect 81898 162810 84330 162838
rect 81898 162798 81904 162810
rect 84324 162798 84330 162810
rect 84382 162798 84388 162850
rect 38 162476 3902 162498
rect 38 162424 2916 162476
rect 2968 162424 2980 162476
rect 3032 162424 3044 162476
rect 3096 162424 3108 162476
rect 3160 162424 3902 162476
rect 38 162402 3902 162424
rect 83298 162476 87806 162498
rect 83298 162424 86916 162476
rect 86968 162424 86980 162476
rect 87032 162424 87044 162476
rect 87096 162424 87108 162476
rect 87160 162424 87806 162476
rect 83298 162402 87806 162424
rect 1892 162118 1898 162170
rect 1950 162158 1956 162170
rect 2260 162158 2266 162170
rect 1950 162130 2266 162158
rect 1950 162118 1956 162130
rect 2260 162118 2266 162130
rect 2318 162118 2324 162170
rect 1892 161982 1898 162034
rect 1950 162022 1956 162034
rect 2260 162022 2266 162034
rect 1950 161994 2266 162022
rect 1950 161982 1956 161994
rect 2260 161982 2266 161994
rect 2318 161982 2324 162034
rect 38 161932 3902 161954
rect 38 161880 916 161932
rect 968 161880 980 161932
rect 1032 161880 1044 161932
rect 1096 161880 1108 161932
rect 1160 161880 3902 161932
rect 38 161858 3902 161880
rect 83298 161932 87806 161954
rect 83298 161880 84916 161932
rect 84968 161880 84980 161932
rect 85032 161880 85044 161932
rect 85096 161880 85108 161932
rect 85160 161880 87806 161932
rect 83298 161858 87806 161880
rect 84324 161778 84330 161830
rect 84382 161818 84388 161830
rect 84600 161818 84606 161830
rect 84382 161790 84606 161818
rect 84382 161778 84388 161790
rect 84600 161778 84606 161790
rect 84658 161778 84664 161830
rect 38 161388 3902 161410
rect 38 161336 2916 161388
rect 2968 161336 2980 161388
rect 3032 161336 3044 161388
rect 3096 161336 3108 161388
rect 3160 161336 3902 161388
rect 38 161314 3902 161336
rect 83298 161388 87806 161410
rect 83298 161336 86916 161388
rect 86968 161336 86980 161388
rect 87032 161336 87044 161388
rect 87096 161336 87108 161388
rect 87160 161336 87806 161388
rect 83298 161314 87806 161336
rect 38 160844 3902 160866
rect 38 160792 916 160844
rect 968 160792 980 160844
rect 1032 160792 1044 160844
rect 1096 160792 1108 160844
rect 1160 160792 3902 160844
rect 38 160770 3902 160792
rect 83298 160844 87806 160866
rect 83298 160792 84916 160844
rect 84968 160792 84980 160844
rect 85032 160792 85044 160844
rect 85096 160792 85108 160844
rect 85160 160792 87806 160844
rect 83298 160770 87806 160792
rect 82576 160690 82582 160742
rect 82634 160730 82640 160742
rect 84600 160730 84606 160742
rect 82634 160702 84606 160730
rect 82634 160690 82640 160702
rect 84600 160690 84606 160702
rect 84658 160690 84664 160742
rect 84416 160622 84422 160674
rect 84474 160662 84480 160674
rect 85336 160662 85342 160674
rect 84474 160634 85342 160662
rect 84474 160622 84480 160634
rect 85336 160622 85342 160634
rect 85394 160622 85400 160674
rect 38 160300 3902 160322
rect 38 160248 2916 160300
rect 2968 160248 2980 160300
rect 3032 160248 3044 160300
rect 3096 160248 3108 160300
rect 3160 160248 3902 160300
rect 38 160226 3902 160248
rect 83298 160300 87806 160322
rect 83298 160248 86916 160300
rect 86968 160248 86980 160300
rect 87032 160248 87044 160300
rect 87096 160248 87108 160300
rect 87160 160248 87806 160300
rect 83298 160226 87806 160248
rect 84508 160146 84514 160198
rect 84566 160146 84572 160198
rect 84526 159994 84554 160146
rect 84508 159942 84514 159994
rect 84566 159942 84572 159994
rect 38 159756 3902 159778
rect 38 159704 916 159756
rect 968 159704 980 159756
rect 1032 159704 1044 159756
rect 1096 159704 1108 159756
rect 1160 159704 3902 159756
rect 38 159682 3902 159704
rect 83298 159756 87806 159778
rect 83298 159704 84916 159756
rect 84968 159704 84980 159756
rect 85032 159704 85044 159756
rect 85096 159704 85108 159756
rect 85160 159704 87806 159756
rect 83298 159682 87806 159704
rect 38 159212 3902 159234
rect 38 159160 2916 159212
rect 2968 159160 2980 159212
rect 3032 159160 3044 159212
rect 3096 159160 3108 159212
rect 3160 159160 3902 159212
rect 38 159138 3902 159160
rect 83298 159212 87806 159234
rect 83298 159160 86916 159212
rect 86968 159160 86980 159212
rect 87032 159160 87044 159212
rect 87096 159160 87108 159212
rect 87160 159160 87806 159212
rect 83298 159138 87806 159160
rect 38 158668 3902 158690
rect 38 158616 916 158668
rect 968 158616 980 158668
rect 1032 158616 1044 158668
rect 1096 158616 1108 158668
rect 1160 158616 3902 158668
rect 38 158594 3902 158616
rect 83298 158668 87806 158690
rect 83298 158616 84916 158668
rect 84968 158616 84980 158668
rect 85032 158616 85044 158668
rect 85096 158616 85108 158668
rect 85160 158616 87806 158668
rect 83298 158594 87806 158616
rect 38 158124 3902 158146
rect 38 158072 2916 158124
rect 2968 158072 2980 158124
rect 3032 158072 3044 158124
rect 3096 158072 3108 158124
rect 3160 158072 3902 158124
rect 38 158050 3902 158072
rect 83298 158124 87806 158146
rect 83298 158072 86916 158124
rect 86968 158072 86980 158124
rect 87032 158072 87044 158124
rect 87096 158072 87108 158124
rect 87160 158072 87806 158124
rect 83298 158050 87806 158072
rect 38 157580 3902 157602
rect 38 157528 916 157580
rect 968 157528 980 157580
rect 1032 157528 1044 157580
rect 1096 157528 1108 157580
rect 1160 157528 3902 157580
rect 38 157506 3902 157528
rect 83298 157580 87806 157602
rect 83298 157528 84916 157580
rect 84968 157528 84980 157580
rect 85032 157528 85044 157580
rect 85096 157528 85108 157580
rect 85160 157528 87806 157580
rect 83298 157506 87806 157528
rect 38 157036 3902 157058
rect 38 156984 2916 157036
rect 2968 156984 2980 157036
rect 3032 156984 3044 157036
rect 3096 156984 3108 157036
rect 3160 156984 3902 157036
rect 38 156962 3902 156984
rect 83298 157036 87806 157058
rect 83298 156984 86916 157036
rect 86968 156984 86980 157036
rect 87032 156984 87044 157036
rect 87096 156984 87108 157036
rect 87160 156984 87806 157036
rect 83298 156962 87806 156984
rect 82484 156882 82490 156934
rect 82542 156922 82548 156934
rect 85060 156922 85066 156934
rect 82542 156894 85066 156922
rect 82542 156882 82548 156894
rect 85060 156882 85066 156894
rect 85118 156882 85124 156934
rect 38 156492 3902 156514
rect 38 156440 916 156492
rect 968 156440 980 156492
rect 1032 156440 1044 156492
rect 1096 156440 1108 156492
rect 1160 156440 3902 156492
rect 38 156418 3902 156440
rect 83298 156492 87806 156514
rect 83298 156440 84916 156492
rect 84968 156440 84980 156492
rect 85032 156440 85044 156492
rect 85096 156440 85108 156492
rect 85160 156440 87806 156492
rect 83298 156418 87806 156440
rect 38 155948 3902 155970
rect 38 155896 2916 155948
rect 2968 155896 2980 155948
rect 3032 155896 3044 155948
rect 3096 155896 3108 155948
rect 3160 155896 3902 155948
rect 38 155874 3902 155896
rect 83298 155948 87806 155970
rect 83298 155896 86916 155948
rect 86968 155896 86980 155948
rect 87032 155896 87044 155948
rect 87096 155896 87108 155948
rect 87160 155896 87806 155948
rect 83298 155874 87806 155896
rect 3456 155658 3462 155710
rect 3514 155698 3520 155710
rect 4011 155701 4069 155707
rect 4011 155698 4023 155701
rect 3514 155670 4023 155698
rect 3514 155658 3520 155670
rect 4011 155667 4023 155670
rect 4057 155667 4069 155701
rect 4011 155661 4069 155667
rect 3548 155590 3554 155642
rect 3606 155630 3612 155642
rect 3732 155630 3738 155642
rect 3606 155602 3738 155630
rect 3606 155590 3612 155602
rect 3732 155590 3738 155602
rect 3790 155590 3796 155642
rect 4008 155562 4014 155574
rect 3750 155534 4014 155562
rect 3750 155506 3778 155534
rect 4008 155522 4014 155534
rect 4066 155522 4072 155574
rect 3732 155454 3738 155506
rect 3790 155454 3796 155506
rect 38 155404 3902 155426
rect 38 155352 916 155404
rect 968 155352 980 155404
rect 1032 155352 1044 155404
rect 1096 155352 1108 155404
rect 1160 155352 3902 155404
rect 83298 155404 87806 155426
rect 4008 155358 4014 155370
rect 38 155330 3902 155352
rect 3969 155330 4014 155358
rect 4008 155318 4014 155330
rect 4066 155318 4072 155370
rect 83298 155352 84916 155404
rect 84968 155352 84980 155404
rect 85032 155352 85044 155404
rect 85096 155352 85108 155404
rect 85160 155352 87806 155404
rect 83298 155330 87806 155352
rect 38 154860 3902 154882
rect 38 154808 2916 154860
rect 2968 154808 2980 154860
rect 3032 154808 3044 154860
rect 3096 154808 3108 154860
rect 3160 154808 3902 154860
rect 38 154786 3902 154808
rect 83298 154860 87806 154882
rect 83298 154808 86916 154860
rect 86968 154808 86980 154860
rect 87032 154808 87044 154860
rect 87096 154808 87108 154860
rect 87160 154808 87806 154860
rect 83298 154786 87806 154808
rect 38 154316 3902 154338
rect 38 154264 916 154316
rect 968 154264 980 154316
rect 1032 154264 1044 154316
rect 1096 154264 1108 154316
rect 1160 154264 3902 154316
rect 38 154242 3902 154264
rect 83298 154316 87806 154338
rect 83298 154264 84916 154316
rect 84968 154264 84980 154316
rect 85032 154264 85044 154316
rect 85096 154264 85108 154316
rect 85160 154264 87806 154316
rect 83298 154242 87806 154264
rect 38 153772 3902 153794
rect 38 153720 2916 153772
rect 2968 153720 2980 153772
rect 3032 153720 3044 153772
rect 3096 153720 3108 153772
rect 3160 153720 3902 153772
rect 38 153698 3902 153720
rect 83298 153772 87806 153794
rect 83298 153720 86916 153772
rect 86968 153720 86980 153772
rect 87032 153720 87044 153772
rect 87096 153720 87108 153772
rect 87160 153720 87806 153772
rect 83298 153698 87806 153720
rect 38 153228 3902 153250
rect 38 153176 916 153228
rect 968 153176 980 153228
rect 1032 153176 1044 153228
rect 1096 153176 1108 153228
rect 1160 153176 3902 153228
rect 38 153154 3902 153176
rect 83298 153228 87806 153250
rect 83298 153176 84916 153228
rect 84968 153176 84980 153228
rect 85032 153176 85044 153228
rect 85096 153176 85108 153228
rect 85160 153176 87806 153228
rect 83298 153154 87806 153176
rect 1892 153074 1898 153126
rect 1950 153114 1956 153126
rect 2260 153114 2266 153126
rect 1950 153086 2266 153114
rect 1950 153074 1956 153086
rect 2260 153074 2266 153086
rect 2318 153074 2324 153126
rect 38 152684 3902 152706
rect 38 152632 2916 152684
rect 2968 152632 2980 152684
rect 3032 152632 3044 152684
rect 3096 152632 3108 152684
rect 3160 152632 3902 152684
rect 38 152610 3902 152632
rect 83298 152684 87806 152706
rect 83298 152632 86916 152684
rect 86968 152632 86980 152684
rect 87032 152632 87044 152684
rect 87096 152632 87108 152684
rect 87160 152632 87806 152684
rect 83298 152610 87806 152632
rect 38 152140 3902 152162
rect 38 152088 916 152140
rect 968 152088 980 152140
rect 1032 152088 1044 152140
rect 1096 152088 1108 152140
rect 1160 152088 3902 152140
rect 38 152066 3902 152088
rect 83298 152140 87806 152162
rect 83298 152088 84916 152140
rect 84968 152088 84980 152140
rect 85032 152088 85044 152140
rect 85096 152088 85108 152140
rect 85160 152088 87806 152140
rect 83298 152066 87806 152088
rect 3456 151782 3462 151834
rect 3514 151822 3520 151834
rect 5572 151822 5578 151834
rect 3514 151794 5578 151822
rect 3514 151782 3520 151794
rect 5572 151782 5578 151794
rect 5630 151782 5636 151834
rect 38 151596 3902 151618
rect 38 151544 2916 151596
rect 2968 151544 2980 151596
rect 3032 151544 3044 151596
rect 3096 151544 3108 151596
rect 3160 151544 3902 151596
rect 38 151522 3902 151544
rect 83298 151596 87806 151618
rect 83298 151544 86916 151596
rect 86968 151544 86980 151596
rect 87032 151544 87044 151596
rect 87096 151544 87108 151596
rect 87160 151544 87806 151596
rect 83298 151522 87806 151544
rect 38 151052 3902 151074
rect 38 151000 916 151052
rect 968 151000 980 151052
rect 1032 151000 1044 151052
rect 1096 151000 1108 151052
rect 1160 151000 3902 151052
rect 38 150978 3902 151000
rect 83298 151052 87806 151074
rect 83298 151000 84916 151052
rect 84968 151000 84980 151052
rect 85032 151000 85044 151052
rect 85096 151000 85108 151052
rect 85160 151000 87806 151052
rect 83298 150978 87806 151000
rect 38 150508 3902 150530
rect 38 150456 2916 150508
rect 2968 150456 2980 150508
rect 3032 150456 3044 150508
rect 3096 150456 3108 150508
rect 3160 150456 3902 150508
rect 38 150434 3902 150456
rect 83298 150508 87806 150530
rect 83298 150456 86916 150508
rect 86968 150456 86980 150508
rect 87032 150456 87044 150508
rect 87096 150456 87108 150508
rect 87160 150456 87806 150508
rect 83298 150434 87806 150456
rect 82392 150082 82398 150134
rect 82450 150122 82456 150134
rect 83956 150122 83962 150134
rect 82450 150094 83962 150122
rect 82450 150082 82456 150094
rect 83956 150082 83962 150094
rect 84014 150082 84020 150134
rect 38 149964 3902 149986
rect 38 149912 916 149964
rect 968 149912 980 149964
rect 1032 149912 1044 149964
rect 1096 149912 1108 149964
rect 1160 149912 3902 149964
rect 38 149890 3902 149912
rect 83298 149964 87806 149986
rect 83298 149912 84916 149964
rect 84968 149912 84980 149964
rect 85032 149912 85044 149964
rect 85096 149912 85108 149964
rect 85160 149912 87806 149964
rect 83298 149890 87806 149912
rect 38 149420 3902 149442
rect 38 149368 2916 149420
rect 2968 149368 2980 149420
rect 3032 149368 3044 149420
rect 3096 149368 3108 149420
rect 3160 149368 3902 149420
rect 38 149346 3902 149368
rect 83298 149420 87806 149442
rect 83298 149368 86916 149420
rect 86968 149368 86980 149420
rect 87032 149368 87044 149420
rect 87096 149368 87108 149420
rect 87160 149368 87806 149420
rect 83298 149346 87806 149368
rect 82300 149130 82306 149182
rect 82358 149170 82364 149182
rect 83956 149170 83962 149182
rect 82358 149142 83962 149170
rect 82358 149130 82364 149142
rect 83956 149130 83962 149142
rect 84014 149130 84020 149182
rect 38 148876 3902 148898
rect 38 148824 916 148876
rect 968 148824 980 148876
rect 1032 148824 1044 148876
rect 1096 148824 1108 148876
rect 1160 148824 3902 148876
rect 38 148802 3902 148824
rect 83298 148876 87806 148898
rect 83298 148824 84916 148876
rect 84968 148824 84980 148876
rect 85032 148824 85044 148876
rect 85096 148824 85108 148876
rect 85160 148824 87806 148876
rect 83298 148802 87806 148824
rect 38 148332 3902 148354
rect 38 148280 2916 148332
rect 2968 148280 2980 148332
rect 3032 148280 3044 148332
rect 3096 148280 3108 148332
rect 3160 148280 3902 148332
rect 38 148258 3902 148280
rect 83298 148332 87806 148354
rect 83298 148280 86916 148332
rect 86968 148280 86980 148332
rect 87032 148280 87044 148332
rect 87096 148280 87108 148332
rect 87160 148280 87806 148332
rect 83298 148258 87806 148280
rect 82208 147838 82214 147890
rect 82266 147878 82272 147890
rect 83956 147878 83962 147890
rect 82266 147850 83962 147878
rect 82266 147838 82272 147850
rect 83956 147838 83962 147850
rect 84014 147838 84020 147890
rect 38 147788 3902 147810
rect 38 147736 916 147788
rect 968 147736 980 147788
rect 1032 147736 1044 147788
rect 1096 147736 1108 147788
rect 1160 147736 3902 147788
rect 38 147714 3902 147736
rect 83298 147788 87806 147810
rect 83298 147736 84916 147788
rect 84968 147736 84980 147788
rect 85032 147736 85044 147788
rect 85096 147736 85108 147788
rect 85160 147736 87806 147788
rect 83298 147714 87806 147736
rect 38 147244 3902 147266
rect 38 147192 2916 147244
rect 2968 147192 2980 147244
rect 3032 147192 3044 147244
rect 3096 147192 3108 147244
rect 3160 147192 3902 147244
rect 38 147170 3902 147192
rect 83298 147244 87806 147266
rect 83298 147192 86916 147244
rect 86968 147192 86980 147244
rect 87032 147192 87044 147244
rect 87096 147192 87108 147244
rect 87160 147192 87806 147244
rect 83298 147170 87806 147192
rect 4008 146858 4014 146870
rect 3969 146830 4014 146858
rect 4008 146818 4014 146830
rect 4066 146818 4072 146870
rect 3548 146750 3554 146802
rect 3606 146790 3612 146802
rect 4103 146793 4161 146799
rect 4103 146790 4115 146793
rect 3606 146762 4115 146790
rect 3606 146750 3612 146762
rect 4103 146759 4115 146762
rect 4149 146759 4161 146793
rect 4103 146753 4161 146759
rect 38 146700 3902 146722
rect 38 146648 916 146700
rect 968 146648 980 146700
rect 1032 146648 1044 146700
rect 1096 146648 1108 146700
rect 1160 146648 3902 146700
rect 38 146626 3902 146648
rect 83298 146700 87806 146722
rect 83298 146648 84916 146700
rect 84968 146648 84980 146700
rect 85032 146648 85044 146700
rect 85096 146648 85108 146700
rect 85160 146648 87806 146700
rect 83298 146626 87806 146648
rect 82116 146546 82122 146598
rect 82174 146586 82180 146598
rect 83956 146586 83962 146598
rect 82174 146558 83962 146586
rect 82174 146546 82180 146558
rect 83956 146546 83962 146558
rect 84014 146546 84020 146598
rect 38 146156 3902 146178
rect 38 146104 2916 146156
rect 2968 146104 2980 146156
rect 3032 146104 3044 146156
rect 3096 146104 3108 146156
rect 3160 146104 3902 146156
rect 38 146082 3902 146104
rect 83298 146156 87806 146178
rect 83298 146104 86916 146156
rect 86968 146104 86980 146156
rect 87032 146104 87044 146156
rect 87096 146104 87108 146156
rect 87160 146104 87806 146156
rect 83298 146082 87806 146104
rect 1892 145934 1898 145986
rect 1950 145974 1956 145986
rect 2260 145974 2266 145986
rect 1950 145946 2266 145974
rect 1950 145934 1956 145946
rect 2260 145934 2266 145946
rect 2318 145934 2324 145986
rect 38 145612 3902 145634
rect 38 145560 916 145612
rect 968 145560 980 145612
rect 1032 145560 1044 145612
rect 1096 145560 1108 145612
rect 1160 145560 3902 145612
rect 38 145538 3902 145560
rect 83298 145612 87806 145634
rect 83298 145560 84916 145612
rect 84968 145560 84980 145612
rect 85032 145560 85044 145612
rect 85096 145560 85108 145612
rect 85160 145560 87806 145612
rect 83298 145538 87806 145560
rect 81932 145254 81938 145306
rect 81990 145294 81996 145306
rect 83956 145294 83962 145306
rect 81990 145266 83962 145294
rect 81990 145254 81996 145266
rect 83956 145254 83962 145266
rect 84014 145254 84020 145306
rect 38 145068 3902 145090
rect 38 145016 2916 145068
rect 2968 145016 2980 145068
rect 3032 145016 3044 145068
rect 3096 145016 3108 145068
rect 3160 145016 3902 145068
rect 38 144994 3902 145016
rect 83298 145068 87806 145090
rect 83298 145016 86916 145068
rect 86968 145016 86980 145068
rect 87032 145016 87044 145068
rect 87096 145016 87108 145068
rect 87160 145016 87806 145068
rect 83298 144994 87806 145016
rect 38 144524 3902 144546
rect 38 144472 916 144524
rect 968 144472 980 144524
rect 1032 144472 1044 144524
rect 1096 144472 1108 144524
rect 1160 144472 3902 144524
rect 38 144450 3902 144472
rect 83298 144524 87806 144546
rect 83298 144472 84916 144524
rect 84968 144472 84980 144524
rect 85032 144472 85044 144524
rect 85096 144472 85108 144524
rect 85160 144472 87806 144524
rect 83298 144450 87806 144472
rect 38 143980 3902 144002
rect 38 143928 2916 143980
rect 2968 143928 2980 143980
rect 3032 143928 3044 143980
rect 3096 143928 3108 143980
rect 3160 143928 3902 143980
rect 38 143906 3902 143928
rect 83298 143980 87806 144002
rect 83298 143928 86916 143980
rect 86968 143928 86980 143980
rect 87032 143928 87044 143980
rect 87096 143928 87108 143980
rect 87160 143928 87806 143980
rect 83298 143906 87806 143928
rect 82024 143826 82030 143878
rect 82082 143866 82088 143878
rect 84232 143866 84238 143878
rect 82082 143838 84238 143866
rect 82082 143826 82088 143838
rect 84232 143826 84238 143838
rect 84290 143826 84296 143878
rect 38 143436 3902 143458
rect 38 143384 916 143436
rect 968 143384 980 143436
rect 1032 143384 1044 143436
rect 1096 143384 1108 143436
rect 1160 143384 3902 143436
rect 38 143362 3902 143384
rect 83298 143436 87806 143458
rect 83298 143384 84916 143436
rect 84968 143384 84980 143436
rect 85032 143384 85044 143436
rect 85096 143384 85108 143436
rect 85160 143384 87806 143436
rect 83298 143362 87806 143384
rect 38 142892 3902 142914
rect 38 142840 2916 142892
rect 2968 142840 2980 142892
rect 3032 142840 3044 142892
rect 3096 142840 3108 142892
rect 3160 142840 3902 142892
rect 38 142818 3902 142840
rect 83298 142892 87806 142914
rect 83298 142840 86916 142892
rect 86968 142840 86980 142892
rect 87032 142840 87044 142892
rect 87096 142840 87108 142892
rect 87160 142840 87806 142892
rect 83298 142818 87806 142840
rect 38 142348 3902 142370
rect 38 142296 916 142348
rect 968 142296 980 142348
rect 1032 142296 1044 142348
rect 1096 142296 1108 142348
rect 1160 142296 3902 142348
rect 38 142274 3902 142296
rect 83298 142348 87806 142370
rect 83298 142296 84916 142348
rect 84968 142296 84980 142348
rect 85032 142296 85044 142348
rect 85096 142296 85108 142348
rect 85160 142296 87806 142348
rect 83298 142274 87806 142296
rect 38 141804 3902 141826
rect 38 141752 2916 141804
rect 2968 141752 2980 141804
rect 3032 141752 3044 141804
rect 3096 141752 3108 141804
rect 3160 141752 3902 141804
rect 38 141730 3902 141752
rect 83298 141804 87806 141826
rect 83298 141752 86916 141804
rect 86968 141752 86980 141804
rect 87032 141752 87044 141804
rect 87096 141752 87108 141804
rect 87160 141752 87806 141804
rect 83298 141730 87806 141752
rect 3732 141582 3738 141634
rect 3790 141622 3796 141634
rect 4103 141625 4161 141631
rect 4103 141622 4115 141625
rect 3790 141594 4115 141622
rect 3790 141582 3796 141594
rect 4103 141591 4115 141594
rect 4149 141591 4161 141625
rect 4103 141585 4161 141591
rect 1892 141514 1898 141566
rect 1950 141554 1956 141566
rect 2168 141554 2174 141566
rect 1950 141526 2174 141554
rect 1950 141514 1956 141526
rect 2168 141514 2174 141526
rect 2226 141514 2232 141566
rect 3548 141514 3554 141566
rect 3606 141554 3612 141566
rect 4011 141557 4069 141563
rect 4011 141554 4023 141557
rect 3606 141526 4023 141554
rect 3606 141514 3612 141526
rect 4011 141523 4023 141526
rect 4057 141523 4069 141557
rect 4011 141517 4069 141523
rect 38 141260 3902 141282
rect 38 141208 916 141260
rect 968 141208 980 141260
rect 1032 141208 1044 141260
rect 1096 141208 1108 141260
rect 1160 141208 3902 141260
rect 38 141186 3902 141208
rect 83298 141260 87806 141282
rect 83298 141208 84916 141260
rect 84968 141208 84980 141260
rect 85032 141208 85044 141260
rect 85096 141208 85108 141260
rect 85160 141208 87806 141260
rect 83298 141186 87806 141208
rect 38 140716 3902 140738
rect 38 140664 2916 140716
rect 2968 140664 2980 140716
rect 3032 140664 3044 140716
rect 3096 140664 3108 140716
rect 3160 140664 3902 140716
rect 38 140642 3902 140664
rect 83298 140716 87806 140738
rect 83298 140664 86916 140716
rect 86968 140664 86980 140716
rect 87032 140664 87044 140716
rect 87096 140664 87108 140716
rect 87160 140664 87806 140716
rect 83298 140642 87806 140664
rect 38 140172 3902 140194
rect 38 140120 916 140172
rect 968 140120 980 140172
rect 1032 140120 1044 140172
rect 1096 140120 1108 140172
rect 1160 140120 3902 140172
rect 38 140098 3902 140120
rect 83298 140172 87806 140194
rect 83298 140120 84916 140172
rect 84968 140120 84980 140172
rect 85032 140120 85044 140172
rect 85096 140120 85108 140172
rect 85160 140120 87806 140172
rect 83298 140098 87806 140120
rect 38 139628 3902 139650
rect 38 139576 2916 139628
rect 2968 139576 2980 139628
rect 3032 139576 3044 139628
rect 3096 139576 3108 139628
rect 3160 139576 3902 139628
rect 38 139554 3902 139576
rect 83298 139628 87806 139650
rect 83298 139576 86916 139628
rect 86968 139576 86980 139628
rect 87032 139576 87044 139628
rect 87096 139576 87108 139628
rect 87160 139576 87806 139628
rect 83298 139554 87806 139576
rect 38 139084 3902 139106
rect 38 139032 916 139084
rect 968 139032 980 139084
rect 1032 139032 1044 139084
rect 1096 139032 1108 139084
rect 1160 139032 3902 139084
rect 38 139010 3902 139032
rect 83298 139084 87806 139106
rect 83298 139032 84916 139084
rect 84968 139032 84980 139084
rect 85032 139032 85044 139084
rect 85096 139032 85108 139084
rect 85160 139032 87806 139084
rect 83298 139010 87806 139032
rect 38 138540 3902 138562
rect 38 138488 2916 138540
rect 2968 138488 2980 138540
rect 3032 138488 3044 138540
rect 3096 138488 3108 138540
rect 3160 138488 3902 138540
rect 38 138466 3902 138488
rect 83298 138540 87806 138562
rect 83298 138488 86916 138540
rect 86968 138488 86980 138540
rect 87032 138488 87044 138540
rect 87096 138488 87108 138540
rect 87160 138488 87806 138540
rect 83298 138466 87806 138488
rect 38 137996 3902 138018
rect 38 137944 916 137996
rect 968 137944 980 137996
rect 1032 137944 1044 137996
rect 1096 137944 1108 137996
rect 1160 137944 3902 137996
rect 38 137922 3902 137944
rect 83298 137996 87806 138018
rect 83298 137944 84916 137996
rect 84968 137944 84980 137996
rect 85032 137944 85044 137996
rect 85096 137944 85108 137996
rect 85160 137944 87806 137996
rect 83298 137922 87806 137944
rect 81932 137638 81938 137690
rect 81990 137678 81996 137690
rect 84232 137678 84238 137690
rect 81990 137650 84238 137678
rect 81990 137638 81996 137650
rect 84232 137638 84238 137650
rect 84290 137638 84296 137690
rect 38 137452 3902 137474
rect 38 137400 2916 137452
rect 2968 137400 2980 137452
rect 3032 137400 3044 137452
rect 3096 137400 3108 137452
rect 3160 137400 3902 137452
rect 38 137378 3902 137400
rect 83298 137452 87806 137474
rect 83298 137400 86916 137452
rect 86968 137400 86980 137452
rect 87032 137400 87044 137452
rect 87096 137400 87108 137452
rect 87160 137400 87806 137452
rect 83298 137378 87806 137400
rect 38 136908 3902 136930
rect 38 136856 916 136908
rect 968 136856 980 136908
rect 1032 136856 1044 136908
rect 1096 136856 1108 136908
rect 1160 136856 3902 136908
rect 38 136834 3902 136856
rect 83298 136908 87806 136930
rect 83298 136856 84916 136908
rect 84968 136856 84980 136908
rect 85032 136856 85044 136908
rect 85096 136856 85108 136908
rect 85160 136856 87806 136908
rect 83298 136834 87806 136856
rect 38 136364 3902 136386
rect 38 136312 2916 136364
rect 2968 136312 2980 136364
rect 3032 136312 3044 136364
rect 3096 136312 3108 136364
rect 3160 136312 3902 136364
rect 38 136290 3902 136312
rect 83298 136364 87806 136386
rect 83298 136312 86916 136364
rect 86968 136312 86980 136364
rect 87032 136312 87044 136364
rect 87096 136312 87108 136364
rect 87160 136312 87806 136364
rect 83298 136290 87806 136312
rect 38 135820 3902 135842
rect 38 135768 916 135820
rect 968 135768 980 135820
rect 1032 135768 1044 135820
rect 1096 135768 1108 135820
rect 1160 135768 3902 135820
rect 38 135746 3902 135768
rect 83298 135820 87806 135842
rect 83298 135768 84916 135820
rect 84968 135768 84980 135820
rect 85032 135768 85044 135820
rect 85096 135768 85108 135820
rect 85160 135768 87806 135820
rect 83298 135746 87806 135768
rect 38 135276 3902 135298
rect 38 135224 2916 135276
rect 2968 135224 2980 135276
rect 3032 135224 3044 135276
rect 3096 135224 3108 135276
rect 3160 135224 3902 135276
rect 38 135202 3902 135224
rect 83298 135276 87806 135298
rect 83298 135224 86916 135276
rect 86968 135224 86980 135276
rect 87032 135224 87044 135276
rect 87096 135224 87108 135276
rect 87160 135224 87806 135276
rect 83298 135202 87806 135224
rect 38 134732 3902 134754
rect 38 134680 916 134732
rect 968 134680 980 134732
rect 1032 134680 1044 134732
rect 1096 134680 1108 134732
rect 1160 134680 3902 134732
rect 38 134658 3902 134680
rect 83298 134732 87806 134754
rect 83298 134680 84916 134732
rect 84968 134680 84980 134732
rect 85032 134680 85044 134732
rect 85096 134680 85108 134732
rect 85160 134680 87806 134732
rect 83298 134658 87806 134680
rect 38 134188 3902 134210
rect 38 134136 2916 134188
rect 2968 134136 2980 134188
rect 3032 134136 3044 134188
rect 3096 134136 3108 134188
rect 3160 134136 3902 134188
rect 38 134114 3902 134136
rect 83298 134188 87806 134210
rect 83298 134136 86916 134188
rect 86968 134136 86980 134188
rect 87032 134136 87044 134188
rect 87096 134136 87108 134188
rect 87160 134136 87806 134188
rect 83298 134114 87806 134136
rect 1892 133694 1898 133746
rect 1950 133734 1956 133746
rect 2260 133734 2266 133746
rect 1950 133706 2266 133734
rect 1950 133694 1956 133706
rect 2260 133694 2266 133706
rect 2318 133694 2324 133746
rect 38 133644 3902 133666
rect 38 133592 916 133644
rect 968 133592 980 133644
rect 1032 133592 1044 133644
rect 1096 133592 1108 133644
rect 1160 133592 3902 133644
rect 38 133570 3902 133592
rect 83298 133644 87806 133666
rect 83298 133592 84916 133644
rect 84968 133592 84980 133644
rect 85032 133592 85044 133644
rect 85096 133592 85108 133644
rect 85160 133592 87806 133644
rect 83298 133570 87806 133592
rect 38 133100 3902 133122
rect 38 133048 2916 133100
rect 2968 133048 2980 133100
rect 3032 133048 3044 133100
rect 3096 133048 3108 133100
rect 3160 133048 3902 133100
rect 38 133026 3902 133048
rect 83298 133100 87806 133122
rect 83298 133048 86916 133100
rect 86968 133048 86980 133100
rect 87032 133048 87044 133100
rect 87096 133048 87108 133100
rect 87160 133048 87806 133100
rect 83298 133026 87806 133048
rect 38 132556 3902 132578
rect 38 132504 916 132556
rect 968 132504 980 132556
rect 1032 132504 1044 132556
rect 1096 132504 1108 132556
rect 1160 132504 3902 132556
rect 38 132482 3902 132504
rect 83298 132556 87806 132578
rect 83298 132504 84916 132556
rect 84968 132504 84980 132556
rect 85032 132504 85044 132556
rect 85096 132504 85108 132556
rect 85160 132504 87806 132556
rect 83298 132482 87806 132504
rect 38 132012 3902 132034
rect 38 131960 2916 132012
rect 2968 131960 2980 132012
rect 3032 131960 3044 132012
rect 3096 131960 3108 132012
rect 3160 131960 3902 132012
rect 38 131938 3902 131960
rect 83298 132012 87806 132034
rect 83298 131960 86916 132012
rect 86968 131960 86980 132012
rect 87032 131960 87044 132012
rect 87096 131960 87108 132012
rect 87160 131960 87806 132012
rect 83298 131938 87806 131960
rect 38 131468 3902 131490
rect 38 131416 916 131468
rect 968 131416 980 131468
rect 1032 131416 1044 131468
rect 1096 131416 1108 131468
rect 1160 131416 3902 131468
rect 38 131394 3902 131416
rect 83298 131468 87806 131490
rect 83298 131416 84916 131468
rect 84968 131416 84980 131468
rect 85032 131416 85044 131468
rect 85096 131416 85108 131468
rect 85160 131416 87806 131468
rect 83298 131394 87806 131416
rect 38 130924 3902 130946
rect 38 130872 2916 130924
rect 2968 130872 2980 130924
rect 3032 130872 3044 130924
rect 3096 130872 3108 130924
rect 3160 130872 3902 130924
rect 38 130850 3902 130872
rect 83298 130924 87806 130946
rect 83298 130872 86916 130924
rect 86968 130872 86980 130924
rect 87032 130872 87044 130924
rect 87096 130872 87108 130924
rect 87160 130872 87806 130924
rect 83298 130850 87806 130872
rect 38 130380 3902 130402
rect 38 130328 916 130380
rect 968 130328 980 130380
rect 1032 130328 1044 130380
rect 1096 130328 1108 130380
rect 1160 130328 3902 130380
rect 38 130306 3902 130328
rect 83298 130380 87806 130402
rect 83298 130328 84916 130380
rect 84968 130328 84980 130380
rect 85032 130328 85044 130380
rect 85096 130328 85108 130380
rect 85160 130328 87806 130380
rect 83298 130306 87806 130328
rect 83220 129886 83226 129938
rect 83278 129926 83284 129938
rect 84508 129926 84514 129938
rect 83278 129898 84514 129926
rect 83278 129886 83284 129898
rect 84508 129886 84514 129898
rect 84566 129886 84572 129938
rect 38 129836 3902 129858
rect 38 129784 2916 129836
rect 2968 129784 2980 129836
rect 3032 129784 3044 129836
rect 3096 129784 3108 129836
rect 3160 129784 3902 129836
rect 38 129762 3902 129784
rect 83298 129836 87806 129858
rect 83298 129784 86916 129836
rect 86968 129784 86980 129836
rect 87032 129784 87044 129836
rect 87096 129784 87108 129836
rect 87160 129784 87806 129836
rect 83298 129762 87806 129784
rect 38 129292 3902 129314
rect 38 129240 916 129292
rect 968 129240 980 129292
rect 1032 129240 1044 129292
rect 1096 129240 1108 129292
rect 1160 129240 3902 129292
rect 38 129218 3902 129240
rect 83298 129292 87806 129314
rect 83298 129240 84916 129292
rect 84968 129240 84980 129292
rect 85032 129240 85044 129292
rect 85096 129240 85108 129292
rect 85160 129240 87806 129292
rect 83298 129218 87806 129240
rect 3548 128798 3554 128850
rect 3606 128838 3612 128850
rect 4011 128841 4069 128847
rect 4011 128838 4023 128841
rect 3606 128810 4023 128838
rect 3606 128798 3612 128810
rect 4011 128807 4023 128810
rect 4057 128807 4069 128841
rect 4011 128801 4069 128807
rect 38 128748 3902 128770
rect 38 128696 2916 128748
rect 2968 128696 2980 128748
rect 3032 128696 3044 128748
rect 3096 128696 3108 128748
rect 3160 128696 3902 128748
rect 38 128674 3902 128696
rect 83298 128748 87806 128770
rect 83298 128696 86916 128748
rect 86968 128696 86980 128748
rect 87032 128696 87044 128748
rect 87096 128696 87108 128748
rect 87160 128696 87806 128748
rect 83298 128674 87806 128696
rect 3732 128594 3738 128646
rect 3790 128634 3796 128646
rect 4103 128637 4161 128643
rect 4103 128634 4115 128637
rect 3790 128606 4115 128634
rect 3790 128594 3796 128606
rect 4103 128603 4115 128606
rect 4149 128603 4161 128637
rect 4103 128597 4161 128603
rect 83128 128594 83134 128646
rect 83186 128634 83192 128646
rect 84416 128634 84422 128646
rect 83186 128606 84422 128634
rect 83186 128594 83192 128606
rect 84416 128594 84422 128606
rect 84474 128594 84480 128646
rect 38 128204 3902 128226
rect 38 128152 916 128204
rect 968 128152 980 128204
rect 1032 128152 1044 128204
rect 1096 128152 1108 128204
rect 1160 128152 3902 128204
rect 38 128130 3902 128152
rect 83298 128204 87806 128226
rect 83298 128152 84916 128204
rect 84968 128152 84980 128204
rect 85032 128152 85044 128204
rect 85096 128152 85108 128204
rect 85160 128152 87806 128204
rect 83298 128130 87806 128152
rect 38 127660 3902 127682
rect 38 127608 2916 127660
rect 2968 127608 2980 127660
rect 3032 127608 3044 127660
rect 3096 127608 3108 127660
rect 3160 127608 3902 127660
rect 38 127586 3902 127608
rect 83298 127660 87806 127682
rect 83298 127608 86916 127660
rect 86968 127608 86980 127660
rect 87032 127608 87044 127660
rect 87096 127608 87108 127660
rect 87160 127608 87806 127660
rect 83298 127586 87806 127608
rect 83404 127370 83410 127422
rect 83462 127410 83468 127422
rect 84232 127410 84238 127422
rect 83462 127382 84238 127410
rect 83462 127370 83468 127382
rect 84232 127370 84238 127382
rect 84290 127370 84296 127422
rect 38 127116 3902 127138
rect 38 127064 916 127116
rect 968 127064 980 127116
rect 1032 127064 1044 127116
rect 1096 127064 1108 127116
rect 1160 127064 3902 127116
rect 38 127042 3902 127064
rect 83298 127116 87806 127138
rect 83298 127064 84916 127116
rect 84968 127064 84980 127116
rect 85032 127064 85044 127116
rect 85096 127064 85108 127116
rect 85160 127064 87806 127116
rect 83298 127042 87806 127064
rect 38 126572 3902 126594
rect 38 126520 2916 126572
rect 2968 126520 2980 126572
rect 3032 126520 3044 126572
rect 3096 126520 3108 126572
rect 3160 126520 3902 126572
rect 38 126498 3902 126520
rect 83298 126572 87806 126594
rect 83298 126520 86916 126572
rect 86968 126520 86980 126572
rect 87032 126520 87044 126572
rect 87096 126520 87108 126572
rect 87160 126520 87806 126572
rect 83298 126498 87806 126520
rect 38 126028 3902 126050
rect 38 125976 916 126028
rect 968 125976 980 126028
rect 1032 125976 1044 126028
rect 1096 125976 1108 126028
rect 1160 125976 3902 126028
rect 38 125954 3902 125976
rect 83298 126028 87806 126050
rect 83298 125976 84916 126028
rect 84968 125976 84980 126028
rect 85032 125976 85044 126028
rect 85096 125976 85108 126028
rect 85160 125976 87806 126028
rect 83298 125954 87806 125976
rect 38 125484 3902 125506
rect 38 125432 2916 125484
rect 2968 125432 2980 125484
rect 3032 125432 3044 125484
rect 3096 125432 3108 125484
rect 3160 125432 3902 125484
rect 38 125410 3902 125432
rect 83298 125484 87806 125506
rect 83298 125432 86916 125484
rect 86968 125432 86980 125484
rect 87032 125432 87044 125484
rect 87096 125432 87108 125484
rect 87160 125432 87806 125484
rect 83298 125410 87806 125432
rect 38 124940 3902 124962
rect 38 124888 916 124940
rect 968 124888 980 124940
rect 1032 124888 1044 124940
rect 1096 124888 1108 124940
rect 1160 124888 3902 124940
rect 38 124866 3902 124888
rect 83298 124940 87806 124962
rect 83298 124888 84916 124940
rect 84968 124888 84980 124940
rect 85032 124888 85044 124940
rect 85096 124888 85108 124940
rect 85160 124888 87806 124940
rect 83298 124866 87806 124888
rect 1892 124718 1898 124770
rect 1950 124758 1956 124770
rect 2168 124758 2174 124770
rect 1950 124730 2174 124758
rect 1950 124718 1956 124730
rect 2168 124718 2174 124730
rect 2226 124718 2232 124770
rect 82024 124718 82030 124770
rect 82082 124758 82088 124770
rect 84232 124758 84238 124770
rect 82082 124730 84238 124758
rect 82082 124718 82088 124730
rect 84232 124718 84238 124730
rect 84290 124718 84296 124770
rect 38 124396 3902 124418
rect 38 124344 2916 124396
rect 2968 124344 2980 124396
rect 3032 124344 3044 124396
rect 3096 124344 3108 124396
rect 3160 124344 3902 124396
rect 38 124322 3902 124344
rect 83298 124396 87806 124418
rect 83298 124344 86916 124396
rect 86968 124344 86980 124396
rect 87032 124344 87044 124396
rect 87096 124344 87108 124396
rect 87160 124344 87806 124396
rect 83298 124322 87806 124344
rect 82116 123902 82122 123954
rect 82174 123942 82180 123954
rect 84416 123942 84422 123954
rect 82174 123914 84422 123942
rect 82174 123902 82180 123914
rect 84416 123902 84422 123914
rect 84474 123902 84480 123954
rect 38 123852 3902 123874
rect 38 123800 916 123852
rect 968 123800 980 123852
rect 1032 123800 1044 123852
rect 1096 123800 1108 123852
rect 1160 123800 3902 123852
rect 38 123778 3902 123800
rect 83298 123852 87806 123874
rect 83298 123800 84916 123852
rect 84968 123800 84980 123852
rect 85032 123800 85044 123852
rect 85096 123800 85108 123852
rect 85160 123800 87806 123852
rect 83298 123778 87806 123800
rect 3732 123494 3738 123546
rect 3790 123534 3796 123546
rect 4103 123537 4161 123543
rect 4103 123534 4115 123537
rect 3790 123506 4115 123534
rect 3790 123494 3796 123506
rect 4103 123503 4115 123506
rect 4149 123503 4161 123537
rect 4103 123497 4161 123503
rect 3548 123426 3554 123478
rect 3606 123466 3612 123478
rect 4011 123469 4069 123475
rect 4011 123466 4023 123469
rect 3606 123438 4023 123466
rect 3606 123426 3612 123438
rect 4011 123435 4023 123438
rect 4057 123435 4069 123469
rect 4011 123429 4069 123435
rect 38 123308 3902 123330
rect 38 123256 2916 123308
rect 2968 123256 2980 123308
rect 3032 123256 3044 123308
rect 3096 123256 3108 123308
rect 3160 123256 3902 123308
rect 38 123234 3902 123256
rect 83298 123308 87806 123330
rect 83298 123256 86916 123308
rect 86968 123256 86980 123308
rect 87032 123256 87044 123308
rect 87096 123256 87108 123308
rect 87160 123256 87806 123308
rect 83298 123234 87806 123256
rect 38 122764 3902 122786
rect 38 122712 916 122764
rect 968 122712 980 122764
rect 1032 122712 1044 122764
rect 1096 122712 1108 122764
rect 1160 122712 3902 122764
rect 38 122690 3902 122712
rect 83298 122764 87806 122786
rect 83298 122712 84916 122764
rect 84968 122712 84980 122764
rect 85032 122712 85044 122764
rect 85096 122712 85108 122764
rect 85160 122712 87806 122764
rect 83298 122690 87806 122712
rect 38 122220 3902 122242
rect 38 122168 2916 122220
rect 2968 122168 2980 122220
rect 3032 122168 3044 122220
rect 3096 122168 3108 122220
rect 3160 122168 3902 122220
rect 38 122146 3902 122168
rect 83298 122220 87806 122242
rect 83298 122168 86916 122220
rect 86968 122168 86980 122220
rect 87032 122168 87044 122220
rect 87096 122168 87108 122220
rect 87160 122168 87806 122220
rect 83298 122146 87806 122168
rect 38 121676 3902 121698
rect 38 121624 916 121676
rect 968 121624 980 121676
rect 1032 121624 1044 121676
rect 1096 121624 1108 121676
rect 1160 121624 3902 121676
rect 38 121602 3902 121624
rect 83298 121676 87806 121698
rect 83298 121624 84916 121676
rect 84968 121624 84980 121676
rect 85032 121624 85044 121676
rect 85096 121624 85108 121676
rect 85160 121624 87806 121676
rect 83298 121602 87806 121624
rect 38 121132 3902 121154
rect 38 121080 2916 121132
rect 2968 121080 2980 121132
rect 3032 121080 3044 121132
rect 3096 121080 3108 121132
rect 3160 121080 3902 121132
rect 38 121058 3902 121080
rect 83298 121132 87806 121154
rect 83298 121080 86916 121132
rect 86968 121080 86980 121132
rect 87032 121080 87044 121132
rect 87096 121080 87108 121132
rect 87160 121080 87806 121132
rect 83298 121058 87806 121080
rect 83036 120842 83042 120894
rect 83094 120882 83100 120894
rect 84324 120882 84330 120894
rect 83094 120854 84330 120882
rect 83094 120842 83100 120854
rect 84324 120842 84330 120854
rect 84382 120842 84388 120894
rect 38 120588 3902 120610
rect 38 120536 916 120588
rect 968 120536 980 120588
rect 1032 120536 1044 120588
rect 1096 120536 1108 120588
rect 1160 120536 3902 120588
rect 38 120514 3902 120536
rect 83298 120588 87806 120610
rect 83298 120536 84916 120588
rect 84968 120536 84980 120588
rect 85032 120536 85044 120588
rect 85096 120536 85108 120588
rect 85160 120536 87806 120588
rect 83298 120514 87806 120536
rect 38 120044 3902 120066
rect 38 119992 2916 120044
rect 2968 119992 2980 120044
rect 3032 119992 3044 120044
rect 3096 119992 3108 120044
rect 3160 119992 3902 120044
rect 38 119970 3902 119992
rect 83298 120044 87806 120066
rect 83298 119992 86916 120044
rect 86968 119992 86980 120044
rect 87032 119992 87044 120044
rect 87096 119992 87108 120044
rect 87160 119992 87806 120044
rect 83298 119970 87806 119992
rect 82208 119618 82214 119670
rect 82266 119658 82272 119670
rect 84232 119658 84238 119670
rect 82266 119630 84238 119658
rect 82266 119618 82272 119630
rect 84232 119618 84238 119630
rect 84290 119618 84296 119670
rect 38 119500 3902 119522
rect 38 119448 916 119500
rect 968 119448 980 119500
rect 1032 119448 1044 119500
rect 1096 119448 1108 119500
rect 1160 119448 3902 119500
rect 38 119426 3902 119448
rect 83298 119500 87806 119522
rect 83298 119448 84916 119500
rect 84968 119448 84980 119500
rect 85032 119448 85044 119500
rect 85096 119448 85108 119500
rect 85160 119448 87806 119500
rect 83298 119426 87806 119448
rect 82484 119346 82490 119398
rect 82542 119386 82548 119398
rect 85336 119386 85342 119398
rect 82542 119358 85342 119386
rect 82542 119346 82548 119358
rect 85336 119346 85342 119358
rect 85394 119346 85400 119398
rect 38 118956 3902 118978
rect 38 118904 2916 118956
rect 2968 118904 2980 118956
rect 3032 118904 3044 118956
rect 3096 118904 3108 118956
rect 3160 118904 3902 118956
rect 38 118882 3902 118904
rect 83298 118956 87806 118978
rect 83298 118904 86916 118956
rect 86968 118904 86980 118956
rect 87032 118904 87044 118956
rect 87096 118904 87108 118956
rect 87160 118904 87806 118956
rect 83298 118882 87806 118904
rect 38 118412 3902 118434
rect 38 118360 916 118412
rect 968 118360 980 118412
rect 1032 118360 1044 118412
rect 1096 118360 1108 118412
rect 1160 118360 3902 118412
rect 38 118338 3902 118360
rect 83298 118412 87806 118434
rect 83298 118360 84916 118412
rect 84968 118360 84980 118412
rect 85032 118360 85044 118412
rect 85096 118360 85108 118412
rect 85160 118360 87806 118412
rect 83298 118338 87806 118360
rect 38 117868 3902 117890
rect 38 117816 2916 117868
rect 2968 117816 2980 117868
rect 3032 117816 3044 117868
rect 3096 117816 3108 117868
rect 3160 117816 3902 117868
rect 38 117794 3902 117816
rect 83298 117868 87806 117890
rect 83298 117816 86916 117868
rect 86968 117816 86980 117868
rect 87032 117816 87044 117868
rect 87096 117816 87108 117868
rect 87160 117816 87806 117868
rect 83298 117794 87806 117816
rect 38 117324 3902 117346
rect 38 117272 916 117324
rect 968 117272 980 117324
rect 1032 117272 1044 117324
rect 1096 117272 1108 117324
rect 1160 117272 3902 117324
rect 38 117250 3902 117272
rect 83298 117324 87806 117346
rect 83298 117272 84916 117324
rect 84968 117272 84980 117324
rect 85032 117272 85044 117324
rect 85096 117272 85108 117324
rect 85160 117272 87806 117324
rect 83298 117250 87806 117272
rect 38 116780 3902 116802
rect 38 116728 2916 116780
rect 2968 116728 2980 116780
rect 3032 116728 3044 116780
rect 3096 116728 3108 116780
rect 3160 116728 3902 116780
rect 38 116706 3902 116728
rect 83298 116780 87806 116802
rect 83298 116728 86916 116780
rect 86968 116728 86980 116780
rect 87032 116728 87044 116780
rect 87096 116728 87108 116780
rect 87160 116728 87806 116780
rect 83298 116706 87806 116728
rect 82392 116626 82398 116678
rect 82450 116666 82456 116678
rect 83956 116666 83962 116678
rect 82450 116638 83962 116666
rect 82450 116626 82456 116638
rect 83956 116626 83962 116638
rect 84014 116626 84020 116678
rect 3551 116465 3609 116471
rect 3551 116431 3563 116465
rect 3597 116462 3609 116465
rect 4100 116462 4106 116474
rect 3597 116434 4106 116462
rect 3597 116431 3609 116434
rect 3551 116425 3609 116431
rect 4100 116422 4106 116434
rect 4158 116462 4164 116474
rect 4284 116462 4290 116474
rect 4158 116434 4290 116462
rect 4158 116422 4164 116434
rect 4284 116422 4290 116434
rect 4342 116422 4348 116474
rect 38 116236 3902 116258
rect 38 116184 916 116236
rect 968 116184 980 116236
rect 1032 116184 1044 116236
rect 1096 116184 1108 116236
rect 1160 116184 3902 116236
rect 38 116162 3902 116184
rect 83298 116236 87806 116258
rect 83298 116184 84916 116236
rect 84968 116184 84980 116236
rect 85032 116184 85044 116236
rect 85096 116184 85108 116236
rect 85160 116184 87806 116236
rect 83298 116162 87806 116184
rect 38 115692 3902 115714
rect 38 115640 2916 115692
rect 2968 115640 2980 115692
rect 3032 115640 3044 115692
rect 3096 115640 3108 115692
rect 3160 115640 3902 115692
rect 38 115618 3902 115640
rect 83298 115692 87806 115714
rect 83298 115640 86916 115692
rect 86968 115640 86980 115692
rect 87032 115640 87044 115692
rect 87096 115640 87108 115692
rect 87160 115640 87806 115692
rect 83298 115618 87806 115640
rect 82944 115538 82950 115590
rect 83002 115578 83008 115590
rect 84324 115578 84330 115590
rect 83002 115550 84330 115578
rect 83002 115538 83008 115550
rect 84324 115538 84330 115550
rect 84382 115538 84388 115590
rect 38 115148 3902 115170
rect 38 115096 916 115148
rect 968 115096 980 115148
rect 1032 115096 1044 115148
rect 1096 115096 1108 115148
rect 1160 115096 3902 115148
rect 38 115074 3902 115096
rect 83298 115148 87806 115170
rect 83298 115096 84916 115148
rect 84968 115096 84980 115148
rect 85032 115096 85044 115148
rect 85096 115096 85108 115148
rect 85160 115096 87806 115148
rect 83298 115074 87806 115096
rect 3456 114858 3462 114910
rect 3514 114898 3520 114910
rect 4284 114898 4290 114910
rect 3514 114870 4290 114898
rect 3514 114858 3520 114870
rect 4284 114858 4290 114870
rect 4342 114858 4348 114910
rect 3456 114762 3462 114774
rect 3417 114734 3462 114762
rect 3456 114722 3462 114734
rect 3514 114722 3520 114774
rect 82300 114654 82306 114706
rect 82358 114694 82364 114706
rect 84324 114694 84330 114706
rect 82358 114666 84330 114694
rect 82358 114654 82364 114666
rect 84324 114654 84330 114666
rect 84382 114654 84388 114706
rect 38 114604 3902 114626
rect 38 114552 2916 114604
rect 2968 114552 2980 114604
rect 3032 114552 3044 114604
rect 3096 114552 3108 114604
rect 3160 114552 3902 114604
rect 38 114530 3902 114552
rect 83298 114604 87806 114626
rect 83298 114552 86916 114604
rect 86968 114552 86980 114604
rect 87032 114552 87044 114604
rect 87096 114552 87108 114604
rect 87160 114552 87806 114604
rect 83298 114530 87806 114552
rect 38 114060 3902 114082
rect 38 114008 916 114060
rect 968 114008 980 114060
rect 1032 114008 1044 114060
rect 1096 114008 1108 114060
rect 1160 114008 3902 114060
rect 38 113986 3902 114008
rect 83298 114060 87806 114082
rect 83298 114008 84916 114060
rect 84968 114008 84980 114060
rect 85032 114008 85044 114060
rect 85096 114008 85108 114060
rect 85160 114008 87806 114060
rect 83298 113986 87806 114008
rect 38 113516 3902 113538
rect 38 113464 2916 113516
rect 2968 113464 2980 113516
rect 3032 113464 3044 113516
rect 3096 113464 3108 113516
rect 3160 113464 3902 113516
rect 38 113442 3902 113464
rect 83298 113516 87806 113538
rect 83298 113464 86916 113516
rect 86968 113464 86980 113516
rect 87032 113464 87044 113516
rect 87096 113464 87108 113516
rect 87160 113464 87806 113516
rect 83298 113442 87806 113464
rect 38 112972 3902 112994
rect 38 112920 916 112972
rect 968 112920 980 112972
rect 1032 112920 1044 112972
rect 1096 112920 1108 112972
rect 1160 112920 3902 112972
rect 38 112898 3902 112920
rect 83298 112972 87806 112994
rect 83298 112920 84916 112972
rect 84968 112920 84980 112972
rect 85032 112920 85044 112972
rect 85096 112920 85108 112972
rect 85160 112920 87806 112972
rect 83298 112898 87806 112920
rect 38 112428 3902 112450
rect 38 112376 2916 112428
rect 2968 112376 2980 112428
rect 3032 112376 3044 112428
rect 3096 112376 3108 112428
rect 3160 112376 3902 112428
rect 38 112354 3902 112376
rect 83298 112428 87806 112450
rect 83298 112376 86916 112428
rect 86968 112376 86980 112428
rect 87032 112376 87044 112428
rect 87096 112376 87108 112428
rect 87160 112376 87806 112428
rect 83298 112354 87806 112376
rect 82484 112002 82490 112054
rect 82542 112042 82548 112054
rect 84876 112042 84882 112054
rect 82542 112014 84882 112042
rect 82542 112002 82548 112014
rect 84876 112002 84882 112014
rect 84934 112002 84940 112054
rect 82852 111934 82858 111986
rect 82910 111974 82916 111986
rect 83956 111974 83962 111986
rect 82910 111946 83962 111974
rect 82910 111934 82916 111946
rect 83956 111934 83962 111946
rect 84014 111934 84020 111986
rect 38 111884 3902 111906
rect 38 111832 916 111884
rect 968 111832 980 111884
rect 1032 111832 1044 111884
rect 1096 111832 1108 111884
rect 1160 111832 3902 111884
rect 38 111810 3902 111832
rect 83298 111884 87806 111906
rect 83298 111832 84916 111884
rect 84968 111832 84980 111884
rect 85032 111832 85044 111884
rect 85096 111832 85108 111884
rect 85160 111832 87806 111884
rect 83298 111810 87806 111832
rect 38 111340 3902 111362
rect 38 111288 2916 111340
rect 2968 111288 2980 111340
rect 3032 111288 3044 111340
rect 3096 111288 3108 111340
rect 3160 111288 3902 111340
rect 38 111266 3902 111288
rect 83298 111340 87806 111362
rect 83298 111288 86916 111340
rect 86968 111288 86980 111340
rect 87032 111288 87044 111340
rect 87096 111288 87108 111340
rect 87160 111288 87806 111340
rect 83298 111266 87806 111288
rect 38 110796 3902 110818
rect 38 110744 916 110796
rect 968 110744 980 110796
rect 1032 110744 1044 110796
rect 1096 110744 1108 110796
rect 1160 110744 3902 110796
rect 38 110722 3902 110744
rect 83298 110796 87806 110818
rect 83298 110744 84916 110796
rect 84968 110744 84980 110796
rect 85032 110744 85044 110796
rect 85096 110744 85108 110796
rect 85160 110744 87806 110796
rect 83298 110722 87806 110744
rect 3548 110642 3554 110694
rect 3606 110682 3612 110694
rect 4011 110685 4069 110691
rect 4011 110682 4023 110685
rect 3606 110654 4023 110682
rect 3606 110642 3612 110654
rect 4011 110651 4023 110654
rect 4057 110651 4069 110685
rect 4011 110645 4069 110651
rect 3732 110574 3738 110626
rect 3790 110614 3796 110626
rect 4103 110617 4161 110623
rect 4103 110614 4115 110617
rect 3790 110586 4115 110614
rect 3790 110574 3796 110586
rect 4103 110583 4115 110586
rect 4149 110583 4161 110617
rect 4103 110577 4161 110583
rect 38 110252 3902 110274
rect 38 110200 2916 110252
rect 2968 110200 2980 110252
rect 3032 110200 3044 110252
rect 3096 110200 3108 110252
rect 3160 110200 3902 110252
rect 38 110178 3902 110200
rect 83298 110252 87806 110274
rect 83298 110200 86916 110252
rect 86968 110200 86980 110252
rect 87032 110200 87044 110252
rect 87096 110200 87108 110252
rect 87160 110200 87806 110252
rect 83298 110178 87806 110200
rect 38 109708 3902 109730
rect 38 109656 916 109708
rect 968 109656 980 109708
rect 1032 109656 1044 109708
rect 1096 109656 1108 109708
rect 1160 109656 3902 109708
rect 38 109634 3902 109656
rect 83298 109708 87806 109730
rect 83298 109656 84916 109708
rect 84968 109656 84980 109708
rect 85032 109656 85044 109708
rect 85096 109656 85108 109708
rect 85160 109656 87806 109708
rect 83298 109634 87806 109656
rect 81840 109282 81846 109334
rect 81898 109322 81904 109334
rect 83956 109322 83962 109334
rect 81898 109294 83962 109322
rect 81898 109282 81904 109294
rect 83956 109282 83962 109294
rect 84014 109282 84020 109334
rect 38 109164 3902 109186
rect 38 109112 2916 109164
rect 2968 109112 2980 109164
rect 3032 109112 3044 109164
rect 3096 109112 3108 109164
rect 3160 109112 3902 109164
rect 38 109090 3902 109112
rect 83298 109164 87806 109186
rect 83298 109112 86916 109164
rect 86968 109112 86980 109164
rect 87032 109112 87044 109164
rect 87096 109112 87108 109164
rect 87160 109112 87806 109164
rect 83298 109090 87806 109112
rect 38 108620 3902 108642
rect 38 108568 916 108620
rect 968 108568 980 108620
rect 1032 108568 1044 108620
rect 1096 108568 1108 108620
rect 1160 108568 3902 108620
rect 38 108546 3902 108568
rect 83298 108620 87806 108642
rect 83298 108568 84916 108620
rect 84968 108568 84980 108620
rect 85032 108568 85044 108620
rect 85096 108568 85108 108620
rect 85160 108568 87806 108620
rect 83298 108546 87806 108568
rect 81656 108126 81662 108178
rect 81714 108166 81720 108178
rect 83956 108166 83962 108178
rect 81714 108138 83962 108166
rect 81714 108126 81720 108138
rect 83956 108126 83962 108138
rect 84014 108126 84020 108178
rect 38 108076 3902 108098
rect 38 108024 2916 108076
rect 2968 108024 2980 108076
rect 3032 108024 3044 108076
rect 3096 108024 3108 108076
rect 3160 108024 3902 108076
rect 38 108002 3902 108024
rect 83298 108076 87806 108098
rect 83298 108024 86916 108076
rect 86968 108024 86980 108076
rect 87032 108024 87044 108076
rect 87096 108024 87108 108076
rect 87160 108024 87806 108076
rect 83298 108002 87806 108024
rect 38 107532 3902 107554
rect 38 107480 916 107532
rect 968 107480 980 107532
rect 1032 107480 1044 107532
rect 1096 107480 1108 107532
rect 1160 107480 3902 107532
rect 38 107458 3902 107480
rect 83298 107532 87806 107554
rect 83298 107480 84916 107532
rect 84968 107480 84980 107532
rect 85032 107480 85044 107532
rect 85096 107480 85108 107532
rect 85160 107480 87806 107532
rect 83298 107458 87806 107480
rect 38 106988 3902 107010
rect 38 106936 2916 106988
rect 2968 106936 2980 106988
rect 3032 106936 3044 106988
rect 3096 106936 3108 106988
rect 3160 106936 3902 106988
rect 38 106914 3902 106936
rect 83298 106988 87806 107010
rect 83298 106936 86916 106988
rect 86968 106936 86980 106988
rect 87032 106936 87044 106988
rect 87096 106936 87108 106988
rect 87160 106936 87806 106988
rect 83298 106914 87806 106936
rect 82576 106562 82582 106614
rect 82634 106602 82640 106614
rect 84232 106602 84238 106614
rect 82634 106574 84238 106602
rect 82634 106562 82640 106574
rect 84232 106562 84238 106574
rect 84290 106562 84296 106614
rect 38 106444 3902 106466
rect 38 106392 916 106444
rect 968 106392 980 106444
rect 1032 106392 1044 106444
rect 1096 106392 1108 106444
rect 1160 106392 3902 106444
rect 38 106370 3902 106392
rect 83298 106444 87806 106466
rect 83298 106392 84916 106444
rect 84968 106392 84980 106444
rect 85032 106392 85044 106444
rect 85096 106392 85108 106444
rect 85160 106392 87806 106444
rect 83298 106370 87806 106392
rect 38 105900 3902 105922
rect 38 105848 2916 105900
rect 2968 105848 2980 105900
rect 3032 105848 3044 105900
rect 3096 105848 3108 105900
rect 3160 105848 3902 105900
rect 38 105826 3902 105848
rect 83298 105900 87806 105922
rect 83298 105848 86916 105900
rect 86968 105848 86980 105900
rect 87032 105848 87044 105900
rect 87096 105848 87108 105900
rect 87160 105848 87806 105900
rect 83298 105826 87806 105848
rect 3732 105474 3738 105526
rect 3790 105514 3796 105526
rect 4103 105517 4161 105523
rect 4103 105514 4115 105517
rect 3790 105486 4115 105514
rect 3790 105474 3796 105486
rect 4103 105483 4115 105486
rect 4149 105483 4161 105517
rect 4103 105477 4161 105483
rect 3548 105406 3554 105458
rect 3606 105446 3612 105458
rect 4011 105449 4069 105455
rect 4011 105446 4023 105449
rect 3606 105418 4023 105446
rect 3606 105406 3612 105418
rect 4011 105415 4023 105418
rect 4057 105415 4069 105449
rect 4011 105409 4069 105415
rect 38 105356 3902 105378
rect 38 105304 916 105356
rect 968 105304 980 105356
rect 1032 105304 1044 105356
rect 1096 105304 1108 105356
rect 1160 105304 3902 105356
rect 38 105282 3902 105304
rect 83298 105356 87806 105378
rect 83298 105304 84916 105356
rect 84968 105304 84980 105356
rect 85032 105304 85044 105356
rect 85096 105304 85108 105356
rect 85160 105304 87806 105356
rect 83298 105282 87806 105304
rect 38 104812 3902 104834
rect 38 104760 2916 104812
rect 2968 104760 2980 104812
rect 3032 104760 3044 104812
rect 3096 104760 3108 104812
rect 3160 104760 3902 104812
rect 38 104738 3902 104760
rect 83298 104812 87806 104834
rect 83298 104760 86916 104812
rect 86968 104760 86980 104812
rect 87032 104760 87044 104812
rect 87096 104760 87108 104812
rect 87160 104760 87806 104812
rect 83298 104738 87806 104760
rect 38 104268 3902 104290
rect 38 104216 916 104268
rect 968 104216 980 104268
rect 1032 104216 1044 104268
rect 1096 104216 1108 104268
rect 1160 104216 3902 104268
rect 38 104194 3902 104216
rect 83298 104268 87806 104290
rect 83298 104216 84916 104268
rect 84968 104216 84980 104268
rect 85032 104216 85044 104268
rect 85096 104216 85108 104268
rect 85160 104216 87806 104268
rect 83298 104194 87806 104216
rect 38 103724 3902 103746
rect 38 103672 2916 103724
rect 2968 103672 2980 103724
rect 3032 103672 3044 103724
rect 3096 103672 3108 103724
rect 3160 103672 3902 103724
rect 38 103650 3902 103672
rect 83298 103724 87806 103746
rect 83298 103672 86916 103724
rect 86968 103672 86980 103724
rect 87032 103672 87044 103724
rect 87096 103672 87108 103724
rect 87160 103672 87806 103724
rect 83298 103650 87806 103672
rect 84784 103434 84790 103486
rect 84842 103474 84848 103486
rect 85244 103474 85250 103486
rect 84842 103446 85250 103474
rect 84842 103434 84848 103446
rect 85244 103434 85250 103446
rect 85302 103434 85308 103486
rect 38 103180 3902 103202
rect 38 103128 916 103180
rect 968 103128 980 103180
rect 1032 103128 1044 103180
rect 1096 103128 1108 103180
rect 1160 103128 3902 103180
rect 38 103106 3902 103128
rect 83298 103180 87806 103202
rect 83298 103128 84916 103180
rect 84968 103128 84980 103180
rect 85032 103128 85044 103180
rect 85096 103128 85108 103180
rect 85160 103128 87806 103180
rect 83298 103106 87806 103128
rect 82760 102822 82766 102874
rect 82818 102862 82824 102874
rect 84508 102862 84514 102874
rect 82818 102834 84514 102862
rect 82818 102822 82824 102834
rect 84508 102822 84514 102834
rect 84566 102822 84572 102874
rect 84048 102686 84054 102738
rect 84106 102726 84112 102738
rect 84508 102726 84514 102738
rect 84106 102698 84514 102726
rect 84106 102686 84112 102698
rect 84508 102686 84514 102698
rect 84566 102686 84572 102738
rect 38 102636 3902 102658
rect 38 102584 2916 102636
rect 2968 102584 2980 102636
rect 3032 102584 3044 102636
rect 3096 102584 3108 102636
rect 3160 102584 3902 102636
rect 38 102562 3902 102584
rect 83298 102636 87806 102658
rect 83298 102584 86916 102636
rect 86968 102584 86980 102636
rect 87032 102584 87044 102636
rect 87096 102584 87108 102636
rect 87160 102584 87806 102636
rect 83298 102562 87806 102584
rect 38 102092 3902 102114
rect 38 102040 916 102092
rect 968 102040 980 102092
rect 1032 102040 1044 102092
rect 1096 102040 1108 102092
rect 1160 102040 3902 102092
rect 38 102018 3902 102040
rect 83298 102092 87806 102114
rect 83298 102040 84916 102092
rect 84968 102040 84980 102092
rect 85032 102040 85044 102092
rect 85096 102040 85108 102092
rect 85160 102040 87806 102092
rect 83298 102018 87806 102040
rect 81748 101598 81754 101650
rect 81806 101638 81812 101650
rect 84324 101638 84330 101650
rect 81806 101610 84330 101638
rect 81806 101598 81812 101610
rect 84324 101598 84330 101610
rect 84382 101598 84388 101650
rect 38 101548 3902 101570
rect 38 101496 2916 101548
rect 2968 101496 2980 101548
rect 3032 101496 3044 101548
rect 3096 101496 3108 101548
rect 3160 101496 3902 101548
rect 38 101474 3902 101496
rect 83298 101548 87806 101570
rect 83298 101496 86916 101548
rect 86968 101496 86980 101548
rect 87032 101496 87044 101548
rect 87096 101496 87108 101548
rect 87160 101496 87806 101548
rect 83298 101474 87806 101496
rect 38 101004 3902 101026
rect 38 100952 916 101004
rect 968 100952 980 101004
rect 1032 100952 1044 101004
rect 1096 100952 1108 101004
rect 1160 100952 3902 101004
rect 38 100930 3902 100952
rect 83298 101004 87806 101026
rect 83298 100952 84916 101004
rect 84968 100952 84980 101004
rect 85032 100952 85044 101004
rect 85096 100952 85108 101004
rect 85160 100952 87806 101004
rect 83298 100930 87806 100952
rect 84048 100510 84054 100562
rect 84106 100550 84112 100562
rect 84324 100550 84330 100562
rect 84106 100522 84330 100550
rect 84106 100510 84112 100522
rect 84324 100510 84330 100522
rect 84382 100510 84388 100562
rect 38 100460 3902 100482
rect 38 100408 2916 100460
rect 2968 100408 2980 100460
rect 3032 100408 3044 100460
rect 3096 100408 3108 100460
rect 3160 100408 3902 100460
rect 38 100386 3902 100408
rect 83298 100460 87806 100482
rect 83298 100408 86916 100460
rect 86968 100408 86980 100460
rect 87032 100408 87044 100460
rect 87096 100408 87108 100460
rect 87160 100408 87806 100460
rect 83298 100386 87806 100408
rect 84048 100306 84054 100358
rect 84106 100346 84112 100358
rect 84692 100346 84698 100358
rect 84106 100318 84698 100346
rect 84106 100306 84112 100318
rect 84692 100306 84698 100318
rect 84750 100306 84756 100358
rect 38 99916 3902 99938
rect 38 99864 916 99916
rect 968 99864 980 99916
rect 1032 99864 1044 99916
rect 1096 99864 1108 99916
rect 1160 99864 3902 99916
rect 38 99842 3902 99864
rect 83298 99916 87806 99938
rect 83298 99864 84916 99916
rect 84968 99864 84980 99916
rect 85032 99864 85044 99916
rect 85096 99864 85108 99916
rect 85160 99864 87806 99916
rect 83298 99842 87806 99864
rect 38 99372 3902 99394
rect 38 99320 2916 99372
rect 2968 99320 2980 99372
rect 3032 99320 3044 99372
rect 3096 99320 3108 99372
rect 3160 99320 3902 99372
rect 38 99298 3902 99320
rect 83298 99372 87806 99394
rect 83298 99320 86916 99372
rect 86968 99320 86980 99372
rect 87032 99320 87044 99372
rect 87096 99320 87108 99372
rect 87160 99320 87806 99372
rect 83298 99298 87806 99320
rect 4011 99125 4069 99131
rect 4011 99091 4023 99125
rect 4057 99122 4069 99125
rect 4560 99122 4566 99134
rect 4057 99094 4566 99122
rect 4057 99091 4069 99094
rect 4011 99085 4069 99091
rect 4560 99082 4566 99094
rect 4618 99082 4624 99134
rect 4376 98946 4382 98998
rect 4434 98986 4440 98998
rect 4744 98986 4750 98998
rect 4434 98958 4750 98986
rect 4434 98946 4440 98958
rect 4744 98946 4750 98958
rect 4802 98946 4808 98998
rect 85244 98986 85250 98998
rect 84894 98958 85250 98986
rect 84894 98918 84922 98958
rect 85244 98946 85250 98958
rect 85302 98946 85308 98998
rect 86532 98918 86538 98930
rect 84894 98890 86538 98918
rect 86532 98878 86538 98890
rect 86590 98878 86596 98930
rect 38 98828 3902 98850
rect 38 98776 916 98828
rect 968 98776 980 98828
rect 1032 98776 1044 98828
rect 1096 98776 1108 98828
rect 1160 98776 3902 98828
rect 38 98754 3902 98776
rect 83298 98828 87806 98850
rect 83298 98776 84916 98828
rect 84968 98776 84980 98828
rect 85032 98776 85044 98828
rect 85096 98776 85108 98828
rect 85160 98776 87806 98828
rect 83298 98754 87806 98776
rect 4652 98674 4658 98726
rect 4710 98714 4716 98726
rect 4928 98714 4934 98726
rect 4710 98686 4934 98714
rect 4710 98674 4716 98686
rect 4928 98674 4934 98686
rect 4986 98674 4992 98726
rect 1892 98334 1898 98386
rect 1950 98374 1956 98386
rect 2812 98374 2818 98386
rect 1950 98346 2818 98374
rect 1950 98334 1956 98346
rect 2812 98334 2818 98346
rect 2870 98374 2876 98386
rect 3091 98377 3149 98383
rect 3091 98374 3103 98377
rect 2870 98346 3103 98374
rect 2870 98334 2876 98346
rect 3091 98343 3103 98346
rect 3137 98343 3149 98377
rect 3091 98337 3149 98343
rect 3551 98377 3609 98383
rect 3551 98343 3563 98377
rect 3597 98374 3609 98377
rect 4100 98374 4106 98386
rect 3597 98346 4106 98374
rect 3597 98343 3609 98346
rect 3551 98337 3609 98343
rect 4100 98334 4106 98346
rect 4158 98334 4164 98386
rect 38 98284 3902 98306
rect 38 98232 2916 98284
rect 2968 98232 2980 98284
rect 3032 98232 3044 98284
rect 3096 98232 3108 98284
rect 3160 98232 3902 98284
rect 38 98210 3902 98232
rect 83298 98284 87806 98306
rect 83298 98232 86916 98284
rect 86968 98232 86980 98284
rect 87032 98232 87044 98284
rect 87096 98232 87108 98284
rect 87160 98232 87806 98284
rect 83298 98210 87806 98232
rect 3551 98173 3609 98179
rect 3551 98139 3563 98173
rect 3597 98170 3609 98173
rect 4100 98170 4106 98182
rect 3597 98142 4106 98170
rect 3597 98139 3609 98142
rect 3551 98133 3609 98139
rect 4100 98130 4106 98142
rect 4158 98170 4164 98182
rect 5112 98170 5118 98182
rect 4158 98142 5118 98170
rect 4158 98130 4164 98142
rect 5112 98130 5118 98142
rect 5170 98130 5176 98182
rect 82668 98130 82674 98182
rect 82726 98170 82732 98182
rect 83864 98170 83870 98182
rect 82726 98142 83870 98170
rect 82726 98130 82732 98142
rect 83864 98130 83870 98142
rect 83922 98130 83928 98182
rect 84324 97994 84330 98046
rect 84382 98034 84388 98046
rect 85152 98034 85158 98046
rect 84382 98006 85158 98034
rect 84382 97994 84388 98006
rect 85152 97994 85158 98006
rect 85210 97994 85216 98046
rect 2260 97790 2266 97842
rect 2318 97830 2324 97842
rect 2355 97833 2413 97839
rect 2355 97830 2367 97833
rect 2318 97802 2367 97830
rect 2318 97790 2324 97802
rect 2355 97799 2367 97802
rect 2401 97830 2413 97833
rect 2444 97830 2450 97842
rect 2401 97802 2450 97830
rect 2401 97799 2413 97802
rect 2355 97793 2413 97799
rect 2444 97790 2450 97802
rect 2502 97790 2508 97842
rect 2815 97833 2873 97839
rect 2815 97799 2827 97833
rect 2861 97830 2873 97833
rect 4011 97833 4069 97839
rect 4011 97830 4023 97833
rect 2861 97802 4023 97830
rect 2861 97799 2873 97802
rect 2815 97793 2873 97799
rect 4011 97799 4023 97802
rect 4057 97799 4069 97833
rect 4011 97793 4069 97799
rect 38 97740 3902 97762
rect 38 97688 916 97740
rect 968 97688 980 97740
rect 1032 97688 1044 97740
rect 1096 97688 1108 97740
rect 1160 97688 3902 97740
rect 38 97666 3902 97688
rect 83298 97740 87806 97762
rect 83298 97688 84916 97740
rect 84968 97688 84980 97740
rect 85032 97688 85044 97740
rect 85096 97688 85108 97740
rect 85160 97688 87806 97740
rect 83298 97666 87806 97688
rect 2812 97626 2818 97638
rect 2773 97598 2818 97626
rect 2812 97586 2818 97598
rect 2870 97586 2876 97638
rect 3183 97629 3241 97635
rect 3183 97595 3195 97629
rect 3229 97626 3241 97629
rect 3364 97626 3370 97638
rect 3229 97598 3370 97626
rect 3229 97595 3241 97598
rect 3183 97589 3241 97595
rect 3364 97586 3370 97598
rect 3422 97626 3428 97638
rect 4376 97626 4382 97638
rect 3422 97598 4382 97626
rect 3422 97586 3428 97598
rect 4376 97586 4382 97598
rect 4434 97586 4440 97638
rect 83039 97629 83097 97635
rect 83039 97595 83051 97629
rect 83085 97626 83097 97629
rect 83956 97626 83962 97638
rect 83085 97598 83962 97626
rect 83085 97595 83097 97598
rect 83039 97589 83097 97595
rect 83956 97586 83962 97598
rect 84014 97586 84020 97638
rect 84235 97629 84293 97635
rect 84235 97595 84247 97629
rect 84281 97626 84293 97629
rect 84508 97626 84514 97638
rect 84281 97598 84514 97626
rect 84281 97595 84293 97598
rect 84235 97589 84293 97595
rect 2076 97518 2082 97570
rect 2134 97558 2140 97570
rect 5759 97561 5817 97567
rect 5759 97558 5771 97561
rect 2134 97530 5771 97558
rect 2134 97518 2140 97530
rect 5759 97527 5771 97530
rect 5805 97527 5817 97561
rect 83772 97558 83778 97570
rect 83733 97530 83778 97558
rect 5759 97521 5817 97527
rect 83772 97518 83778 97530
rect 83830 97518 83836 97570
rect 1711 97493 1769 97499
rect 1711 97459 1723 97493
rect 1757 97490 1769 97493
rect 4100 97490 4106 97502
rect 1757 97462 4106 97490
rect 1757 97459 1769 97462
rect 1711 97453 1769 97459
rect 4100 97450 4106 97462
rect 4158 97450 4164 97502
rect 81472 97450 81478 97502
rect 81530 97490 81536 97502
rect 84250 97490 84278 97589
rect 84508 97586 84514 97598
rect 84566 97586 84572 97638
rect 81530 97462 84278 97490
rect 81530 97450 81536 97462
rect 2812 97382 2818 97434
rect 2870 97422 2876 97434
rect 3916 97422 3922 97434
rect 2870 97394 3922 97422
rect 2870 97382 2876 97394
rect 3916 97382 3922 97394
rect 3974 97382 3980 97434
rect 81291 97425 81349 97431
rect 81291 97391 81303 97425
rect 81337 97422 81349 97425
rect 86072 97422 86078 97434
rect 81337 97394 86078 97422
rect 81337 97391 81349 97394
rect 81291 97385 81349 97391
rect 86072 97382 86078 97394
rect 86130 97382 86136 97434
rect 1340 97314 1346 97366
rect 1398 97354 1404 97366
rect 5759 97357 5817 97363
rect 5759 97354 5771 97357
rect 1398 97326 5771 97354
rect 1398 97314 1404 97326
rect 5759 97323 5771 97326
rect 5805 97323 5817 97357
rect 83128 97354 83134 97366
rect 5759 97317 5817 97323
rect 81306 97326 83134 97354
rect 81306 97298 81334 97326
rect 83128 97314 83134 97326
rect 83186 97314 83192 97366
rect 85796 97354 85802 97366
rect 83698 97326 85802 97354
rect 2076 97286 2082 97298
rect 2037 97258 2082 97286
rect 2076 97246 2082 97258
rect 2134 97246 2140 97298
rect 2352 97246 2358 97298
rect 2410 97286 2416 97298
rect 2447 97289 2505 97295
rect 2447 97286 2459 97289
rect 2410 97258 2459 97286
rect 2410 97246 2416 97258
rect 2447 97255 2459 97258
rect 2493 97286 2505 97289
rect 2536 97286 2542 97298
rect 2493 97258 2542 97286
rect 2493 97255 2505 97258
rect 2447 97249 2505 97255
rect 2536 97246 2542 97258
rect 2594 97246 2600 97298
rect 3364 97246 3370 97298
rect 3422 97286 3428 97298
rect 3459 97289 3517 97295
rect 3459 97286 3471 97289
rect 3422 97258 3471 97286
rect 3422 97246 3428 97258
rect 3459 97255 3471 97258
rect 3505 97255 3517 97289
rect 3459 97249 3517 97255
rect 81288 97246 81294 97298
rect 81346 97246 81352 97298
rect 81383 97289 81441 97295
rect 81383 97255 81395 97289
rect 81429 97286 81441 97289
rect 83698 97286 83726 97326
rect 85796 97314 85802 97326
rect 85854 97314 85860 97366
rect 81429 97258 83726 97286
rect 81429 97255 81441 97258
rect 81383 97249 81441 97255
rect 38 97196 3902 97218
rect 38 97144 2916 97196
rect 2968 97144 2980 97196
rect 3032 97144 3044 97196
rect 3096 97144 3108 97196
rect 3160 97144 3902 97196
rect 83298 97196 87806 97218
rect 83036 97150 83042 97162
rect 38 97122 3902 97144
rect 56650 97122 83042 97150
rect 975 97085 1033 97091
rect 975 97051 987 97085
rect 1021 97082 1033 97085
rect 1021 97054 2030 97082
rect 1021 97051 1033 97054
rect 975 97045 1033 97051
rect 1340 97014 1346 97026
rect 1301 96986 1346 97014
rect 1340 96974 1346 96986
rect 1398 96974 1404 97026
rect 2002 96946 2030 97054
rect 3732 97042 3738 97094
rect 3790 97082 3796 97094
rect 3916 97082 3922 97094
rect 3790 97054 3922 97082
rect 3790 97042 3796 97054
rect 3916 97042 3922 97054
rect 3974 97042 3980 97094
rect 4468 97082 4474 97094
rect 4026 97054 4474 97082
rect 2079 97017 2137 97023
rect 2079 96983 2091 97017
rect 2125 97014 2137 97017
rect 4026 97014 4054 97054
rect 4468 97042 4474 97054
rect 4526 97042 4532 97094
rect 5943 97085 6001 97091
rect 5943 97051 5955 97085
rect 5989 97082 6001 97085
rect 22132 97082 22138 97094
rect 5989 97054 22138 97082
rect 5989 97051 6001 97054
rect 5943 97045 6001 97051
rect 22132 97042 22138 97054
rect 22190 97042 22196 97094
rect 45316 97042 45322 97094
rect 45374 97082 45380 97094
rect 45374 97054 56586 97082
rect 45374 97042 45380 97054
rect 2125 96986 4054 97014
rect 2125 96983 2137 96986
rect 2079 96977 2137 96983
rect 4100 96974 4106 97026
rect 4158 97014 4164 97026
rect 5296 97014 5302 97026
rect 4158 96986 5302 97014
rect 4158 96974 4164 96986
rect 5296 96974 5302 96986
rect 5354 97014 5360 97026
rect 14588 97014 14594 97026
rect 5354 96986 14594 97014
rect 5354 96974 5360 96986
rect 14588 96974 14594 96986
rect 14646 96974 14652 97026
rect 14959 97017 15017 97023
rect 14959 96983 14971 97017
rect 15005 97014 15017 97017
rect 28480 97014 28486 97026
rect 15005 96986 28486 97014
rect 15005 96983 15017 96986
rect 14959 96977 15017 96983
rect 28480 96974 28486 96986
rect 28538 96974 28544 97026
rect 5204 96946 5210 96958
rect 2002 96918 5210 96946
rect 5204 96906 5210 96918
rect 5262 96906 5268 96958
rect 56558 96946 56586 97054
rect 56650 97026 56678 97122
rect 83036 97110 83042 97122
rect 83094 97110 83100 97162
rect 83298 97144 86916 97196
rect 86968 97144 86980 97196
rect 87032 97144 87044 97196
rect 87096 97144 87108 97196
rect 87160 97144 87806 97196
rect 83298 97122 87806 97144
rect 81291 97085 81349 97091
rect 81291 97082 81303 97085
rect 56742 97054 81303 97082
rect 56632 96974 56638 97026
rect 56690 96974 56696 97026
rect 56742 96946 56770 97054
rect 81291 97051 81303 97054
rect 81337 97051 81349 97085
rect 81291 97045 81349 97051
rect 81380 97042 81386 97094
rect 81438 97082 81444 97094
rect 82944 97082 82950 97094
rect 81438 97054 82950 97082
rect 81438 97042 81444 97054
rect 82944 97042 82950 97054
rect 83002 97042 83008 97094
rect 84140 97082 84146 97094
rect 84101 97054 84146 97082
rect 84140 97042 84146 97054
rect 84198 97042 84204 97094
rect 60864 96974 60870 97026
rect 60922 97014 60928 97026
rect 83039 97017 83097 97023
rect 83039 97014 83051 97017
rect 60922 96986 83051 97014
rect 60922 96974 60928 96986
rect 83039 96983 83051 96986
rect 83085 96983 83097 97017
rect 83039 96977 83097 96983
rect 56558 96918 56770 96946
rect 80276 96906 80282 96958
rect 80334 96946 80340 96958
rect 81383 96949 81441 96955
rect 81383 96946 81395 96949
rect 80334 96918 81395 96946
rect 80334 96906 80340 96918
rect 81383 96915 81395 96918
rect 81429 96915 81441 96949
rect 81383 96909 81441 96915
rect 81475 96949 81533 96955
rect 81475 96915 81487 96949
rect 81521 96946 81533 96949
rect 82852 96946 82858 96958
rect 81521 96918 82858 96946
rect 81521 96915 81533 96918
rect 81475 96909 81533 96915
rect 82852 96906 82858 96918
rect 82910 96906 82916 96958
rect 2815 96881 2873 96887
rect 2815 96847 2827 96881
rect 2861 96878 2873 96881
rect 4560 96878 4566 96890
rect 2861 96850 4566 96878
rect 2861 96847 2873 96850
rect 2815 96841 2873 96847
rect 4560 96838 4566 96850
rect 4618 96838 4624 96890
rect 5759 96881 5817 96887
rect 5759 96847 5771 96881
rect 5805 96878 5817 96881
rect 19559 96881 19617 96887
rect 5805 96850 15738 96878
rect 5805 96847 5817 96850
rect 5759 96841 5817 96847
rect 15710 96810 15738 96850
rect 19559 96847 19571 96881
rect 19605 96878 19617 96881
rect 19605 96850 24662 96878
rect 19605 96847 19617 96850
rect 19559 96841 19617 96847
rect 19467 96813 19525 96819
rect 19467 96810 19479 96813
rect 3474 96782 5526 96810
rect 15710 96782 19479 96810
rect 1708 96742 1714 96754
rect 1669 96714 1714 96742
rect 1708 96702 1714 96714
rect 1766 96702 1772 96754
rect 2447 96745 2505 96751
rect 2447 96711 2459 96745
rect 2493 96742 2505 96745
rect 2996 96742 3002 96754
rect 2493 96714 3002 96742
rect 2493 96711 2505 96714
rect 2447 96705 2505 96711
rect 2996 96702 3002 96714
rect 3054 96742 3060 96754
rect 3474 96742 3502 96782
rect 3054 96714 3502 96742
rect 3551 96745 3609 96751
rect 3054 96702 3060 96714
rect 3551 96711 3563 96745
rect 3597 96742 3609 96745
rect 4928 96742 4934 96754
rect 3597 96714 4934 96742
rect 3597 96711 3609 96714
rect 3551 96705 3609 96711
rect 4928 96702 4934 96714
rect 4986 96702 4992 96754
rect 5498 96742 5526 96782
rect 19467 96779 19479 96782
rect 19513 96779 19525 96813
rect 24634 96810 24662 96850
rect 50192 96838 50198 96890
rect 50250 96878 50256 96890
rect 74759 96881 74817 96887
rect 74759 96878 74771 96881
rect 50250 96850 74771 96878
rect 50250 96838 50256 96850
rect 74759 96847 74771 96850
rect 74805 96847 74817 96881
rect 74759 96841 74817 96847
rect 80184 96838 80190 96890
rect 80242 96878 80248 96890
rect 83588 96878 83594 96890
rect 80242 96850 83594 96878
rect 80242 96838 80248 96850
rect 83588 96838 83594 96850
rect 83646 96838 83652 96890
rect 83772 96878 83778 96890
rect 83733 96850 83778 96878
rect 83772 96838 83778 96850
rect 83830 96838 83836 96890
rect 84508 96838 84514 96890
rect 84566 96878 84572 96890
rect 84784 96878 84790 96890
rect 84566 96850 84790 96878
rect 84566 96838 84572 96850
rect 84784 96838 84790 96850
rect 84842 96838 84848 96890
rect 25260 96810 25266 96822
rect 24634 96782 25266 96810
rect 19467 96773 19525 96779
rect 25260 96770 25266 96782
rect 25318 96770 25324 96822
rect 51664 96770 51670 96822
rect 51722 96810 51728 96822
rect 72735 96813 72793 96819
rect 72735 96810 72747 96813
rect 51722 96782 72747 96810
rect 51722 96770 51728 96782
rect 72735 96779 72747 96782
rect 72781 96779 72793 96813
rect 72735 96773 72793 96779
rect 73655 96813 73713 96819
rect 73655 96779 73667 96813
rect 73701 96810 73713 96813
rect 81475 96813 81533 96819
rect 81475 96810 81487 96813
rect 73701 96782 81487 96810
rect 73701 96779 73713 96782
rect 73655 96773 73713 96779
rect 81475 96779 81487 96782
rect 81521 96779 81533 96813
rect 84232 96810 84238 96822
rect 81475 96773 81533 96779
rect 83146 96782 84238 96810
rect 5848 96742 5854 96754
rect 5498 96714 5854 96742
rect 5848 96702 5854 96714
rect 5906 96742 5912 96754
rect 14959 96745 15017 96751
rect 14959 96742 14971 96745
rect 5906 96714 14971 96742
rect 5906 96702 5912 96714
rect 14959 96711 14971 96714
rect 15005 96711 15017 96745
rect 80003 96745 80061 96751
rect 80003 96742 80015 96745
rect 14959 96705 15017 96711
rect 66586 96714 80015 96742
rect 38 96652 3902 96674
rect 38 96600 916 96652
rect 968 96600 980 96652
rect 1032 96600 1044 96652
rect 1096 96600 1108 96652
rect 1160 96600 3902 96652
rect 4560 96634 4566 96686
rect 4618 96674 4624 96686
rect 28940 96674 28946 96686
rect 4618 96646 28946 96674
rect 4618 96634 4624 96646
rect 28940 96634 28946 96646
rect 28998 96634 29004 96686
rect 34920 96634 34926 96686
rect 34978 96674 34984 96686
rect 37036 96674 37042 96686
rect 34978 96646 37042 96674
rect 34978 96634 34984 96646
rect 37036 96634 37042 96646
rect 37094 96634 37100 96686
rect 48904 96634 48910 96686
rect 48962 96674 48968 96686
rect 48962 96646 62106 96674
rect 48962 96634 48968 96646
rect 38 96578 3902 96600
rect 4376 96566 4382 96618
rect 4434 96606 4440 96618
rect 29952 96606 29958 96618
rect 4434 96578 29958 96606
rect 4434 96566 4440 96578
rect 29952 96566 29958 96578
rect 30010 96566 30016 96618
rect 62078 96606 62106 96646
rect 66586 96606 66614 96714
rect 80003 96711 80015 96714
rect 80049 96711 80061 96745
rect 80003 96705 80061 96711
rect 80092 96702 80098 96754
rect 80150 96742 80156 96754
rect 83146 96742 83174 96782
rect 84232 96770 84238 96782
rect 84290 96770 84296 96822
rect 84603 96813 84661 96819
rect 84603 96779 84615 96813
rect 84649 96810 84661 96813
rect 86532 96810 86538 96822
rect 84649 96782 86538 96810
rect 84649 96779 84661 96782
rect 84603 96773 84661 96779
rect 84618 96742 84646 96773
rect 86532 96770 86538 96782
rect 86590 96770 86596 96822
rect 80150 96714 83174 96742
rect 83238 96714 84646 96742
rect 84971 96745 85029 96751
rect 80150 96702 80156 96714
rect 72735 96677 72793 96683
rect 72735 96643 72747 96677
rect 72781 96674 72793 96677
rect 83238 96674 83266 96714
rect 84971 96711 84983 96745
rect 85017 96742 85029 96745
rect 85336 96742 85342 96754
rect 85017 96714 85342 96742
rect 85017 96711 85029 96714
rect 84971 96705 85029 96711
rect 85336 96702 85342 96714
rect 85394 96742 85400 96754
rect 86624 96742 86630 96754
rect 85394 96714 86630 96742
rect 85394 96702 85400 96714
rect 86624 96702 86630 96714
rect 86682 96702 86688 96754
rect 72781 96646 83266 96674
rect 83298 96652 87806 96674
rect 72781 96643 72793 96646
rect 72735 96637 72793 96643
rect 62078 96578 66614 96606
rect 80095 96609 80153 96615
rect 80095 96575 80107 96609
rect 80141 96606 80153 96609
rect 80141 96578 82622 96606
rect 83298 96600 84916 96652
rect 84968 96600 84980 96652
rect 85032 96600 85044 96652
rect 85096 96600 85108 96652
rect 85160 96600 87806 96652
rect 83298 96578 87806 96600
rect 80141 96575 80153 96578
rect 80095 96569 80153 96575
rect 1708 96498 1714 96550
rect 1766 96538 1772 96550
rect 4100 96538 4106 96550
rect 1766 96510 4106 96538
rect 1766 96498 1772 96510
rect 4100 96498 4106 96510
rect 4158 96498 4164 96550
rect 4468 96498 4474 96550
rect 4526 96538 4532 96550
rect 5020 96538 5026 96550
rect 4526 96510 5026 96538
rect 4526 96498 4532 96510
rect 5020 96498 5026 96510
rect 5078 96538 5084 96550
rect 35012 96538 35018 96550
rect 5078 96510 35018 96538
rect 5078 96498 5084 96510
rect 35012 96498 35018 96510
rect 35070 96498 35076 96550
rect 38600 96498 38606 96550
rect 38658 96538 38664 96550
rect 61968 96538 61974 96550
rect 38658 96510 61974 96538
rect 38658 96498 38664 96510
rect 61968 96498 61974 96510
rect 62026 96498 62032 96550
rect 62520 96498 62526 96550
rect 62578 96538 62584 96550
rect 74388 96538 74394 96550
rect 62578 96510 74394 96538
rect 62578 96498 62584 96510
rect 74388 96498 74394 96510
rect 74446 96498 74452 96550
rect 77424 96498 77430 96550
rect 77482 96538 77488 96550
rect 82487 96541 82545 96547
rect 82487 96538 82499 96541
rect 77482 96510 82499 96538
rect 77482 96498 77488 96510
rect 82487 96507 82499 96510
rect 82533 96507 82545 96541
rect 82487 96501 82545 96507
rect 36852 96470 36858 96482
rect 5130 96442 36858 96470
rect 2168 96402 2174 96414
rect 2094 96374 2174 96402
rect 2094 96207 2122 96374
rect 2168 96362 2174 96374
rect 2226 96362 2232 96414
rect 2720 96362 2726 96414
rect 2778 96402 2784 96414
rect 5130 96402 5158 96442
rect 36852 96430 36858 96442
rect 36910 96430 36916 96482
rect 53044 96430 53050 96482
rect 53102 96470 53108 96482
rect 56816 96470 56822 96482
rect 53102 96442 56822 96470
rect 53102 96430 53108 96442
rect 56816 96430 56822 96442
rect 56874 96430 56880 96482
rect 62060 96430 62066 96482
rect 62118 96470 62124 96482
rect 66568 96470 66574 96482
rect 62118 96442 66574 96470
rect 62118 96430 62124 96442
rect 66568 96430 66574 96442
rect 66626 96430 66632 96482
rect 74759 96473 74817 96479
rect 74759 96439 74771 96473
rect 74805 96470 74817 96473
rect 81472 96470 81478 96482
rect 74805 96442 81478 96470
rect 74805 96439 74817 96442
rect 74759 96433 74817 96439
rect 81472 96430 81478 96442
rect 81530 96430 81536 96482
rect 82594 96470 82622 96578
rect 83864 96498 83870 96550
rect 83922 96538 83928 96550
rect 84140 96538 84146 96550
rect 83922 96510 84146 96538
rect 83922 96498 83928 96510
rect 84140 96498 84146 96510
rect 84198 96498 84204 96550
rect 85336 96470 85342 96482
rect 82594 96442 85342 96470
rect 85336 96430 85342 96442
rect 85394 96430 85400 96482
rect 2778 96374 5158 96402
rect 2778 96362 2784 96374
rect 15692 96362 15698 96414
rect 15750 96402 15756 96414
rect 24432 96402 24438 96414
rect 15750 96374 24438 96402
rect 15750 96362 15756 96374
rect 24432 96362 24438 96374
rect 24490 96362 24496 96414
rect 46512 96362 46518 96414
rect 46570 96402 46576 96414
rect 84416 96402 84422 96414
rect 46570 96374 84422 96402
rect 46570 96362 46576 96374
rect 84416 96362 84422 96374
rect 84474 96362 84480 96414
rect 3180 96334 3186 96346
rect 3141 96306 3186 96334
rect 3180 96294 3186 96306
rect 3238 96294 3244 96346
rect 3275 96337 3333 96343
rect 3275 96303 3287 96337
rect 3321 96334 3333 96337
rect 4011 96337 4069 96343
rect 4011 96334 4023 96337
rect 3321 96306 4023 96334
rect 3321 96303 3333 96306
rect 3275 96297 3333 96303
rect 4011 96303 4023 96306
rect 4057 96303 4069 96337
rect 4011 96297 4069 96303
rect 4284 96294 4290 96346
rect 4342 96334 4348 96346
rect 41820 96334 41826 96346
rect 4342 96306 41826 96334
rect 4342 96294 4348 96306
rect 41820 96294 41826 96306
rect 41878 96294 41884 96346
rect 44488 96294 44494 96346
rect 44546 96334 44552 96346
rect 82392 96334 82398 96346
rect 44546 96306 82398 96334
rect 44546 96294 44552 96306
rect 82392 96294 82398 96306
rect 82450 96294 82456 96346
rect 83772 96334 83778 96346
rect 83733 96306 83778 96334
rect 83772 96294 83778 96306
rect 83830 96294 83836 96346
rect 83864 96294 83870 96346
rect 83922 96334 83928 96346
rect 84235 96337 84293 96343
rect 84235 96334 84247 96337
rect 83922 96306 84247 96334
rect 83922 96294 83928 96306
rect 84235 96303 84247 96306
rect 84281 96334 84293 96337
rect 85152 96334 85158 96346
rect 84281 96306 85158 96334
rect 84281 96303 84293 96306
rect 84235 96297 84293 96303
rect 85152 96294 85158 96306
rect 85210 96294 85216 96346
rect 2168 96226 2174 96278
rect 2226 96266 2232 96278
rect 2226 96238 5894 96266
rect 2226 96226 2232 96238
rect 2079 96201 2137 96207
rect 2079 96167 2091 96201
rect 2125 96198 2137 96201
rect 2352 96198 2358 96210
rect 2125 96170 2358 96198
rect 2125 96167 2137 96170
rect 2079 96161 2137 96167
rect 2352 96158 2358 96170
rect 2410 96158 2416 96210
rect 2447 96201 2505 96207
rect 2447 96167 2459 96201
rect 2493 96198 2505 96201
rect 2738 96198 2766 96238
rect 2493 96170 2766 96198
rect 2815 96201 2873 96207
rect 2493 96167 2505 96170
rect 2447 96161 2505 96167
rect 2815 96167 2827 96201
rect 2861 96198 2873 96201
rect 3275 96201 3333 96207
rect 3275 96198 3287 96201
rect 2861 96170 3287 96198
rect 2861 96167 2873 96170
rect 2815 96161 2873 96167
rect 3275 96167 3287 96170
rect 3321 96167 3333 96201
rect 3275 96161 3333 96167
rect 3551 96201 3609 96207
rect 3551 96167 3563 96201
rect 3597 96198 3609 96201
rect 4284 96198 4290 96210
rect 3597 96170 4290 96198
rect 3597 96167 3609 96170
rect 3551 96161 3609 96167
rect 4284 96158 4290 96170
rect 4342 96158 4348 96210
rect 4011 96133 4069 96139
rect 38 96108 3902 96130
rect 38 96056 2916 96108
rect 2968 96056 2980 96108
rect 3032 96056 3044 96108
rect 3096 96056 3108 96108
rect 3160 96056 3902 96108
rect 4011 96099 4023 96133
rect 4057 96130 4069 96133
rect 5480 96130 5486 96142
rect 4057 96102 5486 96130
rect 4057 96099 4069 96102
rect 4011 96093 4069 96099
rect 5480 96090 5486 96102
rect 5538 96130 5544 96142
rect 5756 96130 5762 96142
rect 5538 96102 5762 96130
rect 5538 96090 5544 96102
rect 5756 96090 5762 96102
rect 5814 96090 5820 96142
rect 38 96034 3902 96056
rect 2628 95954 2634 96006
rect 2686 95994 2692 96006
rect 2815 95997 2873 96003
rect 2815 95994 2827 95997
rect 2686 95966 2827 95994
rect 2686 95954 2692 95966
rect 2815 95963 2827 95966
rect 2861 95963 2873 95997
rect 2815 95957 2873 95963
rect 3551 95997 3609 96003
rect 3551 95963 3563 95997
rect 3597 95994 3609 95997
rect 4652 95994 4658 96006
rect 3597 95966 4658 95994
rect 3597 95963 3609 95966
rect 3551 95957 3609 95963
rect 2830 95926 2858 95957
rect 4652 95954 4658 95966
rect 4710 95954 4716 96006
rect 5866 95994 5894 96238
rect 24984 96226 24990 96278
rect 25042 96266 25048 96278
rect 33540 96266 33546 96278
rect 25042 96238 33546 96266
rect 25042 96226 25048 96238
rect 33540 96226 33546 96238
rect 33598 96226 33604 96278
rect 34460 96226 34466 96278
rect 34518 96266 34524 96278
rect 45316 96266 45322 96278
rect 34518 96238 45322 96266
rect 34518 96226 34524 96238
rect 45316 96226 45322 96238
rect 45374 96226 45380 96278
rect 50192 96226 50198 96278
rect 50250 96266 50256 96278
rect 85980 96266 85986 96278
rect 50250 96238 85986 96266
rect 50250 96226 50256 96238
rect 85980 96226 85986 96238
rect 86038 96226 86044 96278
rect 47800 96158 47806 96210
rect 47858 96198 47864 96210
rect 82116 96198 82122 96210
rect 47858 96170 82122 96198
rect 47858 96158 47864 96170
rect 82116 96158 82122 96170
rect 82174 96158 82180 96210
rect 82487 96201 82545 96207
rect 82487 96167 82499 96201
rect 82533 96198 82545 96201
rect 85428 96198 85434 96210
rect 82533 96170 85434 96198
rect 82533 96167 82545 96170
rect 82487 96161 82545 96167
rect 85428 96158 85434 96170
rect 85486 96158 85492 96210
rect 51572 96090 51578 96142
rect 51630 96130 51636 96142
rect 82760 96130 82766 96142
rect 51630 96102 82766 96130
rect 51630 96090 51636 96102
rect 82760 96090 82766 96102
rect 82818 96090 82824 96142
rect 83298 96108 87806 96130
rect 37496 96022 37502 96074
rect 37554 96062 37560 96074
rect 53044 96062 53050 96074
rect 37554 96034 53050 96062
rect 37554 96022 37560 96034
rect 53044 96022 53050 96034
rect 53102 96022 53108 96074
rect 82208 96062 82214 96074
rect 53154 96034 82214 96062
rect 18360 95994 18366 96006
rect 5866 95966 18366 95994
rect 18360 95954 18366 95966
rect 18418 95954 18424 96006
rect 23420 95926 23426 95938
rect 2830 95898 23426 95926
rect 23420 95886 23426 95898
rect 23478 95886 23484 95938
rect 1708 95818 1714 95870
rect 1766 95858 1772 95870
rect 2352 95858 2358 95870
rect 1766 95830 2358 95858
rect 1766 95818 1772 95830
rect 2352 95818 2358 95830
rect 2410 95858 2416 95870
rect 23972 95858 23978 95870
rect 2410 95830 23978 95858
rect 2410 95818 2416 95830
rect 23972 95818 23978 95830
rect 24030 95818 24036 95870
rect 25999 95861 26057 95867
rect 25999 95858 26011 95861
rect 24082 95830 26011 95858
rect 24082 95790 24110 95830
rect 25999 95827 26011 95830
rect 26045 95827 26057 95861
rect 25999 95821 26057 95827
rect 43752 95818 43758 95870
rect 43810 95858 43816 95870
rect 53154 95858 53182 96034
rect 82208 96022 82214 96034
rect 82266 96022 82272 96074
rect 83298 96056 86916 96108
rect 86968 96056 86980 96108
rect 87032 96056 87044 96108
rect 87096 96056 87108 96108
rect 87160 96056 87806 96108
rect 83298 96034 87806 96056
rect 57920 95954 57926 96006
rect 57978 95994 57984 96006
rect 81196 95994 81202 96006
rect 57978 95966 81202 95994
rect 57978 95954 57984 95966
rect 81196 95954 81202 95966
rect 81254 95954 81260 96006
rect 83867 95997 83925 96003
rect 83867 95963 83879 95997
rect 83913 95994 83925 95997
rect 84140 95994 84146 96006
rect 83913 95966 84146 95994
rect 83913 95963 83925 95966
rect 83867 95957 83925 95963
rect 84140 95954 84146 95966
rect 84198 95954 84204 96006
rect 61784 95886 61790 95938
rect 61842 95926 61848 95938
rect 80276 95926 80282 95938
rect 61842 95898 80282 95926
rect 61842 95886 61848 95898
rect 80276 95886 80282 95898
rect 80334 95886 80340 95938
rect 43810 95830 53182 95858
rect 43810 95818 43816 95830
rect 62796 95818 62802 95870
rect 62854 95858 62860 95870
rect 81932 95858 81938 95870
rect 62854 95830 81938 95858
rect 62854 95818 62860 95830
rect 81932 95818 81938 95830
rect 81990 95818 81996 95870
rect 22150 95762 24110 95790
rect 2447 95725 2505 95731
rect 2447 95691 2459 95725
rect 2493 95722 2505 95725
rect 4744 95722 4750 95734
rect 2493 95694 4750 95722
rect 2493 95691 2505 95694
rect 2447 95685 2505 95691
rect 4744 95682 4750 95694
rect 4802 95722 4808 95734
rect 14036 95722 14042 95734
rect 4802 95694 14042 95722
rect 4802 95682 4808 95694
rect 14036 95682 14042 95694
rect 14094 95682 14100 95734
rect 38 95564 3902 95586
rect 38 95512 916 95564
rect 968 95512 980 95564
rect 1032 95512 1044 95564
rect 1096 95512 1108 95564
rect 1160 95512 3902 95564
rect 5480 95546 5486 95598
rect 5538 95586 5544 95598
rect 22150 95586 22178 95762
rect 25720 95750 25726 95802
rect 25778 95790 25784 95802
rect 28299 95793 28357 95799
rect 28299 95790 28311 95793
rect 25778 95762 28311 95790
rect 25778 95750 25784 95762
rect 28299 95759 28311 95762
rect 28345 95759 28357 95793
rect 28299 95753 28357 95759
rect 63440 95750 63446 95802
rect 63498 95790 63504 95802
rect 82576 95790 82582 95802
rect 63498 95762 82582 95790
rect 63498 95750 63504 95762
rect 82576 95750 82582 95762
rect 82634 95750 82640 95802
rect 68960 95682 68966 95734
rect 69018 95722 69024 95734
rect 81288 95722 81294 95734
rect 69018 95694 81294 95722
rect 69018 95682 69024 95694
rect 81288 95682 81294 95694
rect 81346 95682 81352 95734
rect 34920 95654 34926 95666
rect 5538 95558 22178 95586
rect 22242 95626 34926 95654
rect 5538 95546 5544 95558
rect 38 95490 3902 95512
rect 18360 95478 18366 95530
rect 18418 95518 18424 95530
rect 22242 95518 22270 95626
rect 34920 95614 34926 95626
rect 34978 95614 34984 95666
rect 47616 95614 47622 95666
rect 47674 95654 47680 95666
rect 47674 95626 62474 95654
rect 47674 95614 47680 95626
rect 25999 95589 26057 95595
rect 25999 95555 26011 95589
rect 26045 95586 26057 95589
rect 38140 95586 38146 95598
rect 26045 95558 38146 95586
rect 26045 95555 26057 95558
rect 25999 95549 26057 95555
rect 38140 95546 38146 95558
rect 38198 95546 38204 95598
rect 57831 95589 57889 95595
rect 57831 95555 57843 95589
rect 57877 95586 57889 95589
rect 62336 95586 62342 95598
rect 57877 95558 62342 95586
rect 57877 95555 57889 95558
rect 57831 95549 57889 95555
rect 62336 95546 62342 95558
rect 62394 95546 62400 95598
rect 18418 95490 22270 95518
rect 18418 95478 18424 95490
rect 26640 95478 26646 95530
rect 26698 95518 26704 95530
rect 35012 95518 35018 95530
rect 26698 95490 35018 95518
rect 26698 95478 26704 95490
rect 35012 95478 35018 95490
rect 35070 95478 35076 95530
rect 51480 95478 51486 95530
rect 51538 95518 51544 95530
rect 61968 95518 61974 95530
rect 51538 95490 61974 95518
rect 51538 95478 51544 95490
rect 61968 95478 61974 95490
rect 62026 95478 62032 95530
rect 3183 95453 3241 95459
rect 3183 95419 3195 95453
rect 3229 95450 3241 95453
rect 4836 95450 4842 95462
rect 3229 95422 4842 95450
rect 3229 95419 3241 95422
rect 3183 95413 3241 95419
rect 4836 95410 4842 95422
rect 4894 95450 4900 95462
rect 11828 95450 11834 95462
rect 4894 95422 11834 95450
rect 4894 95410 4900 95422
rect 11828 95410 11834 95422
rect 11886 95410 11892 95462
rect 36208 95410 36214 95462
rect 36266 95450 36272 95462
rect 45316 95450 45322 95462
rect 36266 95422 45322 95450
rect 36266 95410 36272 95422
rect 45316 95410 45322 95422
rect 45374 95410 45380 95462
rect 53136 95410 53142 95462
rect 53194 95450 53200 95462
rect 57831 95453 57889 95459
rect 57831 95450 57843 95453
rect 53194 95422 57843 95450
rect 53194 95410 53200 95422
rect 57831 95419 57843 95422
rect 57877 95419 57889 95453
rect 62244 95450 62250 95462
rect 57831 95413 57889 95419
rect 57938 95422 62250 95450
rect 3551 95385 3609 95391
rect 3551 95351 3563 95385
rect 3597 95382 3609 95385
rect 3732 95382 3738 95394
rect 3597 95354 3738 95382
rect 3597 95351 3609 95354
rect 3551 95345 3609 95351
rect 3732 95342 3738 95354
rect 3790 95382 3796 95394
rect 19832 95382 19838 95394
rect 3790 95354 19838 95382
rect 3790 95342 3796 95354
rect 19832 95342 19838 95354
rect 19890 95382 19896 95394
rect 20752 95382 20758 95394
rect 19890 95354 20758 95382
rect 19890 95342 19896 95354
rect 20752 95342 20758 95354
rect 20810 95342 20816 95394
rect 28299 95385 28357 95391
rect 28299 95351 28311 95385
rect 28345 95382 28357 95385
rect 45408 95382 45414 95394
rect 28345 95354 45414 95382
rect 28345 95351 28357 95354
rect 28299 95345 28357 95351
rect 45408 95342 45414 95354
rect 45466 95342 45472 95394
rect 53228 95342 53234 95394
rect 53286 95382 53292 95394
rect 57938 95382 57966 95422
rect 62244 95410 62250 95422
rect 62302 95410 62308 95462
rect 62446 95450 62474 95626
rect 71168 95614 71174 95666
rect 71226 95654 71232 95666
rect 80184 95654 80190 95666
rect 71226 95626 80190 95654
rect 71226 95614 71232 95626
rect 80184 95614 80190 95626
rect 80242 95614 80248 95666
rect 69052 95546 69058 95598
rect 69110 95586 69116 95598
rect 77424 95586 77430 95598
rect 69110 95558 77430 95586
rect 69110 95546 69116 95558
rect 77424 95546 77430 95558
rect 77482 95546 77488 95598
rect 83298 95564 87806 95586
rect 83298 95512 84916 95564
rect 84968 95512 84980 95564
rect 85032 95512 85044 95564
rect 85096 95512 85108 95564
rect 85160 95512 87806 95564
rect 83298 95490 87806 95512
rect 68868 95450 68874 95462
rect 62446 95422 68874 95450
rect 68868 95410 68874 95422
rect 68926 95410 68932 95462
rect 77424 95410 77430 95462
rect 77482 95450 77488 95462
rect 84692 95450 84698 95462
rect 77482 95422 84698 95450
rect 77482 95410 77488 95422
rect 84692 95410 84698 95422
rect 84750 95410 84756 95462
rect 53286 95354 57966 95382
rect 53286 95342 53292 95354
rect 58012 95342 58018 95394
rect 58070 95382 58076 95394
rect 69236 95382 69242 95394
rect 58070 95354 69242 95382
rect 58070 95342 58076 95354
rect 69236 95342 69242 95354
rect 69294 95342 69300 95394
rect 80092 95342 80098 95394
rect 80150 95382 80156 95394
rect 86256 95382 86262 95394
rect 80150 95354 86262 95382
rect 80150 95342 80156 95354
rect 86256 95342 86262 95354
rect 86314 95342 86320 95394
rect 4192 95274 4198 95326
rect 4250 95314 4256 95326
rect 31148 95314 31154 95326
rect 4250 95286 31154 95314
rect 4250 95274 4256 95286
rect 31148 95274 31154 95286
rect 31206 95274 31212 95326
rect 35656 95274 35662 95326
rect 35714 95314 35720 95326
rect 51756 95314 51762 95326
rect 35714 95286 51762 95314
rect 35714 95274 35720 95286
rect 51756 95274 51762 95286
rect 51814 95274 51820 95326
rect 53044 95274 53050 95326
rect 53102 95314 53108 95326
rect 69880 95314 69886 95326
rect 53102 95286 69886 95314
rect 53102 95274 53108 95286
rect 69880 95274 69886 95286
rect 69938 95274 69944 95326
rect 4284 95206 4290 95258
rect 4342 95246 4348 95258
rect 4342 95218 4606 95246
rect 4342 95206 4348 95218
rect 2720 95138 2726 95190
rect 2778 95178 2784 95190
rect 4578 95178 4606 95218
rect 4836 95206 4842 95258
rect 4894 95246 4900 95258
rect 36300 95246 36306 95258
rect 4894 95218 36306 95246
rect 4894 95206 4900 95218
rect 36300 95206 36306 95218
rect 36358 95206 36364 95258
rect 58104 95246 58110 95258
rect 41286 95218 58110 95246
rect 16980 95178 16986 95190
rect 2778 95150 4514 95178
rect 2778 95138 2784 95150
rect 4486 95122 4514 95150
rect 4578 95150 16986 95178
rect 4578 95122 4606 95150
rect 16980 95138 16986 95150
rect 17038 95138 17044 95190
rect 24432 95138 24438 95190
rect 24490 95178 24496 95190
rect 29768 95178 29774 95190
rect 24490 95150 29774 95178
rect 24490 95138 24496 95150
rect 29768 95138 29774 95150
rect 29826 95138 29832 95190
rect 4468 95070 4474 95122
rect 4526 95070 4532 95122
rect 4560 95070 4566 95122
rect 4618 95070 4624 95122
rect 4744 95070 4750 95122
rect 4802 95110 4808 95122
rect 5020 95110 5026 95122
rect 4802 95082 5026 95110
rect 4802 95070 4808 95082
rect 5020 95070 5026 95082
rect 5078 95070 5084 95122
rect 8148 95070 8154 95122
rect 8206 95110 8212 95122
rect 41286 95110 41314 95218
rect 58104 95206 58110 95218
rect 58162 95206 58168 95258
rect 59392 95206 59398 95258
rect 59450 95246 59456 95258
rect 63348 95246 63354 95258
rect 59450 95218 63354 95246
rect 59450 95206 59456 95218
rect 63348 95206 63354 95218
rect 63406 95206 63412 95258
rect 68408 95206 68414 95258
rect 68466 95246 68472 95258
rect 85152 95246 85158 95258
rect 68466 95218 85158 95246
rect 68466 95206 68472 95218
rect 85152 95206 85158 95218
rect 85210 95206 85216 95258
rect 48720 95138 48726 95190
rect 48778 95178 48784 95190
rect 54148 95178 54154 95190
rect 48778 95150 54154 95178
rect 48778 95138 48784 95150
rect 54148 95138 54154 95150
rect 54206 95138 54212 95190
rect 80184 95138 80190 95190
rect 80242 95178 80248 95190
rect 84048 95178 84054 95190
rect 80242 95150 84054 95178
rect 80242 95138 80248 95150
rect 84048 95138 84054 95150
rect 84106 95138 84112 95190
rect 8206 95082 41314 95110
rect 8206 95070 8212 95082
rect 49088 95070 49094 95122
rect 49146 95110 49152 95122
rect 51664 95110 51670 95122
rect 49146 95082 51670 95110
rect 49146 95070 49152 95082
rect 51664 95070 51670 95082
rect 51722 95070 51728 95122
rect 51759 95113 51817 95119
rect 51759 95079 51771 95113
rect 51805 95110 51817 95113
rect 58012 95110 58018 95122
rect 51805 95082 58018 95110
rect 51805 95079 51817 95082
rect 51759 95073 51817 95079
rect 58012 95070 58018 95082
rect 58070 95070 58076 95122
rect 66476 95070 66482 95122
rect 66534 95110 66540 95122
rect 71076 95110 71082 95122
rect 66534 95082 71082 95110
rect 66534 95070 66540 95082
rect 71076 95070 71082 95082
rect 71134 95070 71140 95122
rect 38 95020 3902 95042
rect 38 94968 2916 95020
rect 2968 94968 2980 95020
rect 3032 94968 3044 95020
rect 3096 94968 3108 95020
rect 3160 94968 3902 95020
rect 37312 95002 37318 95054
rect 37370 95042 37376 95054
rect 53044 95042 53050 95054
rect 37370 95014 53050 95042
rect 37370 95002 37376 95014
rect 53044 95002 53050 95014
rect 53102 95002 53108 95054
rect 55807 95045 55865 95051
rect 55807 95011 55819 95045
rect 55853 95042 55865 95045
rect 77424 95042 77430 95054
rect 55853 95014 77430 95042
rect 55853 95011 55865 95014
rect 55807 95005 55865 95011
rect 77424 95002 77430 95014
rect 77482 95002 77488 95054
rect 83298 95020 87806 95042
rect 38 94946 3902 94968
rect 38784 94934 38790 94986
rect 38842 94974 38848 94986
rect 46607 94977 46665 94983
rect 46607 94974 46619 94977
rect 38842 94946 46619 94974
rect 38842 94934 38848 94946
rect 46607 94943 46619 94946
rect 46653 94943 46665 94977
rect 82024 94974 82030 94986
rect 46607 94937 46665 94943
rect 56926 94946 82030 94974
rect 3364 94866 3370 94918
rect 3422 94906 3428 94918
rect 8148 94906 8154 94918
rect 3422 94878 8154 94906
rect 3422 94866 3428 94878
rect 8148 94866 8154 94878
rect 8206 94866 8212 94918
rect 25904 94866 25910 94918
rect 25962 94906 25968 94918
rect 29676 94906 29682 94918
rect 25962 94878 29682 94906
rect 25962 94866 25968 94878
rect 29676 94866 29682 94878
rect 29734 94866 29740 94918
rect 43936 94866 43942 94918
rect 43994 94906 44000 94918
rect 51020 94906 51026 94918
rect 43994 94878 51026 94906
rect 43994 94866 44000 94878
rect 51020 94866 51026 94878
rect 51078 94866 51084 94918
rect 54148 94866 54154 94918
rect 54206 94906 54212 94918
rect 56926 94906 56954 94946
rect 82024 94934 82030 94946
rect 82082 94934 82088 94986
rect 83298 94968 86916 95020
rect 86968 94968 86980 95020
rect 87032 94968 87044 95020
rect 87096 94968 87108 95020
rect 87160 94968 87806 95020
rect 83298 94946 87806 94968
rect 54206 94878 56954 94906
rect 58935 94909 58993 94915
rect 54206 94866 54212 94878
rect 58935 94875 58947 94909
rect 58981 94906 58993 94909
rect 84600 94906 84606 94918
rect 58981 94878 84606 94906
rect 58981 94875 58993 94878
rect 58935 94869 58993 94875
rect 84600 94866 84606 94878
rect 84658 94866 84664 94918
rect 4928 94798 4934 94850
rect 4986 94838 4992 94850
rect 11092 94838 11098 94850
rect 4986 94810 11098 94838
rect 4986 94798 4992 94810
rect 11092 94798 11098 94810
rect 11150 94798 11156 94850
rect 50376 94798 50382 94850
rect 50434 94838 50440 94850
rect 50434 94810 60082 94838
rect 50434 94798 50440 94810
rect 1616 94730 1622 94782
rect 1674 94770 1680 94782
rect 1892 94770 1898 94782
rect 1674 94742 1898 94770
rect 1674 94730 1680 94742
rect 1892 94730 1898 94742
rect 1950 94770 1956 94782
rect 25996 94770 26002 94782
rect 1950 94742 26002 94770
rect 1950 94730 1956 94742
rect 25996 94730 26002 94742
rect 26054 94730 26060 94782
rect 50284 94730 50290 94782
rect 50342 94770 50348 94782
rect 50342 94742 56770 94770
rect 50342 94730 50348 94742
rect 4011 94705 4069 94711
rect 4011 94671 4023 94705
rect 4057 94702 4069 94705
rect 20844 94702 20850 94714
rect 4057 94674 20850 94702
rect 4057 94671 4069 94674
rect 4011 94665 4069 94671
rect 20844 94662 20850 94674
rect 20902 94662 20908 94714
rect 30688 94662 30694 94714
rect 30746 94702 30752 94714
rect 38784 94702 38790 94714
rect 30746 94674 38790 94702
rect 30746 94662 30752 94674
rect 38784 94662 38790 94674
rect 38842 94662 38848 94714
rect 41728 94662 41734 94714
rect 41786 94702 41792 94714
rect 55715 94705 55773 94711
rect 55715 94702 55727 94705
rect 41786 94674 55727 94702
rect 41786 94662 41792 94674
rect 55715 94671 55727 94674
rect 55761 94671 55773 94705
rect 56742 94702 56770 94742
rect 56816 94730 56822 94782
rect 56874 94770 56880 94782
rect 60054 94770 60082 94810
rect 62152 94798 62158 94850
rect 62210 94838 62216 94850
rect 69144 94838 69150 94850
rect 62210 94810 69150 94838
rect 62210 94798 62216 94810
rect 69144 94798 69150 94810
rect 69202 94798 69208 94850
rect 69239 94841 69297 94847
rect 69239 94807 69251 94841
rect 69285 94838 69297 94841
rect 83312 94838 83318 94850
rect 69285 94810 83318 94838
rect 69285 94807 69297 94810
rect 69239 94801 69297 94807
rect 83312 94798 83318 94810
rect 83370 94798 83376 94850
rect 69052 94770 69058 94782
rect 56874 94742 59898 94770
rect 60054 94742 69058 94770
rect 56874 94730 56880 94742
rect 59671 94705 59729 94711
rect 59671 94702 59683 94705
rect 56742 94674 59683 94702
rect 55715 94665 55773 94671
rect 59671 94671 59683 94674
rect 59717 94671 59729 94705
rect 59671 94665 59729 94671
rect 2260 94594 2266 94646
rect 2318 94634 2324 94646
rect 2628 94634 2634 94646
rect 2318 94606 2634 94634
rect 2318 94594 2324 94606
rect 2628 94594 2634 94606
rect 2686 94634 2692 94646
rect 27284 94634 27290 94646
rect 2686 94606 27290 94634
rect 2686 94594 2692 94606
rect 27284 94594 27290 94606
rect 27342 94594 27348 94646
rect 29768 94594 29774 94646
rect 29826 94634 29832 94646
rect 40164 94634 40170 94646
rect 29826 94606 40170 94634
rect 29826 94594 29832 94606
rect 40164 94594 40170 94606
rect 40222 94594 40228 94646
rect 46607 94637 46665 94643
rect 46607 94603 46619 94637
rect 46653 94634 46665 94637
rect 51759 94637 51817 94643
rect 51759 94634 51771 94637
rect 46653 94606 51771 94634
rect 46653 94603 46665 94606
rect 46607 94597 46665 94603
rect 51759 94603 51771 94606
rect 51805 94603 51817 94637
rect 51759 94597 51817 94603
rect 52952 94594 52958 94646
rect 53010 94634 53016 94646
rect 58935 94637 58993 94643
rect 58935 94634 58947 94637
rect 53010 94606 58947 94634
rect 53010 94594 53016 94606
rect 58935 94603 58947 94606
rect 58981 94603 58993 94637
rect 59870 94634 59898 94742
rect 69052 94730 69058 94742
rect 69110 94730 69116 94782
rect 77979 94773 78037 94779
rect 77979 94739 77991 94773
rect 78025 94770 78037 94773
rect 82300 94770 82306 94782
rect 78025 94742 82306 94770
rect 78025 94739 78037 94742
rect 77979 94733 78037 94739
rect 82300 94730 82306 94742
rect 82358 94730 82364 94782
rect 82760 94730 82766 94782
rect 82818 94770 82824 94782
rect 85704 94770 85710 94782
rect 82818 94742 85710 94770
rect 82818 94730 82824 94742
rect 85704 94730 85710 94742
rect 85762 94730 85768 94782
rect 59947 94705 60005 94711
rect 59947 94671 59959 94705
rect 59993 94702 60005 94705
rect 68408 94702 68414 94714
rect 59993 94674 68414 94702
rect 59993 94671 60005 94674
rect 59947 94665 60005 94671
rect 68408 94662 68414 94674
rect 68466 94662 68472 94714
rect 68500 94662 68506 94714
rect 68558 94702 68564 94714
rect 70984 94702 70990 94714
rect 68558 94674 70990 94702
rect 68558 94662 68564 94674
rect 70984 94662 70990 94674
rect 71042 94662 71048 94714
rect 72456 94662 72462 94714
rect 72514 94702 72520 94714
rect 78163 94705 78221 94711
rect 72514 94674 78114 94702
rect 72514 94662 72520 94674
rect 77979 94637 78037 94643
rect 77979 94634 77991 94637
rect 59870 94606 77991 94634
rect 58935 94597 58993 94603
rect 77979 94603 77991 94606
rect 78025 94603 78037 94637
rect 78086 94634 78114 94674
rect 78163 94671 78175 94705
rect 78209 94702 78221 94705
rect 83404 94702 83410 94714
rect 78209 94674 83410 94702
rect 78209 94671 78221 94674
rect 78163 94665 78221 94671
rect 83404 94662 83410 94674
rect 83462 94662 83468 94714
rect 83956 94634 83962 94646
rect 78086 94606 83962 94634
rect 77979 94597 78037 94603
rect 83956 94594 83962 94606
rect 84014 94594 84020 94646
rect 5020 94526 5026 94578
rect 5078 94566 5084 94578
rect 32436 94566 32442 94578
rect 5078 94538 32442 94566
rect 5078 94526 5084 94538
rect 32436 94526 32442 94538
rect 32494 94526 32500 94578
rect 49088 94526 49094 94578
rect 49146 94566 49152 94578
rect 84784 94566 84790 94578
rect 49146 94538 84790 94566
rect 49146 94526 49152 94538
rect 84784 94526 84790 94538
rect 84842 94526 84848 94578
rect 4284 94498 4290 94510
rect 38 94476 3902 94498
rect 38 94424 916 94476
rect 968 94424 980 94476
rect 1032 94424 1044 94476
rect 1096 94424 1108 94476
rect 1160 94424 3902 94476
rect 38 94402 3902 94424
rect 3934 94470 4290 94498
rect 3364 94322 3370 94374
rect 3422 94362 3428 94374
rect 3732 94362 3738 94374
rect 3422 94334 3738 94362
rect 3422 94322 3428 94334
rect 3732 94322 3738 94334
rect 3790 94322 3796 94374
rect 2720 94254 2726 94306
rect 2778 94294 2784 94306
rect 3934 94294 3962 94470
rect 4284 94458 4290 94470
rect 4342 94498 4348 94510
rect 41452 94498 41458 94510
rect 4342 94470 41458 94498
rect 4342 94458 4348 94470
rect 41452 94458 41458 94470
rect 41510 94458 41516 94510
rect 42648 94458 42654 94510
rect 42706 94498 42712 94510
rect 72364 94498 72370 94510
rect 42706 94470 72370 94498
rect 42706 94458 42712 94470
rect 72364 94458 72370 94470
rect 72422 94458 72428 94510
rect 72548 94458 72554 94510
rect 72606 94498 72612 94510
rect 80184 94498 80190 94510
rect 72606 94470 80190 94498
rect 72606 94458 72612 94470
rect 80184 94458 80190 94470
rect 80242 94458 80248 94510
rect 83298 94476 87806 94498
rect 40072 94390 40078 94442
rect 40130 94430 40136 94442
rect 53136 94430 53142 94442
rect 40130 94402 53142 94430
rect 40130 94390 40136 94402
rect 53136 94390 53142 94402
rect 53194 94390 53200 94442
rect 54240 94390 54246 94442
rect 54298 94430 54304 94442
rect 55807 94433 55865 94439
rect 55807 94430 55819 94433
rect 54298 94402 55819 94430
rect 54298 94390 54304 94402
rect 55807 94399 55819 94402
rect 55853 94399 55865 94433
rect 55807 94393 55865 94399
rect 63256 94390 63262 94442
rect 63314 94430 63320 94442
rect 64639 94433 64697 94439
rect 64639 94430 64651 94433
rect 63314 94402 64651 94430
rect 63314 94390 63320 94402
rect 64639 94399 64651 94402
rect 64685 94399 64697 94433
rect 64639 94393 64697 94399
rect 66476 94390 66482 94442
rect 66534 94430 66540 94442
rect 70984 94430 70990 94442
rect 66534 94402 70990 94430
rect 66534 94390 66540 94402
rect 70984 94390 70990 94402
rect 71042 94390 71048 94442
rect 74388 94390 74394 94442
rect 74446 94430 74452 94442
rect 81196 94430 81202 94442
rect 74446 94402 81202 94430
rect 74446 94390 74452 94402
rect 81196 94390 81202 94402
rect 81254 94390 81260 94442
rect 83298 94424 84916 94476
rect 84968 94424 84980 94476
rect 85032 94424 85044 94476
rect 85096 94424 85108 94476
rect 85160 94424 87806 94476
rect 83298 94402 87806 94424
rect 29768 94322 29774 94374
rect 29826 94362 29832 94374
rect 33448 94362 33454 94374
rect 29826 94334 33454 94362
rect 29826 94322 29832 94334
rect 33448 94322 33454 94334
rect 33506 94322 33512 94374
rect 51664 94322 51670 94374
rect 51722 94362 51728 94374
rect 84324 94362 84330 94374
rect 51722 94334 84330 94362
rect 51722 94322 51728 94334
rect 84324 94322 84330 94334
rect 84382 94322 84388 94374
rect 2778 94266 3962 94294
rect 2778 94254 2784 94266
rect 38048 94254 38054 94306
rect 38106 94294 38112 94306
rect 42648 94294 42654 94306
rect 38106 94266 42654 94294
rect 38106 94254 38112 94266
rect 42648 94254 42654 94266
rect 42706 94254 42712 94306
rect 55715 94297 55773 94303
rect 55715 94263 55727 94297
rect 55761 94294 55773 94297
rect 60772 94294 60778 94306
rect 55761 94266 60778 94294
rect 55761 94263 55773 94266
rect 55715 94257 55773 94263
rect 60772 94254 60778 94266
rect 60830 94254 60836 94306
rect 69052 94254 69058 94306
rect 69110 94294 69116 94306
rect 78163 94297 78221 94303
rect 78163 94294 78175 94297
rect 69110 94266 78175 94294
rect 69110 94254 69116 94266
rect 78163 94263 78175 94266
rect 78209 94263 78221 94297
rect 78163 94257 78221 94263
rect 3732 94186 3738 94238
rect 3790 94226 3796 94238
rect 4011 94229 4069 94235
rect 4011 94226 4023 94229
rect 3790 94198 4023 94226
rect 3790 94186 3796 94198
rect 4011 94195 4023 94198
rect 4057 94195 4069 94229
rect 4011 94189 4069 94195
rect 23328 94186 23334 94238
rect 23386 94226 23392 94238
rect 48812 94226 48818 94238
rect 23386 94198 48818 94226
rect 23386 94186 23392 94198
rect 48812 94186 48818 94198
rect 48870 94186 48876 94238
rect 69144 94186 69150 94238
rect 69202 94226 69208 94238
rect 73655 94229 73713 94235
rect 73655 94226 73667 94229
rect 69202 94198 73667 94226
rect 69202 94186 69208 94198
rect 73655 94195 73667 94198
rect 73701 94195 73713 94229
rect 73655 94189 73713 94195
rect 41268 94118 41274 94170
rect 41326 94158 41332 94170
rect 69788 94158 69794 94170
rect 41326 94130 69794 94158
rect 41326 94118 41332 94130
rect 69788 94118 69794 94130
rect 69846 94118 69852 94170
rect 72364 94118 72370 94170
rect 72422 94158 72428 94170
rect 84416 94158 84422 94170
rect 72422 94130 84422 94158
rect 72422 94118 72428 94130
rect 84416 94118 84422 94130
rect 84474 94118 84480 94170
rect 28388 94050 28394 94102
rect 28446 94090 28452 94102
rect 36300 94090 36306 94102
rect 28446 94062 36306 94090
rect 28446 94050 28452 94062
rect 36300 94050 36306 94062
rect 36358 94050 36364 94102
rect 45224 94050 45230 94102
rect 45282 94090 45288 94102
rect 84048 94090 84054 94102
rect 45282 94062 84054 94090
rect 45282 94050 45288 94062
rect 84048 94050 84054 94062
rect 84106 94050 84112 94102
rect 5848 93982 5854 94034
rect 5906 94022 5912 94034
rect 18268 94022 18274 94034
rect 5906 93994 18274 94022
rect 5906 93982 5912 93994
rect 18268 93982 18274 93994
rect 18326 93982 18332 94034
rect 24616 93982 24622 94034
rect 24674 94022 24680 94034
rect 38232 94022 38238 94034
rect 24674 93994 38238 94022
rect 24674 93982 24680 93994
rect 38232 93982 38238 93994
rect 38290 93982 38296 94034
rect 43936 93982 43942 94034
rect 43994 94022 44000 94034
rect 84140 94022 84146 94034
rect 43994 93994 84146 94022
rect 43994 93982 44000 93994
rect 84140 93982 84146 93994
rect 84198 93982 84204 94034
rect 38 93932 3902 93954
rect 38 93880 2916 93932
rect 2968 93880 2980 93932
rect 3032 93880 3044 93932
rect 3096 93880 3108 93932
rect 3160 93880 3902 93932
rect 18176 93914 18182 93966
rect 18234 93954 18240 93966
rect 48444 93954 48450 93966
rect 18234 93926 48450 93954
rect 18234 93914 18240 93926
rect 48444 93914 48450 93926
rect 48502 93914 48508 93966
rect 64639 93957 64697 93963
rect 64639 93923 64651 93957
rect 64685 93954 64697 93957
rect 72548 93954 72554 93966
rect 64685 93926 72554 93954
rect 64685 93923 64697 93926
rect 64639 93917 64697 93923
rect 72548 93914 72554 93926
rect 72606 93914 72612 93966
rect 83298 93932 87806 93954
rect 38 93858 3902 93880
rect 5388 93846 5394 93898
rect 5446 93886 5452 93898
rect 19832 93886 19838 93898
rect 5446 93858 19838 93886
rect 5446 93846 5452 93858
rect 19832 93846 19838 93858
rect 19890 93846 19896 93898
rect 46144 93846 46150 93898
rect 46202 93886 46208 93898
rect 81288 93886 81294 93898
rect 46202 93858 81294 93886
rect 46202 93846 46208 93858
rect 81288 93846 81294 93858
rect 81346 93846 81352 93898
rect 83298 93880 86916 93932
rect 86968 93880 86980 93932
rect 87032 93880 87044 93932
rect 87096 93880 87108 93932
rect 87160 93880 87806 93932
rect 83298 93858 87806 93880
rect 63348 93778 63354 93830
rect 63406 93818 63412 93830
rect 72456 93818 72462 93830
rect 63406 93790 72462 93818
rect 63406 93778 63412 93790
rect 72456 93778 72462 93790
rect 72514 93778 72520 93830
rect 38876 93710 38882 93762
rect 38934 93750 38940 93762
rect 53228 93750 53234 93762
rect 38934 93722 53234 93750
rect 38934 93710 38940 93722
rect 53228 93710 53234 93722
rect 53286 93710 53292 93762
rect 53688 93710 53694 93762
rect 53746 93750 53752 93762
rect 60036 93750 60042 93762
rect 53746 93722 60042 93750
rect 53746 93710 53752 93722
rect 60036 93710 60042 93722
rect 60094 93710 60100 93762
rect 62244 93710 62250 93762
rect 62302 93750 62308 93762
rect 83956 93750 83962 93762
rect 62302 93722 83962 93750
rect 62302 93710 62308 93722
rect 83956 93710 83962 93722
rect 84014 93710 84020 93762
rect 45316 93642 45322 93694
rect 45374 93682 45380 93694
rect 56356 93682 56362 93694
rect 45374 93654 56362 93682
rect 45374 93642 45380 93654
rect 56356 93642 56362 93654
rect 56414 93642 56420 93694
rect 60772 93642 60778 93694
rect 60830 93682 60836 93694
rect 68960 93682 68966 93694
rect 60830 93654 68966 93682
rect 60830 93642 60836 93654
rect 68960 93642 68966 93654
rect 69018 93642 69024 93694
rect 71076 93642 71082 93694
rect 71134 93682 71140 93694
rect 78436 93682 78442 93694
rect 71134 93654 78442 93682
rect 71134 93642 71140 93654
rect 78436 93642 78442 93654
rect 78494 93642 78500 93694
rect 34920 93574 34926 93626
rect 34978 93614 34984 93626
rect 84600 93614 84606 93626
rect 34978 93586 84606 93614
rect 34978 93574 34984 93586
rect 84600 93574 84606 93586
rect 84658 93574 84664 93626
rect 33632 93506 33638 93558
rect 33690 93546 33696 93558
rect 82668 93546 82674 93558
rect 33690 93518 82674 93546
rect 33690 93506 33696 93518
rect 82668 93506 82674 93518
rect 82726 93506 82732 93558
rect 42740 93438 42746 93490
rect 42798 93478 42804 93490
rect 42798 93450 55758 93478
rect 42798 93438 42804 93450
rect 55730 93410 55758 93450
rect 60496 93438 60502 93490
rect 60554 93478 60560 93490
rect 69239 93481 69297 93487
rect 69239 93478 69251 93481
rect 60554 93450 69251 93478
rect 60554 93438 60560 93450
rect 69239 93447 69251 93450
rect 69285 93447 69297 93481
rect 69239 93441 69297 93447
rect 78436 93438 78442 93490
rect 78494 93478 78500 93490
rect 82576 93478 82582 93490
rect 78494 93450 82582 93478
rect 78494 93438 78500 93450
rect 82576 93438 82582 93450
rect 82634 93478 82640 93490
rect 83775 93481 83833 93487
rect 83775 93478 83787 93481
rect 82634 93450 83787 93478
rect 82634 93438 82640 93450
rect 83775 93447 83787 93450
rect 83821 93447 83833 93481
rect 83775 93441 83833 93447
rect 63440 93410 63446 93422
rect 38 93388 3902 93410
rect 38 93336 916 93388
rect 968 93336 980 93388
rect 1032 93336 1044 93388
rect 1096 93336 1108 93388
rect 1160 93336 3902 93388
rect 55730 93382 63446 93410
rect 63440 93370 63446 93382
rect 63498 93370 63504 93422
rect 69880 93370 69886 93422
rect 69938 93410 69944 93422
rect 80184 93410 80190 93422
rect 69938 93382 80190 93410
rect 69938 93370 69944 93382
rect 80184 93370 80190 93382
rect 80242 93370 80248 93422
rect 83298 93388 87806 93410
rect 38 93314 3902 93336
rect 33448 93302 33454 93354
rect 33506 93342 33512 93354
rect 82208 93342 82214 93354
rect 33506 93314 82214 93342
rect 33506 93302 33512 93314
rect 82208 93302 82214 93314
rect 82266 93302 82272 93354
rect 83298 93336 84916 93388
rect 84968 93336 84980 93388
rect 85032 93336 85044 93388
rect 85096 93336 85108 93388
rect 85160 93336 87806 93388
rect 83298 93314 87806 93336
rect 32344 93234 32350 93286
rect 32402 93274 32408 93286
rect 83404 93274 83410 93286
rect 32402 93246 83410 93274
rect 32402 93234 32408 93246
rect 83404 93234 83410 93246
rect 83462 93234 83468 93286
rect 31056 93166 31062 93218
rect 31114 93206 31120 93218
rect 83312 93206 83318 93218
rect 31114 93178 83318 93206
rect 31114 93166 31120 93178
rect 83312 93166 83318 93178
rect 83370 93166 83376 93218
rect 48444 93098 48450 93150
rect 48502 93138 48508 93150
rect 62520 93138 62526 93150
rect 48502 93110 62526 93138
rect 48502 93098 48508 93110
rect 62520 93098 62526 93110
rect 62578 93098 62584 93150
rect 69236 93098 69242 93150
rect 69294 93138 69300 93150
rect 84232 93138 84238 93150
rect 69294 93110 84238 93138
rect 69294 93098 69300 93110
rect 84232 93098 84238 93110
rect 84290 93098 84296 93150
rect 45408 93030 45414 93082
rect 45466 93070 45472 93082
rect 63256 93070 63262 93082
rect 45466 93042 63262 93070
rect 45466 93030 45472 93042
rect 63256 93030 63262 93042
rect 63314 93030 63320 93082
rect 69788 93030 69794 93082
rect 69846 93070 69852 93082
rect 81291 93073 81349 93079
rect 81291 93070 81303 93073
rect 69846 93042 81303 93070
rect 69846 93030 69852 93042
rect 81291 93039 81303 93042
rect 81337 93039 81349 93073
rect 81291 93033 81349 93039
rect 36208 92962 36214 93014
rect 36266 93002 36272 93014
rect 84784 93002 84790 93014
rect 36266 92974 84790 93002
rect 36266 92962 36272 92974
rect 84784 92962 84790 92974
rect 84842 92962 84848 93014
rect 38784 92894 38790 92946
rect 38842 92934 38848 92946
rect 59947 92937 60005 92943
rect 59947 92934 59959 92937
rect 38842 92906 59959 92934
rect 38842 92894 38848 92906
rect 59947 92903 59959 92906
rect 59993 92903 60005 92937
rect 59947 92897 60005 92903
rect 60036 92894 60042 92946
rect 60094 92934 60100 92946
rect 71168 92934 71174 92946
rect 60094 92906 71174 92934
rect 60094 92894 60100 92906
rect 71168 92894 71174 92906
rect 71226 92894 71232 92946
rect 73744 92894 73750 92946
rect 73802 92934 73808 92946
rect 83772 92934 83778 92946
rect 73802 92906 83778 92934
rect 73802 92894 73808 92906
rect 83772 92894 83778 92906
rect 83830 92894 83836 92946
rect 38 92844 3902 92866
rect 38 92792 2916 92844
rect 2968 92792 2980 92844
rect 3032 92792 3044 92844
rect 3096 92792 3108 92844
rect 3160 92792 3902 92844
rect 51756 92826 51762 92878
rect 51814 92866 51820 92878
rect 62428 92866 62434 92878
rect 51814 92838 62434 92866
rect 51814 92826 51820 92838
rect 62428 92826 62434 92838
rect 62486 92826 62492 92878
rect 83298 92844 87806 92866
rect 38 92770 3902 92792
rect 59947 92801 60005 92807
rect 59947 92767 59959 92801
rect 59993 92798 60005 92801
rect 60864 92798 60870 92810
rect 59993 92770 60870 92798
rect 59993 92767 60005 92770
rect 59947 92761 60005 92767
rect 60864 92758 60870 92770
rect 60922 92758 60928 92810
rect 81196 92758 81202 92810
rect 81254 92798 81260 92810
rect 81932 92798 81938 92810
rect 81254 92770 81938 92798
rect 81254 92758 81260 92770
rect 81932 92758 81938 92770
rect 81990 92758 81996 92810
rect 83298 92792 86916 92844
rect 86968 92792 86980 92844
rect 87032 92792 87044 92844
rect 87096 92792 87108 92844
rect 87160 92792 87806 92844
rect 83298 92770 87806 92792
rect 62336 92690 62342 92742
rect 62394 92730 62400 92742
rect 84324 92730 84330 92742
rect 62394 92702 84330 92730
rect 62394 92690 62400 92702
rect 84324 92690 84330 92702
rect 84382 92690 84388 92742
rect 68868 92622 68874 92674
rect 68926 92662 68932 92674
rect 85152 92662 85158 92674
rect 68926 92634 85158 92662
rect 68926 92622 68932 92634
rect 85152 92622 85158 92634
rect 85210 92622 85216 92674
rect 55344 92554 55350 92606
rect 55402 92594 55408 92606
rect 69052 92594 69058 92606
rect 55402 92566 69058 92594
rect 55402 92554 55408 92566
rect 69052 92554 69058 92566
rect 69110 92554 69116 92606
rect 80184 92554 80190 92606
rect 80242 92594 80248 92606
rect 81383 92597 81441 92603
rect 81383 92594 81395 92597
rect 80242 92566 81395 92594
rect 80242 92554 80248 92566
rect 81383 92563 81395 92566
rect 81429 92563 81441 92597
rect 81383 92557 81441 92563
rect 40164 92486 40170 92538
rect 40222 92526 40228 92538
rect 40222 92498 80046 92526
rect 40222 92486 40228 92498
rect 80018 92458 80046 92498
rect 80092 92486 80098 92538
rect 80150 92526 80156 92538
rect 82024 92526 82030 92538
rect 80150 92498 82030 92526
rect 80150 92486 80156 92498
rect 82024 92486 82030 92498
rect 82082 92486 82088 92538
rect 82760 92458 82766 92470
rect 80018 92430 82766 92458
rect 82760 92418 82766 92430
rect 82818 92418 82824 92470
rect 81383 92393 81441 92399
rect 81383 92359 81395 92393
rect 81429 92390 81441 92393
rect 83864 92390 83870 92402
rect 81429 92362 83870 92390
rect 81429 92359 81441 92362
rect 81383 92353 81441 92359
rect 83864 92350 83870 92362
rect 83922 92350 83928 92402
rect 38 92300 3902 92322
rect 38 92248 916 92300
rect 968 92248 980 92300
rect 1032 92248 1044 92300
rect 1096 92248 1108 92300
rect 1160 92248 3902 92300
rect 38 92226 3902 92248
rect 83298 92300 87806 92322
rect 83298 92248 84916 92300
rect 84968 92248 84980 92300
rect 85032 92248 85044 92300
rect 85096 92248 85108 92300
rect 85160 92248 87806 92300
rect 83298 92226 87806 92248
rect 81291 92189 81349 92195
rect 81291 92155 81303 92189
rect 81337 92186 81349 92189
rect 84692 92186 84698 92198
rect 81337 92158 84698 92186
rect 81337 92155 81349 92158
rect 81291 92149 81349 92155
rect 84692 92146 84698 92158
rect 84750 92146 84756 92198
rect 81288 92010 81294 92062
rect 81346 92050 81352 92062
rect 85152 92050 85158 92062
rect 81346 92022 85158 92050
rect 81346 92010 81352 92022
rect 85152 92010 85158 92022
rect 85210 92010 85216 92062
rect 83956 91942 83962 91994
rect 84014 91982 84020 91994
rect 84508 91982 84514 91994
rect 84014 91954 84514 91982
rect 84014 91942 84020 91954
rect 84508 91942 84514 91954
rect 84566 91942 84572 91994
rect 83867 91849 83925 91855
rect 83867 91815 83879 91849
rect 83913 91846 83925 91849
rect 83956 91846 83962 91858
rect 83913 91818 83962 91846
rect 83913 91815 83925 91818
rect 83867 91809 83925 91815
rect 83956 91806 83962 91818
rect 84014 91806 84020 91858
rect 38 91756 3902 91778
rect 38 91704 2916 91756
rect 2968 91704 2980 91756
rect 3032 91704 3044 91756
rect 3096 91704 3108 91756
rect 3160 91704 3902 91756
rect 38 91682 3902 91704
rect 83298 91756 87806 91778
rect 83298 91704 86916 91756
rect 86968 91704 86980 91756
rect 87032 91704 87044 91756
rect 87096 91704 87108 91756
rect 87160 91704 87806 91756
rect 83298 91682 87806 91704
rect 38 91212 3902 91234
rect 38 91160 916 91212
rect 968 91160 980 91212
rect 1032 91160 1044 91212
rect 1096 91160 1108 91212
rect 1160 91160 3902 91212
rect 38 91138 3902 91160
rect 83298 91212 87806 91234
rect 83298 91160 84916 91212
rect 84968 91160 84980 91212
rect 85032 91160 85044 91212
rect 85096 91160 85108 91212
rect 85160 91160 87806 91212
rect 83298 91138 87806 91160
rect 38 90668 3902 90690
rect 38 90616 2916 90668
rect 2968 90616 2980 90668
rect 3032 90616 3044 90668
rect 3096 90616 3108 90668
rect 3160 90616 3902 90668
rect 38 90594 3902 90616
rect 83298 90668 87806 90690
rect 83298 90616 86916 90668
rect 86968 90616 86980 90668
rect 87032 90616 87044 90668
rect 87096 90616 87108 90668
rect 87160 90616 87806 90668
rect 83298 90594 87806 90616
rect 38 90124 3902 90146
rect 38 90072 916 90124
rect 968 90072 980 90124
rect 1032 90072 1044 90124
rect 1096 90072 1108 90124
rect 1160 90072 3902 90124
rect 38 90050 3902 90072
rect 83298 90124 87806 90146
rect 83298 90072 84916 90124
rect 84968 90072 84980 90124
rect 85032 90072 85044 90124
rect 85096 90072 85108 90124
rect 85160 90072 87806 90124
rect 83298 90050 87806 90072
rect 3364 89902 3370 89954
rect 3422 89942 3428 89954
rect 4011 89945 4069 89951
rect 4011 89942 4023 89945
rect 3422 89914 4023 89942
rect 3422 89902 3428 89914
rect 4011 89911 4023 89914
rect 4057 89911 4069 89945
rect 5388 89942 5394 89954
rect 5349 89914 5394 89942
rect 4011 89905 4069 89911
rect 5388 89902 5394 89914
rect 5446 89902 5452 89954
rect 81380 89902 81386 89954
rect 81438 89942 81444 89954
rect 84048 89942 84054 89954
rect 81438 89914 84054 89942
rect 81438 89902 81444 89914
rect 84048 89902 84054 89914
rect 84106 89902 84112 89954
rect 38 89580 3902 89602
rect 38 89528 2916 89580
rect 2968 89528 2980 89580
rect 3032 89528 3044 89580
rect 3096 89528 3108 89580
rect 3160 89528 3902 89580
rect 38 89506 3902 89528
rect 83298 89580 87806 89602
rect 83298 89528 86916 89580
rect 86968 89528 86980 89580
rect 87032 89528 87044 89580
rect 87096 89528 87108 89580
rect 87160 89528 87806 89580
rect 83298 89506 87806 89528
rect 83864 89222 83870 89274
rect 83922 89262 83928 89274
rect 84140 89262 84146 89274
rect 83922 89234 84146 89262
rect 83922 89222 83928 89234
rect 84140 89222 84146 89234
rect 84198 89222 84204 89274
rect 38 89036 3902 89058
rect 38 88984 916 89036
rect 968 88984 980 89036
rect 1032 88984 1044 89036
rect 1096 88984 1108 89036
rect 1160 88984 3902 89036
rect 38 88962 3902 88984
rect 83298 89036 87806 89058
rect 83298 88984 84916 89036
rect 84968 88984 84980 89036
rect 85032 88984 85044 89036
rect 85096 88984 85108 89036
rect 85160 88984 87806 89036
rect 83298 88962 87806 88984
rect 2904 88610 2910 88662
rect 2962 88650 2968 88662
rect 2962 88622 3594 88650
rect 2962 88610 2968 88622
rect 3566 88591 3594 88622
rect 3732 88610 3738 88662
rect 3790 88650 3796 88662
rect 3916 88650 3922 88662
rect 3790 88622 3922 88650
rect 3790 88610 3796 88622
rect 3916 88610 3922 88622
rect 3974 88610 3980 88662
rect 3551 88585 3609 88591
rect 3551 88551 3563 88585
rect 3597 88582 3609 88585
rect 4100 88582 4106 88594
rect 3597 88554 4106 88582
rect 3597 88551 3609 88554
rect 3551 88545 3609 88551
rect 4100 88542 4106 88554
rect 4158 88542 4164 88594
rect 38 88492 3902 88514
rect 38 88440 2916 88492
rect 2968 88440 2980 88492
rect 3032 88440 3044 88492
rect 3096 88440 3108 88492
rect 3160 88440 3902 88492
rect 38 88418 3902 88440
rect 83298 88492 87806 88514
rect 83298 88440 86916 88492
rect 86968 88440 86980 88492
rect 87032 88440 87044 88492
rect 87096 88440 87108 88492
rect 87160 88440 87806 88492
rect 83298 88418 87806 88440
rect 83588 87998 83594 88050
rect 83646 88038 83652 88050
rect 83864 88038 83870 88050
rect 83646 88010 83870 88038
rect 83646 87998 83652 88010
rect 83864 87998 83870 88010
rect 83922 87998 83928 88050
rect 84140 87998 84146 88050
rect 84198 88038 84204 88050
rect 84416 88038 84422 88050
rect 84198 88010 84422 88038
rect 84198 87998 84204 88010
rect 84416 87998 84422 88010
rect 84474 87998 84480 88050
rect 38 87948 3902 87970
rect 38 87896 916 87948
rect 968 87896 980 87948
rect 1032 87896 1044 87948
rect 1096 87896 1108 87948
rect 1160 87896 3902 87948
rect 38 87874 3902 87896
rect 83298 87948 87806 87970
rect 83298 87896 84916 87948
rect 84968 87896 84980 87948
rect 85032 87896 85044 87948
rect 85096 87896 85108 87948
rect 85160 87896 87806 87948
rect 83298 87874 87806 87896
rect 3551 87837 3609 87843
rect 3551 87803 3563 87837
rect 3597 87834 3609 87837
rect 3732 87834 3738 87846
rect 3597 87806 3738 87834
rect 3597 87803 3609 87806
rect 3551 87797 3609 87803
rect 3732 87794 3738 87806
rect 3790 87794 3796 87846
rect 82668 87794 82674 87846
rect 82726 87834 82732 87846
rect 84140 87834 84146 87846
rect 82726 87806 84146 87834
rect 82726 87794 82732 87806
rect 84140 87794 84146 87806
rect 84198 87794 84204 87846
rect 38 87404 3902 87426
rect 38 87352 2916 87404
rect 2968 87352 2980 87404
rect 3032 87352 3044 87404
rect 3096 87352 3108 87404
rect 3160 87352 3902 87404
rect 38 87330 3902 87352
rect 83298 87404 87806 87426
rect 83298 87352 86916 87404
rect 86968 87352 86980 87404
rect 87032 87352 87044 87404
rect 87096 87352 87108 87404
rect 87160 87352 87806 87404
rect 83298 87330 87806 87352
rect 38 86860 3902 86882
rect 38 86808 916 86860
rect 968 86808 980 86860
rect 1032 86808 1044 86860
rect 1096 86808 1108 86860
rect 1160 86808 3902 86860
rect 38 86786 3902 86808
rect 83298 86860 87806 86882
rect 83298 86808 84916 86860
rect 84968 86808 84980 86860
rect 85032 86808 85044 86860
rect 85096 86808 85108 86860
rect 85160 86808 87806 86860
rect 83298 86786 87806 86808
rect 38 86316 3902 86338
rect 38 86264 2916 86316
rect 2968 86264 2980 86316
rect 3032 86264 3044 86316
rect 3096 86264 3108 86316
rect 3160 86264 3902 86316
rect 38 86242 3902 86264
rect 83298 86316 87806 86338
rect 83298 86264 86916 86316
rect 86968 86264 86980 86316
rect 87032 86264 87044 86316
rect 87096 86264 87108 86316
rect 87160 86264 87806 86316
rect 83298 86242 87806 86264
rect 3551 85865 3609 85871
rect 3551 85831 3563 85865
rect 3597 85862 3609 85865
rect 3824 85862 3830 85874
rect 3597 85834 3830 85862
rect 3597 85831 3609 85834
rect 3551 85825 3609 85831
rect 3824 85822 3830 85834
rect 3882 85862 3888 85874
rect 4192 85862 4198 85874
rect 3882 85834 4198 85862
rect 3882 85822 3888 85834
rect 4192 85822 4198 85834
rect 4250 85822 4256 85874
rect 84140 85822 84146 85874
rect 84198 85862 84204 85874
rect 84324 85862 84330 85874
rect 84198 85834 84330 85862
rect 84198 85822 84204 85834
rect 84324 85822 84330 85834
rect 84382 85822 84388 85874
rect 38 85772 3902 85794
rect 38 85720 916 85772
rect 968 85720 980 85772
rect 1032 85720 1044 85772
rect 1096 85720 1108 85772
rect 1160 85720 3902 85772
rect 38 85698 3902 85720
rect 83298 85772 87806 85794
rect 83298 85720 84916 85772
rect 84968 85720 84980 85772
rect 85032 85720 85044 85772
rect 85096 85720 85108 85772
rect 85160 85720 87806 85772
rect 83298 85698 87806 85720
rect 38 85228 3902 85250
rect 38 85176 2916 85228
rect 2968 85176 2980 85228
rect 3032 85176 3044 85228
rect 3096 85176 3108 85228
rect 3160 85176 3902 85228
rect 38 85154 3902 85176
rect 83298 85228 87806 85250
rect 83298 85176 86916 85228
rect 86968 85176 86980 85228
rect 87032 85176 87044 85228
rect 87096 85176 87108 85228
rect 87160 85176 87806 85228
rect 83298 85154 87806 85176
rect 3551 84845 3609 84851
rect 3551 84811 3563 84845
rect 3597 84842 3609 84845
rect 4008 84842 4014 84854
rect 3597 84814 4014 84842
rect 3597 84811 3609 84814
rect 3551 84805 3609 84811
rect 4008 84802 4014 84814
rect 4066 84802 4072 84854
rect 83404 84734 83410 84786
rect 83462 84774 83468 84786
rect 84140 84774 84146 84786
rect 83462 84746 84146 84774
rect 83462 84734 83468 84746
rect 84140 84734 84146 84746
rect 84198 84734 84204 84786
rect 38 84684 3902 84706
rect 38 84632 916 84684
rect 968 84632 980 84684
rect 1032 84632 1044 84684
rect 1096 84632 1108 84684
rect 1160 84632 3902 84684
rect 38 84610 3902 84632
rect 83298 84684 87806 84706
rect 83298 84632 84916 84684
rect 84968 84632 84980 84684
rect 85032 84632 85044 84684
rect 85096 84632 85108 84684
rect 85160 84632 87806 84684
rect 83298 84610 87806 84632
rect 38 84140 3902 84162
rect 38 84088 2916 84140
rect 2968 84088 2980 84140
rect 3032 84088 3044 84140
rect 3096 84088 3108 84140
rect 3160 84088 3902 84140
rect 38 84066 3902 84088
rect 83298 84140 87806 84162
rect 83298 84088 86916 84140
rect 86968 84088 86980 84140
rect 87032 84088 87044 84140
rect 87096 84088 87108 84140
rect 87160 84088 87806 84140
rect 83298 84066 87806 84088
rect 82208 83714 82214 83766
rect 82266 83754 82272 83766
rect 84324 83754 84330 83766
rect 82266 83726 84330 83754
rect 82266 83714 82272 83726
rect 84324 83714 84330 83726
rect 84382 83714 84388 83766
rect 38 83596 3902 83618
rect 38 83544 916 83596
rect 968 83544 980 83596
rect 1032 83544 1044 83596
rect 1096 83544 1108 83596
rect 1160 83544 3902 83596
rect 38 83522 3902 83544
rect 83298 83596 87806 83618
rect 83298 83544 84916 83596
rect 84968 83544 84980 83596
rect 85032 83544 85044 83596
rect 85096 83544 85108 83596
rect 85160 83544 87806 83596
rect 83298 83522 87806 83544
rect 5391 83417 5449 83423
rect 5391 83383 5403 83417
rect 5437 83414 5449 83417
rect 5572 83414 5578 83426
rect 5437 83386 5578 83414
rect 5437 83383 5449 83386
rect 5391 83377 5449 83383
rect 5572 83374 5578 83386
rect 5630 83374 5636 83426
rect 3548 83142 3554 83154
rect 3509 83114 3554 83142
rect 3548 83102 3554 83114
rect 3606 83102 3612 83154
rect 38 83052 3902 83074
rect 38 83000 2916 83052
rect 2968 83000 2980 83052
rect 3032 83000 3044 83052
rect 3096 83000 3108 83052
rect 3160 83000 3902 83052
rect 38 82978 3902 83000
rect 83298 83052 87806 83074
rect 83298 83000 86916 83052
rect 86968 83000 86980 83052
rect 87032 83000 87044 83052
rect 87096 83000 87108 83052
rect 87160 83000 87806 83052
rect 83298 82978 87806 83000
rect 38 82508 3902 82530
rect 38 82456 916 82508
rect 968 82456 980 82508
rect 1032 82456 1044 82508
rect 1096 82456 1108 82508
rect 1160 82456 3902 82508
rect 38 82434 3902 82456
rect 83298 82508 87806 82530
rect 83298 82456 84916 82508
rect 84968 82456 84980 82508
rect 85032 82456 85044 82508
rect 85096 82456 85108 82508
rect 85160 82456 87806 82508
rect 83298 82434 87806 82456
rect 2628 82218 2634 82270
rect 2686 82258 2692 82270
rect 3272 82258 3278 82270
rect 2686 82230 3278 82258
rect 2686 82218 2692 82230
rect 3272 82218 3278 82230
rect 3330 82258 3336 82270
rect 3330 82230 3502 82258
rect 3330 82218 3336 82230
rect 3474 82199 3502 82230
rect 3459 82193 3517 82199
rect 3459 82159 3471 82193
rect 3505 82159 3517 82193
rect 3459 82153 3517 82159
rect 38 81964 3902 81986
rect 38 81912 2916 81964
rect 2968 81912 2980 81964
rect 3032 81912 3044 81964
rect 3096 81912 3108 81964
rect 3160 81912 3902 81964
rect 38 81890 3902 81912
rect 83298 81964 87806 81986
rect 83298 81912 86916 81964
rect 86968 81912 86980 81964
rect 87032 81912 87044 81964
rect 87096 81912 87108 81964
rect 87160 81912 87806 81964
rect 83298 81890 87806 81912
rect 38 81420 3902 81442
rect 38 81368 916 81420
rect 968 81368 980 81420
rect 1032 81368 1044 81420
rect 1096 81368 1108 81420
rect 1160 81368 3902 81420
rect 38 81346 3902 81368
rect 83298 81420 87806 81442
rect 83298 81368 84916 81420
rect 84968 81368 84980 81420
rect 85032 81368 85044 81420
rect 85096 81368 85108 81420
rect 85160 81368 87806 81420
rect 83298 81346 87806 81368
rect 3364 80926 3370 80978
rect 3422 80966 3428 80978
rect 4011 80969 4069 80975
rect 4011 80966 4023 80969
rect 3422 80938 4023 80966
rect 3422 80926 3428 80938
rect 4011 80935 4023 80938
rect 4057 80935 4069 80969
rect 4011 80929 4069 80935
rect 83036 80926 83042 80978
rect 83094 80966 83100 80978
rect 83220 80966 83226 80978
rect 83094 80938 83226 80966
rect 83094 80926 83100 80938
rect 83220 80926 83226 80938
rect 83278 80926 83284 80978
rect 83864 80926 83870 80978
rect 83922 80966 83928 80978
rect 85244 80966 85250 80978
rect 83922 80938 85250 80966
rect 83922 80926 83928 80938
rect 85244 80926 85250 80938
rect 85302 80926 85308 80978
rect 38 80876 3902 80898
rect 38 80824 2916 80876
rect 2968 80824 2980 80876
rect 3032 80824 3044 80876
rect 3096 80824 3108 80876
rect 3160 80824 3902 80876
rect 38 80802 3902 80824
rect 83298 80876 87806 80898
rect 83298 80824 86916 80876
rect 86968 80824 86980 80876
rect 87032 80824 87044 80876
rect 87096 80824 87108 80876
rect 87160 80824 87806 80876
rect 83298 80802 87806 80824
rect 38 80332 3902 80354
rect 38 80280 916 80332
rect 968 80280 980 80332
rect 1032 80280 1044 80332
rect 1096 80280 1108 80332
rect 1160 80280 3902 80332
rect 38 80258 3902 80280
rect 83298 80332 87806 80354
rect 83298 80280 84916 80332
rect 84968 80280 84980 80332
rect 85032 80280 85044 80332
rect 85096 80280 85108 80332
rect 85160 80280 87806 80332
rect 83298 80258 87806 80280
rect 3551 79881 3609 79887
rect 3551 79847 3563 79881
rect 3597 79878 3609 79881
rect 3640 79878 3646 79890
rect 3597 79850 3646 79878
rect 3597 79847 3609 79850
rect 3551 79841 3609 79847
rect 3640 79838 3646 79850
rect 3698 79838 3704 79890
rect 38 79788 3902 79810
rect 38 79736 2916 79788
rect 2968 79736 2980 79788
rect 3032 79736 3044 79788
rect 3096 79736 3108 79788
rect 3160 79736 3902 79788
rect 38 79714 3902 79736
rect 83298 79788 87806 79810
rect 83298 79736 86916 79788
rect 86968 79736 86980 79788
rect 87032 79736 87044 79788
rect 87096 79736 87108 79788
rect 87160 79736 87806 79788
rect 83298 79714 87806 79736
rect 38 79244 3902 79266
rect 38 79192 916 79244
rect 968 79192 980 79244
rect 1032 79192 1044 79244
rect 1096 79192 1108 79244
rect 1160 79192 3902 79244
rect 38 79170 3902 79192
rect 83298 79244 87806 79266
rect 83298 79192 84916 79244
rect 84968 79192 84980 79244
rect 85032 79192 85044 79244
rect 85096 79192 85108 79244
rect 85160 79192 87806 79244
rect 83298 79170 87806 79192
rect 38 78700 3902 78722
rect 38 78648 2916 78700
rect 2968 78648 2980 78700
rect 3032 78648 3044 78700
rect 3096 78648 3108 78700
rect 3160 78648 3902 78700
rect 38 78626 3902 78648
rect 83298 78700 87806 78722
rect 83298 78648 86916 78700
rect 86968 78648 86980 78700
rect 87032 78648 87044 78700
rect 87096 78648 87108 78700
rect 87160 78648 87806 78700
rect 83298 78626 87806 78648
rect 38 78156 3902 78178
rect 38 78104 916 78156
rect 968 78104 980 78156
rect 1032 78104 1044 78156
rect 1096 78104 1108 78156
rect 1160 78104 3902 78156
rect 38 78082 3902 78104
rect 83298 78156 87806 78178
rect 83298 78104 84916 78156
rect 84968 78104 84980 78156
rect 85032 78104 85044 78156
rect 85096 78104 85108 78156
rect 85160 78104 87806 78156
rect 83298 78082 87806 78104
rect 38 77612 3902 77634
rect 38 77560 2916 77612
rect 2968 77560 2980 77612
rect 3032 77560 3044 77612
rect 3096 77560 3108 77612
rect 3160 77560 3902 77612
rect 38 77538 3902 77560
rect 83298 77612 87806 77634
rect 83298 77560 86916 77612
rect 86968 77560 86980 77612
rect 87032 77560 87044 77612
rect 87096 77560 87108 77612
rect 87160 77560 87806 77612
rect 83298 77538 87806 77560
rect 81656 77322 81662 77374
rect 81714 77362 81720 77374
rect 84600 77362 84606 77374
rect 81714 77334 84606 77362
rect 81714 77322 81720 77334
rect 84600 77322 84606 77334
rect 84658 77322 84664 77374
rect 38 77068 3902 77090
rect 38 77016 916 77068
rect 968 77016 980 77068
rect 1032 77016 1044 77068
rect 1096 77016 1108 77068
rect 1160 77016 3902 77068
rect 38 76994 3902 77016
rect 83298 77068 87806 77090
rect 83298 77016 84916 77068
rect 84968 77016 84980 77068
rect 85032 77016 85044 77068
rect 85096 77016 85108 77068
rect 85160 77016 87806 77068
rect 83298 76994 87806 77016
rect 38 76524 3902 76546
rect 38 76472 2916 76524
rect 2968 76472 2980 76524
rect 3032 76472 3044 76524
rect 3096 76472 3108 76524
rect 3160 76472 3902 76524
rect 38 76450 3902 76472
rect 83298 76524 87806 76546
rect 83298 76472 86916 76524
rect 86968 76472 86980 76524
rect 87032 76472 87044 76524
rect 87096 76472 87108 76524
rect 87160 76472 87806 76524
rect 83298 76450 87806 76472
rect 38 75980 3902 76002
rect 38 75928 916 75980
rect 968 75928 980 75980
rect 1032 75928 1044 75980
rect 1096 75928 1108 75980
rect 1160 75928 3902 75980
rect 38 75906 3902 75928
rect 83298 75980 87806 76002
rect 83298 75928 84916 75980
rect 84968 75928 84980 75980
rect 85032 75928 85044 75980
rect 85096 75928 85108 75980
rect 85160 75928 87806 75980
rect 83298 75906 87806 75928
rect 38 75436 3902 75458
rect 38 75384 2916 75436
rect 2968 75384 2980 75436
rect 3032 75384 3044 75436
rect 3096 75384 3108 75436
rect 3160 75384 3902 75436
rect 38 75362 3902 75384
rect 83298 75436 87806 75458
rect 83298 75384 86916 75436
rect 86968 75384 86980 75436
rect 87032 75384 87044 75436
rect 87096 75384 87108 75436
rect 87160 75384 87806 75436
rect 83298 75362 87806 75384
rect 84048 74942 84054 74994
rect 84106 74982 84112 74994
rect 84784 74982 84790 74994
rect 84106 74954 84790 74982
rect 84106 74942 84112 74954
rect 84784 74942 84790 74954
rect 84842 74942 84848 74994
rect 38 74892 3902 74914
rect 38 74840 916 74892
rect 968 74840 980 74892
rect 1032 74840 1044 74892
rect 1096 74840 1108 74892
rect 1160 74840 3902 74892
rect 38 74818 3902 74840
rect 83298 74892 87806 74914
rect 83298 74840 84916 74892
rect 84968 74840 84980 74892
rect 85032 74840 85044 74892
rect 85096 74840 85108 74892
rect 85160 74840 87806 74892
rect 83298 74818 87806 74840
rect 81840 74466 81846 74518
rect 81898 74506 81904 74518
rect 84876 74506 84882 74518
rect 81898 74478 84882 74506
rect 81898 74466 81904 74478
rect 84876 74466 84882 74478
rect 84934 74466 84940 74518
rect 82484 74398 82490 74450
rect 82542 74438 82548 74450
rect 84324 74438 84330 74450
rect 82542 74410 84330 74438
rect 82542 74398 82548 74410
rect 84324 74398 84330 74410
rect 84382 74398 84388 74450
rect 38 74348 3902 74370
rect 38 74296 2916 74348
rect 2968 74296 2980 74348
rect 3032 74296 3044 74348
rect 3096 74296 3108 74348
rect 3160 74296 3902 74348
rect 38 74274 3902 74296
rect 83298 74348 87806 74370
rect 83298 74296 86916 74348
rect 86968 74296 86980 74348
rect 87032 74296 87044 74348
rect 87096 74296 87108 74348
rect 87160 74296 87806 74348
rect 83298 74274 87806 74296
rect 38 73804 3902 73826
rect 38 73752 916 73804
rect 968 73752 980 73804
rect 1032 73752 1044 73804
rect 1096 73752 1108 73804
rect 1160 73752 3902 73804
rect 38 73730 3902 73752
rect 83298 73804 87806 73826
rect 83298 73752 84916 73804
rect 84968 73752 84980 73804
rect 85032 73752 85044 73804
rect 85096 73752 85108 73804
rect 85160 73752 87806 73804
rect 83298 73730 87806 73752
rect 38 73260 3902 73282
rect 38 73208 2916 73260
rect 2968 73208 2980 73260
rect 3032 73208 3044 73260
rect 3096 73208 3108 73260
rect 3160 73208 3902 73260
rect 38 73186 3902 73208
rect 83298 73260 87806 73282
rect 83298 73208 86916 73260
rect 86968 73208 86980 73260
rect 87032 73208 87044 73260
rect 87096 73208 87108 73260
rect 87160 73208 87806 73260
rect 83298 73186 87806 73208
rect 82116 73106 82122 73158
rect 82174 73146 82180 73158
rect 84692 73146 84698 73158
rect 82174 73118 84698 73146
rect 82174 73106 82180 73118
rect 84692 73106 84698 73118
rect 84750 73106 84756 73158
rect 82300 73038 82306 73090
rect 82358 73078 82364 73090
rect 84784 73078 84790 73090
rect 82358 73050 84790 73078
rect 82358 73038 82364 73050
rect 84784 73038 84790 73050
rect 84842 73038 84848 73090
rect 38 72716 3902 72738
rect 38 72664 916 72716
rect 968 72664 980 72716
rect 1032 72664 1044 72716
rect 1096 72664 1108 72716
rect 1160 72664 3902 72716
rect 38 72642 3902 72664
rect 83298 72716 87806 72738
rect 83298 72664 84916 72716
rect 84968 72664 84980 72716
rect 85032 72664 85044 72716
rect 85096 72664 85108 72716
rect 85160 72664 87806 72716
rect 83298 72642 87806 72664
rect 38 72172 3902 72194
rect 38 72120 2916 72172
rect 2968 72120 2980 72172
rect 3032 72120 3044 72172
rect 3096 72120 3108 72172
rect 3160 72120 3902 72172
rect 38 72098 3902 72120
rect 83298 72172 87806 72194
rect 83298 72120 86916 72172
rect 86968 72120 86980 72172
rect 87032 72120 87044 72172
rect 87096 72120 87108 72172
rect 87160 72120 87806 72172
rect 83298 72098 87806 72120
rect 38 71628 3902 71650
rect 38 71576 916 71628
rect 968 71576 980 71628
rect 1032 71576 1044 71628
rect 1096 71576 1108 71628
rect 1160 71576 3902 71628
rect 38 71554 3902 71576
rect 83298 71628 87806 71650
rect 83298 71576 84916 71628
rect 84968 71576 84980 71628
rect 85032 71576 85044 71628
rect 85096 71576 85108 71628
rect 85160 71576 87806 71628
rect 83298 71554 87806 71576
rect 38 71084 3902 71106
rect 38 71032 2916 71084
rect 2968 71032 2980 71084
rect 3032 71032 3044 71084
rect 3096 71032 3108 71084
rect 3160 71032 3902 71084
rect 38 71010 3902 71032
rect 83298 71084 87806 71106
rect 83298 71032 86916 71084
rect 86968 71032 86980 71084
rect 87032 71032 87044 71084
rect 87096 71032 87108 71084
rect 87160 71032 87806 71084
rect 83298 71010 87806 71032
rect 38 70540 3902 70562
rect 38 70488 916 70540
rect 968 70488 980 70540
rect 1032 70488 1044 70540
rect 1096 70488 1108 70540
rect 1160 70488 3902 70540
rect 38 70466 3902 70488
rect 83298 70540 87806 70562
rect 83298 70488 84916 70540
rect 84968 70488 84980 70540
rect 85032 70488 85044 70540
rect 85096 70488 85108 70540
rect 85160 70488 87806 70540
rect 83298 70466 87806 70488
rect 38 69996 3902 70018
rect 38 69944 2916 69996
rect 2968 69944 2980 69996
rect 3032 69944 3044 69996
rect 3096 69944 3108 69996
rect 3160 69944 3902 69996
rect 38 69922 3902 69944
rect 83298 69996 87806 70018
rect 83298 69944 86916 69996
rect 86968 69944 86980 69996
rect 87032 69944 87044 69996
rect 87096 69944 87108 69996
rect 87160 69944 87806 69996
rect 83298 69922 87806 69944
rect 38 69452 3902 69474
rect 38 69400 916 69452
rect 968 69400 980 69452
rect 1032 69400 1044 69452
rect 1096 69400 1108 69452
rect 1160 69400 3902 69452
rect 38 69378 3902 69400
rect 83298 69452 87806 69474
rect 83298 69400 84916 69452
rect 84968 69400 84980 69452
rect 85032 69400 85044 69452
rect 85096 69400 85108 69452
rect 85160 69400 87806 69452
rect 83298 69378 87806 69400
rect 38 68908 3902 68930
rect 38 68856 2916 68908
rect 2968 68856 2980 68908
rect 3032 68856 3044 68908
rect 3096 68856 3108 68908
rect 3160 68856 3902 68908
rect 38 68834 3902 68856
rect 83298 68908 87806 68930
rect 83298 68856 86916 68908
rect 86968 68856 86980 68908
rect 87032 68856 87044 68908
rect 87096 68856 87108 68908
rect 87160 68856 87806 68908
rect 83298 68834 87806 68856
rect 38 68364 3902 68386
rect 38 68312 916 68364
rect 968 68312 980 68364
rect 1032 68312 1044 68364
rect 1096 68312 1108 68364
rect 1160 68312 3902 68364
rect 38 68290 3902 68312
rect 83298 68364 87806 68386
rect 83298 68312 84916 68364
rect 84968 68312 84980 68364
rect 85032 68312 85044 68364
rect 85096 68312 85108 68364
rect 85160 68312 87806 68364
rect 83298 68290 87806 68312
rect 38 67820 3902 67842
rect 38 67768 2916 67820
rect 2968 67768 2980 67820
rect 3032 67768 3044 67820
rect 3096 67768 3108 67820
rect 3160 67768 3902 67820
rect 38 67746 3902 67768
rect 83298 67820 87806 67842
rect 83298 67768 86916 67820
rect 86968 67768 86980 67820
rect 87032 67768 87044 67820
rect 87096 67768 87108 67820
rect 87160 67768 87806 67820
rect 83298 67746 87806 67768
rect 38 67276 3902 67298
rect 38 67224 916 67276
rect 968 67224 980 67276
rect 1032 67224 1044 67276
rect 1096 67224 1108 67276
rect 1160 67224 3902 67276
rect 38 67202 3902 67224
rect 83298 67276 87806 67298
rect 83298 67224 84916 67276
rect 84968 67224 84980 67276
rect 85032 67224 85044 67276
rect 85096 67224 85108 67276
rect 85160 67224 87806 67276
rect 83298 67202 87806 67224
rect 38 66732 3902 66754
rect 38 66680 2916 66732
rect 2968 66680 2980 66732
rect 3032 66680 3044 66732
rect 3096 66680 3108 66732
rect 3160 66680 3902 66732
rect 38 66658 3902 66680
rect 83298 66732 87806 66754
rect 83298 66680 86916 66732
rect 86968 66680 86980 66732
rect 87032 66680 87044 66732
rect 87096 66680 87108 66732
rect 87160 66680 87806 66732
rect 83298 66658 87806 66680
rect 82024 66578 82030 66630
rect 82082 66618 82088 66630
rect 85152 66618 85158 66630
rect 82082 66590 85158 66618
rect 82082 66578 82088 66590
rect 85152 66578 85158 66590
rect 85210 66578 85216 66630
rect 38 66188 3902 66210
rect 38 66136 916 66188
rect 968 66136 980 66188
rect 1032 66136 1044 66188
rect 1096 66136 1108 66188
rect 1160 66136 3902 66188
rect 38 66114 3902 66136
rect 83298 66188 87806 66210
rect 83298 66136 84916 66188
rect 84968 66136 84980 66188
rect 85032 66136 85044 66188
rect 85096 66136 85108 66188
rect 85160 66136 87806 66188
rect 83298 66114 87806 66136
rect 38 65644 3902 65666
rect 38 65592 2916 65644
rect 2968 65592 2980 65644
rect 3032 65592 3044 65644
rect 3096 65592 3108 65644
rect 3160 65592 3902 65644
rect 38 65570 3902 65592
rect 83298 65644 87806 65666
rect 83298 65592 86916 65644
rect 86968 65592 86980 65644
rect 87032 65592 87044 65644
rect 87096 65592 87108 65644
rect 87160 65592 87806 65644
rect 83298 65570 87806 65592
rect 38 65100 3902 65122
rect 38 65048 916 65100
rect 968 65048 980 65100
rect 1032 65048 1044 65100
rect 1096 65048 1108 65100
rect 1160 65048 3902 65100
rect 38 65026 3902 65048
rect 83298 65100 87806 65122
rect 83298 65048 84916 65100
rect 84968 65048 84980 65100
rect 85032 65048 85044 65100
rect 85096 65048 85108 65100
rect 85160 65048 87806 65100
rect 83298 65026 87806 65048
rect 38 64556 3902 64578
rect 38 64504 2916 64556
rect 2968 64504 2980 64556
rect 3032 64504 3044 64556
rect 3096 64504 3108 64556
rect 3160 64504 3902 64556
rect 38 64482 3902 64504
rect 83298 64556 87806 64578
rect 83298 64504 86916 64556
rect 86968 64504 86980 64556
rect 87032 64504 87044 64556
rect 87096 64504 87108 64556
rect 87160 64504 87806 64556
rect 83298 64482 87806 64504
rect 38 64012 3902 64034
rect 38 63960 916 64012
rect 968 63960 980 64012
rect 1032 63960 1044 64012
rect 1096 63960 1108 64012
rect 1160 63960 3902 64012
rect 38 63938 3902 63960
rect 83298 64012 87806 64034
rect 83298 63960 84916 64012
rect 84968 63960 84980 64012
rect 85032 63960 85044 64012
rect 85096 63960 85108 64012
rect 85160 63960 87806 64012
rect 83298 63938 87806 63960
rect 38 63468 3902 63490
rect 38 63416 2916 63468
rect 2968 63416 2980 63468
rect 3032 63416 3044 63468
rect 3096 63416 3108 63468
rect 3160 63416 3902 63468
rect 38 63394 3902 63416
rect 83298 63468 87806 63490
rect 83298 63416 86916 63468
rect 86968 63416 86980 63468
rect 87032 63416 87044 63468
rect 87096 63416 87108 63468
rect 87160 63416 87806 63468
rect 83298 63394 87806 63416
rect 3640 63314 3646 63366
rect 3698 63314 3704 63366
rect 3658 63026 3686 63314
rect 3640 62974 3646 63026
rect 3698 62974 3704 63026
rect 3824 62974 3830 63026
rect 3882 63014 3888 63026
rect 3916 63014 3922 63026
rect 3882 62986 3922 63014
rect 3882 62974 3888 62986
rect 3916 62974 3922 62986
rect 3974 62974 3980 63026
rect 38 62924 3902 62946
rect 38 62872 916 62924
rect 968 62872 980 62924
rect 1032 62872 1044 62924
rect 1096 62872 1108 62924
rect 1160 62872 3902 62924
rect 38 62850 3902 62872
rect 83298 62924 87806 62946
rect 83298 62872 84916 62924
rect 84968 62872 84980 62924
rect 85032 62872 85044 62924
rect 85096 62872 85108 62924
rect 85160 62872 87806 62924
rect 83298 62850 87806 62872
rect 81932 62770 81938 62822
rect 81990 62810 81996 62822
rect 84784 62810 84790 62822
rect 81990 62782 84790 62810
rect 81990 62770 81996 62782
rect 84784 62770 84790 62782
rect 84842 62770 84848 62822
rect 38 62380 3902 62402
rect 38 62328 2916 62380
rect 2968 62328 2980 62380
rect 3032 62328 3044 62380
rect 3096 62328 3108 62380
rect 3160 62328 3902 62380
rect 38 62306 3902 62328
rect 83298 62380 87806 62402
rect 83298 62328 86916 62380
rect 86968 62328 86980 62380
rect 87032 62328 87044 62380
rect 87096 62328 87108 62380
rect 87160 62328 87806 62380
rect 83298 62306 87806 62328
rect 38 61836 3902 61858
rect 38 61784 916 61836
rect 968 61784 980 61836
rect 1032 61784 1044 61836
rect 1096 61784 1108 61836
rect 1160 61784 3902 61836
rect 38 61762 3902 61784
rect 83298 61836 87806 61858
rect 83298 61784 84916 61836
rect 84968 61784 84980 61836
rect 85032 61784 85044 61836
rect 85096 61784 85108 61836
rect 85160 61784 87806 61836
rect 83298 61762 87806 61784
rect 3824 61546 3830 61598
rect 3882 61586 3888 61598
rect 4011 61589 4069 61595
rect 4011 61586 4023 61589
rect 3882 61558 4023 61586
rect 3882 61546 3888 61558
rect 4011 61555 4023 61558
rect 4057 61555 4069 61589
rect 4011 61549 4069 61555
rect 38 61292 3902 61314
rect 38 61240 2916 61292
rect 2968 61240 2980 61292
rect 3032 61240 3044 61292
rect 3096 61240 3108 61292
rect 3160 61240 3902 61292
rect 38 61218 3902 61240
rect 83298 61292 87806 61314
rect 83298 61240 86916 61292
rect 86968 61240 86980 61292
rect 87032 61240 87044 61292
rect 87096 61240 87108 61292
rect 87160 61240 87806 61292
rect 83298 61218 87806 61240
rect 38 60748 3902 60770
rect 38 60696 916 60748
rect 968 60696 980 60748
rect 1032 60696 1044 60748
rect 1096 60696 1108 60748
rect 1160 60696 3902 60748
rect 38 60674 3902 60696
rect 83298 60748 87806 60770
rect 83298 60696 84916 60748
rect 84968 60696 84980 60748
rect 85032 60696 85044 60748
rect 85096 60696 85108 60748
rect 85160 60696 87806 60748
rect 83298 60674 87806 60696
rect 38 60204 3902 60226
rect 38 60152 2916 60204
rect 2968 60152 2980 60204
rect 3032 60152 3044 60204
rect 3096 60152 3108 60204
rect 3160 60152 3902 60204
rect 38 60130 3902 60152
rect 83298 60204 87806 60226
rect 83298 60152 86916 60204
rect 86968 60152 86980 60204
rect 87032 60152 87044 60204
rect 87096 60152 87108 60204
rect 87160 60152 87806 60204
rect 83298 60130 87806 60152
rect 38 59660 3902 59682
rect 38 59608 916 59660
rect 968 59608 980 59660
rect 1032 59608 1044 59660
rect 1096 59608 1108 59660
rect 1160 59608 3902 59660
rect 38 59586 3902 59608
rect 83298 59660 87806 59682
rect 83298 59608 84916 59660
rect 84968 59608 84980 59660
rect 85032 59608 85044 59660
rect 85096 59608 85108 59660
rect 85160 59608 87806 59660
rect 83298 59586 87806 59608
rect 38 59116 3902 59138
rect 38 59064 2916 59116
rect 2968 59064 2980 59116
rect 3032 59064 3044 59116
rect 3096 59064 3108 59116
rect 3160 59064 3902 59116
rect 38 59042 3902 59064
rect 83298 59116 87806 59138
rect 83298 59064 86916 59116
rect 86968 59064 86980 59116
rect 87032 59064 87044 59116
rect 87096 59064 87108 59116
rect 87160 59064 87806 59116
rect 83298 59042 87806 59064
rect 38 58572 3902 58594
rect 38 58520 916 58572
rect 968 58520 980 58572
rect 1032 58520 1044 58572
rect 1096 58520 1108 58572
rect 1160 58520 3902 58572
rect 38 58498 3902 58520
rect 83298 58572 87806 58594
rect 83298 58520 84916 58572
rect 84968 58520 84980 58572
rect 85032 58520 85044 58572
rect 85096 58520 85108 58572
rect 85160 58520 87806 58572
rect 83298 58498 87806 58520
rect 38 58028 3902 58050
rect 38 57976 2916 58028
rect 2968 57976 2980 58028
rect 3032 57976 3044 58028
rect 3096 57976 3108 58028
rect 3160 57976 3902 58028
rect 38 57954 3902 57976
rect 83298 58028 87806 58050
rect 83298 57976 86916 58028
rect 86968 57976 86980 58028
rect 87032 57976 87044 58028
rect 87096 57976 87108 58028
rect 87160 57976 87806 58028
rect 83298 57954 87806 57976
rect 38 57484 3902 57506
rect 38 57432 916 57484
rect 968 57432 980 57484
rect 1032 57432 1044 57484
rect 1096 57432 1108 57484
rect 1160 57432 3902 57484
rect 38 57410 3902 57432
rect 83298 57484 87806 57506
rect 83298 57432 84916 57484
rect 84968 57432 84980 57484
rect 85032 57432 85044 57484
rect 85096 57432 85108 57484
rect 85160 57432 87806 57484
rect 83298 57410 87806 57432
rect 38 56940 3902 56962
rect 38 56888 2916 56940
rect 2968 56888 2980 56940
rect 3032 56888 3044 56940
rect 3096 56888 3108 56940
rect 3160 56888 3902 56940
rect 38 56866 3902 56888
rect 83298 56940 87806 56962
rect 83298 56888 86916 56940
rect 86968 56888 86980 56940
rect 87032 56888 87044 56940
rect 87096 56888 87108 56940
rect 87160 56888 87806 56940
rect 83298 56866 87806 56888
rect 83128 56554 83134 56566
rect 83089 56526 83134 56554
rect 83128 56514 83134 56526
rect 83186 56514 83192 56566
rect 81932 56446 81938 56498
rect 81990 56486 81996 56498
rect 84784 56486 84790 56498
rect 81990 56458 84790 56486
rect 81990 56446 81996 56458
rect 84784 56446 84790 56458
rect 84842 56446 84848 56498
rect 83128 56418 83134 56430
rect 38 56396 3902 56418
rect 38 56344 916 56396
rect 968 56344 980 56396
rect 1032 56344 1044 56396
rect 1096 56344 1108 56396
rect 1160 56344 3902 56396
rect 83089 56390 83134 56418
rect 83128 56378 83134 56390
rect 83186 56378 83192 56430
rect 83298 56396 87806 56418
rect 38 56322 3902 56344
rect 83298 56344 84916 56396
rect 84968 56344 84980 56396
rect 85032 56344 85044 56396
rect 85096 56344 85108 56396
rect 85160 56344 87806 56396
rect 83298 56322 87806 56344
rect 3824 56242 3830 56294
rect 3882 56282 3888 56294
rect 4011 56285 4069 56291
rect 4011 56282 4023 56285
rect 3882 56254 4023 56282
rect 3882 56242 3888 56254
rect 4011 56251 4023 56254
rect 4057 56251 4069 56285
rect 4011 56245 4069 56251
rect 38 55852 3902 55874
rect 38 55800 2916 55852
rect 2968 55800 2980 55852
rect 3032 55800 3044 55852
rect 3096 55800 3108 55852
rect 3160 55800 3902 55852
rect 38 55778 3902 55800
rect 83298 55852 87806 55874
rect 83298 55800 86916 55852
rect 86968 55800 86980 55852
rect 87032 55800 87044 55852
rect 87096 55800 87108 55852
rect 87160 55800 87806 55852
rect 83298 55778 87806 55800
rect 38 55308 3902 55330
rect 38 55256 916 55308
rect 968 55256 980 55308
rect 1032 55256 1044 55308
rect 1096 55256 1108 55308
rect 1160 55256 3902 55308
rect 38 55234 3902 55256
rect 83298 55308 87806 55330
rect 83298 55256 84916 55308
rect 84968 55256 84980 55308
rect 85032 55256 85044 55308
rect 85096 55256 85108 55308
rect 85160 55256 87806 55308
rect 83298 55234 87806 55256
rect 38 54764 3902 54786
rect 38 54712 2916 54764
rect 2968 54712 2980 54764
rect 3032 54712 3044 54764
rect 3096 54712 3108 54764
rect 3160 54712 3902 54764
rect 38 54690 3902 54712
rect 83298 54764 87806 54786
rect 83298 54712 86916 54764
rect 86968 54712 86980 54764
rect 87032 54712 87044 54764
rect 87096 54712 87108 54764
rect 87160 54712 87806 54764
rect 83298 54690 87806 54712
rect 38 54220 3902 54242
rect 38 54168 916 54220
rect 968 54168 980 54220
rect 1032 54168 1044 54220
rect 1096 54168 1108 54220
rect 1160 54168 3902 54220
rect 38 54146 3902 54168
rect 83298 54220 87806 54242
rect 83298 54168 84916 54220
rect 84968 54168 84980 54220
rect 85032 54168 85044 54220
rect 85096 54168 85108 54220
rect 85160 54168 87806 54220
rect 83298 54146 87806 54168
rect 38 53676 3902 53698
rect 38 53624 2916 53676
rect 2968 53624 2980 53676
rect 3032 53624 3044 53676
rect 3096 53624 3108 53676
rect 3160 53624 3902 53676
rect 38 53602 3902 53624
rect 83298 53676 87806 53698
rect 83298 53624 86916 53676
rect 86968 53624 86980 53676
rect 87032 53624 87044 53676
rect 87096 53624 87108 53676
rect 87160 53624 87806 53676
rect 83298 53602 87806 53624
rect 38 53132 3902 53154
rect 38 53080 916 53132
rect 968 53080 980 53132
rect 1032 53080 1044 53132
rect 1096 53080 1108 53132
rect 1160 53080 3902 53132
rect 38 53058 3902 53080
rect 83298 53132 87806 53154
rect 83298 53080 84916 53132
rect 84968 53080 84980 53132
rect 85032 53080 85044 53132
rect 85096 53080 85108 53132
rect 85160 53080 87806 53132
rect 83298 53058 87806 53080
rect 38 52588 3902 52610
rect 38 52536 2916 52588
rect 2968 52536 2980 52588
rect 3032 52536 3044 52588
rect 3096 52536 3108 52588
rect 3160 52536 3902 52588
rect 82852 52570 82858 52622
rect 82910 52610 82916 52622
rect 83128 52610 83134 52622
rect 82910 52582 83134 52610
rect 82910 52570 82916 52582
rect 83128 52570 83134 52582
rect 83186 52570 83192 52622
rect 83298 52588 87806 52610
rect 38 52514 3902 52536
rect 83298 52536 86916 52588
rect 86968 52536 86980 52588
rect 87032 52536 87044 52588
rect 87096 52536 87108 52588
rect 87160 52536 87806 52588
rect 83298 52514 87806 52536
rect 38 52044 3902 52066
rect 38 51992 916 52044
rect 968 51992 980 52044
rect 1032 51992 1044 52044
rect 1096 51992 1108 52044
rect 1160 51992 3902 52044
rect 38 51970 3902 51992
rect 83298 52044 87806 52066
rect 83298 51992 84916 52044
rect 84968 51992 84980 52044
rect 85032 51992 85044 52044
rect 85096 51992 85108 52044
rect 85160 51992 87806 52044
rect 83298 51970 87806 51992
rect 38 51500 3902 51522
rect 38 51448 2916 51500
rect 2968 51448 2980 51500
rect 3032 51448 3044 51500
rect 3096 51448 3108 51500
rect 3160 51448 3902 51500
rect 38 51426 3902 51448
rect 83298 51500 87806 51522
rect 83298 51448 86916 51500
rect 86968 51448 86980 51500
rect 87032 51448 87044 51500
rect 87096 51448 87108 51500
rect 87160 51448 87806 51500
rect 83298 51426 87806 51448
rect 38 50956 3902 50978
rect 38 50904 916 50956
rect 968 50904 980 50956
rect 1032 50904 1044 50956
rect 1096 50904 1108 50956
rect 1160 50904 3902 50956
rect 38 50882 3902 50904
rect 83298 50956 87806 50978
rect 83298 50904 84916 50956
rect 84968 50904 84980 50956
rect 85032 50904 85044 50956
rect 85096 50904 85108 50956
rect 85160 50904 87806 50956
rect 83298 50882 87806 50904
rect 38 50412 3902 50434
rect 38 50360 2916 50412
rect 2968 50360 2980 50412
rect 3032 50360 3044 50412
rect 3096 50360 3108 50412
rect 3160 50360 3902 50412
rect 38 50338 3902 50360
rect 83298 50412 87806 50434
rect 83298 50360 86916 50412
rect 86968 50360 86980 50412
rect 87032 50360 87044 50412
rect 87096 50360 87108 50412
rect 87160 50360 87806 50412
rect 83298 50338 87806 50360
rect 82024 50054 82030 50106
rect 82082 50094 82088 50106
rect 85152 50094 85158 50106
rect 82082 50066 85158 50094
rect 82082 50054 82088 50066
rect 85152 50054 85158 50066
rect 85210 50054 85216 50106
rect 38 49868 3902 49890
rect 38 49816 916 49868
rect 968 49816 980 49868
rect 1032 49816 1044 49868
rect 1096 49816 1108 49868
rect 1160 49816 3902 49868
rect 38 49794 3902 49816
rect 83298 49868 87806 49890
rect 83298 49816 84916 49868
rect 84968 49816 84980 49868
rect 85032 49816 85044 49868
rect 85096 49816 85108 49868
rect 85160 49816 87806 49868
rect 83298 49794 87806 49816
rect 38 49324 3902 49346
rect 38 49272 2916 49324
rect 2968 49272 2980 49324
rect 3032 49272 3044 49324
rect 3096 49272 3108 49324
rect 3160 49272 3902 49324
rect 38 49250 3902 49272
rect 83298 49324 87806 49346
rect 83298 49272 86916 49324
rect 86968 49272 86980 49324
rect 87032 49272 87044 49324
rect 87096 49272 87108 49324
rect 87160 49272 87806 49324
rect 83298 49250 87806 49272
rect 82116 48830 82122 48882
rect 82174 48870 82180 48882
rect 84784 48870 84790 48882
rect 82174 48842 84790 48870
rect 82174 48830 82180 48842
rect 84784 48830 84790 48842
rect 84842 48830 84848 48882
rect 38 48780 3902 48802
rect 38 48728 916 48780
rect 968 48728 980 48780
rect 1032 48728 1044 48780
rect 1096 48728 1108 48780
rect 1160 48728 3902 48780
rect 38 48706 3902 48728
rect 83298 48780 87806 48802
rect 83298 48728 84916 48780
rect 84968 48728 84980 48780
rect 85032 48728 85044 48780
rect 85096 48728 85108 48780
rect 85160 48728 87806 48780
rect 83298 48706 87806 48728
rect 38 48236 3902 48258
rect 38 48184 2916 48236
rect 2968 48184 2980 48236
rect 3032 48184 3044 48236
rect 3096 48184 3108 48236
rect 3160 48184 3902 48236
rect 38 48162 3902 48184
rect 83298 48236 87806 48258
rect 83298 48184 86916 48236
rect 86968 48184 86980 48236
rect 87032 48184 87044 48236
rect 87096 48184 87108 48236
rect 87160 48184 87806 48236
rect 83298 48162 87806 48184
rect 38 47692 3902 47714
rect 38 47640 916 47692
rect 968 47640 980 47692
rect 1032 47640 1044 47692
rect 1096 47640 1108 47692
rect 1160 47640 3902 47692
rect 38 47618 3902 47640
rect 83298 47692 87806 47714
rect 83298 47640 84916 47692
rect 84968 47640 84980 47692
rect 85032 47640 85044 47692
rect 85096 47640 85108 47692
rect 85160 47640 87806 47692
rect 83298 47618 87806 47640
rect 38 47148 3902 47170
rect 38 47096 2916 47148
rect 2968 47096 2980 47148
rect 3032 47096 3044 47148
rect 3096 47096 3108 47148
rect 3160 47096 3902 47148
rect 38 47074 3902 47096
rect 83298 47148 87806 47170
rect 83298 47096 86916 47148
rect 86968 47096 86980 47148
rect 87032 47096 87044 47148
rect 87096 47096 87108 47148
rect 87160 47096 87806 47148
rect 83298 47074 87806 47096
rect 38 46604 3902 46626
rect 38 46552 916 46604
rect 968 46552 980 46604
rect 1032 46552 1044 46604
rect 1096 46552 1108 46604
rect 1160 46552 3902 46604
rect 38 46530 3902 46552
rect 83298 46604 87806 46626
rect 83298 46552 84916 46604
rect 84968 46552 84980 46604
rect 85032 46552 85044 46604
rect 85096 46552 85108 46604
rect 85160 46552 87806 46604
rect 83298 46530 87806 46552
rect 38 46060 3902 46082
rect 38 46008 2916 46060
rect 2968 46008 2980 46060
rect 3032 46008 3044 46060
rect 3096 46008 3108 46060
rect 3160 46008 3902 46060
rect 38 45986 3902 46008
rect 83298 46060 87806 46082
rect 83298 46008 86916 46060
rect 86968 46008 86980 46060
rect 87032 46008 87044 46060
rect 87096 46008 87108 46060
rect 87160 46008 87806 46060
rect 83298 45986 87806 46008
rect 38 45516 3902 45538
rect 38 45464 916 45516
rect 968 45464 980 45516
rect 1032 45464 1044 45516
rect 1096 45464 1108 45516
rect 1160 45464 3902 45516
rect 38 45442 3902 45464
rect 83298 45516 87806 45538
rect 83298 45464 84916 45516
rect 84968 45464 84980 45516
rect 85032 45464 85044 45516
rect 85096 45464 85108 45516
rect 85160 45464 87806 45516
rect 83298 45442 87806 45464
rect 38 44972 3902 44994
rect 38 44920 2916 44972
rect 2968 44920 2980 44972
rect 3032 44920 3044 44972
rect 3096 44920 3108 44972
rect 3160 44920 3902 44972
rect 38 44898 3902 44920
rect 83298 44972 87806 44994
rect 83298 44920 86916 44972
rect 86968 44920 86980 44972
rect 87032 44920 87044 44972
rect 87096 44920 87108 44972
rect 87160 44920 87806 44972
rect 83298 44898 87806 44920
rect 3364 44818 3370 44870
rect 3422 44858 3428 44870
rect 3551 44861 3609 44867
rect 3551 44858 3563 44861
rect 3422 44830 3563 44858
rect 3422 44818 3428 44830
rect 3551 44827 3563 44830
rect 3597 44827 3609 44861
rect 3551 44821 3609 44827
rect 3640 44818 3646 44870
rect 3698 44818 3704 44870
rect 3732 44818 3738 44870
rect 3790 44818 3796 44870
rect 3658 44598 3686 44818
rect 3750 44598 3778 44818
rect 3824 44750 3830 44802
rect 3882 44790 3888 44802
rect 4011 44793 4069 44799
rect 4011 44790 4023 44793
rect 3882 44762 4023 44790
rect 3882 44750 3888 44762
rect 4011 44759 4023 44762
rect 4057 44759 4069 44793
rect 4011 44753 4069 44759
rect 3640 44546 3646 44598
rect 3698 44546 3704 44598
rect 3732 44546 3738 44598
rect 3790 44546 3796 44598
rect 3551 44521 3609 44527
rect 3551 44487 3563 44521
rect 3597 44518 3609 44521
rect 3824 44518 3830 44530
rect 3597 44490 3830 44518
rect 3597 44487 3609 44490
rect 3551 44481 3609 44487
rect 3824 44478 3830 44490
rect 3882 44478 3888 44530
rect 38 44428 3902 44450
rect 38 44376 916 44428
rect 968 44376 980 44428
rect 1032 44376 1044 44428
rect 1096 44376 1108 44428
rect 1160 44376 3902 44428
rect 38 44354 3902 44376
rect 83298 44428 87806 44450
rect 83298 44376 84916 44428
rect 84968 44376 84980 44428
rect 85032 44376 85044 44428
rect 85096 44376 85108 44428
rect 85160 44376 87806 44428
rect 83298 44354 87806 44376
rect 38 43884 3902 43906
rect 38 43832 2916 43884
rect 2968 43832 2980 43884
rect 3032 43832 3044 43884
rect 3096 43832 3108 43884
rect 3160 43832 3902 43884
rect 38 43810 3902 43832
rect 83298 43884 87806 43906
rect 83298 43832 86916 43884
rect 86968 43832 86980 43884
rect 87032 43832 87044 43884
rect 87096 43832 87108 43884
rect 87160 43832 87806 43884
rect 83298 43810 87806 43832
rect 82208 43594 82214 43646
rect 82266 43634 82272 43646
rect 85152 43634 85158 43646
rect 82266 43606 85158 43634
rect 82266 43594 82272 43606
rect 85152 43594 85158 43606
rect 85210 43594 85216 43646
rect 38 43340 3902 43362
rect 38 43288 916 43340
rect 968 43288 980 43340
rect 1032 43288 1044 43340
rect 1096 43288 1108 43340
rect 1160 43288 3902 43340
rect 38 43266 3902 43288
rect 83298 43340 87806 43362
rect 83298 43288 84916 43340
rect 84968 43288 84980 43340
rect 85032 43288 85044 43340
rect 85096 43288 85108 43340
rect 85160 43288 87806 43340
rect 83298 43266 87806 43288
rect 38 42796 3902 42818
rect 38 42744 2916 42796
rect 2968 42744 2980 42796
rect 3032 42744 3044 42796
rect 3096 42744 3108 42796
rect 3160 42744 3902 42796
rect 38 42722 3902 42744
rect 83298 42796 87806 42818
rect 83298 42744 86916 42796
rect 86968 42744 86980 42796
rect 87032 42744 87044 42796
rect 87096 42744 87108 42796
rect 87160 42744 87806 42796
rect 83298 42722 87806 42744
rect 38 42252 3902 42274
rect 38 42200 916 42252
rect 968 42200 980 42252
rect 1032 42200 1044 42252
rect 1096 42200 1108 42252
rect 1160 42200 3902 42252
rect 38 42178 3902 42200
rect 83298 42252 87806 42274
rect 83298 42200 84916 42252
rect 84968 42200 84980 42252
rect 85032 42200 85044 42252
rect 85096 42200 85108 42252
rect 85160 42200 87806 42252
rect 83298 42178 87806 42200
rect 38 41708 3902 41730
rect 38 41656 2916 41708
rect 2968 41656 2980 41708
rect 3032 41656 3044 41708
rect 3096 41656 3108 41708
rect 3160 41656 3902 41708
rect 38 41634 3902 41656
rect 83298 41708 87806 41730
rect 83298 41656 86916 41708
rect 86968 41656 86980 41708
rect 87032 41656 87044 41708
rect 87096 41656 87108 41708
rect 87160 41656 87806 41708
rect 83298 41634 87806 41656
rect 38 41164 3902 41186
rect 38 41112 916 41164
rect 968 41112 980 41164
rect 1032 41112 1044 41164
rect 1096 41112 1108 41164
rect 1160 41112 3902 41164
rect 38 41090 3902 41112
rect 83298 41164 87806 41186
rect 83298 41112 84916 41164
rect 84968 41112 84980 41164
rect 85032 41112 85044 41164
rect 85096 41112 85108 41164
rect 85160 41112 87806 41164
rect 83298 41090 87806 41112
rect 38 40620 3902 40642
rect 38 40568 2916 40620
rect 2968 40568 2980 40620
rect 3032 40568 3044 40620
rect 3096 40568 3108 40620
rect 3160 40568 3902 40620
rect 38 40546 3902 40568
rect 83298 40620 87806 40642
rect 83298 40568 86916 40620
rect 86968 40568 86980 40620
rect 87032 40568 87044 40620
rect 87096 40568 87108 40620
rect 87160 40568 87806 40620
rect 83298 40546 87806 40568
rect 38 40076 3902 40098
rect 38 40024 916 40076
rect 968 40024 980 40076
rect 1032 40024 1044 40076
rect 1096 40024 1108 40076
rect 1160 40024 3902 40076
rect 38 40002 3902 40024
rect 83298 40076 87806 40098
rect 83298 40024 84916 40076
rect 84968 40024 84980 40076
rect 85032 40024 85044 40076
rect 85096 40024 85108 40076
rect 85160 40024 87806 40076
rect 83298 40002 87806 40024
rect 82300 39922 82306 39974
rect 82358 39962 82364 39974
rect 84784 39962 84790 39974
rect 82358 39934 84790 39962
rect 82358 39922 82364 39934
rect 84784 39922 84790 39934
rect 84842 39922 84848 39974
rect 38 39532 3902 39554
rect 38 39480 2916 39532
rect 2968 39480 2980 39532
rect 3032 39480 3044 39532
rect 3096 39480 3108 39532
rect 3160 39480 3902 39532
rect 38 39458 3902 39480
rect 83298 39532 87806 39554
rect 83298 39480 86916 39532
rect 86968 39480 86980 39532
rect 87032 39480 87044 39532
rect 87096 39480 87108 39532
rect 87160 39480 87806 39532
rect 83298 39458 87806 39480
rect 38 38988 3902 39010
rect 38 38936 916 38988
rect 968 38936 980 38988
rect 1032 38936 1044 38988
rect 1096 38936 1108 38988
rect 1160 38936 3902 38988
rect 38 38914 3902 38936
rect 83298 38988 87806 39010
rect 83298 38936 84916 38988
rect 84968 38936 84980 38988
rect 85032 38936 85044 38988
rect 85096 38936 85108 38988
rect 85160 38936 87806 38988
rect 83298 38914 87806 38936
rect 38 38444 3902 38466
rect 38 38392 2916 38444
rect 2968 38392 2980 38444
rect 3032 38392 3044 38444
rect 3096 38392 3108 38444
rect 3160 38392 3902 38444
rect 38 38370 3902 38392
rect 83298 38444 87806 38466
rect 83298 38392 86916 38444
rect 86968 38392 86980 38444
rect 87032 38392 87044 38444
rect 87096 38392 87108 38444
rect 87160 38392 87806 38444
rect 83298 38370 87806 38392
rect 3916 38290 3922 38342
rect 3974 38330 3980 38342
rect 4011 38333 4069 38339
rect 4011 38330 4023 38333
rect 3974 38302 4023 38330
rect 3974 38290 3980 38302
rect 4011 38299 4023 38302
rect 4057 38299 4069 38333
rect 4011 38293 4069 38299
rect 38 37900 3902 37922
rect 38 37848 916 37900
rect 968 37848 980 37900
rect 1032 37848 1044 37900
rect 1096 37848 1108 37900
rect 1160 37848 3902 37900
rect 38 37826 3902 37848
rect 83298 37900 87806 37922
rect 83298 37848 84916 37900
rect 84968 37848 84980 37900
rect 85032 37848 85044 37900
rect 85096 37848 85108 37900
rect 85160 37848 87806 37900
rect 83298 37826 87806 37848
rect 38 37356 3902 37378
rect 38 37304 2916 37356
rect 2968 37304 2980 37356
rect 3032 37304 3044 37356
rect 3096 37304 3108 37356
rect 3160 37304 3902 37356
rect 38 37282 3902 37304
rect 83298 37356 87806 37378
rect 83298 37304 86916 37356
rect 86968 37304 86980 37356
rect 87032 37304 87044 37356
rect 87096 37304 87108 37356
rect 87160 37304 87806 37356
rect 83298 37282 87806 37304
rect 38 36812 3902 36834
rect 38 36760 916 36812
rect 968 36760 980 36812
rect 1032 36760 1044 36812
rect 1096 36760 1108 36812
rect 1160 36760 3902 36812
rect 38 36738 3902 36760
rect 83298 36812 87806 36834
rect 83298 36760 84916 36812
rect 84968 36760 84980 36812
rect 85032 36760 85044 36812
rect 85096 36760 85108 36812
rect 85160 36760 87806 36812
rect 83298 36738 87806 36760
rect 38 36268 3902 36290
rect 38 36216 2916 36268
rect 2968 36216 2980 36268
rect 3032 36216 3044 36268
rect 3096 36216 3108 36268
rect 3160 36216 3902 36268
rect 38 36194 3902 36216
rect 83298 36268 87806 36290
rect 83298 36216 86916 36268
rect 86968 36216 86980 36268
rect 87032 36216 87044 36268
rect 87096 36216 87108 36268
rect 87160 36216 87806 36268
rect 83298 36194 87806 36216
rect 3272 35842 3278 35894
rect 3330 35882 3336 35894
rect 3824 35882 3830 35894
rect 3330 35854 3830 35882
rect 3330 35842 3336 35854
rect 3824 35842 3830 35854
rect 3882 35842 3888 35894
rect 38 35724 3902 35746
rect 38 35672 916 35724
rect 968 35672 980 35724
rect 1032 35672 1044 35724
rect 1096 35672 1108 35724
rect 1160 35672 3902 35724
rect 38 35650 3902 35672
rect 83298 35724 87806 35746
rect 83298 35672 84916 35724
rect 84968 35672 84980 35724
rect 85032 35672 85044 35724
rect 85096 35672 85108 35724
rect 85160 35672 87806 35724
rect 83298 35650 87806 35672
rect 82392 35434 82398 35486
rect 82450 35474 82456 35486
rect 84140 35474 84146 35486
rect 82450 35446 84146 35474
rect 82450 35434 82456 35446
rect 84140 35434 84146 35446
rect 84198 35434 84204 35486
rect 38 35180 3902 35202
rect 38 35128 2916 35180
rect 2968 35128 2980 35180
rect 3032 35128 3044 35180
rect 3096 35128 3108 35180
rect 3160 35128 3902 35180
rect 38 35106 3902 35128
rect 83298 35180 87806 35202
rect 83298 35128 86916 35180
rect 86968 35128 86980 35180
rect 87032 35128 87044 35180
rect 87096 35128 87108 35180
rect 87160 35128 87806 35180
rect 83298 35106 87806 35128
rect 38 34636 3902 34658
rect 38 34584 916 34636
rect 968 34584 980 34636
rect 1032 34584 1044 34636
rect 1096 34584 1108 34636
rect 1160 34584 3902 34636
rect 38 34562 3902 34584
rect 83298 34636 87806 34658
rect 83298 34584 84916 34636
rect 84968 34584 84980 34636
rect 85032 34584 85044 34636
rect 85096 34584 85108 34636
rect 85160 34584 87806 34636
rect 83298 34562 87806 34584
rect 38 34092 3902 34114
rect 38 34040 2916 34092
rect 2968 34040 2980 34092
rect 3032 34040 3044 34092
rect 3096 34040 3108 34092
rect 3160 34040 3902 34092
rect 38 34018 3902 34040
rect 83298 34092 87806 34114
rect 83298 34040 86916 34092
rect 86968 34040 86980 34092
rect 87032 34040 87044 34092
rect 87096 34040 87108 34092
rect 87160 34040 87806 34092
rect 83298 34018 87806 34040
rect 38 33548 3902 33570
rect 38 33496 916 33548
rect 968 33496 980 33548
rect 1032 33496 1044 33548
rect 1096 33496 1108 33548
rect 1160 33496 3902 33548
rect 38 33474 3902 33496
rect 83298 33548 87806 33570
rect 83298 33496 84916 33548
rect 84968 33496 84980 33548
rect 85032 33496 85044 33548
rect 85096 33496 85108 33548
rect 85160 33496 87806 33548
rect 83298 33474 87806 33496
rect 38 33004 3902 33026
rect 38 32952 2916 33004
rect 2968 32952 2980 33004
rect 3032 32952 3044 33004
rect 3096 32952 3108 33004
rect 3160 32952 3902 33004
rect 38 32930 3902 32952
rect 83298 33004 87806 33026
rect 83298 32952 86916 33004
rect 86968 32952 86980 33004
rect 87032 32952 87044 33004
rect 87096 32952 87108 33004
rect 87160 32952 87806 33004
rect 83298 32930 87806 32952
rect 38 32460 3902 32482
rect 38 32408 916 32460
rect 968 32408 980 32460
rect 1032 32408 1044 32460
rect 1096 32408 1108 32460
rect 1160 32408 3902 32460
rect 38 32386 3902 32408
rect 83298 32460 87806 32482
rect 83298 32408 84916 32460
rect 84968 32408 84980 32460
rect 85032 32408 85044 32460
rect 85096 32408 85108 32460
rect 85160 32408 87806 32460
rect 83298 32386 87806 32408
rect 82484 32034 82490 32086
rect 82542 32074 82548 32086
rect 84232 32074 84238 32086
rect 82542 32046 84238 32074
rect 82542 32034 82548 32046
rect 84232 32034 84238 32046
rect 84290 32034 84296 32086
rect 83680 31966 83686 32018
rect 83738 32006 83744 32018
rect 85336 32006 85342 32018
rect 83738 31978 85342 32006
rect 83738 31966 83744 31978
rect 85336 31966 85342 31978
rect 85394 31966 85400 32018
rect 38 31916 3902 31938
rect 38 31864 2916 31916
rect 2968 31864 2980 31916
rect 3032 31864 3044 31916
rect 3096 31864 3108 31916
rect 3160 31864 3902 31916
rect 38 31842 3902 31864
rect 83298 31916 87806 31938
rect 83298 31864 86916 31916
rect 86968 31864 86980 31916
rect 87032 31864 87044 31916
rect 87096 31864 87108 31916
rect 87160 31864 87806 31916
rect 83298 31842 87806 31864
rect 83867 31465 83925 31471
rect 83867 31431 83879 31465
rect 83913 31462 83925 31465
rect 84048 31462 84054 31474
rect 83913 31434 84054 31462
rect 83913 31431 83925 31434
rect 83867 31425 83925 31431
rect 84048 31422 84054 31434
rect 84106 31462 84112 31474
rect 85980 31462 85986 31474
rect 84106 31434 85986 31462
rect 84106 31422 84112 31434
rect 85980 31422 85986 31434
rect 86038 31422 86044 31474
rect 38 31372 3902 31394
rect 38 31320 916 31372
rect 968 31320 980 31372
rect 1032 31320 1044 31372
rect 1096 31320 1108 31372
rect 1160 31320 3902 31372
rect 38 31298 3902 31320
rect 83298 31372 87806 31394
rect 83298 31320 84916 31372
rect 84968 31320 84980 31372
rect 85032 31320 85044 31372
rect 85096 31320 85108 31372
rect 85160 31320 87806 31372
rect 83298 31298 87806 31320
rect 82944 30878 82950 30930
rect 83002 30918 83008 30930
rect 84140 30918 84146 30930
rect 83002 30890 84146 30918
rect 83002 30878 83008 30890
rect 84140 30878 84146 30890
rect 84198 30878 84204 30930
rect 38 30828 3902 30850
rect 38 30776 2916 30828
rect 2968 30776 2980 30828
rect 3032 30776 3044 30828
rect 3096 30776 3108 30828
rect 3160 30776 3902 30828
rect 38 30754 3902 30776
rect 83298 30828 87806 30850
rect 83298 30776 86916 30828
rect 86968 30776 86980 30828
rect 87032 30776 87044 30828
rect 87096 30776 87108 30828
rect 87160 30776 87806 30828
rect 83298 30754 87806 30776
rect 38 30284 3902 30306
rect 38 30232 916 30284
rect 968 30232 980 30284
rect 1032 30232 1044 30284
rect 1096 30232 1108 30284
rect 1160 30232 3902 30284
rect 38 30210 3902 30232
rect 83298 30284 87806 30306
rect 83298 30232 84916 30284
rect 84968 30232 84980 30284
rect 85032 30232 85044 30284
rect 85096 30232 85108 30284
rect 85160 30232 87806 30284
rect 83298 30210 87806 30232
rect 83867 29901 83925 29907
rect 83867 29867 83879 29901
rect 83913 29898 83925 29901
rect 84048 29898 84054 29910
rect 83913 29870 84054 29898
rect 83913 29867 83925 29870
rect 83867 29861 83925 29867
rect 84048 29858 84054 29870
rect 84106 29858 84112 29910
rect 38 29740 3902 29762
rect 38 29688 2916 29740
rect 2968 29688 2980 29740
rect 3032 29688 3044 29740
rect 3096 29688 3108 29740
rect 3160 29688 3902 29740
rect 38 29666 3902 29688
rect 83298 29740 87806 29762
rect 83298 29688 86916 29740
rect 86968 29688 86980 29740
rect 87032 29688 87044 29740
rect 87096 29688 87108 29740
rect 87160 29688 87806 29740
rect 83298 29666 87806 29688
rect 3824 29450 3830 29502
rect 3882 29450 3888 29502
rect 81840 29450 81846 29502
rect 81898 29490 81904 29502
rect 84324 29490 84330 29502
rect 81898 29462 84330 29490
rect 81898 29450 81904 29462
rect 84324 29450 84330 29462
rect 84382 29450 84388 29502
rect 3842 29366 3870 29450
rect 84784 29422 84790 29434
rect 84342 29394 84790 29422
rect 84342 29366 84370 29394
rect 84784 29382 84790 29394
rect 84842 29382 84848 29434
rect 3824 29314 3830 29366
rect 3882 29314 3888 29366
rect 84324 29314 84330 29366
rect 84382 29314 84388 29366
rect 38 29196 3902 29218
rect 38 29144 916 29196
rect 968 29144 980 29196
rect 1032 29144 1044 29196
rect 1096 29144 1108 29196
rect 1160 29144 3902 29196
rect 38 29122 3902 29144
rect 83298 29196 87806 29218
rect 83298 29144 84916 29196
rect 84968 29144 84980 29196
rect 85032 29144 85044 29196
rect 85096 29144 85108 29196
rect 85160 29144 87806 29196
rect 83298 29122 87806 29144
rect 83867 28745 83925 28751
rect 83867 28711 83879 28745
rect 83913 28742 83925 28745
rect 84140 28742 84146 28754
rect 83913 28714 84146 28742
rect 83913 28711 83925 28714
rect 83867 28705 83925 28711
rect 84140 28702 84146 28714
rect 84198 28702 84204 28754
rect 38 28652 3902 28674
rect 38 28600 2916 28652
rect 2968 28600 2980 28652
rect 3032 28600 3044 28652
rect 3096 28600 3108 28652
rect 3160 28600 3902 28652
rect 38 28578 3902 28600
rect 83298 28652 87806 28674
rect 83298 28600 86916 28652
rect 86968 28600 86980 28652
rect 87032 28600 87044 28652
rect 87096 28600 87108 28652
rect 87160 28600 87806 28652
rect 83298 28578 87806 28600
rect 81748 28498 81754 28550
rect 81806 28538 81812 28550
rect 84416 28538 84422 28550
rect 81806 28510 84422 28538
rect 81806 28498 81812 28510
rect 84416 28498 84422 28510
rect 84474 28498 84480 28550
rect 83220 28226 83226 28278
rect 83278 28266 83284 28278
rect 85428 28266 85434 28278
rect 83278 28238 85434 28266
rect 83278 28226 83284 28238
rect 85428 28226 85434 28238
rect 85486 28226 85492 28278
rect 82852 28158 82858 28210
rect 82910 28198 82916 28210
rect 84692 28198 84698 28210
rect 82910 28170 84698 28198
rect 82910 28158 82916 28170
rect 84692 28158 84698 28170
rect 84750 28158 84756 28210
rect 38 28108 3902 28130
rect 38 28056 916 28108
rect 968 28056 980 28108
rect 1032 28056 1044 28108
rect 1096 28056 1108 28108
rect 1160 28056 3902 28108
rect 38 28034 3902 28056
rect 83298 28108 87806 28130
rect 83298 28056 84916 28108
rect 84968 28056 84980 28108
rect 85032 28056 85044 28108
rect 85096 28056 85108 28108
rect 85160 28056 87806 28108
rect 83298 28034 87806 28056
rect 38 27564 3902 27586
rect 38 27512 2916 27564
rect 2968 27512 2980 27564
rect 3032 27512 3044 27564
rect 3096 27512 3108 27564
rect 3160 27512 3902 27564
rect 38 27490 3902 27512
rect 83298 27564 87806 27586
rect 83298 27512 86916 27564
rect 86968 27512 86980 27564
rect 87032 27512 87044 27564
rect 87096 27512 87108 27564
rect 87160 27512 87806 27564
rect 83298 27490 87806 27512
rect 83867 27113 83925 27119
rect 83867 27079 83879 27113
rect 83913 27110 83925 27113
rect 84232 27110 84238 27122
rect 83913 27082 84238 27110
rect 83913 27079 83925 27082
rect 83867 27073 83925 27079
rect 84232 27070 84238 27082
rect 84290 27110 84296 27122
rect 84692 27110 84698 27122
rect 84290 27082 84698 27110
rect 84290 27070 84296 27082
rect 84692 27070 84698 27082
rect 84750 27070 84756 27122
rect 38 27020 3902 27042
rect 38 26968 916 27020
rect 968 26968 980 27020
rect 1032 26968 1044 27020
rect 1096 26968 1108 27020
rect 1160 26968 3902 27020
rect 38 26946 3902 26968
rect 83298 27020 87806 27042
rect 83298 26968 84916 27020
rect 84968 26968 84980 27020
rect 85032 26968 85044 27020
rect 85096 26968 85108 27020
rect 85160 26968 87806 27020
rect 83298 26946 87806 26968
rect 38 26476 3902 26498
rect 38 26424 2916 26476
rect 2968 26424 2980 26476
rect 3032 26424 3044 26476
rect 3096 26424 3108 26476
rect 3160 26424 3902 26476
rect 38 26402 3902 26424
rect 83298 26476 87806 26498
rect 83298 26424 86916 26476
rect 86968 26424 86980 26476
rect 87032 26424 87044 26476
rect 87096 26424 87108 26476
rect 87160 26424 87806 26476
rect 83298 26402 87806 26424
rect 83496 25982 83502 26034
rect 83554 26022 83560 26034
rect 83775 26025 83833 26031
rect 83775 26022 83787 26025
rect 83554 25994 83787 26022
rect 83554 25982 83560 25994
rect 83775 25991 83787 25994
rect 83821 25991 83833 26025
rect 83775 25985 83833 25991
rect 38 25932 3902 25954
rect 38 25880 916 25932
rect 968 25880 980 25932
rect 1032 25880 1044 25932
rect 1096 25880 1108 25932
rect 1160 25880 3902 25932
rect 38 25858 3902 25880
rect 83298 25932 87806 25954
rect 83298 25880 84916 25932
rect 84968 25880 84980 25932
rect 85032 25880 85044 25932
rect 85096 25880 85108 25932
rect 85160 25880 87806 25932
rect 83298 25858 87806 25880
rect 81656 25574 81662 25626
rect 81714 25614 81720 25626
rect 84876 25614 84882 25626
rect 81714 25586 84882 25614
rect 81714 25574 81720 25586
rect 84876 25574 84882 25586
rect 84934 25574 84940 25626
rect 3272 25506 3278 25558
rect 3330 25546 3336 25558
rect 3364 25546 3370 25558
rect 3330 25518 3370 25546
rect 3330 25506 3336 25518
rect 3364 25506 3370 25518
rect 3422 25506 3428 25558
rect 38 25388 3902 25410
rect 38 25336 2916 25388
rect 2968 25336 2980 25388
rect 3032 25336 3044 25388
rect 3096 25336 3108 25388
rect 3160 25336 3902 25388
rect 38 25314 3902 25336
rect 83298 25388 87806 25410
rect 83298 25336 86916 25388
rect 86968 25336 86980 25388
rect 87032 25336 87044 25388
rect 87096 25336 87108 25388
rect 87160 25336 87806 25388
rect 83298 25314 87806 25336
rect 38 24844 3902 24866
rect 38 24792 916 24844
rect 968 24792 980 24844
rect 1032 24792 1044 24844
rect 1096 24792 1108 24844
rect 1160 24792 3902 24844
rect 38 24770 3902 24792
rect 83298 24844 87806 24866
rect 83298 24792 84916 24844
rect 84968 24792 84980 24844
rect 85032 24792 85044 24844
rect 85096 24792 85108 24844
rect 85160 24792 87806 24844
rect 83298 24770 87806 24792
rect 38 24300 3902 24322
rect 38 24248 2916 24300
rect 2968 24248 2980 24300
rect 3032 24248 3044 24300
rect 3096 24248 3108 24300
rect 3160 24248 3902 24300
rect 38 24226 3902 24248
rect 83298 24300 87806 24322
rect 83298 24248 86916 24300
rect 86968 24248 86980 24300
rect 87032 24248 87044 24300
rect 87096 24248 87108 24300
rect 87160 24248 87806 24300
rect 83298 24226 87806 24248
rect 3272 24146 3278 24198
rect 3330 24186 3336 24198
rect 4103 24189 4161 24195
rect 4103 24186 4115 24189
rect 3330 24158 4115 24186
rect 3330 24146 3336 24158
rect 4103 24155 4115 24158
rect 4149 24155 4161 24189
rect 4103 24149 4161 24155
rect 84232 24010 84238 24062
rect 84290 24050 84296 24062
rect 84692 24050 84698 24062
rect 84290 24022 84698 24050
rect 84290 24010 84296 24022
rect 84692 24010 84698 24022
rect 84750 24010 84756 24062
rect 83867 23849 83925 23855
rect 83867 23815 83879 23849
rect 83913 23846 83925 23849
rect 84232 23846 84238 23858
rect 83913 23818 84238 23846
rect 83913 23815 83925 23818
rect 83867 23809 83925 23815
rect 84232 23806 84238 23818
rect 84290 23806 84296 23858
rect 38 23756 3902 23778
rect 38 23704 916 23756
rect 968 23704 980 23756
rect 1032 23704 1044 23756
rect 1096 23704 1108 23756
rect 1160 23704 3902 23756
rect 38 23682 3902 23704
rect 83298 23756 87806 23778
rect 83298 23704 84916 23756
rect 84968 23704 84980 23756
rect 85032 23704 85044 23756
rect 85096 23704 85108 23756
rect 85160 23704 87806 23756
rect 83298 23682 87806 23704
rect 38 23212 3902 23234
rect 38 23160 2916 23212
rect 2968 23160 2980 23212
rect 3032 23160 3044 23212
rect 3096 23160 3108 23212
rect 3160 23160 3902 23212
rect 38 23138 3902 23160
rect 83298 23212 87806 23234
rect 83298 23160 86916 23212
rect 86968 23160 86980 23212
rect 87032 23160 87044 23212
rect 87096 23160 87108 23212
rect 87160 23160 87806 23212
rect 83298 23138 87806 23160
rect 3824 22922 3830 22974
rect 3882 22962 3888 22974
rect 4011 22965 4069 22971
rect 4011 22962 4023 22965
rect 3882 22934 4023 22962
rect 3882 22922 3888 22934
rect 4011 22931 4023 22934
rect 4057 22931 4069 22965
rect 4011 22925 4069 22931
rect 83867 22965 83925 22971
rect 83867 22931 83879 22965
rect 83913 22962 83925 22965
rect 83956 22962 83962 22974
rect 83913 22934 83962 22962
rect 83913 22931 83925 22934
rect 83867 22925 83925 22931
rect 83956 22922 83962 22934
rect 84014 22922 84020 22974
rect 38 22668 3902 22690
rect 38 22616 916 22668
rect 968 22616 980 22668
rect 1032 22616 1044 22668
rect 1096 22616 1108 22668
rect 1160 22616 3902 22668
rect 38 22594 3902 22616
rect 83298 22668 87806 22690
rect 83298 22616 84916 22668
rect 84968 22616 84980 22668
rect 85032 22616 85044 22668
rect 85096 22616 85108 22668
rect 85160 22616 87806 22668
rect 83298 22594 87806 22616
rect 3551 22557 3609 22563
rect 3551 22523 3563 22557
rect 3597 22554 3609 22557
rect 3824 22554 3830 22566
rect 3597 22526 3830 22554
rect 3597 22523 3609 22526
rect 3551 22517 3609 22523
rect 3824 22514 3830 22526
rect 3882 22514 3888 22566
rect 38 22124 3902 22146
rect 38 22072 2916 22124
rect 2968 22072 2980 22124
rect 3032 22072 3044 22124
rect 3096 22072 3108 22124
rect 3160 22072 3902 22124
rect 38 22050 3902 22072
rect 83298 22124 87806 22146
rect 83298 22072 86916 22124
rect 86968 22072 86980 22124
rect 87032 22072 87044 22124
rect 87096 22072 87108 22124
rect 87160 22072 87806 22124
rect 83298 22050 87806 22072
rect 38 21580 3902 21602
rect 38 21528 916 21580
rect 968 21528 980 21580
rect 1032 21528 1044 21580
rect 1096 21528 1108 21580
rect 1160 21528 3902 21580
rect 38 21506 3902 21528
rect 83298 21580 87806 21602
rect 83298 21528 84916 21580
rect 84968 21528 84980 21580
rect 85032 21528 85044 21580
rect 85096 21528 85108 21580
rect 85160 21528 87806 21580
rect 83298 21506 87806 21528
rect 38 21036 3902 21058
rect 38 20984 2916 21036
rect 2968 20984 2980 21036
rect 3032 20984 3044 21036
rect 3096 20984 3108 21036
rect 3160 20984 3902 21036
rect 38 20962 3902 20984
rect 83298 21036 87806 21058
rect 83298 20984 86916 21036
rect 86968 20984 86980 21036
rect 87032 20984 87044 21036
rect 87096 20984 87108 21036
rect 87160 20984 87806 21036
rect 83298 20962 87806 20984
rect 3551 20585 3609 20591
rect 3551 20551 3563 20585
rect 3597 20582 3609 20585
rect 4284 20582 4290 20594
rect 3597 20554 4290 20582
rect 3597 20551 3609 20554
rect 3551 20545 3609 20551
rect 4284 20542 4290 20554
rect 4342 20542 4348 20594
rect 38 20492 3902 20514
rect 38 20440 916 20492
rect 968 20440 980 20492
rect 1032 20440 1044 20492
rect 1096 20440 1108 20492
rect 1160 20440 3902 20492
rect 38 20418 3902 20440
rect 83298 20492 87806 20514
rect 83298 20440 84916 20492
rect 84968 20440 84980 20492
rect 85032 20440 85044 20492
rect 85096 20440 85108 20492
rect 85160 20440 87806 20492
rect 83298 20418 87806 20440
rect 83496 20202 83502 20254
rect 83554 20242 83560 20254
rect 84784 20242 84790 20254
rect 83554 20214 84790 20242
rect 83554 20202 83560 20214
rect 84784 20202 84790 20214
rect 84842 20202 84848 20254
rect 83496 19998 83502 20050
rect 83554 20038 83560 20050
rect 84048 20038 84054 20050
rect 83554 20010 84054 20038
rect 83554 19998 83560 20010
rect 84048 19998 84054 20010
rect 84106 19998 84112 20050
rect 38 19948 3902 19970
rect 38 19896 2916 19948
rect 2968 19896 2980 19948
rect 3032 19896 3044 19948
rect 3096 19896 3108 19948
rect 3160 19896 3902 19948
rect 38 19874 3902 19896
rect 83298 19948 87806 19970
rect 83298 19896 86916 19948
rect 86968 19896 86980 19948
rect 87032 19896 87044 19948
rect 87096 19896 87108 19948
rect 87160 19896 87806 19948
rect 83298 19874 87806 19896
rect 82576 19590 82582 19642
rect 82634 19630 82640 19642
rect 85520 19630 85526 19642
rect 82634 19602 85526 19630
rect 82634 19590 82640 19602
rect 85520 19590 85526 19602
rect 85578 19590 85584 19642
rect 38 19404 3902 19426
rect 38 19352 916 19404
rect 968 19352 980 19404
rect 1032 19352 1044 19404
rect 1096 19352 1108 19404
rect 1160 19352 3902 19404
rect 38 19330 3902 19352
rect 83298 19404 87806 19426
rect 83298 19352 84916 19404
rect 84968 19352 84980 19404
rect 85032 19352 85044 19404
rect 85096 19352 85108 19404
rect 85160 19352 87806 19404
rect 83298 19330 87806 19352
rect 38 18860 3902 18882
rect 38 18808 2916 18860
rect 2968 18808 2980 18860
rect 3032 18808 3044 18860
rect 3096 18808 3108 18860
rect 3160 18808 3902 18860
rect 38 18786 3902 18808
rect 83298 18860 87806 18882
rect 83298 18808 86916 18860
rect 86968 18808 86980 18860
rect 87032 18808 87044 18860
rect 87096 18808 87108 18860
rect 87160 18808 87806 18860
rect 83298 18786 87806 18808
rect 83496 18366 83502 18418
rect 83554 18406 83560 18418
rect 83956 18406 83962 18418
rect 83554 18378 83962 18406
rect 83554 18366 83560 18378
rect 83956 18366 83962 18378
rect 84014 18366 84020 18418
rect 38 18316 3902 18338
rect 38 18264 916 18316
rect 968 18264 980 18316
rect 1032 18264 1044 18316
rect 1096 18264 1108 18316
rect 1160 18264 3902 18316
rect 38 18242 3902 18264
rect 83298 18316 87806 18338
rect 83298 18264 84916 18316
rect 84968 18264 84980 18316
rect 85032 18264 85044 18316
rect 85096 18264 85108 18316
rect 85160 18264 87806 18316
rect 83298 18242 87806 18264
rect 38 17772 3902 17794
rect 38 17720 2916 17772
rect 2968 17720 2980 17772
rect 3032 17720 3044 17772
rect 3096 17720 3108 17772
rect 3160 17720 3902 17772
rect 38 17698 3902 17720
rect 83298 17772 87806 17794
rect 83298 17720 86916 17772
rect 86968 17720 86980 17772
rect 87032 17720 87044 17772
rect 87096 17720 87108 17772
rect 87160 17720 87806 17772
rect 83298 17698 87806 17720
rect 38 17228 3902 17250
rect 38 17176 916 17228
rect 968 17176 980 17228
rect 1032 17176 1044 17228
rect 1096 17176 1108 17228
rect 1160 17176 3902 17228
rect 38 17154 3902 17176
rect 83298 17228 87806 17250
rect 83298 17176 84916 17228
rect 84968 17176 84980 17228
rect 85032 17176 85044 17228
rect 85096 17176 85108 17228
rect 85160 17176 87806 17228
rect 83298 17154 87806 17176
rect 38 16684 3902 16706
rect 38 16632 2916 16684
rect 2968 16632 2980 16684
rect 3032 16632 3044 16684
rect 3096 16632 3108 16684
rect 3160 16632 3902 16684
rect 38 16610 3902 16632
rect 83298 16684 87806 16706
rect 83298 16632 86916 16684
rect 86968 16632 86980 16684
rect 87032 16632 87044 16684
rect 87096 16632 87108 16684
rect 87160 16632 87806 16684
rect 83298 16610 87806 16632
rect 3916 16530 3922 16582
rect 3974 16570 3980 16582
rect 4011 16573 4069 16579
rect 4011 16570 4023 16573
rect 3974 16542 4023 16570
rect 3974 16530 3980 16542
rect 4011 16539 4023 16542
rect 4057 16539 4069 16573
rect 4011 16533 4069 16539
rect 38 16140 3902 16162
rect 38 16088 916 16140
rect 968 16088 980 16140
rect 1032 16088 1044 16140
rect 1096 16088 1108 16140
rect 1160 16088 3902 16140
rect 38 16066 3902 16088
rect 83298 16140 87806 16162
rect 83298 16088 84916 16140
rect 84968 16088 84980 16140
rect 85032 16088 85044 16140
rect 85096 16088 85108 16140
rect 85160 16088 87806 16140
rect 83298 16066 87806 16088
rect 84324 15850 84330 15902
rect 84382 15890 84388 15902
rect 84600 15890 84606 15902
rect 84382 15862 84606 15890
rect 84382 15850 84388 15862
rect 84600 15850 84606 15862
rect 84658 15850 84664 15902
rect 38 15596 3902 15618
rect 38 15544 2916 15596
rect 2968 15544 2980 15596
rect 3032 15544 3044 15596
rect 3096 15544 3108 15596
rect 3160 15544 3902 15596
rect 38 15522 3902 15544
rect 83298 15596 87806 15618
rect 83298 15544 86916 15596
rect 86968 15544 86980 15596
rect 87032 15544 87044 15596
rect 87096 15544 87108 15596
rect 87160 15544 87806 15596
rect 83298 15522 87806 15544
rect 3272 15238 3278 15290
rect 3330 15278 3336 15290
rect 4103 15281 4161 15287
rect 4103 15278 4115 15281
rect 3330 15250 4115 15278
rect 3330 15238 3336 15250
rect 4103 15247 4115 15250
rect 4149 15247 4161 15281
rect 4103 15241 4161 15247
rect 38 15052 3902 15074
rect 38 15000 916 15052
rect 968 15000 980 15052
rect 1032 15000 1044 15052
rect 1096 15000 1108 15052
rect 1160 15000 3902 15052
rect 38 14978 3902 15000
rect 83298 15052 87806 15074
rect 83298 15000 84916 15052
rect 84968 15000 84980 15052
rect 85032 15000 85044 15052
rect 85096 15000 85108 15052
rect 85160 15000 87806 15052
rect 83298 14978 87806 15000
rect 38 14508 3902 14530
rect 38 14456 2916 14508
rect 2968 14456 2980 14508
rect 3032 14456 3044 14508
rect 3096 14456 3108 14508
rect 3160 14456 3902 14508
rect 38 14434 3902 14456
rect 83298 14508 87806 14530
rect 83298 14456 86916 14508
rect 86968 14456 86980 14508
rect 87032 14456 87044 14508
rect 87096 14456 87108 14508
rect 87160 14456 87806 14508
rect 83298 14434 87806 14456
rect 38 13964 3902 13986
rect 38 13912 916 13964
rect 968 13912 980 13964
rect 1032 13912 1044 13964
rect 1096 13912 1108 13964
rect 1160 13912 3902 13964
rect 38 13890 3902 13912
rect 83298 13964 87806 13986
rect 83298 13912 84916 13964
rect 84968 13912 84980 13964
rect 85032 13912 85044 13964
rect 85096 13912 85108 13964
rect 85160 13912 87806 13964
rect 83298 13890 87806 13912
rect 83772 13810 83778 13862
rect 83830 13850 83836 13862
rect 84140 13850 84146 13862
rect 83830 13822 84146 13850
rect 83830 13810 83836 13822
rect 84140 13810 84146 13822
rect 84198 13810 84204 13862
rect 3272 13606 3278 13658
rect 3330 13646 3336 13658
rect 4011 13649 4069 13655
rect 4011 13646 4023 13649
rect 3330 13618 4023 13646
rect 3330 13606 3336 13618
rect 4011 13615 4023 13618
rect 4057 13615 4069 13649
rect 4011 13609 4069 13615
rect 38 13420 3902 13442
rect 38 13368 2916 13420
rect 2968 13368 2980 13420
rect 3032 13368 3044 13420
rect 3096 13368 3108 13420
rect 3160 13368 3902 13420
rect 38 13346 3902 13368
rect 83298 13420 87806 13442
rect 83298 13368 86916 13420
rect 86968 13368 86980 13420
rect 87032 13368 87044 13420
rect 87096 13368 87108 13420
rect 87160 13368 87806 13420
rect 83298 13346 87806 13368
rect 38 12876 3902 12898
rect 38 12824 916 12876
rect 968 12824 980 12876
rect 1032 12824 1044 12876
rect 1096 12824 1108 12876
rect 1160 12824 3902 12876
rect 38 12802 3902 12824
rect 83298 12876 87806 12898
rect 83298 12824 84916 12876
rect 84968 12824 84980 12876
rect 85032 12824 85044 12876
rect 85096 12824 85108 12876
rect 85160 12824 87806 12876
rect 83298 12802 87806 12824
rect 38 12332 3902 12354
rect 38 12280 2916 12332
rect 2968 12280 2980 12332
rect 3032 12280 3044 12332
rect 3096 12280 3108 12332
rect 3160 12280 3902 12332
rect 38 12258 3902 12280
rect 83298 12332 87806 12354
rect 83298 12280 86916 12332
rect 86968 12280 86980 12332
rect 87032 12280 87044 12332
rect 87096 12280 87108 12332
rect 87160 12280 87806 12332
rect 83298 12258 87806 12280
rect 38 11788 3902 11810
rect 38 11736 916 11788
rect 968 11736 980 11788
rect 1032 11736 1044 11788
rect 1096 11736 1108 11788
rect 1160 11736 3902 11788
rect 38 11714 3902 11736
rect 83298 11788 87806 11810
rect 83298 11736 84916 11788
rect 84968 11736 84980 11788
rect 85032 11736 85044 11788
rect 85096 11736 85108 11788
rect 85160 11736 87806 11788
rect 83298 11714 87806 11736
rect 3916 11470 3922 11482
rect 3842 11442 3922 11470
rect 3842 11414 3870 11442
rect 3916 11430 3922 11442
rect 3974 11430 3980 11482
rect 5572 11470 5578 11482
rect 5498 11442 5578 11470
rect 5498 11414 5526 11442
rect 5572 11430 5578 11442
rect 5630 11430 5636 11482
rect 3824 11362 3830 11414
rect 3882 11362 3888 11414
rect 5480 11362 5486 11414
rect 5538 11362 5544 11414
rect 38 11244 3902 11266
rect 38 11192 2916 11244
rect 2968 11192 2980 11244
rect 3032 11192 3044 11244
rect 3096 11192 3108 11244
rect 3160 11192 3902 11244
rect 38 11170 3902 11192
rect 83298 11244 87806 11266
rect 83298 11192 86916 11244
rect 86968 11192 86980 11244
rect 87032 11192 87044 11244
rect 87096 11192 87108 11244
rect 87160 11192 87806 11244
rect 83298 11170 87806 11192
rect 38 10700 3902 10722
rect 38 10648 916 10700
rect 968 10648 980 10700
rect 1032 10648 1044 10700
rect 1096 10648 1108 10700
rect 1160 10648 3902 10700
rect 38 10626 3902 10648
rect 83298 10700 87806 10722
rect 83298 10648 84916 10700
rect 84968 10648 84980 10700
rect 85032 10648 85044 10700
rect 85096 10648 85108 10700
rect 85160 10648 87806 10700
rect 83298 10626 87806 10648
rect 38 10156 3902 10178
rect 38 10104 2916 10156
rect 2968 10104 2980 10156
rect 3032 10104 3044 10156
rect 3096 10104 3108 10156
rect 3160 10104 3902 10156
rect 38 10082 3902 10104
rect 83298 10156 87806 10178
rect 83298 10104 86916 10156
rect 86968 10104 86980 10156
rect 87032 10104 87044 10156
rect 87096 10104 87108 10156
rect 87160 10104 87806 10156
rect 83298 10082 87806 10104
rect 38 9612 3902 9634
rect 38 9560 916 9612
rect 968 9560 980 9612
rect 1032 9560 1044 9612
rect 1096 9560 1108 9612
rect 1160 9560 3902 9612
rect 38 9538 3902 9560
rect 83298 9612 87806 9634
rect 83298 9560 84916 9612
rect 84968 9560 84980 9612
rect 85032 9560 85044 9612
rect 85096 9560 85108 9612
rect 85160 9560 87806 9612
rect 83298 9538 87806 9560
rect 38 9068 3902 9090
rect 38 9016 2916 9068
rect 2968 9016 2980 9068
rect 3032 9016 3044 9068
rect 3096 9016 3108 9068
rect 3160 9016 3902 9068
rect 38 8994 3902 9016
rect 83298 9068 87806 9090
rect 83298 9016 86916 9068
rect 86968 9016 86980 9068
rect 87032 9016 87044 9068
rect 87096 9016 87108 9068
rect 87160 9016 87806 9068
rect 83298 8994 87806 9016
rect 82576 8818 82582 8830
rect 82537 8790 82582 8818
rect 82576 8778 82582 8790
rect 82634 8778 82640 8830
rect 38 8524 3902 8546
rect 38 8472 916 8524
rect 968 8472 980 8524
rect 1032 8472 1044 8524
rect 1096 8472 1108 8524
rect 1160 8472 3902 8524
rect 38 8450 3902 8472
rect 83298 8524 87806 8546
rect 83298 8472 84916 8524
rect 84968 8472 84980 8524
rect 85032 8472 85044 8524
rect 85096 8472 85108 8524
rect 85160 8472 87806 8524
rect 83298 8450 87806 8472
rect 38 7980 3902 8002
rect 38 7928 2916 7980
rect 2968 7928 2980 7980
rect 3032 7928 3044 7980
rect 3096 7928 3108 7980
rect 3160 7928 3902 7980
rect 38 7906 3902 7928
rect 83298 7980 87806 8002
rect 83298 7928 86916 7980
rect 86968 7928 86980 7980
rect 87032 7928 87044 7980
rect 87096 7928 87108 7980
rect 87160 7928 87806 7980
rect 83298 7906 87806 7928
rect 82576 7554 82582 7606
rect 82634 7594 82640 7606
rect 85060 7594 85066 7606
rect 82634 7566 85066 7594
rect 82634 7554 82640 7566
rect 85060 7554 85066 7566
rect 85118 7554 85124 7606
rect 38 7436 3902 7458
rect 38 7384 916 7436
rect 968 7384 980 7436
rect 1032 7384 1044 7436
rect 1096 7384 1108 7436
rect 1160 7384 3902 7436
rect 38 7362 3902 7384
rect 83298 7436 87806 7458
rect 83298 7384 84916 7436
rect 84968 7384 84980 7436
rect 85032 7384 85044 7436
rect 85096 7384 85108 7436
rect 85160 7384 87806 7436
rect 83298 7362 87806 7384
rect 84324 7146 84330 7198
rect 84382 7186 84388 7198
rect 84784 7186 84790 7198
rect 84382 7158 84790 7186
rect 84382 7146 84388 7158
rect 84784 7146 84790 7158
rect 84842 7146 84848 7198
rect 81564 7010 81570 7062
rect 81622 7050 81628 7062
rect 82024 7050 82030 7062
rect 81622 7022 82030 7050
rect 81622 7010 81628 7022
rect 82024 7010 82030 7022
rect 82082 7010 82088 7062
rect 38 6892 3902 6914
rect 38 6840 2916 6892
rect 2968 6840 2980 6892
rect 3032 6840 3044 6892
rect 3096 6840 3108 6892
rect 3160 6840 3902 6892
rect 82024 6874 82030 6926
rect 82082 6914 82088 6926
rect 82392 6914 82398 6926
rect 82082 6886 82398 6914
rect 82082 6874 82088 6886
rect 82392 6874 82398 6886
rect 82450 6874 82456 6926
rect 83298 6892 87806 6914
rect 38 6818 3902 6840
rect 83298 6840 86916 6892
rect 86968 6840 86980 6892
rect 87032 6840 87044 6892
rect 87096 6840 87108 6892
rect 87160 6840 87806 6892
rect 83298 6818 87806 6840
rect 38 6348 3902 6370
rect 38 6296 916 6348
rect 968 6296 980 6348
rect 1032 6296 1044 6348
rect 1096 6296 1108 6348
rect 1160 6296 3902 6348
rect 38 6274 3902 6296
rect 83298 6348 87806 6370
rect 83298 6296 84916 6348
rect 84968 6296 84980 6348
rect 85032 6296 85044 6348
rect 85096 6296 85108 6348
rect 85160 6296 87806 6348
rect 83298 6274 87806 6296
rect 3640 6194 3646 6246
rect 3698 6234 3704 6246
rect 5756 6234 5762 6246
rect 3698 6206 5762 6234
rect 3698 6194 3704 6206
rect 5756 6194 5762 6206
rect 5814 6194 5820 6246
rect 38 5804 3902 5826
rect 38 5752 2916 5804
rect 2968 5752 2980 5804
rect 3032 5752 3044 5804
rect 3096 5752 3108 5804
rect 3160 5752 3902 5804
rect 38 5730 3902 5752
rect 83298 5804 87806 5826
rect 83298 5752 86916 5804
rect 86968 5752 86980 5804
rect 87032 5752 87044 5804
rect 87096 5752 87108 5804
rect 87160 5752 87806 5804
rect 83298 5730 87806 5752
rect 38 5260 3902 5282
rect 38 5208 916 5260
rect 968 5208 980 5260
rect 1032 5208 1044 5260
rect 1096 5208 1108 5260
rect 1160 5208 3902 5260
rect 38 5186 3902 5208
rect 83298 5260 87806 5282
rect 83298 5208 84916 5260
rect 84968 5208 84980 5260
rect 85032 5208 85044 5260
rect 85096 5208 85108 5260
rect 85160 5208 87806 5260
rect 83298 5186 87806 5208
rect 3551 5149 3609 5155
rect 3551 5115 3563 5149
rect 3597 5146 3609 5149
rect 3640 5146 3646 5158
rect 3597 5118 3646 5146
rect 3597 5115 3609 5118
rect 3551 5109 3609 5115
rect 3640 5106 3646 5118
rect 3698 5106 3704 5158
rect 4468 4834 4474 4886
rect 4526 4834 4532 4886
rect 38 4716 3902 4738
rect 38 4664 2916 4716
rect 2968 4664 2980 4716
rect 3032 4664 3044 4716
rect 3096 4664 3108 4716
rect 3160 4664 3902 4716
rect 38 4642 3902 4664
rect 3551 4605 3609 4611
rect 3551 4571 3563 4605
rect 3597 4602 3609 4605
rect 4376 4602 4382 4614
rect 3597 4574 4382 4602
rect 3597 4571 3609 4574
rect 3551 4565 3609 4571
rect 4376 4562 4382 4574
rect 4434 4562 4440 4614
rect 4486 4534 4514 4834
rect 83298 4716 87806 4738
rect 83298 4664 86916 4716
rect 86968 4664 86980 4716
rect 87032 4664 87044 4716
rect 87096 4664 87108 4716
rect 87160 4664 87806 4716
rect 83298 4642 87806 4664
rect 4394 4506 4514 4534
rect 4394 4478 4422 4506
rect 4376 4426 4382 4478
rect 4434 4426 4440 4478
rect 1524 4222 1530 4274
rect 1582 4262 1588 4274
rect 2815 4265 2873 4271
rect 2815 4262 2827 4265
rect 1582 4234 2827 4262
rect 1582 4222 1588 4234
rect 2815 4231 2827 4234
rect 2861 4262 2873 4265
rect 2904 4262 2910 4274
rect 2861 4234 2910 4262
rect 2861 4231 2873 4234
rect 2815 4225 2873 4231
rect 2904 4222 2910 4234
rect 2962 4222 2968 4274
rect 38 4172 3902 4194
rect 38 4120 916 4172
rect 968 4120 980 4172
rect 1032 4120 1044 4172
rect 1096 4120 1108 4172
rect 1160 4120 3902 4172
rect 38 4098 3902 4120
rect 83298 4172 87806 4194
rect 83298 4120 84916 4172
rect 84968 4120 84980 4172
rect 85032 4120 85044 4172
rect 85096 4120 85108 4172
rect 85160 4120 87806 4172
rect 83298 4098 87806 4120
rect 1984 4058 1990 4070
rect 1945 4030 1990 4058
rect 1984 4018 1990 4030
rect 2042 4058 2048 4070
rect 2260 4058 2266 4070
rect 2042 4030 2266 4058
rect 2042 4018 2048 4030
rect 2260 4018 2266 4030
rect 2318 4018 2324 4070
rect 2447 4061 2505 4067
rect 2447 4027 2459 4061
rect 2493 4058 2505 4061
rect 2536 4058 2542 4070
rect 2493 4030 2542 4058
rect 2493 4027 2505 4030
rect 2447 4021 2505 4027
rect 2536 4018 2542 4030
rect 2594 4018 2600 4070
rect 2812 4058 2818 4070
rect 2773 4030 2818 4058
rect 2812 4018 2818 4030
rect 2870 4058 2876 4070
rect 3916 4058 3922 4070
rect 2870 4030 3922 4058
rect 2870 4018 2876 4030
rect 3916 4018 3922 4030
rect 3974 4018 3980 4070
rect 82763 4061 82821 4067
rect 82763 4027 82775 4061
rect 82809 4058 82821 4061
rect 83772 4058 83778 4070
rect 82809 4030 83778 4058
rect 82809 4027 82821 4030
rect 82763 4021 82821 4027
rect 83772 4018 83778 4030
rect 83830 4018 83836 4070
rect 3364 3950 3370 4002
rect 3422 3990 3428 4002
rect 3551 3993 3609 3999
rect 3551 3990 3563 3993
rect 3422 3962 3563 3990
rect 3422 3950 3428 3962
rect 3551 3959 3563 3962
rect 3597 3990 3609 3993
rect 5020 3990 5026 4002
rect 3597 3962 5026 3990
rect 3597 3959 3609 3962
rect 3551 3953 3609 3959
rect 5020 3950 5026 3962
rect 5078 3950 5084 4002
rect 3183 3925 3241 3931
rect 3183 3891 3195 3925
rect 3229 3922 3241 3925
rect 5296 3922 5302 3934
rect 3229 3894 5302 3922
rect 3229 3891 3241 3894
rect 3183 3885 3241 3891
rect 5296 3882 5302 3894
rect 5354 3882 5360 3934
rect 81383 3721 81441 3727
rect 81383 3687 81395 3721
rect 81429 3718 81441 3721
rect 83588 3718 83594 3730
rect 81429 3690 83594 3718
rect 81429 3687 81441 3690
rect 81383 3681 81441 3687
rect 83588 3678 83594 3690
rect 83646 3678 83652 3730
rect 38 3628 3902 3650
rect 38 3576 2916 3628
rect 2968 3576 2980 3628
rect 3032 3576 3044 3628
rect 3096 3576 3108 3628
rect 3160 3576 3902 3628
rect 82392 3610 82398 3662
rect 82450 3650 82456 3662
rect 82760 3650 82766 3662
rect 82450 3622 82766 3650
rect 82450 3610 82456 3622
rect 82760 3610 82766 3622
rect 82818 3610 82824 3662
rect 83298 3628 87806 3650
rect 38 3554 3902 3576
rect 83298 3576 86916 3628
rect 86968 3576 86980 3628
rect 87032 3576 87044 3628
rect 87096 3576 87108 3628
rect 87160 3576 87806 3628
rect 83298 3554 87806 3576
rect 2815 3517 2873 3523
rect 2815 3483 2827 3517
rect 2861 3514 2873 3517
rect 3272 3514 3278 3526
rect 2861 3486 3278 3514
rect 2861 3483 2873 3486
rect 2815 3477 2873 3483
rect 3272 3474 3278 3486
rect 3330 3474 3336 3526
rect 82760 3514 82766 3526
rect 82721 3486 82766 3514
rect 82760 3474 82766 3486
rect 82818 3474 82824 3526
rect 84051 3517 84109 3523
rect 84051 3483 84063 3517
rect 84097 3514 84109 3517
rect 84603 3517 84661 3523
rect 84603 3514 84615 3517
rect 84097 3486 84615 3514
rect 84097 3483 84109 3486
rect 84051 3477 84109 3483
rect 84603 3483 84615 3486
rect 84649 3514 84661 3517
rect 85428 3514 85434 3526
rect 84649 3486 85434 3514
rect 84649 3483 84661 3486
rect 84603 3477 84661 3483
rect 85428 3474 85434 3486
rect 85486 3474 85492 3526
rect 2076 3406 2082 3458
rect 2134 3446 2140 3458
rect 2352 3446 2358 3458
rect 2134 3418 2358 3446
rect 2134 3406 2140 3418
rect 2352 3406 2358 3418
rect 2410 3446 2416 3458
rect 5759 3449 5817 3455
rect 5759 3446 5771 3449
rect 2410 3418 5771 3446
rect 2410 3406 2416 3418
rect 5759 3415 5771 3418
rect 5805 3415 5817 3449
rect 5759 3409 5817 3415
rect 2812 3338 2818 3390
rect 2870 3378 2876 3390
rect 4468 3378 4474 3390
rect 2870 3350 4474 3378
rect 2870 3338 2876 3350
rect 4468 3338 4474 3350
rect 4526 3338 4532 3390
rect 81291 3381 81349 3387
rect 81291 3347 81303 3381
rect 81337 3378 81349 3381
rect 85796 3378 85802 3390
rect 81337 3350 85802 3378
rect 81337 3347 81349 3350
rect 81291 3341 81349 3347
rect 85796 3338 85802 3350
rect 85854 3338 85860 3390
rect 2079 3313 2137 3319
rect 2079 3279 2091 3313
rect 2125 3310 2137 3313
rect 4011 3313 4069 3319
rect 4011 3310 4023 3313
rect 2125 3282 4023 3310
rect 2125 3279 2137 3282
rect 2079 3273 2137 3279
rect 4011 3279 4023 3282
rect 4057 3279 4069 3313
rect 84051 3313 84109 3319
rect 84051 3310 84063 3313
rect 4011 3273 4069 3279
rect 82318 3282 84063 3310
rect 1708 3242 1714 3254
rect 1621 3214 1714 3242
rect 1708 3202 1714 3214
rect 1766 3242 1772 3254
rect 4655 3245 4713 3251
rect 4655 3242 4667 3245
rect 1766 3214 2950 3242
rect 1766 3202 1772 3214
rect 1340 3174 1346 3186
rect 1301 3146 1346 3174
rect 1340 3134 1346 3146
rect 1398 3134 1404 3186
rect 2444 3174 2450 3186
rect 2405 3146 2450 3174
rect 2444 3134 2450 3146
rect 2502 3134 2508 3186
rect 2922 3174 2950 3214
rect 3474 3214 4667 3242
rect 3474 3174 3502 3214
rect 4655 3211 4667 3214
rect 4701 3211 4713 3245
rect 4655 3205 4713 3211
rect 2922 3146 3502 3174
rect 3551 3177 3609 3183
rect 3551 3143 3563 3177
rect 3597 3174 3609 3177
rect 3597 3146 5894 3174
rect 3597 3143 3609 3146
rect 3551 3137 3609 3143
rect 38 3084 3902 3106
rect 38 3032 916 3084
rect 968 3032 980 3084
rect 1032 3032 1044 3084
rect 1096 3032 1108 3084
rect 1160 3032 3902 3084
rect 38 3010 3902 3032
rect 5866 3038 5894 3146
rect 8700 3038 8706 3050
rect 5866 3010 8706 3038
rect 8700 2998 8706 3010
rect 8758 2998 8764 3050
rect 36944 2998 36950 3050
rect 37002 3038 37008 3050
rect 82208 3038 82214 3050
rect 37002 3010 82214 3038
rect 37002 2998 37008 3010
rect 82208 2998 82214 3010
rect 82266 2998 82272 3050
rect 1343 2973 1401 2979
rect 1343 2939 1355 2973
rect 1389 2970 1401 2973
rect 2352 2970 2358 2982
rect 1389 2942 2358 2970
rect 1389 2939 1401 2942
rect 1343 2933 1401 2939
rect 2352 2930 2358 2942
rect 2410 2930 2416 2982
rect 2812 2970 2818 2982
rect 2773 2942 2818 2970
rect 2812 2930 2818 2942
rect 2870 2930 2876 2982
rect 3272 2930 3278 2982
rect 3330 2970 3336 2982
rect 33724 2970 33730 2982
rect 3330 2942 33730 2970
rect 3330 2930 3336 2942
rect 33724 2930 33730 2942
rect 33782 2930 33788 2982
rect 53688 2930 53694 2982
rect 53746 2970 53752 2982
rect 82318 2970 82346 3282
rect 84051 3279 84063 3282
rect 84097 3279 84109 3313
rect 84051 3273 84109 3279
rect 82392 3202 82398 3254
rect 82450 3242 82456 3254
rect 84143 3245 84201 3251
rect 84143 3242 84155 3245
rect 82450 3214 84155 3242
rect 82450 3202 82456 3214
rect 84143 3211 84155 3214
rect 84189 3211 84201 3245
rect 84143 3205 84201 3211
rect 83772 3174 83778 3186
rect 83733 3146 83778 3174
rect 83772 3134 83778 3146
rect 83830 3134 83836 3186
rect 83298 3084 87806 3106
rect 83298 3032 84916 3084
rect 84968 3032 84980 3084
rect 85032 3032 85044 3084
rect 85096 3032 85108 3084
rect 85160 3032 87806 3084
rect 83298 3010 87806 3032
rect 53746 2942 82346 2970
rect 53746 2930 53752 2942
rect 82668 2930 82674 2982
rect 82726 2970 82732 2982
rect 83775 2973 83833 2979
rect 83775 2970 83787 2973
rect 82726 2942 83787 2970
rect 82726 2930 82732 2942
rect 83775 2939 83787 2942
rect 83821 2939 83833 2973
rect 84232 2970 84238 2982
rect 84145 2942 84238 2970
rect 83775 2933 83833 2939
rect 84232 2930 84238 2942
rect 84290 2970 84296 2982
rect 85336 2970 85342 2982
rect 84290 2942 85342 2970
rect 84290 2930 84296 2942
rect 85336 2930 85342 2942
rect 85394 2930 85400 2982
rect 1711 2905 1769 2911
rect 1711 2871 1723 2905
rect 1757 2902 1769 2905
rect 1800 2902 1806 2914
rect 1757 2874 1806 2902
rect 1757 2871 1769 2874
rect 1711 2865 1769 2871
rect 1800 2862 1806 2874
rect 1858 2862 1864 2914
rect 2447 2905 2505 2911
rect 2447 2871 2459 2905
rect 2493 2902 2505 2905
rect 2996 2902 3002 2914
rect 2493 2874 3002 2902
rect 2493 2871 2505 2874
rect 2447 2865 2505 2871
rect 2996 2862 3002 2874
rect 3054 2862 3060 2914
rect 3183 2905 3241 2911
rect 3183 2871 3195 2905
rect 3229 2902 3241 2905
rect 4560 2902 4566 2914
rect 3229 2874 4566 2902
rect 3229 2871 3241 2874
rect 3183 2865 3241 2871
rect 4560 2862 4566 2874
rect 4618 2862 4624 2914
rect 4655 2905 4713 2911
rect 4655 2871 4667 2905
rect 4701 2902 4713 2905
rect 23972 2902 23978 2914
rect 4701 2874 23978 2902
rect 4701 2871 4713 2874
rect 4655 2865 4713 2871
rect 23972 2862 23978 2874
rect 24030 2862 24036 2914
rect 34828 2862 34834 2914
rect 34886 2902 34892 2914
rect 61603 2905 61661 2911
rect 61603 2902 61615 2905
rect 34886 2874 61615 2902
rect 34886 2862 34892 2874
rect 61603 2871 61615 2874
rect 61649 2871 61661 2905
rect 61603 2865 61661 2871
rect 61879 2905 61937 2911
rect 61879 2871 61891 2905
rect 61925 2902 61937 2905
rect 84784 2902 84790 2914
rect 61925 2874 84790 2902
rect 61925 2871 61937 2874
rect 61879 2865 61937 2871
rect 84784 2862 84790 2874
rect 84842 2862 84848 2914
rect 84968 2902 84974 2914
rect 84881 2874 84974 2902
rect 84968 2862 84974 2874
rect 85026 2902 85032 2914
rect 86624 2902 86630 2914
rect 85026 2874 86630 2902
rect 85026 2862 85032 2874
rect 86624 2862 86630 2874
rect 86682 2862 86688 2914
rect 2720 2794 2726 2846
rect 2778 2834 2784 2846
rect 2778 2806 2858 2834
rect 2778 2794 2784 2806
rect 607 2701 665 2707
rect 607 2667 619 2701
rect 653 2698 665 2701
rect 2079 2701 2137 2707
rect 653 2670 2030 2698
rect 653 2667 665 2670
rect 607 2661 665 2667
rect 972 2630 978 2642
rect 933 2602 978 2630
rect 972 2590 978 2602
rect 1030 2590 1036 2642
rect 2002 2630 2030 2670
rect 2079 2667 2091 2701
rect 2125 2698 2137 2701
rect 2720 2698 2726 2710
rect 2125 2670 2726 2698
rect 2125 2667 2137 2670
rect 2079 2661 2137 2667
rect 2720 2658 2726 2670
rect 2778 2658 2784 2710
rect 2830 2630 2858 2806
rect 3014 2766 3042 2862
rect 3551 2837 3609 2843
rect 3551 2803 3563 2837
rect 3597 2834 3609 2837
rect 4928 2834 4934 2846
rect 3597 2806 4934 2834
rect 3597 2803 3609 2806
rect 3551 2797 3609 2803
rect 4928 2794 4934 2806
rect 4986 2794 4992 2846
rect 5023 2837 5081 2843
rect 5023 2803 5035 2837
rect 5069 2834 5081 2837
rect 27468 2834 27474 2846
rect 5069 2806 27474 2834
rect 5069 2803 5081 2806
rect 5023 2797 5081 2803
rect 27468 2794 27474 2806
rect 27526 2794 27532 2846
rect 38784 2794 38790 2846
rect 38842 2834 38848 2846
rect 57463 2837 57521 2843
rect 57463 2834 57475 2837
rect 38842 2806 57475 2834
rect 38842 2794 38848 2806
rect 57463 2803 57475 2806
rect 57509 2803 57521 2837
rect 57463 2797 57521 2803
rect 61968 2794 61974 2846
rect 62026 2834 62032 2846
rect 85888 2834 85894 2846
rect 62026 2806 85894 2834
rect 62026 2794 62032 2806
rect 85888 2794 85894 2806
rect 85946 2794 85952 2846
rect 5575 2769 5633 2775
rect 5575 2766 5587 2769
rect 3014 2738 5587 2766
rect 5575 2735 5587 2738
rect 5621 2735 5633 2769
rect 5575 2729 5633 2735
rect 5759 2769 5817 2775
rect 5759 2735 5771 2769
rect 5805 2766 5817 2769
rect 22132 2766 22138 2778
rect 5805 2738 22138 2766
rect 5805 2735 5817 2738
rect 5759 2729 5817 2735
rect 22132 2726 22138 2738
rect 22190 2726 22196 2778
rect 37588 2726 37594 2778
rect 37646 2766 37652 2778
rect 61787 2769 61845 2775
rect 61787 2766 61799 2769
rect 37646 2738 61799 2766
rect 37646 2726 37652 2738
rect 61787 2735 61799 2738
rect 61833 2735 61845 2769
rect 61787 2729 61845 2735
rect 61879 2769 61937 2775
rect 61879 2735 61891 2769
rect 61925 2766 61937 2769
rect 84324 2766 84330 2778
rect 61925 2738 84330 2766
rect 61925 2735 61937 2738
rect 61879 2729 61937 2735
rect 84324 2726 84330 2738
rect 84382 2726 84388 2778
rect 84603 2769 84661 2775
rect 84603 2735 84615 2769
rect 84649 2766 84661 2769
rect 86532 2766 86538 2778
rect 84649 2738 86538 2766
rect 84649 2735 84661 2738
rect 84603 2729 84661 2735
rect 4011 2701 4069 2707
rect 4011 2667 4023 2701
rect 4057 2698 4069 2701
rect 19740 2698 19746 2710
rect 4057 2670 19746 2698
rect 4057 2667 4069 2670
rect 4011 2661 4069 2667
rect 19740 2658 19746 2670
rect 19798 2658 19804 2710
rect 41360 2658 41366 2710
rect 41418 2698 41424 2710
rect 81291 2701 81349 2707
rect 81291 2698 81303 2701
rect 41418 2670 81303 2698
rect 41418 2658 41424 2670
rect 81291 2667 81303 2670
rect 81337 2667 81349 2701
rect 81291 2661 81349 2667
rect 81380 2658 81386 2710
rect 81438 2698 81444 2710
rect 82392 2698 82398 2710
rect 81438 2670 82398 2698
rect 81438 2658 81444 2670
rect 82392 2658 82398 2670
rect 82450 2658 82456 2710
rect 84618 2698 84646 2729
rect 86532 2726 86538 2738
rect 86590 2726 86596 2778
rect 82502 2670 84646 2698
rect 5023 2633 5081 2639
rect 5023 2630 5035 2633
rect 2002 2602 5035 2630
rect 5023 2599 5035 2602
rect 5069 2599 5081 2633
rect 5023 2593 5081 2599
rect 19464 2590 19470 2642
rect 19522 2630 19528 2642
rect 24616 2630 24622 2642
rect 19522 2602 24622 2630
rect 19522 2590 19528 2602
rect 24616 2590 24622 2602
rect 24674 2590 24680 2642
rect 82502 2630 82530 2670
rect 57386 2602 64498 2630
rect 25076 2562 25082 2574
rect 38 2540 3902 2562
rect 38 2488 2916 2540
rect 2968 2488 2980 2540
rect 3032 2488 3044 2540
rect 3096 2488 3108 2540
rect 3160 2488 3902 2540
rect 38 2466 3902 2488
rect 3934 2534 25082 2562
rect 972 2386 978 2438
rect 1030 2426 1036 2438
rect 1432 2426 1438 2438
rect 1030 2398 1438 2426
rect 1030 2386 1036 2398
rect 1432 2386 1438 2398
rect 1490 2426 1496 2438
rect 3934 2426 3962 2534
rect 25076 2522 25082 2534
rect 25134 2522 25140 2574
rect 50468 2522 50474 2574
rect 50526 2562 50532 2574
rect 50526 2534 55482 2562
rect 50526 2522 50532 2534
rect 4100 2454 4106 2506
rect 4158 2494 4164 2506
rect 7872 2494 7878 2506
rect 4158 2466 7878 2494
rect 4158 2454 4164 2466
rect 7872 2454 7878 2466
rect 7930 2454 7936 2506
rect 25996 2454 26002 2506
rect 26054 2494 26060 2506
rect 28388 2494 28394 2506
rect 26054 2466 28394 2494
rect 26054 2454 26060 2466
rect 28388 2454 28394 2466
rect 28446 2454 28452 2506
rect 55454 2494 55482 2534
rect 57386 2494 57414 2602
rect 57463 2565 57521 2571
rect 57463 2531 57475 2565
rect 57509 2562 57521 2565
rect 61968 2562 61974 2574
rect 57509 2534 61974 2562
rect 57509 2531 57521 2534
rect 57463 2525 57521 2531
rect 61968 2522 61974 2534
rect 62026 2522 62032 2574
rect 55454 2466 57414 2494
rect 64470 2494 64498 2602
rect 80110 2602 82530 2630
rect 78715 2565 78773 2571
rect 78715 2531 78727 2565
rect 78761 2562 78773 2565
rect 80110 2562 80138 2602
rect 83496 2590 83502 2642
rect 83554 2630 83560 2642
rect 84968 2630 84974 2642
rect 83554 2602 84974 2630
rect 83554 2590 83560 2602
rect 84968 2590 84974 2602
rect 85026 2590 85032 2642
rect 78761 2534 80138 2562
rect 83298 2540 87806 2562
rect 78761 2531 78773 2534
rect 78715 2525 78773 2531
rect 69791 2497 69849 2503
rect 69791 2494 69803 2497
rect 64470 2466 69803 2494
rect 69791 2463 69803 2466
rect 69837 2463 69849 2497
rect 83298 2488 86916 2540
rect 86968 2488 86980 2540
rect 87032 2488 87044 2540
rect 87096 2488 87108 2540
rect 87160 2488 87806 2540
rect 83298 2466 87806 2488
rect 69791 2457 69849 2463
rect 1490 2398 3962 2426
rect 5575 2429 5633 2435
rect 1490 2386 1496 2398
rect 5575 2395 5587 2429
rect 5621 2426 5633 2429
rect 31056 2426 31062 2438
rect 5621 2398 31062 2426
rect 5621 2395 5633 2398
rect 5575 2389 5633 2395
rect 31056 2386 31062 2398
rect 31114 2386 31120 2438
rect 50192 2386 50198 2438
rect 50250 2426 50256 2438
rect 81380 2426 81386 2438
rect 50250 2398 81386 2426
rect 50250 2386 50256 2398
rect 81380 2386 81386 2398
rect 81438 2386 81444 2438
rect 3548 2318 3554 2370
rect 3606 2358 3612 2370
rect 84048 2358 84054 2370
rect 3606 2330 84054 2358
rect 3606 2318 3612 2330
rect 84048 2318 84054 2330
rect 84106 2318 84112 2370
rect 2815 2293 2873 2299
rect 2815 2259 2827 2293
rect 2861 2290 2873 2293
rect 4836 2290 4842 2302
rect 2861 2262 4842 2290
rect 2861 2259 2873 2262
rect 2815 2253 2873 2259
rect 4836 2250 4842 2262
rect 4894 2250 4900 2302
rect 5756 2250 5762 2302
rect 5814 2290 5820 2302
rect 83956 2290 83962 2302
rect 5814 2262 83962 2290
rect 5814 2250 5820 2262
rect 83956 2250 83962 2262
rect 84014 2250 84020 2302
rect 2628 2182 2634 2234
rect 2686 2222 2692 2234
rect 81288 2222 81294 2234
rect 2686 2194 81294 2222
rect 2686 2182 2692 2194
rect 81288 2182 81294 2194
rect 81346 2182 81352 2234
rect 83867 2225 83925 2231
rect 83867 2222 83879 2225
rect 82134 2194 83879 2222
rect 2168 2114 2174 2166
rect 2226 2154 2232 2166
rect 2447 2157 2505 2163
rect 2447 2154 2459 2157
rect 2226 2126 2459 2154
rect 2226 2114 2232 2126
rect 2447 2123 2459 2126
rect 2493 2154 2505 2157
rect 18268 2154 18274 2166
rect 2493 2126 18274 2154
rect 2493 2123 2505 2126
rect 2447 2117 2505 2123
rect 18268 2114 18274 2126
rect 18326 2114 18332 2166
rect 35012 2114 35018 2166
rect 35070 2154 35076 2166
rect 42464 2154 42470 2166
rect 35070 2126 42470 2154
rect 35070 2114 35076 2126
rect 42464 2114 42470 2126
rect 42522 2114 42528 2166
rect 69791 2157 69849 2163
rect 69791 2123 69803 2157
rect 69837 2154 69849 2157
rect 78715 2157 78773 2163
rect 78715 2154 78727 2157
rect 69837 2126 78727 2154
rect 69837 2123 69849 2126
rect 69791 2117 69849 2123
rect 78715 2123 78727 2126
rect 78761 2123 78773 2157
rect 78715 2117 78773 2123
rect 1708 2086 1714 2098
rect 1669 2058 1714 2086
rect 1708 2046 1714 2058
rect 1766 2046 1772 2098
rect 2079 2089 2137 2095
rect 2079 2055 2091 2089
rect 2125 2086 2137 2089
rect 2812 2086 2818 2098
rect 2125 2058 2818 2086
rect 2125 2055 2137 2058
rect 2079 2049 2137 2055
rect 2812 2046 2818 2058
rect 2870 2046 2876 2098
rect 3551 2089 3609 2095
rect 3551 2055 3563 2089
rect 3597 2086 3609 2089
rect 4652 2086 4658 2098
rect 3597 2058 4658 2086
rect 3597 2055 3609 2058
rect 3551 2049 3609 2055
rect 4652 2046 4658 2058
rect 4710 2046 4716 2098
rect 46696 2046 46702 2098
rect 46754 2086 46760 2098
rect 82134 2086 82162 2194
rect 83867 2191 83879 2194
rect 83913 2222 83925 2225
rect 85244 2222 85250 2234
rect 83913 2194 85250 2222
rect 83913 2191 83925 2194
rect 83867 2185 83925 2191
rect 85244 2182 85250 2194
rect 85302 2182 85308 2234
rect 83496 2114 83502 2166
rect 83554 2154 83560 2166
rect 84143 2157 84201 2163
rect 84143 2154 84155 2157
rect 83554 2126 84155 2154
rect 83554 2114 83560 2126
rect 84143 2123 84155 2126
rect 84189 2123 84201 2157
rect 84143 2117 84201 2123
rect 46754 2058 82162 2086
rect 46754 2046 46760 2058
rect 38 1996 3902 2018
rect 38 1944 916 1996
rect 968 1944 980 1996
rect 1032 1944 1044 1996
rect 1096 1944 1108 1996
rect 1160 1944 3902 1996
rect 38 1922 3902 1944
rect 83298 1996 87806 2018
rect 83298 1944 84916 1996
rect 84968 1944 84980 1996
rect 85032 1944 85044 1996
rect 85096 1944 85108 1996
rect 85160 1944 87806 1996
rect 83298 1922 87806 1944
rect 1708 1842 1714 1894
rect 1766 1882 1772 1894
rect 26364 1882 26370 1894
rect 1766 1854 26370 1882
rect 1766 1842 1772 1854
rect 26364 1842 26370 1854
rect 26422 1842 26428 1894
rect 2812 1774 2818 1826
rect 2870 1814 2876 1826
rect 3824 1814 3830 1826
rect 2870 1786 3830 1814
rect 2870 1774 2876 1786
rect 3824 1774 3830 1786
rect 3882 1774 3888 1826
rect 47892 1774 47898 1826
rect 47950 1814 47956 1826
rect 84600 1814 84606 1826
rect 47950 1786 84606 1814
rect 47950 1774 47956 1786
rect 84600 1774 84606 1786
rect 84658 1774 84664 1826
rect 39980 1706 39986 1758
rect 40038 1746 40044 1758
rect 84692 1746 84698 1758
rect 40038 1718 84698 1746
rect 40038 1706 40044 1718
rect 84692 1706 84698 1718
rect 84750 1706 84756 1758
rect 54240 1570 54246 1622
rect 54298 1610 54304 1622
rect 83312 1610 83318 1622
rect 54298 1582 83318 1610
rect 54298 1570 54304 1582
rect 83312 1570 83318 1582
rect 83370 1570 83376 1622
rect 3916 1502 3922 1554
rect 3974 1542 3980 1554
rect 41820 1542 41826 1554
rect 3974 1514 41826 1542
rect 3974 1502 3980 1514
rect 41820 1502 41826 1514
rect 41878 1502 41884 1554
rect 49824 1502 49830 1554
rect 49882 1542 49888 1554
rect 81932 1542 81938 1554
rect 49882 1514 81938 1542
rect 49882 1502 49888 1514
rect 81932 1502 81938 1514
rect 81990 1502 81996 1554
rect 4652 1434 4658 1486
rect 4710 1474 4716 1486
rect 29216 1474 29222 1486
rect 4710 1446 29222 1474
rect 4710 1434 4716 1446
rect 29216 1434 29222 1446
rect 29274 1434 29280 1486
rect 51480 1434 51486 1486
rect 51538 1474 51544 1486
rect 83496 1474 83502 1486
rect 51538 1446 83502 1474
rect 51538 1434 51544 1446
rect 83496 1434 83502 1446
rect 83554 1434 83560 1486
rect 4836 1366 4842 1418
rect 4894 1406 4900 1418
rect 36300 1406 36306 1418
rect 4894 1378 36306 1406
rect 4894 1366 4900 1378
rect 36300 1366 36306 1378
rect 36358 1366 36364 1418
rect 45224 1366 45230 1418
rect 45282 1406 45288 1418
rect 81383 1409 81441 1415
rect 81383 1406 81395 1409
rect 45282 1378 81395 1406
rect 45282 1366 45288 1378
rect 81383 1375 81395 1378
rect 81429 1375 81441 1409
rect 81383 1369 81441 1375
rect 42280 1298 42286 1350
rect 42338 1338 42344 1350
rect 82116 1338 82122 1350
rect 42338 1310 82122 1338
rect 42338 1298 42344 1310
rect 82116 1298 82122 1310
rect 82174 1298 82180 1350
rect 24708 1230 24714 1282
rect 24766 1270 24772 1282
rect 82944 1270 82950 1282
rect 24766 1242 82950 1270
rect 24766 1230 24772 1242
rect 82944 1230 82950 1242
rect 83002 1230 83008 1282
rect 3824 1162 3830 1214
rect 3882 1202 3888 1214
rect 20844 1202 20850 1214
rect 3882 1174 20850 1202
rect 3882 1162 3888 1174
rect 20844 1162 20850 1174
rect 20902 1162 20908 1214
rect 22408 1162 22414 1214
rect 22466 1202 22472 1214
rect 82852 1202 82858 1214
rect 22466 1174 82858 1202
rect 22466 1162 22472 1174
rect 82852 1162 82858 1174
rect 82910 1162 82916 1214
rect 18912 1094 18918 1146
rect 18970 1134 18976 1146
rect 81656 1134 81662 1146
rect 18970 1106 81662 1134
rect 18970 1094 18976 1106
rect 81656 1094 81662 1106
rect 81714 1094 81720 1146
rect 2260 1026 2266 1078
rect 2318 1066 2324 1078
rect 11828 1066 11834 1078
rect 2318 1038 11834 1066
rect 2318 1026 2324 1038
rect 11828 1026 11834 1038
rect 11886 1026 11892 1078
rect 28296 1026 28302 1078
rect 28354 1066 28360 1078
rect 33080 1066 33086 1078
rect 28354 1038 33086 1066
rect 28354 1026 28360 1038
rect 33080 1026 33086 1038
rect 33138 1026 33144 1078
rect 3640 958 3646 1010
rect 3698 998 3704 1010
rect 14404 998 14410 1010
rect 3698 970 14410 998
rect 3698 958 3704 970
rect 14404 958 14410 970
rect 14462 958 14468 1010
rect 29400 958 29406 1010
rect 29458 998 29464 1010
rect 37588 998 37594 1010
rect 29458 970 37594 998
rect 29458 958 29464 970
rect 37588 958 37594 970
rect 37646 958 37652 1010
rect 4928 890 4934 942
rect 4986 930 4992 942
rect 11736 930 11742 942
rect 4986 902 11742 930
rect 4986 890 4992 902
rect 11736 890 11742 902
rect 11794 890 11800 942
rect 21304 890 21310 942
rect 21362 930 21368 942
rect 83220 930 83226 942
rect 21362 902 83226 930
rect 21362 890 21368 902
rect 83220 890 83226 902
rect 83278 890 83284 942
rect 2536 822 2542 874
rect 2594 862 2600 874
rect 23420 862 23426 874
rect 2594 834 23426 862
rect 2594 822 2600 834
rect 23420 822 23426 834
rect 23478 822 23484 874
rect 24248 822 24254 874
rect 24306 862 24312 874
rect 83680 862 83686 874
rect 24306 834 83686 862
rect 24306 822 24312 834
rect 83680 822 83686 834
rect 83738 822 83744 874
rect 4560 754 4566 806
rect 4618 794 4624 806
rect 16980 794 16986 806
rect 4618 766 16986 794
rect 4618 754 4624 766
rect 16980 754 16986 766
rect 17038 754 17044 806
rect 31056 754 31062 806
rect 31114 794 31120 806
rect 83036 794 83042 806
rect 31114 766 83042 794
rect 31114 754 31120 766
rect 83036 754 83042 766
rect 83094 754 83100 806
rect 31884 686 31890 738
rect 31942 726 31948 738
rect 83128 726 83134 738
rect 31942 698 83134 726
rect 31942 686 31948 698
rect 83128 686 83134 698
rect 83186 686 83192 738
rect 2904 618 2910 670
rect 2962 658 2968 670
rect 29860 658 29866 670
rect 2962 630 29866 658
rect 2962 618 2968 630
rect 29860 618 29866 630
rect 29918 618 29924 670
rect 32896 618 32902 670
rect 32954 658 32960 670
rect 82300 658 82306 670
rect 32954 630 82306 658
rect 32954 618 32960 630
rect 82300 618 82306 630
rect 82358 618 82364 670
rect 18084 550 18090 602
rect 18142 590 18148 602
rect 18142 562 32574 590
rect 18142 550 18148 562
rect 3272 482 3278 534
rect 3330 522 3336 534
rect 32436 522 32442 534
rect 3330 494 32442 522
rect 3330 482 3336 494
rect 32436 482 32442 494
rect 32494 482 32500 534
rect 32546 522 32574 562
rect 34736 550 34742 602
rect 34794 590 34800 602
rect 82579 593 82637 599
rect 82579 590 82591 593
rect 34794 562 82591 590
rect 34794 550 34800 562
rect 82579 559 82591 562
rect 82625 559 82637 593
rect 82579 553 82637 559
rect 34828 522 34834 534
rect 32546 494 34834 522
rect 34828 482 34834 494
rect 34886 482 34892 534
rect 35288 482 35294 534
rect 35346 522 35352 534
rect 82024 522 82030 534
rect 35346 494 82030 522
rect 35346 482 35352 494
rect 82024 482 82030 494
rect 82082 482 82088 534
rect 11736 414 11742 466
rect 11794 454 11800 466
rect 83956 454 83962 466
rect 11794 426 83962 454
rect 11794 414 11800 426
rect 83956 414 83962 426
rect 84014 414 84020 466
rect 20752 346 20758 398
rect 20810 386 20816 398
rect 39980 386 39986 398
rect 20810 358 39986 386
rect 20810 346 20816 358
rect 39980 346 39986 358
rect 40038 346 40044 398
rect 40072 346 40078 398
rect 40130 386 40136 398
rect 82484 386 82490 398
rect 40130 358 82490 386
rect 40130 346 40136 358
rect 82484 346 82490 358
rect 82542 346 82548 398
rect 5296 278 5302 330
rect 5354 318 5360 330
rect 38048 318 38054 330
rect 5354 290 38054 318
rect 5354 278 5360 290
rect 38048 278 38054 290
rect 38106 278 38112 330
rect 38324 278 38330 330
rect 38382 318 38388 330
rect 81840 318 81846 330
rect 38382 290 81846 318
rect 38382 278 38388 290
rect 81840 278 81846 290
rect 81898 278 81904 330
rect 43936 210 43942 262
rect 43994 250 44000 262
rect 81564 250 81570 262
rect 43994 222 81570 250
rect 43994 210 44000 222
rect 81564 210 81570 222
rect 81622 210 81628 262
rect 46144 142 46150 194
rect 46202 182 46208 194
rect 83404 182 83410 194
rect 46202 154 83410 182
rect 46202 142 46208 154
rect 83404 142 83410 154
rect 83462 142 83468 194
rect 4284 74 4290 126
rect 4342 114 4348 126
rect 84416 114 84422 126
rect 4342 86 84422 114
rect 4342 74 4348 86
rect 84416 74 84422 86
rect 84474 74 84480 126
rect 8700 6 8706 58
rect 8758 46 8764 58
rect 85520 46 85526 58
rect 8758 18 85526 46
rect 8758 6 8764 18
rect 85520 6 85526 18
rect 85578 6 85584 58
<< via1 >>
rect 5854 188502 5906 188554
rect 82490 188502 82542 188554
rect 5210 188434 5262 188486
rect 84330 188434 84382 188486
rect 5302 188366 5354 188418
rect 85158 188366 85210 188418
rect 2634 188298 2686 188350
rect 82122 188298 82174 188350
rect 2358 188230 2410 188282
rect 81846 188230 81898 188282
rect 2818 188162 2870 188214
rect 82398 188162 82450 188214
rect 2082 188094 2134 188146
rect 81938 188094 81990 188146
rect 2726 188026 2778 188078
rect 82582 188026 82634 188078
rect 82214 187958 82266 188010
rect 2450 187890 2502 187942
rect 83226 187890 83278 187942
rect 1346 187822 1398 187874
rect 82306 187822 82358 187874
rect 4750 187550 4802 187602
rect 2916 187448 2968 187500
rect 2980 187448 3032 187500
rect 3044 187448 3096 187500
rect 3108 187448 3160 187500
rect 86916 187448 86968 187500
rect 86980 187448 87032 187500
rect 87044 187448 87096 187500
rect 87108 187448 87160 187500
rect 5118 187346 5170 187398
rect 84790 187346 84842 187398
rect 4566 187278 4618 187330
rect 82030 187278 82082 187330
rect 5762 187210 5814 187262
rect 84054 187210 84106 187262
rect 4474 187142 4526 187194
rect 83318 187142 83370 187194
rect 4934 187074 4986 187126
rect 84422 187074 84474 187126
rect 4198 187006 4250 187058
rect 84330 187006 84382 187058
rect 916 186904 968 186956
rect 980 186904 1032 186956
rect 1044 186904 1096 186956
rect 1108 186904 1160 186956
rect 84916 186904 84968 186956
rect 84980 186904 85032 186956
rect 85044 186904 85096 186956
rect 85108 186904 85160 186956
rect 4658 186802 4710 186854
rect 84698 186802 84750 186854
rect 4106 186734 4158 186786
rect 84146 186734 84198 186786
rect 4842 186666 4894 186718
rect 85158 186666 85210 186718
rect 3370 186598 3422 186650
rect 84514 186598 84566 186650
rect 1990 186530 2042 186582
rect 83962 186530 84014 186582
rect 2916 186360 2968 186412
rect 2980 186360 3032 186412
rect 3044 186360 3096 186412
rect 3108 186360 3160 186412
rect 86916 186360 86968 186412
rect 86980 186360 87032 186412
rect 87044 186360 87096 186412
rect 87108 186360 87160 186412
rect 916 185816 968 185868
rect 980 185816 1032 185868
rect 1044 185816 1096 185868
rect 1108 185816 1160 185868
rect 84916 185816 84968 185868
rect 84980 185816 85032 185868
rect 85044 185816 85096 185868
rect 85108 185816 85160 185868
rect 84330 185374 84382 185426
rect 84790 185374 84842 185426
rect 2916 185272 2968 185324
rect 2980 185272 3032 185324
rect 3044 185272 3096 185324
rect 3108 185272 3160 185324
rect 86916 185272 86968 185324
rect 86980 185272 87032 185324
rect 87044 185272 87096 185324
rect 87108 185272 87160 185324
rect 916 184728 968 184780
rect 980 184728 1032 184780
rect 1044 184728 1096 184780
rect 1108 184728 1160 184780
rect 84916 184728 84968 184780
rect 84980 184728 85032 184780
rect 85044 184728 85096 184780
rect 85108 184728 85160 184780
rect 2916 184184 2968 184236
rect 2980 184184 3032 184236
rect 3044 184184 3096 184236
rect 3108 184184 3160 184236
rect 86916 184184 86968 184236
rect 86980 184184 87032 184236
rect 87044 184184 87096 184236
rect 87108 184184 87160 184236
rect 916 183640 968 183692
rect 980 183640 1032 183692
rect 1044 183640 1096 183692
rect 1108 183640 1160 183692
rect 84916 183640 84968 183692
rect 84980 183640 85032 183692
rect 85044 183640 85096 183692
rect 85108 183640 85160 183692
rect 2916 183096 2968 183148
rect 2980 183096 3032 183148
rect 3044 183096 3096 183148
rect 3108 183096 3160 183148
rect 86916 183096 86968 183148
rect 86980 183096 87032 183148
rect 87044 183096 87096 183148
rect 87108 183096 87160 183148
rect 3922 182722 3974 182774
rect 916 182552 968 182604
rect 980 182552 1032 182604
rect 1044 182552 1096 182604
rect 1108 182552 1160 182604
rect 84916 182552 84968 182604
rect 84980 182552 85032 182604
rect 85044 182552 85096 182604
rect 85108 182552 85160 182604
rect 84238 182246 84290 182298
rect 84422 182246 84474 182298
rect 84422 182110 84474 182162
rect 84606 182110 84658 182162
rect 2916 182008 2968 182060
rect 2980 182008 3032 182060
rect 3044 182008 3096 182060
rect 3108 182008 3160 182060
rect 86916 182008 86968 182060
rect 86980 182008 87032 182060
rect 87044 182008 87096 182060
rect 87108 182008 87160 182060
rect 3554 181677 3606 181686
rect 3554 181643 3563 181677
rect 3563 181643 3597 181677
rect 3597 181643 3606 181677
rect 3554 181634 3606 181643
rect 916 181464 968 181516
rect 980 181464 1032 181516
rect 1044 181464 1096 181516
rect 1108 181464 1160 181516
rect 84916 181464 84968 181516
rect 84980 181464 85032 181516
rect 85044 181464 85096 181516
rect 85108 181464 85160 181516
rect 2916 180920 2968 180972
rect 2980 180920 3032 180972
rect 3044 180920 3096 180972
rect 3108 180920 3160 180972
rect 86916 180920 86968 180972
rect 86980 180920 87032 180972
rect 87044 180920 87096 180972
rect 87108 180920 87160 180972
rect 916 180376 968 180428
rect 980 180376 1032 180428
rect 1044 180376 1096 180428
rect 1108 180376 1160 180428
rect 84916 180376 84968 180428
rect 84980 180376 85032 180428
rect 85044 180376 85096 180428
rect 85108 180376 85160 180428
rect 2174 180138 2226 180190
rect 3554 180181 3606 180190
rect 3554 180147 3563 180181
rect 3563 180147 3597 180181
rect 3597 180147 3606 180181
rect 3554 180138 3606 180147
rect 84330 180138 84382 180190
rect 2916 179832 2968 179884
rect 2980 179832 3032 179884
rect 3044 179832 3096 179884
rect 3108 179832 3160 179884
rect 86916 179832 86968 179884
rect 86980 179832 87032 179884
rect 87044 179832 87096 179884
rect 87108 179832 87160 179884
rect 916 179288 968 179340
rect 980 179288 1032 179340
rect 1044 179288 1096 179340
rect 1108 179288 1160 179340
rect 84916 179288 84968 179340
rect 84980 179288 85032 179340
rect 85044 179288 85096 179340
rect 85108 179288 85160 179340
rect 4014 178846 4066 178898
rect 2916 178744 2968 178796
rect 2980 178744 3032 178796
rect 3044 178744 3096 178796
rect 3108 178744 3160 178796
rect 86916 178744 86968 178796
rect 86980 178744 87032 178796
rect 87044 178744 87096 178796
rect 87108 178744 87160 178796
rect 84698 178506 84750 178558
rect 84698 178302 84750 178354
rect 916 178200 968 178252
rect 980 178200 1032 178252
rect 1044 178200 1096 178252
rect 1108 178200 1160 178252
rect 84916 178200 84968 178252
rect 84980 178200 85032 178252
rect 85044 178200 85096 178252
rect 85108 178200 85160 178252
rect 2916 177656 2968 177708
rect 2980 177656 3032 177708
rect 3044 177656 3096 177708
rect 3108 177656 3160 177708
rect 86916 177656 86968 177708
rect 86980 177656 87032 177708
rect 87044 177656 87096 177708
rect 87108 177656 87160 177708
rect 916 177112 968 177164
rect 980 177112 1032 177164
rect 1044 177112 1096 177164
rect 1108 177112 1160 177164
rect 84916 177112 84968 177164
rect 84980 177112 85032 177164
rect 85044 177112 85096 177164
rect 85108 177112 85160 177164
rect 3646 176670 3698 176722
rect 2916 176568 2968 176620
rect 2980 176568 3032 176620
rect 3044 176568 3096 176620
rect 3108 176568 3160 176620
rect 86916 176568 86968 176620
rect 86980 176568 87032 176620
rect 87044 176568 87096 176620
rect 87108 176568 87160 176620
rect 916 176024 968 176076
rect 980 176024 1032 176076
rect 1044 176024 1096 176076
rect 1108 176024 1160 176076
rect 84916 176024 84968 176076
rect 84980 176024 85032 176076
rect 85044 176024 85096 176076
rect 85108 176024 85160 176076
rect 3278 175582 3330 175634
rect 84606 175582 84658 175634
rect 84790 175582 84842 175634
rect 2916 175480 2968 175532
rect 2980 175480 3032 175532
rect 3044 175480 3096 175532
rect 3108 175480 3160 175532
rect 86916 175480 86968 175532
rect 86980 175480 87032 175532
rect 87044 175480 87096 175532
rect 87108 175480 87160 175532
rect 916 174936 968 174988
rect 980 174936 1032 174988
rect 1044 174936 1096 174988
rect 1108 174936 1160 174988
rect 84916 174936 84968 174988
rect 84980 174936 85032 174988
rect 85044 174936 85096 174988
rect 85108 174936 85160 174988
rect 2916 174392 2968 174444
rect 2980 174392 3032 174444
rect 3044 174392 3096 174444
rect 3108 174392 3160 174444
rect 86916 174392 86968 174444
rect 86980 174392 87032 174444
rect 87044 174392 87096 174444
rect 87108 174392 87160 174444
rect 3646 174154 3698 174206
rect 3646 173950 3698 174002
rect 916 173848 968 173900
rect 980 173848 1032 173900
rect 1044 173848 1096 173900
rect 1108 173848 1160 173900
rect 84916 173848 84968 173900
rect 84980 173848 85032 173900
rect 85044 173848 85096 173900
rect 85108 173848 85160 173900
rect 2174 173610 2226 173662
rect 3462 173610 3514 173662
rect 84330 173610 84382 173662
rect 84790 173610 84842 173662
rect 2266 173542 2318 173594
rect 2916 173304 2968 173356
rect 2980 173304 3032 173356
rect 3044 173304 3096 173356
rect 3108 173304 3160 173356
rect 86916 173304 86968 173356
rect 86980 173304 87032 173356
rect 87044 173304 87096 173356
rect 87108 173304 87160 173356
rect 916 172760 968 172812
rect 980 172760 1032 172812
rect 1044 172760 1096 172812
rect 1108 172760 1160 172812
rect 84916 172760 84968 172812
rect 84980 172760 85032 172812
rect 85044 172760 85096 172812
rect 85108 172760 85160 172812
rect 2916 172216 2968 172268
rect 2980 172216 3032 172268
rect 3044 172216 3096 172268
rect 3108 172216 3160 172268
rect 86916 172216 86968 172268
rect 86980 172216 87032 172268
rect 87044 172216 87096 172268
rect 87108 172216 87160 172268
rect 916 171672 968 171724
rect 980 171672 1032 171724
rect 1044 171672 1096 171724
rect 1108 171672 1160 171724
rect 84916 171672 84968 171724
rect 84980 171672 85032 171724
rect 85044 171672 85096 171724
rect 85108 171672 85160 171724
rect 2916 171128 2968 171180
rect 2980 171128 3032 171180
rect 3044 171128 3096 171180
rect 3108 171128 3160 171180
rect 86916 171128 86968 171180
rect 86980 171128 87032 171180
rect 87044 171128 87096 171180
rect 87108 171128 87160 171180
rect 84330 171026 84382 171078
rect 84790 171026 84842 171078
rect 916 170584 968 170636
rect 980 170584 1032 170636
rect 1044 170584 1096 170636
rect 1108 170584 1160 170636
rect 84916 170584 84968 170636
rect 84980 170584 85032 170636
rect 85044 170584 85096 170636
rect 85108 170584 85160 170636
rect 2916 170040 2968 170092
rect 2980 170040 3032 170092
rect 3044 170040 3096 170092
rect 3108 170040 3160 170092
rect 86916 170040 86968 170092
rect 86980 170040 87032 170092
rect 87044 170040 87096 170092
rect 87108 170040 87160 170092
rect 916 169496 968 169548
rect 980 169496 1032 169548
rect 1044 169496 1096 169548
rect 1108 169496 1160 169548
rect 84916 169496 84968 169548
rect 84980 169496 85032 169548
rect 85044 169496 85096 169548
rect 85108 169496 85160 169548
rect 2916 168952 2968 169004
rect 2980 168952 3032 169004
rect 3044 168952 3096 169004
rect 3108 168952 3160 169004
rect 86916 168952 86968 169004
rect 86980 168952 87032 169004
rect 87044 168952 87096 169004
rect 87108 168952 87160 169004
rect 916 168408 968 168460
rect 980 168408 1032 168460
rect 1044 168408 1096 168460
rect 1108 168408 1160 168460
rect 84916 168408 84968 168460
rect 84980 168408 85032 168460
rect 85044 168408 85096 168460
rect 85108 168408 85160 168460
rect 2916 167864 2968 167916
rect 2980 167864 3032 167916
rect 3044 167864 3096 167916
rect 3108 167864 3160 167916
rect 86916 167864 86968 167916
rect 86980 167864 87032 167916
rect 87044 167864 87096 167916
rect 87108 167864 87160 167916
rect 916 167320 968 167372
rect 980 167320 1032 167372
rect 1044 167320 1096 167372
rect 1108 167320 1160 167372
rect 84916 167320 84968 167372
rect 84980 167320 85032 167372
rect 85044 167320 85096 167372
rect 85108 167320 85160 167372
rect 2916 166776 2968 166828
rect 2980 166776 3032 166828
rect 3044 166776 3096 166828
rect 3108 166776 3160 166828
rect 86916 166776 86968 166828
rect 86980 166776 87032 166828
rect 87044 166776 87096 166828
rect 87108 166776 87160 166828
rect 916 166232 968 166284
rect 980 166232 1032 166284
rect 1044 166232 1096 166284
rect 1108 166232 1160 166284
rect 84916 166232 84968 166284
rect 84980 166232 85032 166284
rect 85044 166232 85096 166284
rect 85108 166232 85160 166284
rect 2916 165688 2968 165740
rect 2980 165688 3032 165740
rect 3044 165688 3096 165740
rect 3108 165688 3160 165740
rect 86916 165688 86968 165740
rect 86980 165688 87032 165740
rect 87044 165688 87096 165740
rect 87108 165688 87160 165740
rect 916 165144 968 165196
rect 980 165144 1032 165196
rect 1044 165144 1096 165196
rect 1108 165144 1160 165196
rect 84916 165144 84968 165196
rect 84980 165144 85032 165196
rect 85044 165144 85096 165196
rect 85108 165144 85160 165196
rect 83962 164838 84014 164890
rect 84422 164838 84474 164890
rect 84238 164770 84290 164822
rect 3738 164702 3790 164754
rect 84606 164702 84658 164754
rect 2916 164600 2968 164652
rect 2980 164600 3032 164652
rect 3044 164600 3096 164652
rect 3108 164600 3160 164652
rect 86916 164600 86968 164652
rect 86980 164600 87032 164652
rect 87044 164600 87096 164652
rect 87108 164600 87160 164652
rect 3738 164498 3790 164550
rect 83962 164498 84014 164550
rect 84238 164498 84290 164550
rect 84330 164498 84382 164550
rect 85158 164498 85210 164550
rect 916 164056 968 164108
rect 980 164056 1032 164108
rect 1044 164056 1096 164108
rect 1108 164056 1160 164108
rect 84916 164056 84968 164108
rect 84980 164056 85032 164108
rect 85044 164056 85096 164108
rect 85108 164056 85160 164108
rect 81754 163886 81806 163938
rect 85158 163886 85210 163938
rect 2916 163512 2968 163564
rect 2980 163512 3032 163564
rect 3044 163512 3096 163564
rect 3108 163512 3160 163564
rect 86916 163512 86968 163564
rect 86980 163512 87032 163564
rect 87044 163512 87096 163564
rect 87108 163512 87160 163564
rect 916 162968 968 163020
rect 980 162968 1032 163020
rect 1044 162968 1096 163020
rect 1108 162968 1160 163020
rect 84916 162968 84968 163020
rect 84980 162968 85032 163020
rect 85044 162968 85096 163020
rect 85108 162968 85160 163020
rect 81846 162798 81898 162850
rect 84330 162798 84382 162850
rect 2916 162424 2968 162476
rect 2980 162424 3032 162476
rect 3044 162424 3096 162476
rect 3108 162424 3160 162476
rect 86916 162424 86968 162476
rect 86980 162424 87032 162476
rect 87044 162424 87096 162476
rect 87108 162424 87160 162476
rect 1898 162118 1950 162170
rect 2266 162118 2318 162170
rect 1898 161982 1950 162034
rect 2266 161982 2318 162034
rect 916 161880 968 161932
rect 980 161880 1032 161932
rect 1044 161880 1096 161932
rect 1108 161880 1160 161932
rect 84916 161880 84968 161932
rect 84980 161880 85032 161932
rect 85044 161880 85096 161932
rect 85108 161880 85160 161932
rect 84330 161778 84382 161830
rect 84606 161778 84658 161830
rect 2916 161336 2968 161388
rect 2980 161336 3032 161388
rect 3044 161336 3096 161388
rect 3108 161336 3160 161388
rect 86916 161336 86968 161388
rect 86980 161336 87032 161388
rect 87044 161336 87096 161388
rect 87108 161336 87160 161388
rect 916 160792 968 160844
rect 980 160792 1032 160844
rect 1044 160792 1096 160844
rect 1108 160792 1160 160844
rect 84916 160792 84968 160844
rect 84980 160792 85032 160844
rect 85044 160792 85096 160844
rect 85108 160792 85160 160844
rect 82582 160690 82634 160742
rect 84606 160690 84658 160742
rect 84422 160622 84474 160674
rect 85342 160622 85394 160674
rect 2916 160248 2968 160300
rect 2980 160248 3032 160300
rect 3044 160248 3096 160300
rect 3108 160248 3160 160300
rect 86916 160248 86968 160300
rect 86980 160248 87032 160300
rect 87044 160248 87096 160300
rect 87108 160248 87160 160300
rect 84514 160146 84566 160198
rect 84514 159942 84566 159994
rect 916 159704 968 159756
rect 980 159704 1032 159756
rect 1044 159704 1096 159756
rect 1108 159704 1160 159756
rect 84916 159704 84968 159756
rect 84980 159704 85032 159756
rect 85044 159704 85096 159756
rect 85108 159704 85160 159756
rect 2916 159160 2968 159212
rect 2980 159160 3032 159212
rect 3044 159160 3096 159212
rect 3108 159160 3160 159212
rect 86916 159160 86968 159212
rect 86980 159160 87032 159212
rect 87044 159160 87096 159212
rect 87108 159160 87160 159212
rect 916 158616 968 158668
rect 980 158616 1032 158668
rect 1044 158616 1096 158668
rect 1108 158616 1160 158668
rect 84916 158616 84968 158668
rect 84980 158616 85032 158668
rect 85044 158616 85096 158668
rect 85108 158616 85160 158668
rect 2916 158072 2968 158124
rect 2980 158072 3032 158124
rect 3044 158072 3096 158124
rect 3108 158072 3160 158124
rect 86916 158072 86968 158124
rect 86980 158072 87032 158124
rect 87044 158072 87096 158124
rect 87108 158072 87160 158124
rect 916 157528 968 157580
rect 980 157528 1032 157580
rect 1044 157528 1096 157580
rect 1108 157528 1160 157580
rect 84916 157528 84968 157580
rect 84980 157528 85032 157580
rect 85044 157528 85096 157580
rect 85108 157528 85160 157580
rect 2916 156984 2968 157036
rect 2980 156984 3032 157036
rect 3044 156984 3096 157036
rect 3108 156984 3160 157036
rect 86916 156984 86968 157036
rect 86980 156984 87032 157036
rect 87044 156984 87096 157036
rect 87108 156984 87160 157036
rect 82490 156882 82542 156934
rect 85066 156882 85118 156934
rect 916 156440 968 156492
rect 980 156440 1032 156492
rect 1044 156440 1096 156492
rect 1108 156440 1160 156492
rect 84916 156440 84968 156492
rect 84980 156440 85032 156492
rect 85044 156440 85096 156492
rect 85108 156440 85160 156492
rect 2916 155896 2968 155948
rect 2980 155896 3032 155948
rect 3044 155896 3096 155948
rect 3108 155896 3160 155948
rect 86916 155896 86968 155948
rect 86980 155896 87032 155948
rect 87044 155896 87096 155948
rect 87108 155896 87160 155948
rect 3462 155658 3514 155710
rect 3554 155590 3606 155642
rect 3738 155590 3790 155642
rect 4014 155522 4066 155574
rect 3738 155454 3790 155506
rect 916 155352 968 155404
rect 980 155352 1032 155404
rect 1044 155352 1096 155404
rect 1108 155352 1160 155404
rect 4014 155361 4066 155370
rect 4014 155327 4023 155361
rect 4023 155327 4057 155361
rect 4057 155327 4066 155361
rect 4014 155318 4066 155327
rect 84916 155352 84968 155404
rect 84980 155352 85032 155404
rect 85044 155352 85096 155404
rect 85108 155352 85160 155404
rect 2916 154808 2968 154860
rect 2980 154808 3032 154860
rect 3044 154808 3096 154860
rect 3108 154808 3160 154860
rect 86916 154808 86968 154860
rect 86980 154808 87032 154860
rect 87044 154808 87096 154860
rect 87108 154808 87160 154860
rect 916 154264 968 154316
rect 980 154264 1032 154316
rect 1044 154264 1096 154316
rect 1108 154264 1160 154316
rect 84916 154264 84968 154316
rect 84980 154264 85032 154316
rect 85044 154264 85096 154316
rect 85108 154264 85160 154316
rect 2916 153720 2968 153772
rect 2980 153720 3032 153772
rect 3044 153720 3096 153772
rect 3108 153720 3160 153772
rect 86916 153720 86968 153772
rect 86980 153720 87032 153772
rect 87044 153720 87096 153772
rect 87108 153720 87160 153772
rect 916 153176 968 153228
rect 980 153176 1032 153228
rect 1044 153176 1096 153228
rect 1108 153176 1160 153228
rect 84916 153176 84968 153228
rect 84980 153176 85032 153228
rect 85044 153176 85096 153228
rect 85108 153176 85160 153228
rect 1898 153074 1950 153126
rect 2266 153074 2318 153126
rect 2916 152632 2968 152684
rect 2980 152632 3032 152684
rect 3044 152632 3096 152684
rect 3108 152632 3160 152684
rect 86916 152632 86968 152684
rect 86980 152632 87032 152684
rect 87044 152632 87096 152684
rect 87108 152632 87160 152684
rect 916 152088 968 152140
rect 980 152088 1032 152140
rect 1044 152088 1096 152140
rect 1108 152088 1160 152140
rect 84916 152088 84968 152140
rect 84980 152088 85032 152140
rect 85044 152088 85096 152140
rect 85108 152088 85160 152140
rect 3462 151782 3514 151834
rect 5578 151782 5630 151834
rect 2916 151544 2968 151596
rect 2980 151544 3032 151596
rect 3044 151544 3096 151596
rect 3108 151544 3160 151596
rect 86916 151544 86968 151596
rect 86980 151544 87032 151596
rect 87044 151544 87096 151596
rect 87108 151544 87160 151596
rect 916 151000 968 151052
rect 980 151000 1032 151052
rect 1044 151000 1096 151052
rect 1108 151000 1160 151052
rect 84916 151000 84968 151052
rect 84980 151000 85032 151052
rect 85044 151000 85096 151052
rect 85108 151000 85160 151052
rect 2916 150456 2968 150508
rect 2980 150456 3032 150508
rect 3044 150456 3096 150508
rect 3108 150456 3160 150508
rect 86916 150456 86968 150508
rect 86980 150456 87032 150508
rect 87044 150456 87096 150508
rect 87108 150456 87160 150508
rect 82398 150082 82450 150134
rect 83962 150082 84014 150134
rect 916 149912 968 149964
rect 980 149912 1032 149964
rect 1044 149912 1096 149964
rect 1108 149912 1160 149964
rect 84916 149912 84968 149964
rect 84980 149912 85032 149964
rect 85044 149912 85096 149964
rect 85108 149912 85160 149964
rect 2916 149368 2968 149420
rect 2980 149368 3032 149420
rect 3044 149368 3096 149420
rect 3108 149368 3160 149420
rect 86916 149368 86968 149420
rect 86980 149368 87032 149420
rect 87044 149368 87096 149420
rect 87108 149368 87160 149420
rect 82306 149130 82358 149182
rect 83962 149130 84014 149182
rect 916 148824 968 148876
rect 980 148824 1032 148876
rect 1044 148824 1096 148876
rect 1108 148824 1160 148876
rect 84916 148824 84968 148876
rect 84980 148824 85032 148876
rect 85044 148824 85096 148876
rect 85108 148824 85160 148876
rect 2916 148280 2968 148332
rect 2980 148280 3032 148332
rect 3044 148280 3096 148332
rect 3108 148280 3160 148332
rect 86916 148280 86968 148332
rect 86980 148280 87032 148332
rect 87044 148280 87096 148332
rect 87108 148280 87160 148332
rect 82214 147838 82266 147890
rect 83962 147838 84014 147890
rect 916 147736 968 147788
rect 980 147736 1032 147788
rect 1044 147736 1096 147788
rect 1108 147736 1160 147788
rect 84916 147736 84968 147788
rect 84980 147736 85032 147788
rect 85044 147736 85096 147788
rect 85108 147736 85160 147788
rect 2916 147192 2968 147244
rect 2980 147192 3032 147244
rect 3044 147192 3096 147244
rect 3108 147192 3160 147244
rect 86916 147192 86968 147244
rect 86980 147192 87032 147244
rect 87044 147192 87096 147244
rect 87108 147192 87160 147244
rect 4014 146861 4066 146870
rect 4014 146827 4023 146861
rect 4023 146827 4057 146861
rect 4057 146827 4066 146861
rect 4014 146818 4066 146827
rect 3554 146750 3606 146802
rect 916 146648 968 146700
rect 980 146648 1032 146700
rect 1044 146648 1096 146700
rect 1108 146648 1160 146700
rect 84916 146648 84968 146700
rect 84980 146648 85032 146700
rect 85044 146648 85096 146700
rect 85108 146648 85160 146700
rect 82122 146546 82174 146598
rect 83962 146546 84014 146598
rect 2916 146104 2968 146156
rect 2980 146104 3032 146156
rect 3044 146104 3096 146156
rect 3108 146104 3160 146156
rect 86916 146104 86968 146156
rect 86980 146104 87032 146156
rect 87044 146104 87096 146156
rect 87108 146104 87160 146156
rect 1898 145934 1950 145986
rect 2266 145934 2318 145986
rect 916 145560 968 145612
rect 980 145560 1032 145612
rect 1044 145560 1096 145612
rect 1108 145560 1160 145612
rect 84916 145560 84968 145612
rect 84980 145560 85032 145612
rect 85044 145560 85096 145612
rect 85108 145560 85160 145612
rect 81938 145254 81990 145306
rect 83962 145254 84014 145306
rect 2916 145016 2968 145068
rect 2980 145016 3032 145068
rect 3044 145016 3096 145068
rect 3108 145016 3160 145068
rect 86916 145016 86968 145068
rect 86980 145016 87032 145068
rect 87044 145016 87096 145068
rect 87108 145016 87160 145068
rect 916 144472 968 144524
rect 980 144472 1032 144524
rect 1044 144472 1096 144524
rect 1108 144472 1160 144524
rect 84916 144472 84968 144524
rect 84980 144472 85032 144524
rect 85044 144472 85096 144524
rect 85108 144472 85160 144524
rect 2916 143928 2968 143980
rect 2980 143928 3032 143980
rect 3044 143928 3096 143980
rect 3108 143928 3160 143980
rect 86916 143928 86968 143980
rect 86980 143928 87032 143980
rect 87044 143928 87096 143980
rect 87108 143928 87160 143980
rect 82030 143826 82082 143878
rect 84238 143826 84290 143878
rect 916 143384 968 143436
rect 980 143384 1032 143436
rect 1044 143384 1096 143436
rect 1108 143384 1160 143436
rect 84916 143384 84968 143436
rect 84980 143384 85032 143436
rect 85044 143384 85096 143436
rect 85108 143384 85160 143436
rect 2916 142840 2968 142892
rect 2980 142840 3032 142892
rect 3044 142840 3096 142892
rect 3108 142840 3160 142892
rect 86916 142840 86968 142892
rect 86980 142840 87032 142892
rect 87044 142840 87096 142892
rect 87108 142840 87160 142892
rect 916 142296 968 142348
rect 980 142296 1032 142348
rect 1044 142296 1096 142348
rect 1108 142296 1160 142348
rect 84916 142296 84968 142348
rect 84980 142296 85032 142348
rect 85044 142296 85096 142348
rect 85108 142296 85160 142348
rect 2916 141752 2968 141804
rect 2980 141752 3032 141804
rect 3044 141752 3096 141804
rect 3108 141752 3160 141804
rect 86916 141752 86968 141804
rect 86980 141752 87032 141804
rect 87044 141752 87096 141804
rect 87108 141752 87160 141804
rect 3738 141582 3790 141634
rect 1898 141514 1950 141566
rect 2174 141514 2226 141566
rect 3554 141514 3606 141566
rect 916 141208 968 141260
rect 980 141208 1032 141260
rect 1044 141208 1096 141260
rect 1108 141208 1160 141260
rect 84916 141208 84968 141260
rect 84980 141208 85032 141260
rect 85044 141208 85096 141260
rect 85108 141208 85160 141260
rect 2916 140664 2968 140716
rect 2980 140664 3032 140716
rect 3044 140664 3096 140716
rect 3108 140664 3160 140716
rect 86916 140664 86968 140716
rect 86980 140664 87032 140716
rect 87044 140664 87096 140716
rect 87108 140664 87160 140716
rect 916 140120 968 140172
rect 980 140120 1032 140172
rect 1044 140120 1096 140172
rect 1108 140120 1160 140172
rect 84916 140120 84968 140172
rect 84980 140120 85032 140172
rect 85044 140120 85096 140172
rect 85108 140120 85160 140172
rect 2916 139576 2968 139628
rect 2980 139576 3032 139628
rect 3044 139576 3096 139628
rect 3108 139576 3160 139628
rect 86916 139576 86968 139628
rect 86980 139576 87032 139628
rect 87044 139576 87096 139628
rect 87108 139576 87160 139628
rect 916 139032 968 139084
rect 980 139032 1032 139084
rect 1044 139032 1096 139084
rect 1108 139032 1160 139084
rect 84916 139032 84968 139084
rect 84980 139032 85032 139084
rect 85044 139032 85096 139084
rect 85108 139032 85160 139084
rect 2916 138488 2968 138540
rect 2980 138488 3032 138540
rect 3044 138488 3096 138540
rect 3108 138488 3160 138540
rect 86916 138488 86968 138540
rect 86980 138488 87032 138540
rect 87044 138488 87096 138540
rect 87108 138488 87160 138540
rect 916 137944 968 137996
rect 980 137944 1032 137996
rect 1044 137944 1096 137996
rect 1108 137944 1160 137996
rect 84916 137944 84968 137996
rect 84980 137944 85032 137996
rect 85044 137944 85096 137996
rect 85108 137944 85160 137996
rect 81938 137638 81990 137690
rect 84238 137638 84290 137690
rect 2916 137400 2968 137452
rect 2980 137400 3032 137452
rect 3044 137400 3096 137452
rect 3108 137400 3160 137452
rect 86916 137400 86968 137452
rect 86980 137400 87032 137452
rect 87044 137400 87096 137452
rect 87108 137400 87160 137452
rect 916 136856 968 136908
rect 980 136856 1032 136908
rect 1044 136856 1096 136908
rect 1108 136856 1160 136908
rect 84916 136856 84968 136908
rect 84980 136856 85032 136908
rect 85044 136856 85096 136908
rect 85108 136856 85160 136908
rect 2916 136312 2968 136364
rect 2980 136312 3032 136364
rect 3044 136312 3096 136364
rect 3108 136312 3160 136364
rect 86916 136312 86968 136364
rect 86980 136312 87032 136364
rect 87044 136312 87096 136364
rect 87108 136312 87160 136364
rect 916 135768 968 135820
rect 980 135768 1032 135820
rect 1044 135768 1096 135820
rect 1108 135768 1160 135820
rect 84916 135768 84968 135820
rect 84980 135768 85032 135820
rect 85044 135768 85096 135820
rect 85108 135768 85160 135820
rect 2916 135224 2968 135276
rect 2980 135224 3032 135276
rect 3044 135224 3096 135276
rect 3108 135224 3160 135276
rect 86916 135224 86968 135276
rect 86980 135224 87032 135276
rect 87044 135224 87096 135276
rect 87108 135224 87160 135276
rect 916 134680 968 134732
rect 980 134680 1032 134732
rect 1044 134680 1096 134732
rect 1108 134680 1160 134732
rect 84916 134680 84968 134732
rect 84980 134680 85032 134732
rect 85044 134680 85096 134732
rect 85108 134680 85160 134732
rect 2916 134136 2968 134188
rect 2980 134136 3032 134188
rect 3044 134136 3096 134188
rect 3108 134136 3160 134188
rect 86916 134136 86968 134188
rect 86980 134136 87032 134188
rect 87044 134136 87096 134188
rect 87108 134136 87160 134188
rect 1898 133694 1950 133746
rect 2266 133694 2318 133746
rect 916 133592 968 133644
rect 980 133592 1032 133644
rect 1044 133592 1096 133644
rect 1108 133592 1160 133644
rect 84916 133592 84968 133644
rect 84980 133592 85032 133644
rect 85044 133592 85096 133644
rect 85108 133592 85160 133644
rect 2916 133048 2968 133100
rect 2980 133048 3032 133100
rect 3044 133048 3096 133100
rect 3108 133048 3160 133100
rect 86916 133048 86968 133100
rect 86980 133048 87032 133100
rect 87044 133048 87096 133100
rect 87108 133048 87160 133100
rect 916 132504 968 132556
rect 980 132504 1032 132556
rect 1044 132504 1096 132556
rect 1108 132504 1160 132556
rect 84916 132504 84968 132556
rect 84980 132504 85032 132556
rect 85044 132504 85096 132556
rect 85108 132504 85160 132556
rect 2916 131960 2968 132012
rect 2980 131960 3032 132012
rect 3044 131960 3096 132012
rect 3108 131960 3160 132012
rect 86916 131960 86968 132012
rect 86980 131960 87032 132012
rect 87044 131960 87096 132012
rect 87108 131960 87160 132012
rect 916 131416 968 131468
rect 980 131416 1032 131468
rect 1044 131416 1096 131468
rect 1108 131416 1160 131468
rect 84916 131416 84968 131468
rect 84980 131416 85032 131468
rect 85044 131416 85096 131468
rect 85108 131416 85160 131468
rect 2916 130872 2968 130924
rect 2980 130872 3032 130924
rect 3044 130872 3096 130924
rect 3108 130872 3160 130924
rect 86916 130872 86968 130924
rect 86980 130872 87032 130924
rect 87044 130872 87096 130924
rect 87108 130872 87160 130924
rect 916 130328 968 130380
rect 980 130328 1032 130380
rect 1044 130328 1096 130380
rect 1108 130328 1160 130380
rect 84916 130328 84968 130380
rect 84980 130328 85032 130380
rect 85044 130328 85096 130380
rect 85108 130328 85160 130380
rect 83226 129886 83278 129938
rect 84514 129886 84566 129938
rect 2916 129784 2968 129836
rect 2980 129784 3032 129836
rect 3044 129784 3096 129836
rect 3108 129784 3160 129836
rect 86916 129784 86968 129836
rect 86980 129784 87032 129836
rect 87044 129784 87096 129836
rect 87108 129784 87160 129836
rect 916 129240 968 129292
rect 980 129240 1032 129292
rect 1044 129240 1096 129292
rect 1108 129240 1160 129292
rect 84916 129240 84968 129292
rect 84980 129240 85032 129292
rect 85044 129240 85096 129292
rect 85108 129240 85160 129292
rect 3554 128798 3606 128850
rect 2916 128696 2968 128748
rect 2980 128696 3032 128748
rect 3044 128696 3096 128748
rect 3108 128696 3160 128748
rect 86916 128696 86968 128748
rect 86980 128696 87032 128748
rect 87044 128696 87096 128748
rect 87108 128696 87160 128748
rect 3738 128594 3790 128646
rect 83134 128594 83186 128646
rect 84422 128594 84474 128646
rect 916 128152 968 128204
rect 980 128152 1032 128204
rect 1044 128152 1096 128204
rect 1108 128152 1160 128204
rect 84916 128152 84968 128204
rect 84980 128152 85032 128204
rect 85044 128152 85096 128204
rect 85108 128152 85160 128204
rect 2916 127608 2968 127660
rect 2980 127608 3032 127660
rect 3044 127608 3096 127660
rect 3108 127608 3160 127660
rect 86916 127608 86968 127660
rect 86980 127608 87032 127660
rect 87044 127608 87096 127660
rect 87108 127608 87160 127660
rect 83410 127370 83462 127422
rect 84238 127370 84290 127422
rect 916 127064 968 127116
rect 980 127064 1032 127116
rect 1044 127064 1096 127116
rect 1108 127064 1160 127116
rect 84916 127064 84968 127116
rect 84980 127064 85032 127116
rect 85044 127064 85096 127116
rect 85108 127064 85160 127116
rect 2916 126520 2968 126572
rect 2980 126520 3032 126572
rect 3044 126520 3096 126572
rect 3108 126520 3160 126572
rect 86916 126520 86968 126572
rect 86980 126520 87032 126572
rect 87044 126520 87096 126572
rect 87108 126520 87160 126572
rect 916 125976 968 126028
rect 980 125976 1032 126028
rect 1044 125976 1096 126028
rect 1108 125976 1160 126028
rect 84916 125976 84968 126028
rect 84980 125976 85032 126028
rect 85044 125976 85096 126028
rect 85108 125976 85160 126028
rect 2916 125432 2968 125484
rect 2980 125432 3032 125484
rect 3044 125432 3096 125484
rect 3108 125432 3160 125484
rect 86916 125432 86968 125484
rect 86980 125432 87032 125484
rect 87044 125432 87096 125484
rect 87108 125432 87160 125484
rect 916 124888 968 124940
rect 980 124888 1032 124940
rect 1044 124888 1096 124940
rect 1108 124888 1160 124940
rect 84916 124888 84968 124940
rect 84980 124888 85032 124940
rect 85044 124888 85096 124940
rect 85108 124888 85160 124940
rect 1898 124718 1950 124770
rect 2174 124718 2226 124770
rect 82030 124718 82082 124770
rect 84238 124718 84290 124770
rect 2916 124344 2968 124396
rect 2980 124344 3032 124396
rect 3044 124344 3096 124396
rect 3108 124344 3160 124396
rect 86916 124344 86968 124396
rect 86980 124344 87032 124396
rect 87044 124344 87096 124396
rect 87108 124344 87160 124396
rect 82122 123902 82174 123954
rect 84422 123902 84474 123954
rect 916 123800 968 123852
rect 980 123800 1032 123852
rect 1044 123800 1096 123852
rect 1108 123800 1160 123852
rect 84916 123800 84968 123852
rect 84980 123800 85032 123852
rect 85044 123800 85096 123852
rect 85108 123800 85160 123852
rect 3738 123494 3790 123546
rect 3554 123426 3606 123478
rect 2916 123256 2968 123308
rect 2980 123256 3032 123308
rect 3044 123256 3096 123308
rect 3108 123256 3160 123308
rect 86916 123256 86968 123308
rect 86980 123256 87032 123308
rect 87044 123256 87096 123308
rect 87108 123256 87160 123308
rect 916 122712 968 122764
rect 980 122712 1032 122764
rect 1044 122712 1096 122764
rect 1108 122712 1160 122764
rect 84916 122712 84968 122764
rect 84980 122712 85032 122764
rect 85044 122712 85096 122764
rect 85108 122712 85160 122764
rect 2916 122168 2968 122220
rect 2980 122168 3032 122220
rect 3044 122168 3096 122220
rect 3108 122168 3160 122220
rect 86916 122168 86968 122220
rect 86980 122168 87032 122220
rect 87044 122168 87096 122220
rect 87108 122168 87160 122220
rect 916 121624 968 121676
rect 980 121624 1032 121676
rect 1044 121624 1096 121676
rect 1108 121624 1160 121676
rect 84916 121624 84968 121676
rect 84980 121624 85032 121676
rect 85044 121624 85096 121676
rect 85108 121624 85160 121676
rect 2916 121080 2968 121132
rect 2980 121080 3032 121132
rect 3044 121080 3096 121132
rect 3108 121080 3160 121132
rect 86916 121080 86968 121132
rect 86980 121080 87032 121132
rect 87044 121080 87096 121132
rect 87108 121080 87160 121132
rect 83042 120842 83094 120894
rect 84330 120842 84382 120894
rect 916 120536 968 120588
rect 980 120536 1032 120588
rect 1044 120536 1096 120588
rect 1108 120536 1160 120588
rect 84916 120536 84968 120588
rect 84980 120536 85032 120588
rect 85044 120536 85096 120588
rect 85108 120536 85160 120588
rect 2916 119992 2968 120044
rect 2980 119992 3032 120044
rect 3044 119992 3096 120044
rect 3108 119992 3160 120044
rect 86916 119992 86968 120044
rect 86980 119992 87032 120044
rect 87044 119992 87096 120044
rect 87108 119992 87160 120044
rect 82214 119618 82266 119670
rect 84238 119618 84290 119670
rect 916 119448 968 119500
rect 980 119448 1032 119500
rect 1044 119448 1096 119500
rect 1108 119448 1160 119500
rect 84916 119448 84968 119500
rect 84980 119448 85032 119500
rect 85044 119448 85096 119500
rect 85108 119448 85160 119500
rect 82490 119346 82542 119398
rect 85342 119346 85394 119398
rect 2916 118904 2968 118956
rect 2980 118904 3032 118956
rect 3044 118904 3096 118956
rect 3108 118904 3160 118956
rect 86916 118904 86968 118956
rect 86980 118904 87032 118956
rect 87044 118904 87096 118956
rect 87108 118904 87160 118956
rect 916 118360 968 118412
rect 980 118360 1032 118412
rect 1044 118360 1096 118412
rect 1108 118360 1160 118412
rect 84916 118360 84968 118412
rect 84980 118360 85032 118412
rect 85044 118360 85096 118412
rect 85108 118360 85160 118412
rect 2916 117816 2968 117868
rect 2980 117816 3032 117868
rect 3044 117816 3096 117868
rect 3108 117816 3160 117868
rect 86916 117816 86968 117868
rect 86980 117816 87032 117868
rect 87044 117816 87096 117868
rect 87108 117816 87160 117868
rect 916 117272 968 117324
rect 980 117272 1032 117324
rect 1044 117272 1096 117324
rect 1108 117272 1160 117324
rect 84916 117272 84968 117324
rect 84980 117272 85032 117324
rect 85044 117272 85096 117324
rect 85108 117272 85160 117324
rect 2916 116728 2968 116780
rect 2980 116728 3032 116780
rect 3044 116728 3096 116780
rect 3108 116728 3160 116780
rect 86916 116728 86968 116780
rect 86980 116728 87032 116780
rect 87044 116728 87096 116780
rect 87108 116728 87160 116780
rect 82398 116626 82450 116678
rect 83962 116626 84014 116678
rect 4106 116422 4158 116474
rect 4290 116422 4342 116474
rect 916 116184 968 116236
rect 980 116184 1032 116236
rect 1044 116184 1096 116236
rect 1108 116184 1160 116236
rect 84916 116184 84968 116236
rect 84980 116184 85032 116236
rect 85044 116184 85096 116236
rect 85108 116184 85160 116236
rect 2916 115640 2968 115692
rect 2980 115640 3032 115692
rect 3044 115640 3096 115692
rect 3108 115640 3160 115692
rect 86916 115640 86968 115692
rect 86980 115640 87032 115692
rect 87044 115640 87096 115692
rect 87108 115640 87160 115692
rect 82950 115538 83002 115590
rect 84330 115538 84382 115590
rect 916 115096 968 115148
rect 980 115096 1032 115148
rect 1044 115096 1096 115148
rect 1108 115096 1160 115148
rect 84916 115096 84968 115148
rect 84980 115096 85032 115148
rect 85044 115096 85096 115148
rect 85108 115096 85160 115148
rect 3462 114858 3514 114910
rect 4290 114858 4342 114910
rect 3462 114765 3514 114774
rect 3462 114731 3471 114765
rect 3471 114731 3505 114765
rect 3505 114731 3514 114765
rect 3462 114722 3514 114731
rect 82306 114654 82358 114706
rect 84330 114654 84382 114706
rect 2916 114552 2968 114604
rect 2980 114552 3032 114604
rect 3044 114552 3096 114604
rect 3108 114552 3160 114604
rect 86916 114552 86968 114604
rect 86980 114552 87032 114604
rect 87044 114552 87096 114604
rect 87108 114552 87160 114604
rect 916 114008 968 114060
rect 980 114008 1032 114060
rect 1044 114008 1096 114060
rect 1108 114008 1160 114060
rect 84916 114008 84968 114060
rect 84980 114008 85032 114060
rect 85044 114008 85096 114060
rect 85108 114008 85160 114060
rect 2916 113464 2968 113516
rect 2980 113464 3032 113516
rect 3044 113464 3096 113516
rect 3108 113464 3160 113516
rect 86916 113464 86968 113516
rect 86980 113464 87032 113516
rect 87044 113464 87096 113516
rect 87108 113464 87160 113516
rect 916 112920 968 112972
rect 980 112920 1032 112972
rect 1044 112920 1096 112972
rect 1108 112920 1160 112972
rect 84916 112920 84968 112972
rect 84980 112920 85032 112972
rect 85044 112920 85096 112972
rect 85108 112920 85160 112972
rect 2916 112376 2968 112428
rect 2980 112376 3032 112428
rect 3044 112376 3096 112428
rect 3108 112376 3160 112428
rect 86916 112376 86968 112428
rect 86980 112376 87032 112428
rect 87044 112376 87096 112428
rect 87108 112376 87160 112428
rect 82490 112002 82542 112054
rect 84882 112002 84934 112054
rect 82858 111934 82910 111986
rect 83962 111934 84014 111986
rect 916 111832 968 111884
rect 980 111832 1032 111884
rect 1044 111832 1096 111884
rect 1108 111832 1160 111884
rect 84916 111832 84968 111884
rect 84980 111832 85032 111884
rect 85044 111832 85096 111884
rect 85108 111832 85160 111884
rect 2916 111288 2968 111340
rect 2980 111288 3032 111340
rect 3044 111288 3096 111340
rect 3108 111288 3160 111340
rect 86916 111288 86968 111340
rect 86980 111288 87032 111340
rect 87044 111288 87096 111340
rect 87108 111288 87160 111340
rect 916 110744 968 110796
rect 980 110744 1032 110796
rect 1044 110744 1096 110796
rect 1108 110744 1160 110796
rect 84916 110744 84968 110796
rect 84980 110744 85032 110796
rect 85044 110744 85096 110796
rect 85108 110744 85160 110796
rect 3554 110642 3606 110694
rect 3738 110574 3790 110626
rect 2916 110200 2968 110252
rect 2980 110200 3032 110252
rect 3044 110200 3096 110252
rect 3108 110200 3160 110252
rect 86916 110200 86968 110252
rect 86980 110200 87032 110252
rect 87044 110200 87096 110252
rect 87108 110200 87160 110252
rect 916 109656 968 109708
rect 980 109656 1032 109708
rect 1044 109656 1096 109708
rect 1108 109656 1160 109708
rect 84916 109656 84968 109708
rect 84980 109656 85032 109708
rect 85044 109656 85096 109708
rect 85108 109656 85160 109708
rect 81846 109282 81898 109334
rect 83962 109282 84014 109334
rect 2916 109112 2968 109164
rect 2980 109112 3032 109164
rect 3044 109112 3096 109164
rect 3108 109112 3160 109164
rect 86916 109112 86968 109164
rect 86980 109112 87032 109164
rect 87044 109112 87096 109164
rect 87108 109112 87160 109164
rect 916 108568 968 108620
rect 980 108568 1032 108620
rect 1044 108568 1096 108620
rect 1108 108568 1160 108620
rect 84916 108568 84968 108620
rect 84980 108568 85032 108620
rect 85044 108568 85096 108620
rect 85108 108568 85160 108620
rect 81662 108126 81714 108178
rect 83962 108126 84014 108178
rect 2916 108024 2968 108076
rect 2980 108024 3032 108076
rect 3044 108024 3096 108076
rect 3108 108024 3160 108076
rect 86916 108024 86968 108076
rect 86980 108024 87032 108076
rect 87044 108024 87096 108076
rect 87108 108024 87160 108076
rect 916 107480 968 107532
rect 980 107480 1032 107532
rect 1044 107480 1096 107532
rect 1108 107480 1160 107532
rect 84916 107480 84968 107532
rect 84980 107480 85032 107532
rect 85044 107480 85096 107532
rect 85108 107480 85160 107532
rect 2916 106936 2968 106988
rect 2980 106936 3032 106988
rect 3044 106936 3096 106988
rect 3108 106936 3160 106988
rect 86916 106936 86968 106988
rect 86980 106936 87032 106988
rect 87044 106936 87096 106988
rect 87108 106936 87160 106988
rect 82582 106562 82634 106614
rect 84238 106562 84290 106614
rect 916 106392 968 106444
rect 980 106392 1032 106444
rect 1044 106392 1096 106444
rect 1108 106392 1160 106444
rect 84916 106392 84968 106444
rect 84980 106392 85032 106444
rect 85044 106392 85096 106444
rect 85108 106392 85160 106444
rect 2916 105848 2968 105900
rect 2980 105848 3032 105900
rect 3044 105848 3096 105900
rect 3108 105848 3160 105900
rect 86916 105848 86968 105900
rect 86980 105848 87032 105900
rect 87044 105848 87096 105900
rect 87108 105848 87160 105900
rect 3738 105474 3790 105526
rect 3554 105406 3606 105458
rect 916 105304 968 105356
rect 980 105304 1032 105356
rect 1044 105304 1096 105356
rect 1108 105304 1160 105356
rect 84916 105304 84968 105356
rect 84980 105304 85032 105356
rect 85044 105304 85096 105356
rect 85108 105304 85160 105356
rect 2916 104760 2968 104812
rect 2980 104760 3032 104812
rect 3044 104760 3096 104812
rect 3108 104760 3160 104812
rect 86916 104760 86968 104812
rect 86980 104760 87032 104812
rect 87044 104760 87096 104812
rect 87108 104760 87160 104812
rect 916 104216 968 104268
rect 980 104216 1032 104268
rect 1044 104216 1096 104268
rect 1108 104216 1160 104268
rect 84916 104216 84968 104268
rect 84980 104216 85032 104268
rect 85044 104216 85096 104268
rect 85108 104216 85160 104268
rect 2916 103672 2968 103724
rect 2980 103672 3032 103724
rect 3044 103672 3096 103724
rect 3108 103672 3160 103724
rect 86916 103672 86968 103724
rect 86980 103672 87032 103724
rect 87044 103672 87096 103724
rect 87108 103672 87160 103724
rect 84790 103434 84842 103486
rect 85250 103434 85302 103486
rect 916 103128 968 103180
rect 980 103128 1032 103180
rect 1044 103128 1096 103180
rect 1108 103128 1160 103180
rect 84916 103128 84968 103180
rect 84980 103128 85032 103180
rect 85044 103128 85096 103180
rect 85108 103128 85160 103180
rect 82766 102822 82818 102874
rect 84514 102822 84566 102874
rect 84054 102686 84106 102738
rect 84514 102686 84566 102738
rect 2916 102584 2968 102636
rect 2980 102584 3032 102636
rect 3044 102584 3096 102636
rect 3108 102584 3160 102636
rect 86916 102584 86968 102636
rect 86980 102584 87032 102636
rect 87044 102584 87096 102636
rect 87108 102584 87160 102636
rect 916 102040 968 102092
rect 980 102040 1032 102092
rect 1044 102040 1096 102092
rect 1108 102040 1160 102092
rect 84916 102040 84968 102092
rect 84980 102040 85032 102092
rect 85044 102040 85096 102092
rect 85108 102040 85160 102092
rect 81754 101598 81806 101650
rect 84330 101598 84382 101650
rect 2916 101496 2968 101548
rect 2980 101496 3032 101548
rect 3044 101496 3096 101548
rect 3108 101496 3160 101548
rect 86916 101496 86968 101548
rect 86980 101496 87032 101548
rect 87044 101496 87096 101548
rect 87108 101496 87160 101548
rect 916 100952 968 101004
rect 980 100952 1032 101004
rect 1044 100952 1096 101004
rect 1108 100952 1160 101004
rect 84916 100952 84968 101004
rect 84980 100952 85032 101004
rect 85044 100952 85096 101004
rect 85108 100952 85160 101004
rect 84054 100510 84106 100562
rect 84330 100510 84382 100562
rect 2916 100408 2968 100460
rect 2980 100408 3032 100460
rect 3044 100408 3096 100460
rect 3108 100408 3160 100460
rect 86916 100408 86968 100460
rect 86980 100408 87032 100460
rect 87044 100408 87096 100460
rect 87108 100408 87160 100460
rect 84054 100306 84106 100358
rect 84698 100306 84750 100358
rect 916 99864 968 99916
rect 980 99864 1032 99916
rect 1044 99864 1096 99916
rect 1108 99864 1160 99916
rect 84916 99864 84968 99916
rect 84980 99864 85032 99916
rect 85044 99864 85096 99916
rect 85108 99864 85160 99916
rect 2916 99320 2968 99372
rect 2980 99320 3032 99372
rect 3044 99320 3096 99372
rect 3108 99320 3160 99372
rect 86916 99320 86968 99372
rect 86980 99320 87032 99372
rect 87044 99320 87096 99372
rect 87108 99320 87160 99372
rect 4566 99082 4618 99134
rect 4382 98946 4434 98998
rect 4750 98946 4802 98998
rect 85250 98946 85302 98998
rect 86538 98878 86590 98930
rect 916 98776 968 98828
rect 980 98776 1032 98828
rect 1044 98776 1096 98828
rect 1108 98776 1160 98828
rect 84916 98776 84968 98828
rect 84980 98776 85032 98828
rect 85044 98776 85096 98828
rect 85108 98776 85160 98828
rect 4658 98674 4710 98726
rect 4934 98674 4986 98726
rect 1898 98334 1950 98386
rect 2818 98334 2870 98386
rect 4106 98334 4158 98386
rect 2916 98232 2968 98284
rect 2980 98232 3032 98284
rect 3044 98232 3096 98284
rect 3108 98232 3160 98284
rect 86916 98232 86968 98284
rect 86980 98232 87032 98284
rect 87044 98232 87096 98284
rect 87108 98232 87160 98284
rect 4106 98130 4158 98182
rect 5118 98130 5170 98182
rect 82674 98130 82726 98182
rect 83870 98173 83922 98182
rect 83870 98139 83879 98173
rect 83879 98139 83913 98173
rect 83913 98139 83922 98173
rect 83870 98130 83922 98139
rect 84330 97994 84382 98046
rect 85158 97994 85210 98046
rect 2266 97790 2318 97842
rect 2450 97790 2502 97842
rect 916 97688 968 97740
rect 980 97688 1032 97740
rect 1044 97688 1096 97740
rect 1108 97688 1160 97740
rect 84916 97688 84968 97740
rect 84980 97688 85032 97740
rect 85044 97688 85096 97740
rect 85108 97688 85160 97740
rect 2818 97629 2870 97638
rect 2818 97595 2827 97629
rect 2827 97595 2861 97629
rect 2861 97595 2870 97629
rect 2818 97586 2870 97595
rect 3370 97586 3422 97638
rect 4382 97586 4434 97638
rect 83962 97586 84014 97638
rect 2082 97518 2134 97570
rect 83778 97561 83830 97570
rect 83778 97527 83787 97561
rect 83787 97527 83821 97561
rect 83821 97527 83830 97561
rect 83778 97518 83830 97527
rect 4106 97450 4158 97502
rect 81478 97450 81530 97502
rect 84514 97586 84566 97638
rect 2818 97382 2870 97434
rect 3922 97382 3974 97434
rect 86078 97382 86130 97434
rect 1346 97314 1398 97366
rect 83134 97314 83186 97366
rect 2082 97289 2134 97298
rect 2082 97255 2091 97289
rect 2091 97255 2125 97289
rect 2125 97255 2134 97289
rect 2082 97246 2134 97255
rect 2358 97246 2410 97298
rect 2542 97246 2594 97298
rect 3370 97246 3422 97298
rect 81294 97246 81346 97298
rect 85802 97314 85854 97366
rect 2916 97144 2968 97196
rect 2980 97144 3032 97196
rect 3044 97144 3096 97196
rect 3108 97144 3160 97196
rect 1346 97017 1398 97026
rect 1346 96983 1355 97017
rect 1355 96983 1389 97017
rect 1389 96983 1398 97017
rect 1346 96974 1398 96983
rect 3738 97042 3790 97094
rect 3922 97042 3974 97094
rect 4474 97042 4526 97094
rect 22138 97042 22190 97094
rect 45322 97042 45374 97094
rect 4106 96974 4158 97026
rect 5302 96974 5354 97026
rect 14594 96974 14646 97026
rect 28486 96974 28538 97026
rect 5210 96906 5262 96958
rect 83042 97110 83094 97162
rect 86916 97144 86968 97196
rect 86980 97144 87032 97196
rect 87044 97144 87096 97196
rect 87108 97144 87160 97196
rect 56638 96974 56690 97026
rect 81386 97042 81438 97094
rect 82950 97042 83002 97094
rect 84146 97085 84198 97094
rect 84146 97051 84155 97085
rect 84155 97051 84189 97085
rect 84189 97051 84198 97085
rect 84146 97042 84198 97051
rect 60870 96974 60922 97026
rect 80282 96906 80334 96958
rect 82858 96906 82910 96958
rect 4566 96838 4618 96890
rect 1714 96745 1766 96754
rect 1714 96711 1723 96745
rect 1723 96711 1757 96745
rect 1757 96711 1766 96745
rect 1714 96702 1766 96711
rect 3002 96702 3054 96754
rect 4934 96702 4986 96754
rect 50198 96838 50250 96890
rect 80190 96838 80242 96890
rect 83594 96838 83646 96890
rect 83778 96881 83830 96890
rect 83778 96847 83787 96881
rect 83787 96847 83821 96881
rect 83821 96847 83830 96881
rect 83778 96838 83830 96847
rect 84514 96838 84566 96890
rect 84790 96838 84842 96890
rect 25266 96770 25318 96822
rect 51670 96770 51722 96822
rect 5854 96702 5906 96754
rect 916 96600 968 96652
rect 980 96600 1032 96652
rect 1044 96600 1096 96652
rect 1108 96600 1160 96652
rect 4566 96634 4618 96686
rect 28946 96634 28998 96686
rect 34926 96634 34978 96686
rect 37042 96634 37094 96686
rect 48910 96634 48962 96686
rect 4382 96566 4434 96618
rect 29958 96566 30010 96618
rect 80098 96702 80150 96754
rect 84238 96770 84290 96822
rect 86538 96770 86590 96822
rect 85342 96702 85394 96754
rect 86630 96702 86682 96754
rect 84916 96600 84968 96652
rect 84980 96600 85032 96652
rect 85044 96600 85096 96652
rect 85108 96600 85160 96652
rect 1714 96498 1766 96550
rect 4106 96498 4158 96550
rect 4474 96498 4526 96550
rect 5026 96498 5078 96550
rect 35018 96498 35070 96550
rect 38606 96498 38658 96550
rect 61974 96498 62026 96550
rect 62526 96498 62578 96550
rect 74394 96498 74446 96550
rect 77430 96498 77482 96550
rect 2174 96362 2226 96414
rect 2726 96362 2778 96414
rect 36858 96430 36910 96482
rect 53050 96430 53102 96482
rect 56822 96430 56874 96482
rect 62066 96430 62118 96482
rect 66574 96430 66626 96482
rect 81478 96430 81530 96482
rect 83870 96498 83922 96550
rect 84146 96498 84198 96550
rect 85342 96430 85394 96482
rect 15698 96362 15750 96414
rect 24438 96362 24490 96414
rect 46518 96362 46570 96414
rect 84422 96362 84474 96414
rect 3186 96337 3238 96346
rect 3186 96303 3195 96337
rect 3195 96303 3229 96337
rect 3229 96303 3238 96337
rect 3186 96294 3238 96303
rect 4290 96294 4342 96346
rect 41826 96294 41878 96346
rect 44494 96294 44546 96346
rect 82398 96294 82450 96346
rect 83778 96337 83830 96346
rect 83778 96303 83787 96337
rect 83787 96303 83821 96337
rect 83821 96303 83830 96337
rect 83778 96294 83830 96303
rect 83870 96294 83922 96346
rect 85158 96294 85210 96346
rect 2174 96226 2226 96278
rect 2358 96158 2410 96210
rect 4290 96158 4342 96210
rect 2916 96056 2968 96108
rect 2980 96056 3032 96108
rect 3044 96056 3096 96108
rect 3108 96056 3160 96108
rect 5486 96090 5538 96142
rect 5762 96090 5814 96142
rect 2634 95954 2686 96006
rect 4658 95954 4710 96006
rect 24990 96226 25042 96278
rect 33546 96226 33598 96278
rect 34466 96226 34518 96278
rect 45322 96226 45374 96278
rect 50198 96226 50250 96278
rect 85986 96226 86038 96278
rect 47806 96158 47858 96210
rect 82122 96158 82174 96210
rect 85434 96158 85486 96210
rect 51578 96090 51630 96142
rect 82766 96090 82818 96142
rect 37502 96022 37554 96074
rect 53050 96022 53102 96074
rect 18366 95954 18418 96006
rect 23426 95886 23478 95938
rect 1714 95818 1766 95870
rect 2358 95818 2410 95870
rect 23978 95818 24030 95870
rect 43758 95818 43810 95870
rect 82214 96022 82266 96074
rect 86916 96056 86968 96108
rect 86980 96056 87032 96108
rect 87044 96056 87096 96108
rect 87108 96056 87160 96108
rect 57926 95954 57978 96006
rect 81202 95954 81254 96006
rect 84146 95954 84198 96006
rect 61790 95886 61842 95938
rect 80282 95886 80334 95938
rect 62802 95818 62854 95870
rect 81938 95818 81990 95870
rect 4750 95682 4802 95734
rect 14042 95682 14094 95734
rect 916 95512 968 95564
rect 980 95512 1032 95564
rect 1044 95512 1096 95564
rect 1108 95512 1160 95564
rect 5486 95546 5538 95598
rect 25726 95750 25778 95802
rect 63446 95750 63498 95802
rect 82582 95750 82634 95802
rect 68966 95682 69018 95734
rect 81294 95682 81346 95734
rect 18366 95478 18418 95530
rect 34926 95614 34978 95666
rect 47622 95614 47674 95666
rect 38146 95546 38198 95598
rect 62342 95546 62394 95598
rect 26646 95478 26698 95530
rect 35018 95478 35070 95530
rect 51486 95478 51538 95530
rect 61974 95478 62026 95530
rect 4842 95410 4894 95462
rect 11834 95410 11886 95462
rect 36214 95410 36266 95462
rect 45322 95410 45374 95462
rect 53142 95410 53194 95462
rect 3738 95342 3790 95394
rect 19838 95342 19890 95394
rect 20758 95342 20810 95394
rect 45414 95342 45466 95394
rect 53234 95342 53286 95394
rect 62250 95410 62302 95462
rect 71174 95614 71226 95666
rect 80190 95614 80242 95666
rect 69058 95546 69110 95598
rect 77430 95546 77482 95598
rect 84916 95512 84968 95564
rect 84980 95512 85032 95564
rect 85044 95512 85096 95564
rect 85108 95512 85160 95564
rect 68874 95410 68926 95462
rect 77430 95410 77482 95462
rect 84698 95410 84750 95462
rect 58018 95342 58070 95394
rect 69242 95342 69294 95394
rect 80098 95342 80150 95394
rect 86262 95342 86314 95394
rect 4198 95274 4250 95326
rect 31154 95274 31206 95326
rect 35662 95274 35714 95326
rect 51762 95274 51814 95326
rect 53050 95274 53102 95326
rect 69886 95274 69938 95326
rect 4290 95206 4342 95258
rect 2726 95138 2778 95190
rect 4842 95206 4894 95258
rect 36306 95206 36358 95258
rect 16986 95138 17038 95190
rect 24438 95138 24490 95190
rect 29774 95138 29826 95190
rect 4474 95070 4526 95122
rect 4566 95070 4618 95122
rect 4750 95070 4802 95122
rect 5026 95070 5078 95122
rect 8154 95070 8206 95122
rect 58110 95206 58162 95258
rect 59398 95206 59450 95258
rect 63354 95206 63406 95258
rect 68414 95206 68466 95258
rect 85158 95206 85210 95258
rect 48726 95138 48778 95190
rect 54154 95138 54206 95190
rect 80190 95138 80242 95190
rect 84054 95138 84106 95190
rect 49094 95070 49146 95122
rect 51670 95070 51722 95122
rect 58018 95070 58070 95122
rect 66482 95070 66534 95122
rect 71082 95070 71134 95122
rect 2916 94968 2968 95020
rect 2980 94968 3032 95020
rect 3044 94968 3096 95020
rect 3108 94968 3160 95020
rect 37318 95002 37370 95054
rect 53050 95002 53102 95054
rect 77430 95002 77482 95054
rect 38790 94934 38842 94986
rect 3370 94866 3422 94918
rect 8154 94866 8206 94918
rect 25910 94866 25962 94918
rect 29682 94866 29734 94918
rect 43942 94866 43994 94918
rect 51026 94866 51078 94918
rect 54154 94866 54206 94918
rect 82030 94934 82082 94986
rect 86916 94968 86968 95020
rect 86980 94968 87032 95020
rect 87044 94968 87096 95020
rect 87108 94968 87160 95020
rect 84606 94866 84658 94918
rect 4934 94798 4986 94850
rect 11098 94798 11150 94850
rect 50382 94798 50434 94850
rect 1622 94730 1674 94782
rect 1898 94730 1950 94782
rect 26002 94730 26054 94782
rect 50290 94730 50342 94782
rect 20850 94662 20902 94714
rect 30694 94662 30746 94714
rect 38790 94662 38842 94714
rect 41734 94662 41786 94714
rect 56822 94730 56874 94782
rect 62158 94798 62210 94850
rect 69150 94798 69202 94850
rect 83318 94798 83370 94850
rect 2266 94594 2318 94646
rect 2634 94594 2686 94646
rect 27290 94594 27342 94646
rect 29774 94594 29826 94646
rect 40170 94594 40222 94646
rect 52958 94594 53010 94646
rect 69058 94730 69110 94782
rect 82306 94730 82358 94782
rect 82766 94730 82818 94782
rect 85710 94730 85762 94782
rect 68414 94662 68466 94714
rect 68506 94662 68558 94714
rect 70990 94662 71042 94714
rect 72462 94662 72514 94714
rect 83410 94662 83462 94714
rect 83962 94594 84014 94646
rect 5026 94526 5078 94578
rect 32442 94526 32494 94578
rect 49094 94526 49146 94578
rect 84790 94526 84842 94578
rect 916 94424 968 94476
rect 980 94424 1032 94476
rect 1044 94424 1096 94476
rect 1108 94424 1160 94476
rect 3370 94322 3422 94374
rect 3738 94322 3790 94374
rect 2726 94254 2778 94306
rect 4290 94458 4342 94510
rect 41458 94458 41510 94510
rect 42654 94458 42706 94510
rect 72370 94458 72422 94510
rect 72554 94458 72606 94510
rect 80190 94458 80242 94510
rect 40078 94390 40130 94442
rect 53142 94390 53194 94442
rect 54246 94390 54298 94442
rect 63262 94390 63314 94442
rect 66482 94390 66534 94442
rect 70990 94390 71042 94442
rect 74394 94390 74446 94442
rect 81202 94390 81254 94442
rect 84916 94424 84968 94476
rect 84980 94424 85032 94476
rect 85044 94424 85096 94476
rect 85108 94424 85160 94476
rect 29774 94322 29826 94374
rect 33454 94322 33506 94374
rect 51670 94322 51722 94374
rect 84330 94322 84382 94374
rect 38054 94254 38106 94306
rect 42654 94254 42706 94306
rect 60778 94254 60830 94306
rect 69058 94254 69110 94306
rect 3738 94186 3790 94238
rect 23334 94186 23386 94238
rect 48818 94186 48870 94238
rect 69150 94186 69202 94238
rect 41274 94118 41326 94170
rect 69794 94118 69846 94170
rect 72370 94118 72422 94170
rect 84422 94118 84474 94170
rect 28394 94050 28446 94102
rect 36306 94050 36358 94102
rect 45230 94050 45282 94102
rect 84054 94050 84106 94102
rect 5854 93982 5906 94034
rect 18274 93982 18326 94034
rect 24622 93982 24674 94034
rect 38238 93982 38290 94034
rect 43942 93982 43994 94034
rect 84146 93982 84198 94034
rect 2916 93880 2968 93932
rect 2980 93880 3032 93932
rect 3044 93880 3096 93932
rect 3108 93880 3160 93932
rect 18182 93914 18234 93966
rect 48450 93914 48502 93966
rect 72554 93914 72606 93966
rect 5394 93846 5446 93898
rect 19838 93846 19890 93898
rect 46150 93846 46202 93898
rect 81294 93846 81346 93898
rect 86916 93880 86968 93932
rect 86980 93880 87032 93932
rect 87044 93880 87096 93932
rect 87108 93880 87160 93932
rect 63354 93778 63406 93830
rect 72462 93778 72514 93830
rect 38882 93710 38934 93762
rect 53234 93710 53286 93762
rect 53694 93710 53746 93762
rect 60042 93710 60094 93762
rect 62250 93710 62302 93762
rect 83962 93710 84014 93762
rect 45322 93642 45374 93694
rect 56362 93642 56414 93694
rect 60778 93642 60830 93694
rect 68966 93642 69018 93694
rect 71082 93642 71134 93694
rect 78442 93642 78494 93694
rect 34926 93574 34978 93626
rect 84606 93574 84658 93626
rect 33638 93506 33690 93558
rect 82674 93506 82726 93558
rect 42746 93438 42798 93490
rect 60502 93438 60554 93490
rect 78442 93438 78494 93490
rect 82582 93438 82634 93490
rect 916 93336 968 93388
rect 980 93336 1032 93388
rect 1044 93336 1096 93388
rect 1108 93336 1160 93388
rect 63446 93370 63498 93422
rect 69886 93370 69938 93422
rect 80190 93370 80242 93422
rect 33454 93302 33506 93354
rect 82214 93302 82266 93354
rect 84916 93336 84968 93388
rect 84980 93336 85032 93388
rect 85044 93336 85096 93388
rect 85108 93336 85160 93388
rect 32350 93234 32402 93286
rect 83410 93234 83462 93286
rect 31062 93166 31114 93218
rect 83318 93166 83370 93218
rect 48450 93098 48502 93150
rect 62526 93098 62578 93150
rect 69242 93098 69294 93150
rect 84238 93098 84290 93150
rect 45414 93030 45466 93082
rect 63262 93030 63314 93082
rect 69794 93030 69846 93082
rect 36214 92962 36266 93014
rect 84790 92962 84842 93014
rect 38790 92894 38842 92946
rect 60042 92894 60094 92946
rect 71174 92894 71226 92946
rect 73750 92894 73802 92946
rect 83778 92937 83830 92946
rect 83778 92903 83787 92937
rect 83787 92903 83821 92937
rect 83821 92903 83830 92937
rect 83778 92894 83830 92903
rect 2916 92792 2968 92844
rect 2980 92792 3032 92844
rect 3044 92792 3096 92844
rect 3108 92792 3160 92844
rect 51762 92826 51814 92878
rect 62434 92826 62486 92878
rect 60870 92758 60922 92810
rect 81202 92758 81254 92810
rect 81938 92758 81990 92810
rect 86916 92792 86968 92844
rect 86980 92792 87032 92844
rect 87044 92792 87096 92844
rect 87108 92792 87160 92844
rect 62342 92690 62394 92742
rect 84330 92690 84382 92742
rect 68874 92622 68926 92674
rect 85158 92622 85210 92674
rect 55350 92554 55402 92606
rect 69058 92554 69110 92606
rect 80190 92554 80242 92606
rect 40170 92486 40222 92538
rect 80098 92486 80150 92538
rect 82030 92486 82082 92538
rect 82766 92418 82818 92470
rect 83870 92350 83922 92402
rect 916 92248 968 92300
rect 980 92248 1032 92300
rect 1044 92248 1096 92300
rect 1108 92248 1160 92300
rect 84916 92248 84968 92300
rect 84980 92248 85032 92300
rect 85044 92248 85096 92300
rect 85108 92248 85160 92300
rect 84698 92146 84750 92198
rect 81294 92010 81346 92062
rect 85158 92010 85210 92062
rect 83962 91942 84014 91994
rect 84514 91942 84566 91994
rect 83962 91806 84014 91858
rect 2916 91704 2968 91756
rect 2980 91704 3032 91756
rect 3044 91704 3096 91756
rect 3108 91704 3160 91756
rect 86916 91704 86968 91756
rect 86980 91704 87032 91756
rect 87044 91704 87096 91756
rect 87108 91704 87160 91756
rect 916 91160 968 91212
rect 980 91160 1032 91212
rect 1044 91160 1096 91212
rect 1108 91160 1160 91212
rect 84916 91160 84968 91212
rect 84980 91160 85032 91212
rect 85044 91160 85096 91212
rect 85108 91160 85160 91212
rect 2916 90616 2968 90668
rect 2980 90616 3032 90668
rect 3044 90616 3096 90668
rect 3108 90616 3160 90668
rect 86916 90616 86968 90668
rect 86980 90616 87032 90668
rect 87044 90616 87096 90668
rect 87108 90616 87160 90668
rect 916 90072 968 90124
rect 980 90072 1032 90124
rect 1044 90072 1096 90124
rect 1108 90072 1160 90124
rect 84916 90072 84968 90124
rect 84980 90072 85032 90124
rect 85044 90072 85096 90124
rect 85108 90072 85160 90124
rect 3370 89902 3422 89954
rect 5394 89945 5446 89954
rect 5394 89911 5403 89945
rect 5403 89911 5437 89945
rect 5437 89911 5446 89945
rect 5394 89902 5446 89911
rect 81386 89902 81438 89954
rect 84054 89902 84106 89954
rect 2916 89528 2968 89580
rect 2980 89528 3032 89580
rect 3044 89528 3096 89580
rect 3108 89528 3160 89580
rect 86916 89528 86968 89580
rect 86980 89528 87032 89580
rect 87044 89528 87096 89580
rect 87108 89528 87160 89580
rect 83870 89222 83922 89274
rect 84146 89222 84198 89274
rect 916 88984 968 89036
rect 980 88984 1032 89036
rect 1044 88984 1096 89036
rect 1108 88984 1160 89036
rect 84916 88984 84968 89036
rect 84980 88984 85032 89036
rect 85044 88984 85096 89036
rect 85108 88984 85160 89036
rect 2910 88610 2962 88662
rect 3738 88610 3790 88662
rect 3922 88610 3974 88662
rect 4106 88542 4158 88594
rect 2916 88440 2968 88492
rect 2980 88440 3032 88492
rect 3044 88440 3096 88492
rect 3108 88440 3160 88492
rect 86916 88440 86968 88492
rect 86980 88440 87032 88492
rect 87044 88440 87096 88492
rect 87108 88440 87160 88492
rect 83594 87998 83646 88050
rect 83870 87998 83922 88050
rect 84146 87998 84198 88050
rect 84422 87998 84474 88050
rect 916 87896 968 87948
rect 980 87896 1032 87948
rect 1044 87896 1096 87948
rect 1108 87896 1160 87948
rect 84916 87896 84968 87948
rect 84980 87896 85032 87948
rect 85044 87896 85096 87948
rect 85108 87896 85160 87948
rect 3738 87794 3790 87846
rect 82674 87794 82726 87846
rect 84146 87794 84198 87846
rect 2916 87352 2968 87404
rect 2980 87352 3032 87404
rect 3044 87352 3096 87404
rect 3108 87352 3160 87404
rect 86916 87352 86968 87404
rect 86980 87352 87032 87404
rect 87044 87352 87096 87404
rect 87108 87352 87160 87404
rect 916 86808 968 86860
rect 980 86808 1032 86860
rect 1044 86808 1096 86860
rect 1108 86808 1160 86860
rect 84916 86808 84968 86860
rect 84980 86808 85032 86860
rect 85044 86808 85096 86860
rect 85108 86808 85160 86860
rect 2916 86264 2968 86316
rect 2980 86264 3032 86316
rect 3044 86264 3096 86316
rect 3108 86264 3160 86316
rect 86916 86264 86968 86316
rect 86980 86264 87032 86316
rect 87044 86264 87096 86316
rect 87108 86264 87160 86316
rect 3830 85822 3882 85874
rect 4198 85822 4250 85874
rect 84146 85822 84198 85874
rect 84330 85822 84382 85874
rect 916 85720 968 85772
rect 980 85720 1032 85772
rect 1044 85720 1096 85772
rect 1108 85720 1160 85772
rect 84916 85720 84968 85772
rect 84980 85720 85032 85772
rect 85044 85720 85096 85772
rect 85108 85720 85160 85772
rect 2916 85176 2968 85228
rect 2980 85176 3032 85228
rect 3044 85176 3096 85228
rect 3108 85176 3160 85228
rect 86916 85176 86968 85228
rect 86980 85176 87032 85228
rect 87044 85176 87096 85228
rect 87108 85176 87160 85228
rect 4014 84802 4066 84854
rect 83410 84734 83462 84786
rect 84146 84734 84198 84786
rect 916 84632 968 84684
rect 980 84632 1032 84684
rect 1044 84632 1096 84684
rect 1108 84632 1160 84684
rect 84916 84632 84968 84684
rect 84980 84632 85032 84684
rect 85044 84632 85096 84684
rect 85108 84632 85160 84684
rect 2916 84088 2968 84140
rect 2980 84088 3032 84140
rect 3044 84088 3096 84140
rect 3108 84088 3160 84140
rect 86916 84088 86968 84140
rect 86980 84088 87032 84140
rect 87044 84088 87096 84140
rect 87108 84088 87160 84140
rect 82214 83714 82266 83766
rect 84330 83714 84382 83766
rect 916 83544 968 83596
rect 980 83544 1032 83596
rect 1044 83544 1096 83596
rect 1108 83544 1160 83596
rect 84916 83544 84968 83596
rect 84980 83544 85032 83596
rect 85044 83544 85096 83596
rect 85108 83544 85160 83596
rect 5578 83374 5630 83426
rect 3554 83145 3606 83154
rect 3554 83111 3563 83145
rect 3563 83111 3597 83145
rect 3597 83111 3606 83145
rect 3554 83102 3606 83111
rect 2916 83000 2968 83052
rect 2980 83000 3032 83052
rect 3044 83000 3096 83052
rect 3108 83000 3160 83052
rect 86916 83000 86968 83052
rect 86980 83000 87032 83052
rect 87044 83000 87096 83052
rect 87108 83000 87160 83052
rect 916 82456 968 82508
rect 980 82456 1032 82508
rect 1044 82456 1096 82508
rect 1108 82456 1160 82508
rect 84916 82456 84968 82508
rect 84980 82456 85032 82508
rect 85044 82456 85096 82508
rect 85108 82456 85160 82508
rect 2634 82218 2686 82270
rect 3278 82218 3330 82270
rect 2916 81912 2968 81964
rect 2980 81912 3032 81964
rect 3044 81912 3096 81964
rect 3108 81912 3160 81964
rect 86916 81912 86968 81964
rect 86980 81912 87032 81964
rect 87044 81912 87096 81964
rect 87108 81912 87160 81964
rect 916 81368 968 81420
rect 980 81368 1032 81420
rect 1044 81368 1096 81420
rect 1108 81368 1160 81420
rect 84916 81368 84968 81420
rect 84980 81368 85032 81420
rect 85044 81368 85096 81420
rect 85108 81368 85160 81420
rect 3370 80926 3422 80978
rect 83042 80926 83094 80978
rect 83226 80926 83278 80978
rect 83870 80926 83922 80978
rect 85250 80926 85302 80978
rect 2916 80824 2968 80876
rect 2980 80824 3032 80876
rect 3044 80824 3096 80876
rect 3108 80824 3160 80876
rect 86916 80824 86968 80876
rect 86980 80824 87032 80876
rect 87044 80824 87096 80876
rect 87108 80824 87160 80876
rect 916 80280 968 80332
rect 980 80280 1032 80332
rect 1044 80280 1096 80332
rect 1108 80280 1160 80332
rect 84916 80280 84968 80332
rect 84980 80280 85032 80332
rect 85044 80280 85096 80332
rect 85108 80280 85160 80332
rect 3646 79838 3698 79890
rect 2916 79736 2968 79788
rect 2980 79736 3032 79788
rect 3044 79736 3096 79788
rect 3108 79736 3160 79788
rect 86916 79736 86968 79788
rect 86980 79736 87032 79788
rect 87044 79736 87096 79788
rect 87108 79736 87160 79788
rect 916 79192 968 79244
rect 980 79192 1032 79244
rect 1044 79192 1096 79244
rect 1108 79192 1160 79244
rect 84916 79192 84968 79244
rect 84980 79192 85032 79244
rect 85044 79192 85096 79244
rect 85108 79192 85160 79244
rect 2916 78648 2968 78700
rect 2980 78648 3032 78700
rect 3044 78648 3096 78700
rect 3108 78648 3160 78700
rect 86916 78648 86968 78700
rect 86980 78648 87032 78700
rect 87044 78648 87096 78700
rect 87108 78648 87160 78700
rect 916 78104 968 78156
rect 980 78104 1032 78156
rect 1044 78104 1096 78156
rect 1108 78104 1160 78156
rect 84916 78104 84968 78156
rect 84980 78104 85032 78156
rect 85044 78104 85096 78156
rect 85108 78104 85160 78156
rect 2916 77560 2968 77612
rect 2980 77560 3032 77612
rect 3044 77560 3096 77612
rect 3108 77560 3160 77612
rect 86916 77560 86968 77612
rect 86980 77560 87032 77612
rect 87044 77560 87096 77612
rect 87108 77560 87160 77612
rect 81662 77322 81714 77374
rect 84606 77322 84658 77374
rect 916 77016 968 77068
rect 980 77016 1032 77068
rect 1044 77016 1096 77068
rect 1108 77016 1160 77068
rect 84916 77016 84968 77068
rect 84980 77016 85032 77068
rect 85044 77016 85096 77068
rect 85108 77016 85160 77068
rect 2916 76472 2968 76524
rect 2980 76472 3032 76524
rect 3044 76472 3096 76524
rect 3108 76472 3160 76524
rect 86916 76472 86968 76524
rect 86980 76472 87032 76524
rect 87044 76472 87096 76524
rect 87108 76472 87160 76524
rect 916 75928 968 75980
rect 980 75928 1032 75980
rect 1044 75928 1096 75980
rect 1108 75928 1160 75980
rect 84916 75928 84968 75980
rect 84980 75928 85032 75980
rect 85044 75928 85096 75980
rect 85108 75928 85160 75980
rect 2916 75384 2968 75436
rect 2980 75384 3032 75436
rect 3044 75384 3096 75436
rect 3108 75384 3160 75436
rect 86916 75384 86968 75436
rect 86980 75384 87032 75436
rect 87044 75384 87096 75436
rect 87108 75384 87160 75436
rect 84054 74942 84106 74994
rect 84790 74942 84842 74994
rect 916 74840 968 74892
rect 980 74840 1032 74892
rect 1044 74840 1096 74892
rect 1108 74840 1160 74892
rect 84916 74840 84968 74892
rect 84980 74840 85032 74892
rect 85044 74840 85096 74892
rect 85108 74840 85160 74892
rect 81846 74466 81898 74518
rect 84882 74466 84934 74518
rect 82490 74398 82542 74450
rect 84330 74398 84382 74450
rect 2916 74296 2968 74348
rect 2980 74296 3032 74348
rect 3044 74296 3096 74348
rect 3108 74296 3160 74348
rect 86916 74296 86968 74348
rect 86980 74296 87032 74348
rect 87044 74296 87096 74348
rect 87108 74296 87160 74348
rect 916 73752 968 73804
rect 980 73752 1032 73804
rect 1044 73752 1096 73804
rect 1108 73752 1160 73804
rect 84916 73752 84968 73804
rect 84980 73752 85032 73804
rect 85044 73752 85096 73804
rect 85108 73752 85160 73804
rect 2916 73208 2968 73260
rect 2980 73208 3032 73260
rect 3044 73208 3096 73260
rect 3108 73208 3160 73260
rect 86916 73208 86968 73260
rect 86980 73208 87032 73260
rect 87044 73208 87096 73260
rect 87108 73208 87160 73260
rect 82122 73106 82174 73158
rect 84698 73106 84750 73158
rect 82306 73038 82358 73090
rect 84790 73038 84842 73090
rect 916 72664 968 72716
rect 980 72664 1032 72716
rect 1044 72664 1096 72716
rect 1108 72664 1160 72716
rect 84916 72664 84968 72716
rect 84980 72664 85032 72716
rect 85044 72664 85096 72716
rect 85108 72664 85160 72716
rect 2916 72120 2968 72172
rect 2980 72120 3032 72172
rect 3044 72120 3096 72172
rect 3108 72120 3160 72172
rect 86916 72120 86968 72172
rect 86980 72120 87032 72172
rect 87044 72120 87096 72172
rect 87108 72120 87160 72172
rect 916 71576 968 71628
rect 980 71576 1032 71628
rect 1044 71576 1096 71628
rect 1108 71576 1160 71628
rect 84916 71576 84968 71628
rect 84980 71576 85032 71628
rect 85044 71576 85096 71628
rect 85108 71576 85160 71628
rect 2916 71032 2968 71084
rect 2980 71032 3032 71084
rect 3044 71032 3096 71084
rect 3108 71032 3160 71084
rect 86916 71032 86968 71084
rect 86980 71032 87032 71084
rect 87044 71032 87096 71084
rect 87108 71032 87160 71084
rect 916 70488 968 70540
rect 980 70488 1032 70540
rect 1044 70488 1096 70540
rect 1108 70488 1160 70540
rect 84916 70488 84968 70540
rect 84980 70488 85032 70540
rect 85044 70488 85096 70540
rect 85108 70488 85160 70540
rect 2916 69944 2968 69996
rect 2980 69944 3032 69996
rect 3044 69944 3096 69996
rect 3108 69944 3160 69996
rect 86916 69944 86968 69996
rect 86980 69944 87032 69996
rect 87044 69944 87096 69996
rect 87108 69944 87160 69996
rect 916 69400 968 69452
rect 980 69400 1032 69452
rect 1044 69400 1096 69452
rect 1108 69400 1160 69452
rect 84916 69400 84968 69452
rect 84980 69400 85032 69452
rect 85044 69400 85096 69452
rect 85108 69400 85160 69452
rect 2916 68856 2968 68908
rect 2980 68856 3032 68908
rect 3044 68856 3096 68908
rect 3108 68856 3160 68908
rect 86916 68856 86968 68908
rect 86980 68856 87032 68908
rect 87044 68856 87096 68908
rect 87108 68856 87160 68908
rect 916 68312 968 68364
rect 980 68312 1032 68364
rect 1044 68312 1096 68364
rect 1108 68312 1160 68364
rect 84916 68312 84968 68364
rect 84980 68312 85032 68364
rect 85044 68312 85096 68364
rect 85108 68312 85160 68364
rect 2916 67768 2968 67820
rect 2980 67768 3032 67820
rect 3044 67768 3096 67820
rect 3108 67768 3160 67820
rect 86916 67768 86968 67820
rect 86980 67768 87032 67820
rect 87044 67768 87096 67820
rect 87108 67768 87160 67820
rect 916 67224 968 67276
rect 980 67224 1032 67276
rect 1044 67224 1096 67276
rect 1108 67224 1160 67276
rect 84916 67224 84968 67276
rect 84980 67224 85032 67276
rect 85044 67224 85096 67276
rect 85108 67224 85160 67276
rect 2916 66680 2968 66732
rect 2980 66680 3032 66732
rect 3044 66680 3096 66732
rect 3108 66680 3160 66732
rect 86916 66680 86968 66732
rect 86980 66680 87032 66732
rect 87044 66680 87096 66732
rect 87108 66680 87160 66732
rect 82030 66578 82082 66630
rect 85158 66578 85210 66630
rect 916 66136 968 66188
rect 980 66136 1032 66188
rect 1044 66136 1096 66188
rect 1108 66136 1160 66188
rect 84916 66136 84968 66188
rect 84980 66136 85032 66188
rect 85044 66136 85096 66188
rect 85108 66136 85160 66188
rect 2916 65592 2968 65644
rect 2980 65592 3032 65644
rect 3044 65592 3096 65644
rect 3108 65592 3160 65644
rect 86916 65592 86968 65644
rect 86980 65592 87032 65644
rect 87044 65592 87096 65644
rect 87108 65592 87160 65644
rect 916 65048 968 65100
rect 980 65048 1032 65100
rect 1044 65048 1096 65100
rect 1108 65048 1160 65100
rect 84916 65048 84968 65100
rect 84980 65048 85032 65100
rect 85044 65048 85096 65100
rect 85108 65048 85160 65100
rect 2916 64504 2968 64556
rect 2980 64504 3032 64556
rect 3044 64504 3096 64556
rect 3108 64504 3160 64556
rect 86916 64504 86968 64556
rect 86980 64504 87032 64556
rect 87044 64504 87096 64556
rect 87108 64504 87160 64556
rect 916 63960 968 64012
rect 980 63960 1032 64012
rect 1044 63960 1096 64012
rect 1108 63960 1160 64012
rect 84916 63960 84968 64012
rect 84980 63960 85032 64012
rect 85044 63960 85096 64012
rect 85108 63960 85160 64012
rect 2916 63416 2968 63468
rect 2980 63416 3032 63468
rect 3044 63416 3096 63468
rect 3108 63416 3160 63468
rect 86916 63416 86968 63468
rect 86980 63416 87032 63468
rect 87044 63416 87096 63468
rect 87108 63416 87160 63468
rect 3646 63314 3698 63366
rect 3646 62974 3698 63026
rect 3830 62974 3882 63026
rect 3922 62974 3974 63026
rect 916 62872 968 62924
rect 980 62872 1032 62924
rect 1044 62872 1096 62924
rect 1108 62872 1160 62924
rect 84916 62872 84968 62924
rect 84980 62872 85032 62924
rect 85044 62872 85096 62924
rect 85108 62872 85160 62924
rect 81938 62770 81990 62822
rect 84790 62770 84842 62822
rect 2916 62328 2968 62380
rect 2980 62328 3032 62380
rect 3044 62328 3096 62380
rect 3108 62328 3160 62380
rect 86916 62328 86968 62380
rect 86980 62328 87032 62380
rect 87044 62328 87096 62380
rect 87108 62328 87160 62380
rect 916 61784 968 61836
rect 980 61784 1032 61836
rect 1044 61784 1096 61836
rect 1108 61784 1160 61836
rect 84916 61784 84968 61836
rect 84980 61784 85032 61836
rect 85044 61784 85096 61836
rect 85108 61784 85160 61836
rect 3830 61546 3882 61598
rect 2916 61240 2968 61292
rect 2980 61240 3032 61292
rect 3044 61240 3096 61292
rect 3108 61240 3160 61292
rect 86916 61240 86968 61292
rect 86980 61240 87032 61292
rect 87044 61240 87096 61292
rect 87108 61240 87160 61292
rect 916 60696 968 60748
rect 980 60696 1032 60748
rect 1044 60696 1096 60748
rect 1108 60696 1160 60748
rect 84916 60696 84968 60748
rect 84980 60696 85032 60748
rect 85044 60696 85096 60748
rect 85108 60696 85160 60748
rect 2916 60152 2968 60204
rect 2980 60152 3032 60204
rect 3044 60152 3096 60204
rect 3108 60152 3160 60204
rect 86916 60152 86968 60204
rect 86980 60152 87032 60204
rect 87044 60152 87096 60204
rect 87108 60152 87160 60204
rect 916 59608 968 59660
rect 980 59608 1032 59660
rect 1044 59608 1096 59660
rect 1108 59608 1160 59660
rect 84916 59608 84968 59660
rect 84980 59608 85032 59660
rect 85044 59608 85096 59660
rect 85108 59608 85160 59660
rect 2916 59064 2968 59116
rect 2980 59064 3032 59116
rect 3044 59064 3096 59116
rect 3108 59064 3160 59116
rect 86916 59064 86968 59116
rect 86980 59064 87032 59116
rect 87044 59064 87096 59116
rect 87108 59064 87160 59116
rect 916 58520 968 58572
rect 980 58520 1032 58572
rect 1044 58520 1096 58572
rect 1108 58520 1160 58572
rect 84916 58520 84968 58572
rect 84980 58520 85032 58572
rect 85044 58520 85096 58572
rect 85108 58520 85160 58572
rect 2916 57976 2968 58028
rect 2980 57976 3032 58028
rect 3044 57976 3096 58028
rect 3108 57976 3160 58028
rect 86916 57976 86968 58028
rect 86980 57976 87032 58028
rect 87044 57976 87096 58028
rect 87108 57976 87160 58028
rect 916 57432 968 57484
rect 980 57432 1032 57484
rect 1044 57432 1096 57484
rect 1108 57432 1160 57484
rect 84916 57432 84968 57484
rect 84980 57432 85032 57484
rect 85044 57432 85096 57484
rect 85108 57432 85160 57484
rect 2916 56888 2968 56940
rect 2980 56888 3032 56940
rect 3044 56888 3096 56940
rect 3108 56888 3160 56940
rect 86916 56888 86968 56940
rect 86980 56888 87032 56940
rect 87044 56888 87096 56940
rect 87108 56888 87160 56940
rect 83134 56557 83186 56566
rect 83134 56523 83143 56557
rect 83143 56523 83177 56557
rect 83177 56523 83186 56557
rect 83134 56514 83186 56523
rect 81938 56446 81990 56498
rect 84790 56446 84842 56498
rect 83134 56421 83186 56430
rect 916 56344 968 56396
rect 980 56344 1032 56396
rect 1044 56344 1096 56396
rect 1108 56344 1160 56396
rect 83134 56387 83143 56421
rect 83143 56387 83177 56421
rect 83177 56387 83186 56421
rect 83134 56378 83186 56387
rect 84916 56344 84968 56396
rect 84980 56344 85032 56396
rect 85044 56344 85096 56396
rect 85108 56344 85160 56396
rect 3830 56242 3882 56294
rect 2916 55800 2968 55852
rect 2980 55800 3032 55852
rect 3044 55800 3096 55852
rect 3108 55800 3160 55852
rect 86916 55800 86968 55852
rect 86980 55800 87032 55852
rect 87044 55800 87096 55852
rect 87108 55800 87160 55852
rect 916 55256 968 55308
rect 980 55256 1032 55308
rect 1044 55256 1096 55308
rect 1108 55256 1160 55308
rect 84916 55256 84968 55308
rect 84980 55256 85032 55308
rect 85044 55256 85096 55308
rect 85108 55256 85160 55308
rect 2916 54712 2968 54764
rect 2980 54712 3032 54764
rect 3044 54712 3096 54764
rect 3108 54712 3160 54764
rect 86916 54712 86968 54764
rect 86980 54712 87032 54764
rect 87044 54712 87096 54764
rect 87108 54712 87160 54764
rect 916 54168 968 54220
rect 980 54168 1032 54220
rect 1044 54168 1096 54220
rect 1108 54168 1160 54220
rect 84916 54168 84968 54220
rect 84980 54168 85032 54220
rect 85044 54168 85096 54220
rect 85108 54168 85160 54220
rect 2916 53624 2968 53676
rect 2980 53624 3032 53676
rect 3044 53624 3096 53676
rect 3108 53624 3160 53676
rect 86916 53624 86968 53676
rect 86980 53624 87032 53676
rect 87044 53624 87096 53676
rect 87108 53624 87160 53676
rect 916 53080 968 53132
rect 980 53080 1032 53132
rect 1044 53080 1096 53132
rect 1108 53080 1160 53132
rect 84916 53080 84968 53132
rect 84980 53080 85032 53132
rect 85044 53080 85096 53132
rect 85108 53080 85160 53132
rect 2916 52536 2968 52588
rect 2980 52536 3032 52588
rect 3044 52536 3096 52588
rect 3108 52536 3160 52588
rect 82858 52570 82910 52622
rect 83134 52570 83186 52622
rect 86916 52536 86968 52588
rect 86980 52536 87032 52588
rect 87044 52536 87096 52588
rect 87108 52536 87160 52588
rect 916 51992 968 52044
rect 980 51992 1032 52044
rect 1044 51992 1096 52044
rect 1108 51992 1160 52044
rect 84916 51992 84968 52044
rect 84980 51992 85032 52044
rect 85044 51992 85096 52044
rect 85108 51992 85160 52044
rect 2916 51448 2968 51500
rect 2980 51448 3032 51500
rect 3044 51448 3096 51500
rect 3108 51448 3160 51500
rect 86916 51448 86968 51500
rect 86980 51448 87032 51500
rect 87044 51448 87096 51500
rect 87108 51448 87160 51500
rect 916 50904 968 50956
rect 980 50904 1032 50956
rect 1044 50904 1096 50956
rect 1108 50904 1160 50956
rect 84916 50904 84968 50956
rect 84980 50904 85032 50956
rect 85044 50904 85096 50956
rect 85108 50904 85160 50956
rect 2916 50360 2968 50412
rect 2980 50360 3032 50412
rect 3044 50360 3096 50412
rect 3108 50360 3160 50412
rect 86916 50360 86968 50412
rect 86980 50360 87032 50412
rect 87044 50360 87096 50412
rect 87108 50360 87160 50412
rect 82030 50054 82082 50106
rect 85158 50054 85210 50106
rect 916 49816 968 49868
rect 980 49816 1032 49868
rect 1044 49816 1096 49868
rect 1108 49816 1160 49868
rect 84916 49816 84968 49868
rect 84980 49816 85032 49868
rect 85044 49816 85096 49868
rect 85108 49816 85160 49868
rect 2916 49272 2968 49324
rect 2980 49272 3032 49324
rect 3044 49272 3096 49324
rect 3108 49272 3160 49324
rect 86916 49272 86968 49324
rect 86980 49272 87032 49324
rect 87044 49272 87096 49324
rect 87108 49272 87160 49324
rect 82122 48830 82174 48882
rect 84790 48830 84842 48882
rect 916 48728 968 48780
rect 980 48728 1032 48780
rect 1044 48728 1096 48780
rect 1108 48728 1160 48780
rect 84916 48728 84968 48780
rect 84980 48728 85032 48780
rect 85044 48728 85096 48780
rect 85108 48728 85160 48780
rect 2916 48184 2968 48236
rect 2980 48184 3032 48236
rect 3044 48184 3096 48236
rect 3108 48184 3160 48236
rect 86916 48184 86968 48236
rect 86980 48184 87032 48236
rect 87044 48184 87096 48236
rect 87108 48184 87160 48236
rect 916 47640 968 47692
rect 980 47640 1032 47692
rect 1044 47640 1096 47692
rect 1108 47640 1160 47692
rect 84916 47640 84968 47692
rect 84980 47640 85032 47692
rect 85044 47640 85096 47692
rect 85108 47640 85160 47692
rect 2916 47096 2968 47148
rect 2980 47096 3032 47148
rect 3044 47096 3096 47148
rect 3108 47096 3160 47148
rect 86916 47096 86968 47148
rect 86980 47096 87032 47148
rect 87044 47096 87096 47148
rect 87108 47096 87160 47148
rect 916 46552 968 46604
rect 980 46552 1032 46604
rect 1044 46552 1096 46604
rect 1108 46552 1160 46604
rect 84916 46552 84968 46604
rect 84980 46552 85032 46604
rect 85044 46552 85096 46604
rect 85108 46552 85160 46604
rect 2916 46008 2968 46060
rect 2980 46008 3032 46060
rect 3044 46008 3096 46060
rect 3108 46008 3160 46060
rect 86916 46008 86968 46060
rect 86980 46008 87032 46060
rect 87044 46008 87096 46060
rect 87108 46008 87160 46060
rect 916 45464 968 45516
rect 980 45464 1032 45516
rect 1044 45464 1096 45516
rect 1108 45464 1160 45516
rect 84916 45464 84968 45516
rect 84980 45464 85032 45516
rect 85044 45464 85096 45516
rect 85108 45464 85160 45516
rect 2916 44920 2968 44972
rect 2980 44920 3032 44972
rect 3044 44920 3096 44972
rect 3108 44920 3160 44972
rect 86916 44920 86968 44972
rect 86980 44920 87032 44972
rect 87044 44920 87096 44972
rect 87108 44920 87160 44972
rect 3370 44818 3422 44870
rect 3646 44818 3698 44870
rect 3738 44818 3790 44870
rect 3830 44750 3882 44802
rect 3646 44546 3698 44598
rect 3738 44546 3790 44598
rect 3830 44478 3882 44530
rect 916 44376 968 44428
rect 980 44376 1032 44428
rect 1044 44376 1096 44428
rect 1108 44376 1160 44428
rect 84916 44376 84968 44428
rect 84980 44376 85032 44428
rect 85044 44376 85096 44428
rect 85108 44376 85160 44428
rect 2916 43832 2968 43884
rect 2980 43832 3032 43884
rect 3044 43832 3096 43884
rect 3108 43832 3160 43884
rect 86916 43832 86968 43884
rect 86980 43832 87032 43884
rect 87044 43832 87096 43884
rect 87108 43832 87160 43884
rect 82214 43594 82266 43646
rect 85158 43594 85210 43646
rect 916 43288 968 43340
rect 980 43288 1032 43340
rect 1044 43288 1096 43340
rect 1108 43288 1160 43340
rect 84916 43288 84968 43340
rect 84980 43288 85032 43340
rect 85044 43288 85096 43340
rect 85108 43288 85160 43340
rect 2916 42744 2968 42796
rect 2980 42744 3032 42796
rect 3044 42744 3096 42796
rect 3108 42744 3160 42796
rect 86916 42744 86968 42796
rect 86980 42744 87032 42796
rect 87044 42744 87096 42796
rect 87108 42744 87160 42796
rect 916 42200 968 42252
rect 980 42200 1032 42252
rect 1044 42200 1096 42252
rect 1108 42200 1160 42252
rect 84916 42200 84968 42252
rect 84980 42200 85032 42252
rect 85044 42200 85096 42252
rect 85108 42200 85160 42252
rect 2916 41656 2968 41708
rect 2980 41656 3032 41708
rect 3044 41656 3096 41708
rect 3108 41656 3160 41708
rect 86916 41656 86968 41708
rect 86980 41656 87032 41708
rect 87044 41656 87096 41708
rect 87108 41656 87160 41708
rect 916 41112 968 41164
rect 980 41112 1032 41164
rect 1044 41112 1096 41164
rect 1108 41112 1160 41164
rect 84916 41112 84968 41164
rect 84980 41112 85032 41164
rect 85044 41112 85096 41164
rect 85108 41112 85160 41164
rect 2916 40568 2968 40620
rect 2980 40568 3032 40620
rect 3044 40568 3096 40620
rect 3108 40568 3160 40620
rect 86916 40568 86968 40620
rect 86980 40568 87032 40620
rect 87044 40568 87096 40620
rect 87108 40568 87160 40620
rect 916 40024 968 40076
rect 980 40024 1032 40076
rect 1044 40024 1096 40076
rect 1108 40024 1160 40076
rect 84916 40024 84968 40076
rect 84980 40024 85032 40076
rect 85044 40024 85096 40076
rect 85108 40024 85160 40076
rect 82306 39922 82358 39974
rect 84790 39922 84842 39974
rect 2916 39480 2968 39532
rect 2980 39480 3032 39532
rect 3044 39480 3096 39532
rect 3108 39480 3160 39532
rect 86916 39480 86968 39532
rect 86980 39480 87032 39532
rect 87044 39480 87096 39532
rect 87108 39480 87160 39532
rect 916 38936 968 38988
rect 980 38936 1032 38988
rect 1044 38936 1096 38988
rect 1108 38936 1160 38988
rect 84916 38936 84968 38988
rect 84980 38936 85032 38988
rect 85044 38936 85096 38988
rect 85108 38936 85160 38988
rect 2916 38392 2968 38444
rect 2980 38392 3032 38444
rect 3044 38392 3096 38444
rect 3108 38392 3160 38444
rect 86916 38392 86968 38444
rect 86980 38392 87032 38444
rect 87044 38392 87096 38444
rect 87108 38392 87160 38444
rect 3922 38290 3974 38342
rect 916 37848 968 37900
rect 980 37848 1032 37900
rect 1044 37848 1096 37900
rect 1108 37848 1160 37900
rect 84916 37848 84968 37900
rect 84980 37848 85032 37900
rect 85044 37848 85096 37900
rect 85108 37848 85160 37900
rect 2916 37304 2968 37356
rect 2980 37304 3032 37356
rect 3044 37304 3096 37356
rect 3108 37304 3160 37356
rect 86916 37304 86968 37356
rect 86980 37304 87032 37356
rect 87044 37304 87096 37356
rect 87108 37304 87160 37356
rect 916 36760 968 36812
rect 980 36760 1032 36812
rect 1044 36760 1096 36812
rect 1108 36760 1160 36812
rect 84916 36760 84968 36812
rect 84980 36760 85032 36812
rect 85044 36760 85096 36812
rect 85108 36760 85160 36812
rect 2916 36216 2968 36268
rect 2980 36216 3032 36268
rect 3044 36216 3096 36268
rect 3108 36216 3160 36268
rect 86916 36216 86968 36268
rect 86980 36216 87032 36268
rect 87044 36216 87096 36268
rect 87108 36216 87160 36268
rect 3278 35842 3330 35894
rect 3830 35842 3882 35894
rect 916 35672 968 35724
rect 980 35672 1032 35724
rect 1044 35672 1096 35724
rect 1108 35672 1160 35724
rect 84916 35672 84968 35724
rect 84980 35672 85032 35724
rect 85044 35672 85096 35724
rect 85108 35672 85160 35724
rect 82398 35434 82450 35486
rect 84146 35434 84198 35486
rect 2916 35128 2968 35180
rect 2980 35128 3032 35180
rect 3044 35128 3096 35180
rect 3108 35128 3160 35180
rect 86916 35128 86968 35180
rect 86980 35128 87032 35180
rect 87044 35128 87096 35180
rect 87108 35128 87160 35180
rect 916 34584 968 34636
rect 980 34584 1032 34636
rect 1044 34584 1096 34636
rect 1108 34584 1160 34636
rect 84916 34584 84968 34636
rect 84980 34584 85032 34636
rect 85044 34584 85096 34636
rect 85108 34584 85160 34636
rect 2916 34040 2968 34092
rect 2980 34040 3032 34092
rect 3044 34040 3096 34092
rect 3108 34040 3160 34092
rect 86916 34040 86968 34092
rect 86980 34040 87032 34092
rect 87044 34040 87096 34092
rect 87108 34040 87160 34092
rect 916 33496 968 33548
rect 980 33496 1032 33548
rect 1044 33496 1096 33548
rect 1108 33496 1160 33548
rect 84916 33496 84968 33548
rect 84980 33496 85032 33548
rect 85044 33496 85096 33548
rect 85108 33496 85160 33548
rect 2916 32952 2968 33004
rect 2980 32952 3032 33004
rect 3044 32952 3096 33004
rect 3108 32952 3160 33004
rect 86916 32952 86968 33004
rect 86980 32952 87032 33004
rect 87044 32952 87096 33004
rect 87108 32952 87160 33004
rect 916 32408 968 32460
rect 980 32408 1032 32460
rect 1044 32408 1096 32460
rect 1108 32408 1160 32460
rect 84916 32408 84968 32460
rect 84980 32408 85032 32460
rect 85044 32408 85096 32460
rect 85108 32408 85160 32460
rect 82490 32034 82542 32086
rect 84238 32034 84290 32086
rect 83686 31966 83738 32018
rect 85342 31966 85394 32018
rect 2916 31864 2968 31916
rect 2980 31864 3032 31916
rect 3044 31864 3096 31916
rect 3108 31864 3160 31916
rect 86916 31864 86968 31916
rect 86980 31864 87032 31916
rect 87044 31864 87096 31916
rect 87108 31864 87160 31916
rect 84054 31422 84106 31474
rect 85986 31422 86038 31474
rect 916 31320 968 31372
rect 980 31320 1032 31372
rect 1044 31320 1096 31372
rect 1108 31320 1160 31372
rect 84916 31320 84968 31372
rect 84980 31320 85032 31372
rect 85044 31320 85096 31372
rect 85108 31320 85160 31372
rect 82950 30878 83002 30930
rect 84146 30878 84198 30930
rect 2916 30776 2968 30828
rect 2980 30776 3032 30828
rect 3044 30776 3096 30828
rect 3108 30776 3160 30828
rect 86916 30776 86968 30828
rect 86980 30776 87032 30828
rect 87044 30776 87096 30828
rect 87108 30776 87160 30828
rect 916 30232 968 30284
rect 980 30232 1032 30284
rect 1044 30232 1096 30284
rect 1108 30232 1160 30284
rect 84916 30232 84968 30284
rect 84980 30232 85032 30284
rect 85044 30232 85096 30284
rect 85108 30232 85160 30284
rect 84054 29858 84106 29910
rect 2916 29688 2968 29740
rect 2980 29688 3032 29740
rect 3044 29688 3096 29740
rect 3108 29688 3160 29740
rect 86916 29688 86968 29740
rect 86980 29688 87032 29740
rect 87044 29688 87096 29740
rect 87108 29688 87160 29740
rect 3830 29450 3882 29502
rect 81846 29450 81898 29502
rect 84330 29450 84382 29502
rect 84790 29382 84842 29434
rect 3830 29314 3882 29366
rect 84330 29314 84382 29366
rect 916 29144 968 29196
rect 980 29144 1032 29196
rect 1044 29144 1096 29196
rect 1108 29144 1160 29196
rect 84916 29144 84968 29196
rect 84980 29144 85032 29196
rect 85044 29144 85096 29196
rect 85108 29144 85160 29196
rect 84146 28702 84198 28754
rect 2916 28600 2968 28652
rect 2980 28600 3032 28652
rect 3044 28600 3096 28652
rect 3108 28600 3160 28652
rect 86916 28600 86968 28652
rect 86980 28600 87032 28652
rect 87044 28600 87096 28652
rect 87108 28600 87160 28652
rect 81754 28498 81806 28550
rect 84422 28498 84474 28550
rect 83226 28226 83278 28278
rect 85434 28226 85486 28278
rect 82858 28158 82910 28210
rect 84698 28158 84750 28210
rect 916 28056 968 28108
rect 980 28056 1032 28108
rect 1044 28056 1096 28108
rect 1108 28056 1160 28108
rect 84916 28056 84968 28108
rect 84980 28056 85032 28108
rect 85044 28056 85096 28108
rect 85108 28056 85160 28108
rect 2916 27512 2968 27564
rect 2980 27512 3032 27564
rect 3044 27512 3096 27564
rect 3108 27512 3160 27564
rect 86916 27512 86968 27564
rect 86980 27512 87032 27564
rect 87044 27512 87096 27564
rect 87108 27512 87160 27564
rect 84238 27070 84290 27122
rect 84698 27070 84750 27122
rect 916 26968 968 27020
rect 980 26968 1032 27020
rect 1044 26968 1096 27020
rect 1108 26968 1160 27020
rect 84916 26968 84968 27020
rect 84980 26968 85032 27020
rect 85044 26968 85096 27020
rect 85108 26968 85160 27020
rect 2916 26424 2968 26476
rect 2980 26424 3032 26476
rect 3044 26424 3096 26476
rect 3108 26424 3160 26476
rect 86916 26424 86968 26476
rect 86980 26424 87032 26476
rect 87044 26424 87096 26476
rect 87108 26424 87160 26476
rect 83502 25982 83554 26034
rect 916 25880 968 25932
rect 980 25880 1032 25932
rect 1044 25880 1096 25932
rect 1108 25880 1160 25932
rect 84916 25880 84968 25932
rect 84980 25880 85032 25932
rect 85044 25880 85096 25932
rect 85108 25880 85160 25932
rect 81662 25574 81714 25626
rect 84882 25574 84934 25626
rect 3278 25506 3330 25558
rect 3370 25506 3422 25558
rect 2916 25336 2968 25388
rect 2980 25336 3032 25388
rect 3044 25336 3096 25388
rect 3108 25336 3160 25388
rect 86916 25336 86968 25388
rect 86980 25336 87032 25388
rect 87044 25336 87096 25388
rect 87108 25336 87160 25388
rect 916 24792 968 24844
rect 980 24792 1032 24844
rect 1044 24792 1096 24844
rect 1108 24792 1160 24844
rect 84916 24792 84968 24844
rect 84980 24792 85032 24844
rect 85044 24792 85096 24844
rect 85108 24792 85160 24844
rect 2916 24248 2968 24300
rect 2980 24248 3032 24300
rect 3044 24248 3096 24300
rect 3108 24248 3160 24300
rect 86916 24248 86968 24300
rect 86980 24248 87032 24300
rect 87044 24248 87096 24300
rect 87108 24248 87160 24300
rect 3278 24146 3330 24198
rect 84238 24010 84290 24062
rect 84698 24010 84750 24062
rect 84238 23806 84290 23858
rect 916 23704 968 23756
rect 980 23704 1032 23756
rect 1044 23704 1096 23756
rect 1108 23704 1160 23756
rect 84916 23704 84968 23756
rect 84980 23704 85032 23756
rect 85044 23704 85096 23756
rect 85108 23704 85160 23756
rect 2916 23160 2968 23212
rect 2980 23160 3032 23212
rect 3044 23160 3096 23212
rect 3108 23160 3160 23212
rect 86916 23160 86968 23212
rect 86980 23160 87032 23212
rect 87044 23160 87096 23212
rect 87108 23160 87160 23212
rect 3830 22922 3882 22974
rect 83962 22922 84014 22974
rect 916 22616 968 22668
rect 980 22616 1032 22668
rect 1044 22616 1096 22668
rect 1108 22616 1160 22668
rect 84916 22616 84968 22668
rect 84980 22616 85032 22668
rect 85044 22616 85096 22668
rect 85108 22616 85160 22668
rect 3830 22514 3882 22566
rect 2916 22072 2968 22124
rect 2980 22072 3032 22124
rect 3044 22072 3096 22124
rect 3108 22072 3160 22124
rect 86916 22072 86968 22124
rect 86980 22072 87032 22124
rect 87044 22072 87096 22124
rect 87108 22072 87160 22124
rect 916 21528 968 21580
rect 980 21528 1032 21580
rect 1044 21528 1096 21580
rect 1108 21528 1160 21580
rect 84916 21528 84968 21580
rect 84980 21528 85032 21580
rect 85044 21528 85096 21580
rect 85108 21528 85160 21580
rect 2916 20984 2968 21036
rect 2980 20984 3032 21036
rect 3044 20984 3096 21036
rect 3108 20984 3160 21036
rect 86916 20984 86968 21036
rect 86980 20984 87032 21036
rect 87044 20984 87096 21036
rect 87108 20984 87160 21036
rect 4290 20542 4342 20594
rect 916 20440 968 20492
rect 980 20440 1032 20492
rect 1044 20440 1096 20492
rect 1108 20440 1160 20492
rect 84916 20440 84968 20492
rect 84980 20440 85032 20492
rect 85044 20440 85096 20492
rect 85108 20440 85160 20492
rect 83502 20202 83554 20254
rect 84790 20202 84842 20254
rect 83502 19998 83554 20050
rect 84054 19998 84106 20050
rect 2916 19896 2968 19948
rect 2980 19896 3032 19948
rect 3044 19896 3096 19948
rect 3108 19896 3160 19948
rect 86916 19896 86968 19948
rect 86980 19896 87032 19948
rect 87044 19896 87096 19948
rect 87108 19896 87160 19948
rect 82582 19590 82634 19642
rect 85526 19590 85578 19642
rect 916 19352 968 19404
rect 980 19352 1032 19404
rect 1044 19352 1096 19404
rect 1108 19352 1160 19404
rect 84916 19352 84968 19404
rect 84980 19352 85032 19404
rect 85044 19352 85096 19404
rect 85108 19352 85160 19404
rect 2916 18808 2968 18860
rect 2980 18808 3032 18860
rect 3044 18808 3096 18860
rect 3108 18808 3160 18860
rect 86916 18808 86968 18860
rect 86980 18808 87032 18860
rect 87044 18808 87096 18860
rect 87108 18808 87160 18860
rect 83502 18366 83554 18418
rect 83962 18366 84014 18418
rect 916 18264 968 18316
rect 980 18264 1032 18316
rect 1044 18264 1096 18316
rect 1108 18264 1160 18316
rect 84916 18264 84968 18316
rect 84980 18264 85032 18316
rect 85044 18264 85096 18316
rect 85108 18264 85160 18316
rect 2916 17720 2968 17772
rect 2980 17720 3032 17772
rect 3044 17720 3096 17772
rect 3108 17720 3160 17772
rect 86916 17720 86968 17772
rect 86980 17720 87032 17772
rect 87044 17720 87096 17772
rect 87108 17720 87160 17772
rect 916 17176 968 17228
rect 980 17176 1032 17228
rect 1044 17176 1096 17228
rect 1108 17176 1160 17228
rect 84916 17176 84968 17228
rect 84980 17176 85032 17228
rect 85044 17176 85096 17228
rect 85108 17176 85160 17228
rect 2916 16632 2968 16684
rect 2980 16632 3032 16684
rect 3044 16632 3096 16684
rect 3108 16632 3160 16684
rect 86916 16632 86968 16684
rect 86980 16632 87032 16684
rect 87044 16632 87096 16684
rect 87108 16632 87160 16684
rect 3922 16530 3974 16582
rect 916 16088 968 16140
rect 980 16088 1032 16140
rect 1044 16088 1096 16140
rect 1108 16088 1160 16140
rect 84916 16088 84968 16140
rect 84980 16088 85032 16140
rect 85044 16088 85096 16140
rect 85108 16088 85160 16140
rect 84330 15850 84382 15902
rect 84606 15850 84658 15902
rect 2916 15544 2968 15596
rect 2980 15544 3032 15596
rect 3044 15544 3096 15596
rect 3108 15544 3160 15596
rect 86916 15544 86968 15596
rect 86980 15544 87032 15596
rect 87044 15544 87096 15596
rect 87108 15544 87160 15596
rect 3278 15238 3330 15290
rect 916 15000 968 15052
rect 980 15000 1032 15052
rect 1044 15000 1096 15052
rect 1108 15000 1160 15052
rect 84916 15000 84968 15052
rect 84980 15000 85032 15052
rect 85044 15000 85096 15052
rect 85108 15000 85160 15052
rect 2916 14456 2968 14508
rect 2980 14456 3032 14508
rect 3044 14456 3096 14508
rect 3108 14456 3160 14508
rect 86916 14456 86968 14508
rect 86980 14456 87032 14508
rect 87044 14456 87096 14508
rect 87108 14456 87160 14508
rect 916 13912 968 13964
rect 980 13912 1032 13964
rect 1044 13912 1096 13964
rect 1108 13912 1160 13964
rect 84916 13912 84968 13964
rect 84980 13912 85032 13964
rect 85044 13912 85096 13964
rect 85108 13912 85160 13964
rect 83778 13810 83830 13862
rect 84146 13810 84198 13862
rect 3278 13606 3330 13658
rect 2916 13368 2968 13420
rect 2980 13368 3032 13420
rect 3044 13368 3096 13420
rect 3108 13368 3160 13420
rect 86916 13368 86968 13420
rect 86980 13368 87032 13420
rect 87044 13368 87096 13420
rect 87108 13368 87160 13420
rect 916 12824 968 12876
rect 980 12824 1032 12876
rect 1044 12824 1096 12876
rect 1108 12824 1160 12876
rect 84916 12824 84968 12876
rect 84980 12824 85032 12876
rect 85044 12824 85096 12876
rect 85108 12824 85160 12876
rect 2916 12280 2968 12332
rect 2980 12280 3032 12332
rect 3044 12280 3096 12332
rect 3108 12280 3160 12332
rect 86916 12280 86968 12332
rect 86980 12280 87032 12332
rect 87044 12280 87096 12332
rect 87108 12280 87160 12332
rect 916 11736 968 11788
rect 980 11736 1032 11788
rect 1044 11736 1096 11788
rect 1108 11736 1160 11788
rect 84916 11736 84968 11788
rect 84980 11736 85032 11788
rect 85044 11736 85096 11788
rect 85108 11736 85160 11788
rect 3922 11430 3974 11482
rect 5578 11430 5630 11482
rect 3830 11362 3882 11414
rect 5486 11362 5538 11414
rect 2916 11192 2968 11244
rect 2980 11192 3032 11244
rect 3044 11192 3096 11244
rect 3108 11192 3160 11244
rect 86916 11192 86968 11244
rect 86980 11192 87032 11244
rect 87044 11192 87096 11244
rect 87108 11192 87160 11244
rect 916 10648 968 10700
rect 980 10648 1032 10700
rect 1044 10648 1096 10700
rect 1108 10648 1160 10700
rect 84916 10648 84968 10700
rect 84980 10648 85032 10700
rect 85044 10648 85096 10700
rect 85108 10648 85160 10700
rect 2916 10104 2968 10156
rect 2980 10104 3032 10156
rect 3044 10104 3096 10156
rect 3108 10104 3160 10156
rect 86916 10104 86968 10156
rect 86980 10104 87032 10156
rect 87044 10104 87096 10156
rect 87108 10104 87160 10156
rect 916 9560 968 9612
rect 980 9560 1032 9612
rect 1044 9560 1096 9612
rect 1108 9560 1160 9612
rect 84916 9560 84968 9612
rect 84980 9560 85032 9612
rect 85044 9560 85096 9612
rect 85108 9560 85160 9612
rect 2916 9016 2968 9068
rect 2980 9016 3032 9068
rect 3044 9016 3096 9068
rect 3108 9016 3160 9068
rect 86916 9016 86968 9068
rect 86980 9016 87032 9068
rect 87044 9016 87096 9068
rect 87108 9016 87160 9068
rect 82582 8821 82634 8830
rect 82582 8787 82591 8821
rect 82591 8787 82625 8821
rect 82625 8787 82634 8821
rect 82582 8778 82634 8787
rect 916 8472 968 8524
rect 980 8472 1032 8524
rect 1044 8472 1096 8524
rect 1108 8472 1160 8524
rect 84916 8472 84968 8524
rect 84980 8472 85032 8524
rect 85044 8472 85096 8524
rect 85108 8472 85160 8524
rect 2916 7928 2968 7980
rect 2980 7928 3032 7980
rect 3044 7928 3096 7980
rect 3108 7928 3160 7980
rect 86916 7928 86968 7980
rect 86980 7928 87032 7980
rect 87044 7928 87096 7980
rect 87108 7928 87160 7980
rect 82582 7554 82634 7606
rect 85066 7554 85118 7606
rect 916 7384 968 7436
rect 980 7384 1032 7436
rect 1044 7384 1096 7436
rect 1108 7384 1160 7436
rect 84916 7384 84968 7436
rect 84980 7384 85032 7436
rect 85044 7384 85096 7436
rect 85108 7384 85160 7436
rect 84330 7146 84382 7198
rect 84790 7146 84842 7198
rect 81570 7010 81622 7062
rect 82030 7010 82082 7062
rect 2916 6840 2968 6892
rect 2980 6840 3032 6892
rect 3044 6840 3096 6892
rect 3108 6840 3160 6892
rect 82030 6874 82082 6926
rect 82398 6874 82450 6926
rect 86916 6840 86968 6892
rect 86980 6840 87032 6892
rect 87044 6840 87096 6892
rect 87108 6840 87160 6892
rect 916 6296 968 6348
rect 980 6296 1032 6348
rect 1044 6296 1096 6348
rect 1108 6296 1160 6348
rect 84916 6296 84968 6348
rect 84980 6296 85032 6348
rect 85044 6296 85096 6348
rect 85108 6296 85160 6348
rect 3646 6194 3698 6246
rect 5762 6194 5814 6246
rect 2916 5752 2968 5804
rect 2980 5752 3032 5804
rect 3044 5752 3096 5804
rect 3108 5752 3160 5804
rect 86916 5752 86968 5804
rect 86980 5752 87032 5804
rect 87044 5752 87096 5804
rect 87108 5752 87160 5804
rect 916 5208 968 5260
rect 980 5208 1032 5260
rect 1044 5208 1096 5260
rect 1108 5208 1160 5260
rect 84916 5208 84968 5260
rect 84980 5208 85032 5260
rect 85044 5208 85096 5260
rect 85108 5208 85160 5260
rect 3646 5106 3698 5158
rect 4474 4834 4526 4886
rect 2916 4664 2968 4716
rect 2980 4664 3032 4716
rect 3044 4664 3096 4716
rect 3108 4664 3160 4716
rect 4382 4562 4434 4614
rect 86916 4664 86968 4716
rect 86980 4664 87032 4716
rect 87044 4664 87096 4716
rect 87108 4664 87160 4716
rect 4382 4426 4434 4478
rect 1530 4222 1582 4274
rect 2910 4222 2962 4274
rect 916 4120 968 4172
rect 980 4120 1032 4172
rect 1044 4120 1096 4172
rect 1108 4120 1160 4172
rect 84916 4120 84968 4172
rect 84980 4120 85032 4172
rect 85044 4120 85096 4172
rect 85108 4120 85160 4172
rect 1990 4061 2042 4070
rect 1990 4027 1999 4061
rect 1999 4027 2033 4061
rect 2033 4027 2042 4061
rect 1990 4018 2042 4027
rect 2266 4018 2318 4070
rect 2542 4018 2594 4070
rect 2818 4061 2870 4070
rect 2818 4027 2827 4061
rect 2827 4027 2861 4061
rect 2861 4027 2870 4061
rect 2818 4018 2870 4027
rect 3922 4018 3974 4070
rect 83778 4061 83830 4070
rect 83778 4027 83787 4061
rect 83787 4027 83821 4061
rect 83821 4027 83830 4061
rect 83778 4018 83830 4027
rect 3370 3950 3422 4002
rect 5026 3950 5078 4002
rect 5302 3882 5354 3934
rect 83594 3678 83646 3730
rect 2916 3576 2968 3628
rect 2980 3576 3032 3628
rect 3044 3576 3096 3628
rect 3108 3576 3160 3628
rect 82398 3610 82450 3662
rect 82766 3610 82818 3662
rect 86916 3576 86968 3628
rect 86980 3576 87032 3628
rect 87044 3576 87096 3628
rect 87108 3576 87160 3628
rect 3278 3474 3330 3526
rect 82766 3517 82818 3526
rect 82766 3483 82775 3517
rect 82775 3483 82809 3517
rect 82809 3483 82818 3517
rect 82766 3474 82818 3483
rect 85434 3474 85486 3526
rect 2082 3406 2134 3458
rect 2358 3406 2410 3458
rect 2818 3338 2870 3390
rect 4474 3338 4526 3390
rect 85802 3338 85854 3390
rect 1714 3245 1766 3254
rect 1714 3211 1723 3245
rect 1723 3211 1757 3245
rect 1757 3211 1766 3245
rect 1714 3202 1766 3211
rect 1346 3177 1398 3186
rect 1346 3143 1355 3177
rect 1355 3143 1389 3177
rect 1389 3143 1398 3177
rect 1346 3134 1398 3143
rect 2450 3177 2502 3186
rect 2450 3143 2459 3177
rect 2459 3143 2493 3177
rect 2493 3143 2502 3177
rect 2450 3134 2502 3143
rect 916 3032 968 3084
rect 980 3032 1032 3084
rect 1044 3032 1096 3084
rect 1108 3032 1160 3084
rect 8706 2998 8758 3050
rect 36950 2998 37002 3050
rect 82214 2998 82266 3050
rect 2358 2930 2410 2982
rect 2818 2973 2870 2982
rect 2818 2939 2827 2973
rect 2827 2939 2861 2973
rect 2861 2939 2870 2973
rect 2818 2930 2870 2939
rect 3278 2930 3330 2982
rect 33730 2930 33782 2982
rect 53694 2930 53746 2982
rect 82398 3202 82450 3254
rect 83778 3177 83830 3186
rect 83778 3143 83787 3177
rect 83787 3143 83821 3177
rect 83821 3143 83830 3177
rect 83778 3134 83830 3143
rect 84916 3032 84968 3084
rect 84980 3032 85032 3084
rect 85044 3032 85096 3084
rect 85108 3032 85160 3084
rect 82674 2930 82726 2982
rect 84238 2973 84290 2982
rect 84238 2939 84247 2973
rect 84247 2939 84281 2973
rect 84281 2939 84290 2973
rect 84238 2930 84290 2939
rect 85342 2930 85394 2982
rect 1806 2862 1858 2914
rect 3002 2862 3054 2914
rect 4566 2862 4618 2914
rect 23978 2862 24030 2914
rect 34834 2862 34886 2914
rect 84790 2862 84842 2914
rect 84974 2905 85026 2914
rect 84974 2871 84983 2905
rect 84983 2871 85017 2905
rect 85017 2871 85026 2905
rect 84974 2862 85026 2871
rect 86630 2862 86682 2914
rect 2726 2794 2778 2846
rect 978 2633 1030 2642
rect 978 2599 987 2633
rect 987 2599 1021 2633
rect 1021 2599 1030 2633
rect 978 2590 1030 2599
rect 2726 2658 2778 2710
rect 4934 2794 4986 2846
rect 27474 2794 27526 2846
rect 38790 2794 38842 2846
rect 61974 2794 62026 2846
rect 85894 2794 85946 2846
rect 22138 2726 22190 2778
rect 37594 2726 37646 2778
rect 84330 2726 84382 2778
rect 19746 2658 19798 2710
rect 41366 2658 41418 2710
rect 81386 2658 81438 2710
rect 82398 2658 82450 2710
rect 86538 2726 86590 2778
rect 19470 2590 19522 2642
rect 24622 2590 24674 2642
rect 2916 2488 2968 2540
rect 2980 2488 3032 2540
rect 3044 2488 3096 2540
rect 3108 2488 3160 2540
rect 978 2386 1030 2438
rect 1438 2386 1490 2438
rect 25082 2522 25134 2574
rect 50474 2522 50526 2574
rect 4106 2454 4158 2506
rect 7878 2454 7930 2506
rect 26002 2454 26054 2506
rect 28394 2454 28446 2506
rect 61974 2522 62026 2574
rect 83502 2590 83554 2642
rect 84974 2590 85026 2642
rect 86916 2488 86968 2540
rect 86980 2488 87032 2540
rect 87044 2488 87096 2540
rect 87108 2488 87160 2540
rect 31062 2386 31114 2438
rect 50198 2386 50250 2438
rect 81386 2386 81438 2438
rect 3554 2318 3606 2370
rect 84054 2318 84106 2370
rect 4842 2250 4894 2302
rect 5762 2250 5814 2302
rect 83962 2250 84014 2302
rect 2634 2182 2686 2234
rect 81294 2182 81346 2234
rect 2174 2114 2226 2166
rect 18274 2114 18326 2166
rect 35018 2114 35070 2166
rect 42470 2114 42522 2166
rect 1714 2089 1766 2098
rect 1714 2055 1723 2089
rect 1723 2055 1757 2089
rect 1757 2055 1766 2089
rect 1714 2046 1766 2055
rect 2818 2046 2870 2098
rect 4658 2046 4710 2098
rect 46702 2046 46754 2098
rect 85250 2182 85302 2234
rect 83502 2114 83554 2166
rect 916 1944 968 1996
rect 980 1944 1032 1996
rect 1044 1944 1096 1996
rect 1108 1944 1160 1996
rect 84916 1944 84968 1996
rect 84980 1944 85032 1996
rect 85044 1944 85096 1996
rect 85108 1944 85160 1996
rect 1714 1842 1766 1894
rect 26370 1842 26422 1894
rect 2818 1774 2870 1826
rect 3830 1774 3882 1826
rect 47898 1774 47950 1826
rect 84606 1774 84658 1826
rect 39986 1706 40038 1758
rect 84698 1706 84750 1758
rect 54246 1570 54298 1622
rect 83318 1570 83370 1622
rect 3922 1502 3974 1554
rect 41826 1502 41878 1554
rect 49830 1502 49882 1554
rect 81938 1502 81990 1554
rect 4658 1434 4710 1486
rect 29222 1434 29274 1486
rect 51486 1434 51538 1486
rect 83502 1434 83554 1486
rect 4842 1366 4894 1418
rect 36306 1366 36358 1418
rect 45230 1366 45282 1418
rect 42286 1298 42338 1350
rect 82122 1298 82174 1350
rect 24714 1230 24766 1282
rect 82950 1230 83002 1282
rect 3830 1162 3882 1214
rect 20850 1162 20902 1214
rect 22414 1162 22466 1214
rect 82858 1162 82910 1214
rect 18918 1094 18970 1146
rect 81662 1094 81714 1146
rect 2266 1026 2318 1078
rect 11834 1026 11886 1078
rect 28302 1026 28354 1078
rect 33086 1026 33138 1078
rect 3646 958 3698 1010
rect 14410 958 14462 1010
rect 29406 958 29458 1010
rect 37594 958 37646 1010
rect 4934 890 4986 942
rect 11742 890 11794 942
rect 21310 890 21362 942
rect 83226 890 83278 942
rect 2542 822 2594 874
rect 23426 822 23478 874
rect 24254 822 24306 874
rect 83686 822 83738 874
rect 4566 754 4618 806
rect 16986 754 17038 806
rect 31062 754 31114 806
rect 83042 754 83094 806
rect 31890 686 31942 738
rect 83134 686 83186 738
rect 2910 618 2962 670
rect 29866 618 29918 670
rect 32902 618 32954 670
rect 82306 618 82358 670
rect 18090 550 18142 602
rect 3278 482 3330 534
rect 32442 482 32494 534
rect 34742 550 34794 602
rect 34834 482 34886 534
rect 35294 482 35346 534
rect 82030 482 82082 534
rect 11742 414 11794 466
rect 83962 414 84014 466
rect 20758 346 20810 398
rect 39986 346 40038 398
rect 40078 346 40130 398
rect 82490 346 82542 398
rect 5302 278 5354 330
rect 38054 278 38106 330
rect 38330 278 38382 330
rect 81846 278 81898 330
rect 43942 210 43994 262
rect 81570 210 81622 262
rect 46150 142 46202 194
rect 83410 142 83462 194
rect 4290 74 4342 126
rect 84422 74 84474 126
rect 8706 6 8758 58
rect 85526 6 85578 58
<< metal2 >>
rect 84328 189202 84384 189211
rect 84328 189137 84384 189146
rect 5854 188554 5906 188560
rect 5854 188496 5906 188502
rect 82490 188554 82542 188560
rect 82490 188496 82542 188502
rect 5210 188486 5262 188492
rect 5210 188428 5262 188434
rect 2634 188350 2686 188356
rect 2634 188292 2686 188298
rect 2358 188282 2410 188288
rect 2358 188224 2410 188230
rect 2082 188146 2134 188152
rect 2082 188088 2134 188094
rect 1346 187874 1398 187880
rect 1346 187816 1398 187822
rect 1252 187298 1308 187307
rect 1252 187233 1308 187242
rect 890 186958 1186 186978
rect 946 186956 970 186958
rect 1026 186956 1050 186958
rect 1106 186956 1130 186958
rect 968 186904 970 186956
rect 1032 186904 1044 186956
rect 1106 186904 1108 186956
rect 946 186902 970 186904
rect 1026 186902 1050 186904
rect 1106 186902 1130 186904
rect 890 186882 1186 186902
rect 890 185870 1186 185890
rect 946 185868 970 185870
rect 1026 185868 1050 185870
rect 1106 185868 1130 185870
rect 968 185816 970 185868
rect 1032 185816 1044 185868
rect 1106 185816 1108 185868
rect 946 185814 970 185816
rect 1026 185814 1050 185816
rect 1106 185814 1130 185816
rect 890 185794 1186 185814
rect 890 184782 1186 184802
rect 946 184780 970 184782
rect 1026 184780 1050 184782
rect 1106 184780 1130 184782
rect 968 184728 970 184780
rect 1032 184728 1044 184780
rect 1106 184728 1108 184780
rect 946 184726 970 184728
rect 1026 184726 1050 184728
rect 1106 184726 1130 184728
rect 890 184706 1186 184726
rect 890 183694 1186 183714
rect 946 183692 970 183694
rect 1026 183692 1050 183694
rect 1106 183692 1130 183694
rect 968 183640 970 183692
rect 1032 183640 1044 183692
rect 1106 183640 1108 183692
rect 946 183638 970 183640
rect 1026 183638 1050 183640
rect 1106 183638 1130 183640
rect 890 183618 1186 183638
rect 890 182606 1186 182626
rect 946 182604 970 182606
rect 1026 182604 1050 182606
rect 1106 182604 1130 182606
rect 968 182552 970 182604
rect 1032 182552 1044 182604
rect 1106 182552 1108 182604
rect 946 182550 970 182552
rect 1026 182550 1050 182552
rect 1106 182550 1130 182552
rect 890 182530 1186 182550
rect 890 181518 1186 181538
rect 946 181516 970 181518
rect 1026 181516 1050 181518
rect 1106 181516 1130 181518
rect 968 181464 970 181516
rect 1032 181464 1044 181516
rect 1106 181464 1108 181516
rect 946 181462 970 181464
rect 1026 181462 1050 181464
rect 1106 181462 1130 181464
rect 890 181442 1186 181462
rect 890 180430 1186 180450
rect 946 180428 970 180430
rect 1026 180428 1050 180430
rect 1106 180428 1130 180430
rect 968 180376 970 180428
rect 1032 180376 1044 180428
rect 1106 180376 1108 180428
rect 946 180374 970 180376
rect 1026 180374 1050 180376
rect 1106 180374 1130 180376
rect 890 180354 1186 180374
rect 890 179342 1186 179362
rect 946 179340 970 179342
rect 1026 179340 1050 179342
rect 1106 179340 1130 179342
rect 968 179288 970 179340
rect 1032 179288 1044 179340
rect 1106 179288 1108 179340
rect 946 179286 970 179288
rect 1026 179286 1050 179288
rect 1106 179286 1130 179288
rect 890 179266 1186 179286
rect 890 178254 1186 178274
rect 946 178252 970 178254
rect 1026 178252 1050 178254
rect 1106 178252 1130 178254
rect 968 178200 970 178252
rect 1032 178200 1044 178252
rect 1106 178200 1108 178252
rect 946 178198 970 178200
rect 1026 178198 1050 178200
rect 1106 178198 1130 178200
rect 890 178178 1186 178198
rect 890 177166 1186 177186
rect 946 177164 970 177166
rect 1026 177164 1050 177166
rect 1106 177164 1130 177166
rect 968 177112 970 177164
rect 1032 177112 1044 177164
rect 1106 177112 1108 177164
rect 946 177110 970 177112
rect 1026 177110 1050 177112
rect 1106 177110 1130 177112
rect 890 177090 1186 177110
rect 890 176078 1186 176098
rect 946 176076 970 176078
rect 1026 176076 1050 176078
rect 1106 176076 1130 176078
rect 968 176024 970 176076
rect 1032 176024 1044 176076
rect 1106 176024 1108 176076
rect 946 176022 970 176024
rect 1026 176022 1050 176024
rect 1106 176022 1130 176024
rect 890 176002 1186 176022
rect 890 174990 1186 175010
rect 946 174988 970 174990
rect 1026 174988 1050 174990
rect 1106 174988 1130 174990
rect 968 174936 970 174988
rect 1032 174936 1044 174988
rect 1106 174936 1108 174988
rect 946 174934 970 174936
rect 1026 174934 1050 174936
rect 1106 174934 1130 174936
rect 890 174914 1186 174934
rect 890 173902 1186 173922
rect 946 173900 970 173902
rect 1026 173900 1050 173902
rect 1106 173900 1130 173902
rect 968 173848 970 173900
rect 1032 173848 1044 173900
rect 1106 173848 1108 173900
rect 946 173846 970 173848
rect 1026 173846 1050 173848
rect 1106 173846 1130 173848
rect 890 173826 1186 173846
rect 890 172814 1186 172834
rect 946 172812 970 172814
rect 1026 172812 1050 172814
rect 1106 172812 1130 172814
rect 968 172760 970 172812
rect 1032 172760 1044 172812
rect 1106 172760 1108 172812
rect 946 172758 970 172760
rect 1026 172758 1050 172760
rect 1106 172758 1130 172760
rect 890 172738 1186 172758
rect 890 171726 1186 171746
rect 946 171724 970 171726
rect 1026 171724 1050 171726
rect 1106 171724 1130 171726
rect 968 171672 970 171724
rect 1032 171672 1044 171724
rect 1106 171672 1108 171724
rect 946 171670 970 171672
rect 1026 171670 1050 171672
rect 1106 171670 1130 171672
rect 890 171650 1186 171670
rect 890 170638 1186 170658
rect 946 170636 970 170638
rect 1026 170636 1050 170638
rect 1106 170636 1130 170638
rect 968 170584 970 170636
rect 1032 170584 1044 170636
rect 1106 170584 1108 170636
rect 946 170582 970 170584
rect 1026 170582 1050 170584
rect 1106 170582 1130 170584
rect 890 170562 1186 170582
rect 890 169550 1186 169570
rect 946 169548 970 169550
rect 1026 169548 1050 169550
rect 1106 169548 1130 169550
rect 968 169496 970 169548
rect 1032 169496 1044 169548
rect 1106 169496 1108 169548
rect 946 169494 970 169496
rect 1026 169494 1050 169496
rect 1106 169494 1130 169496
rect 890 169474 1186 169494
rect 890 168462 1186 168482
rect 946 168460 970 168462
rect 1026 168460 1050 168462
rect 1106 168460 1130 168462
rect 968 168408 970 168460
rect 1032 168408 1044 168460
rect 1106 168408 1108 168460
rect 946 168406 970 168408
rect 1026 168406 1050 168408
rect 1106 168406 1130 168408
rect 890 168386 1186 168406
rect 890 167374 1186 167394
rect 946 167372 970 167374
rect 1026 167372 1050 167374
rect 1106 167372 1130 167374
rect 968 167320 970 167372
rect 1032 167320 1044 167372
rect 1106 167320 1108 167372
rect 946 167318 970 167320
rect 1026 167318 1050 167320
rect 1106 167318 1130 167320
rect 890 167298 1186 167318
rect 890 166286 1186 166306
rect 946 166284 970 166286
rect 1026 166284 1050 166286
rect 1106 166284 1130 166286
rect 968 166232 970 166284
rect 1032 166232 1044 166284
rect 1106 166232 1108 166284
rect 946 166230 970 166232
rect 1026 166230 1050 166232
rect 1106 166230 1130 166232
rect 890 166210 1186 166230
rect 890 165198 1186 165218
rect 946 165196 970 165198
rect 1026 165196 1050 165198
rect 1106 165196 1130 165198
rect 968 165144 970 165196
rect 1032 165144 1044 165196
rect 1106 165144 1108 165196
rect 946 165142 970 165144
rect 1026 165142 1050 165144
rect 1106 165142 1130 165144
rect 890 165122 1186 165142
rect 890 164110 1186 164130
rect 946 164108 970 164110
rect 1026 164108 1050 164110
rect 1106 164108 1130 164110
rect 968 164056 970 164108
rect 1032 164056 1044 164108
rect 1106 164056 1108 164108
rect 946 164054 970 164056
rect 1026 164054 1050 164056
rect 1106 164054 1130 164056
rect 890 164034 1186 164054
rect 890 163022 1186 163042
rect 946 163020 970 163022
rect 1026 163020 1050 163022
rect 1106 163020 1130 163022
rect 968 162968 970 163020
rect 1032 162968 1044 163020
rect 1106 162968 1108 163020
rect 946 162966 970 162968
rect 1026 162966 1050 162968
rect 1106 162966 1130 162968
rect 890 162946 1186 162966
rect 890 161934 1186 161954
rect 946 161932 970 161934
rect 1026 161932 1050 161934
rect 1106 161932 1130 161934
rect 968 161880 970 161932
rect 1032 161880 1044 161932
rect 1106 161880 1108 161932
rect 946 161878 970 161880
rect 1026 161878 1050 161880
rect 1106 161878 1130 161880
rect 890 161858 1186 161878
rect 890 160846 1186 160866
rect 946 160844 970 160846
rect 1026 160844 1050 160846
rect 1106 160844 1130 160846
rect 968 160792 970 160844
rect 1032 160792 1044 160844
rect 1106 160792 1108 160844
rect 946 160790 970 160792
rect 1026 160790 1050 160792
rect 1106 160790 1130 160792
rect 890 160770 1186 160790
rect 890 159758 1186 159778
rect 946 159756 970 159758
rect 1026 159756 1050 159758
rect 1106 159756 1130 159758
rect 968 159704 970 159756
rect 1032 159704 1044 159756
rect 1106 159704 1108 159756
rect 946 159702 970 159704
rect 1026 159702 1050 159704
rect 1106 159702 1130 159704
rect 890 159682 1186 159702
rect 890 158670 1186 158690
rect 946 158668 970 158670
rect 1026 158668 1050 158670
rect 1106 158668 1130 158670
rect 968 158616 970 158668
rect 1032 158616 1044 158668
rect 1106 158616 1108 158668
rect 946 158614 970 158616
rect 1026 158614 1050 158616
rect 1106 158614 1130 158616
rect 890 158594 1186 158614
rect 890 157582 1186 157602
rect 946 157580 970 157582
rect 1026 157580 1050 157582
rect 1106 157580 1130 157582
rect 968 157528 970 157580
rect 1032 157528 1044 157580
rect 1106 157528 1108 157580
rect 946 157526 970 157528
rect 1026 157526 1050 157528
rect 1106 157526 1130 157528
rect 890 157506 1186 157526
rect 890 156494 1186 156514
rect 946 156492 970 156494
rect 1026 156492 1050 156494
rect 1106 156492 1130 156494
rect 968 156440 970 156492
rect 1032 156440 1044 156492
rect 1106 156440 1108 156492
rect 946 156438 970 156440
rect 1026 156438 1050 156440
rect 1106 156438 1130 156440
rect 890 156418 1186 156438
rect 890 155406 1186 155426
rect 946 155404 970 155406
rect 1026 155404 1050 155406
rect 1106 155404 1130 155406
rect 968 155352 970 155404
rect 1032 155352 1044 155404
rect 1106 155352 1108 155404
rect 946 155350 970 155352
rect 1026 155350 1050 155352
rect 1106 155350 1130 155352
rect 890 155330 1186 155350
rect 890 154318 1186 154338
rect 946 154316 970 154318
rect 1026 154316 1050 154318
rect 1106 154316 1130 154318
rect 968 154264 970 154316
rect 1032 154264 1044 154316
rect 1106 154264 1108 154316
rect 946 154262 970 154264
rect 1026 154262 1050 154264
rect 1106 154262 1130 154264
rect 890 154242 1186 154262
rect 890 153230 1186 153250
rect 946 153228 970 153230
rect 1026 153228 1050 153230
rect 1106 153228 1130 153230
rect 968 153176 970 153228
rect 1032 153176 1044 153228
rect 1106 153176 1108 153228
rect 946 153174 970 153176
rect 1026 153174 1050 153176
rect 1106 153174 1130 153176
rect 890 153154 1186 153174
rect 890 152142 1186 152162
rect 946 152140 970 152142
rect 1026 152140 1050 152142
rect 1106 152140 1130 152142
rect 968 152088 970 152140
rect 1032 152088 1044 152140
rect 1106 152088 1108 152140
rect 946 152086 970 152088
rect 1026 152086 1050 152088
rect 1106 152086 1130 152088
rect 890 152066 1186 152086
rect 890 151054 1186 151074
rect 946 151052 970 151054
rect 1026 151052 1050 151054
rect 1106 151052 1130 151054
rect 968 151000 970 151052
rect 1032 151000 1044 151052
rect 1106 151000 1108 151052
rect 946 150998 970 151000
rect 1026 150998 1050 151000
rect 1106 150998 1130 151000
rect 890 150978 1186 150998
rect 890 149966 1186 149986
rect 946 149964 970 149966
rect 1026 149964 1050 149966
rect 1106 149964 1130 149966
rect 968 149912 970 149964
rect 1032 149912 1044 149964
rect 1106 149912 1108 149964
rect 946 149910 970 149912
rect 1026 149910 1050 149912
rect 1106 149910 1130 149912
rect 890 149890 1186 149910
rect 890 148878 1186 148898
rect 946 148876 970 148878
rect 1026 148876 1050 148878
rect 1106 148876 1130 148878
rect 968 148824 970 148876
rect 1032 148824 1044 148876
rect 1106 148824 1108 148876
rect 946 148822 970 148824
rect 1026 148822 1050 148824
rect 1106 148822 1130 148824
rect 890 148802 1186 148822
rect 890 147790 1186 147810
rect 946 147788 970 147790
rect 1026 147788 1050 147790
rect 1106 147788 1130 147790
rect 968 147736 970 147788
rect 1032 147736 1044 147788
rect 1106 147736 1108 147788
rect 946 147734 970 147736
rect 1026 147734 1050 147736
rect 1106 147734 1130 147736
rect 890 147714 1186 147734
rect 890 146702 1186 146722
rect 946 146700 970 146702
rect 1026 146700 1050 146702
rect 1106 146700 1130 146702
rect 968 146648 970 146700
rect 1032 146648 1044 146700
rect 1106 146648 1108 146700
rect 946 146646 970 146648
rect 1026 146646 1050 146648
rect 1106 146646 1130 146648
rect 890 146626 1186 146646
rect 890 145614 1186 145634
rect 946 145612 970 145614
rect 1026 145612 1050 145614
rect 1106 145612 1130 145614
rect 968 145560 970 145612
rect 1032 145560 1044 145612
rect 1106 145560 1108 145612
rect 946 145558 970 145560
rect 1026 145558 1050 145560
rect 1106 145558 1130 145560
rect 890 145538 1186 145558
rect 890 144526 1186 144546
rect 946 144524 970 144526
rect 1026 144524 1050 144526
rect 1106 144524 1130 144526
rect 968 144472 970 144524
rect 1032 144472 1044 144524
rect 1106 144472 1108 144524
rect 946 144470 970 144472
rect 1026 144470 1050 144472
rect 1106 144470 1130 144472
rect 890 144450 1186 144470
rect 890 143438 1186 143458
rect 946 143436 970 143438
rect 1026 143436 1050 143438
rect 1106 143436 1130 143438
rect 968 143384 970 143436
rect 1032 143384 1044 143436
rect 1106 143384 1108 143436
rect 946 143382 970 143384
rect 1026 143382 1050 143384
rect 1106 143382 1130 143384
rect 890 143362 1186 143382
rect 890 142350 1186 142370
rect 946 142348 970 142350
rect 1026 142348 1050 142350
rect 1106 142348 1130 142350
rect 968 142296 970 142348
rect 1032 142296 1044 142348
rect 1106 142296 1108 142348
rect 946 142294 970 142296
rect 1026 142294 1050 142296
rect 1106 142294 1130 142296
rect 890 142274 1186 142294
rect 890 141262 1186 141282
rect 946 141260 970 141262
rect 1026 141260 1050 141262
rect 1106 141260 1130 141262
rect 968 141208 970 141260
rect 1032 141208 1044 141260
rect 1106 141208 1108 141260
rect 946 141206 970 141208
rect 1026 141206 1050 141208
rect 1106 141206 1130 141208
rect 890 141186 1186 141206
rect 890 140174 1186 140194
rect 946 140172 970 140174
rect 1026 140172 1050 140174
rect 1106 140172 1130 140174
rect 968 140120 970 140172
rect 1032 140120 1044 140172
rect 1106 140120 1108 140172
rect 946 140118 970 140120
rect 1026 140118 1050 140120
rect 1106 140118 1130 140120
rect 890 140098 1186 140118
rect 890 139086 1186 139106
rect 946 139084 970 139086
rect 1026 139084 1050 139086
rect 1106 139084 1130 139086
rect 968 139032 970 139084
rect 1032 139032 1044 139084
rect 1106 139032 1108 139084
rect 946 139030 970 139032
rect 1026 139030 1050 139032
rect 1106 139030 1130 139032
rect 890 139010 1186 139030
rect 890 137998 1186 138018
rect 946 137996 970 137998
rect 1026 137996 1050 137998
rect 1106 137996 1130 137998
rect 968 137944 970 137996
rect 1032 137944 1044 137996
rect 1106 137944 1108 137996
rect 946 137942 970 137944
rect 1026 137942 1050 137944
rect 1106 137942 1130 137944
rect 890 137922 1186 137942
rect 890 136910 1186 136930
rect 946 136908 970 136910
rect 1026 136908 1050 136910
rect 1106 136908 1130 136910
rect 968 136856 970 136908
rect 1032 136856 1044 136908
rect 1106 136856 1108 136908
rect 946 136854 970 136856
rect 1026 136854 1050 136856
rect 1106 136854 1130 136856
rect 890 136834 1186 136854
rect 890 135822 1186 135842
rect 946 135820 970 135822
rect 1026 135820 1050 135822
rect 1106 135820 1130 135822
rect 968 135768 970 135820
rect 1032 135768 1044 135820
rect 1106 135768 1108 135820
rect 946 135766 970 135768
rect 1026 135766 1050 135768
rect 1106 135766 1130 135768
rect 890 135746 1186 135766
rect 890 134734 1186 134754
rect 946 134732 970 134734
rect 1026 134732 1050 134734
rect 1106 134732 1130 134734
rect 968 134680 970 134732
rect 1032 134680 1044 134732
rect 1106 134680 1108 134732
rect 946 134678 970 134680
rect 1026 134678 1050 134680
rect 1106 134678 1130 134680
rect 890 134658 1186 134678
rect 890 133646 1186 133666
rect 946 133644 970 133646
rect 1026 133644 1050 133646
rect 1106 133644 1130 133646
rect 968 133592 970 133644
rect 1032 133592 1044 133644
rect 1106 133592 1108 133644
rect 946 133590 970 133592
rect 1026 133590 1050 133592
rect 1106 133590 1130 133592
rect 890 133570 1186 133590
rect 890 132558 1186 132578
rect 946 132556 970 132558
rect 1026 132556 1050 132558
rect 1106 132556 1130 132558
rect 968 132504 970 132556
rect 1032 132504 1044 132556
rect 1106 132504 1108 132556
rect 946 132502 970 132504
rect 1026 132502 1050 132504
rect 1106 132502 1130 132504
rect 890 132482 1186 132502
rect 890 131470 1186 131490
rect 946 131468 970 131470
rect 1026 131468 1050 131470
rect 1106 131468 1130 131470
rect 968 131416 970 131468
rect 1032 131416 1044 131468
rect 1106 131416 1108 131468
rect 946 131414 970 131416
rect 1026 131414 1050 131416
rect 1106 131414 1130 131416
rect 890 131394 1186 131414
rect 890 130382 1186 130402
rect 946 130380 970 130382
rect 1026 130380 1050 130382
rect 1106 130380 1130 130382
rect 968 130328 970 130380
rect 1032 130328 1044 130380
rect 1106 130328 1108 130380
rect 946 130326 970 130328
rect 1026 130326 1050 130328
rect 1106 130326 1130 130328
rect 890 130306 1186 130326
rect 890 129294 1186 129314
rect 946 129292 970 129294
rect 1026 129292 1050 129294
rect 1106 129292 1130 129294
rect 968 129240 970 129292
rect 1032 129240 1044 129292
rect 1106 129240 1108 129292
rect 946 129238 970 129240
rect 1026 129238 1050 129240
rect 1106 129238 1130 129240
rect 890 129218 1186 129238
rect 890 128206 1186 128226
rect 946 128204 970 128206
rect 1026 128204 1050 128206
rect 1106 128204 1130 128206
rect 968 128152 970 128204
rect 1032 128152 1044 128204
rect 1106 128152 1108 128204
rect 946 128150 970 128152
rect 1026 128150 1050 128152
rect 1106 128150 1130 128152
rect 890 128130 1186 128150
rect 890 127118 1186 127138
rect 946 127116 970 127118
rect 1026 127116 1050 127118
rect 1106 127116 1130 127118
rect 968 127064 970 127116
rect 1032 127064 1044 127116
rect 1106 127064 1108 127116
rect 946 127062 970 127064
rect 1026 127062 1050 127064
rect 1106 127062 1130 127064
rect 890 127042 1186 127062
rect 890 126030 1186 126050
rect 946 126028 970 126030
rect 1026 126028 1050 126030
rect 1106 126028 1130 126030
rect 968 125976 970 126028
rect 1032 125976 1044 126028
rect 1106 125976 1108 126028
rect 946 125974 970 125976
rect 1026 125974 1050 125976
rect 1106 125974 1130 125976
rect 890 125954 1186 125974
rect 890 124942 1186 124962
rect 946 124940 970 124942
rect 1026 124940 1050 124942
rect 1106 124940 1130 124942
rect 968 124888 970 124940
rect 1032 124888 1044 124940
rect 1106 124888 1108 124940
rect 946 124886 970 124888
rect 1026 124886 1050 124888
rect 1106 124886 1130 124888
rect 890 124866 1186 124886
rect 890 123854 1186 123874
rect 946 123852 970 123854
rect 1026 123852 1050 123854
rect 1106 123852 1130 123854
rect 968 123800 970 123852
rect 1032 123800 1044 123852
rect 1106 123800 1108 123852
rect 946 123798 970 123800
rect 1026 123798 1050 123800
rect 1106 123798 1130 123800
rect 890 123778 1186 123798
rect 890 122766 1186 122786
rect 946 122764 970 122766
rect 1026 122764 1050 122766
rect 1106 122764 1130 122766
rect 968 122712 970 122764
rect 1032 122712 1044 122764
rect 1106 122712 1108 122764
rect 946 122710 970 122712
rect 1026 122710 1050 122712
rect 1106 122710 1130 122712
rect 890 122690 1186 122710
rect 890 121678 1186 121698
rect 946 121676 970 121678
rect 1026 121676 1050 121678
rect 1106 121676 1130 121678
rect 968 121624 970 121676
rect 1032 121624 1044 121676
rect 1106 121624 1108 121676
rect 946 121622 970 121624
rect 1026 121622 1050 121624
rect 1106 121622 1130 121624
rect 890 121602 1186 121622
rect 890 120590 1186 120610
rect 946 120588 970 120590
rect 1026 120588 1050 120590
rect 1106 120588 1130 120590
rect 968 120536 970 120588
rect 1032 120536 1044 120588
rect 1106 120536 1108 120588
rect 946 120534 970 120536
rect 1026 120534 1050 120536
rect 1106 120534 1130 120536
rect 890 120514 1186 120534
rect 890 119502 1186 119522
rect 946 119500 970 119502
rect 1026 119500 1050 119502
rect 1106 119500 1130 119502
rect 968 119448 970 119500
rect 1032 119448 1044 119500
rect 1106 119448 1108 119500
rect 946 119446 970 119448
rect 1026 119446 1050 119448
rect 1106 119446 1130 119448
rect 890 119426 1186 119446
rect 890 118414 1186 118434
rect 946 118412 970 118414
rect 1026 118412 1050 118414
rect 1106 118412 1130 118414
rect 968 118360 970 118412
rect 1032 118360 1044 118412
rect 1106 118360 1108 118412
rect 946 118358 970 118360
rect 1026 118358 1050 118360
rect 1106 118358 1130 118360
rect 890 118338 1186 118358
rect 890 117326 1186 117346
rect 946 117324 970 117326
rect 1026 117324 1050 117326
rect 1106 117324 1130 117326
rect 968 117272 970 117324
rect 1032 117272 1044 117324
rect 1106 117272 1108 117324
rect 946 117270 970 117272
rect 1026 117270 1050 117272
rect 1106 117270 1130 117272
rect 890 117250 1186 117270
rect 890 116238 1186 116258
rect 946 116236 970 116238
rect 1026 116236 1050 116238
rect 1106 116236 1130 116238
rect 968 116184 970 116236
rect 1032 116184 1044 116236
rect 1106 116184 1108 116236
rect 946 116182 970 116184
rect 1026 116182 1050 116184
rect 1106 116182 1130 116184
rect 890 116162 1186 116182
rect 890 115150 1186 115170
rect 946 115148 970 115150
rect 1026 115148 1050 115150
rect 1106 115148 1130 115150
rect 968 115096 970 115148
rect 1032 115096 1044 115148
rect 1106 115096 1108 115148
rect 946 115094 970 115096
rect 1026 115094 1050 115096
rect 1106 115094 1130 115096
rect 890 115074 1186 115094
rect 890 114062 1186 114082
rect 946 114060 970 114062
rect 1026 114060 1050 114062
rect 1106 114060 1130 114062
rect 968 114008 970 114060
rect 1032 114008 1044 114060
rect 1106 114008 1108 114060
rect 946 114006 970 114008
rect 1026 114006 1050 114008
rect 1106 114006 1130 114008
rect 890 113986 1186 114006
rect 890 112974 1186 112994
rect 946 112972 970 112974
rect 1026 112972 1050 112974
rect 1106 112972 1130 112974
rect 968 112920 970 112972
rect 1032 112920 1044 112972
rect 1106 112920 1108 112972
rect 946 112918 970 112920
rect 1026 112918 1050 112920
rect 1106 112918 1130 112920
rect 890 112898 1186 112918
rect 890 111886 1186 111906
rect 946 111884 970 111886
rect 1026 111884 1050 111886
rect 1106 111884 1130 111886
rect 968 111832 970 111884
rect 1032 111832 1044 111884
rect 1106 111832 1108 111884
rect 946 111830 970 111832
rect 1026 111830 1050 111832
rect 1106 111830 1130 111832
rect 890 111810 1186 111830
rect 890 110798 1186 110818
rect 946 110796 970 110798
rect 1026 110796 1050 110798
rect 1106 110796 1130 110798
rect 968 110744 970 110796
rect 1032 110744 1044 110796
rect 1106 110744 1108 110796
rect 946 110742 970 110744
rect 1026 110742 1050 110744
rect 1106 110742 1130 110744
rect 890 110722 1186 110742
rect 890 109710 1186 109730
rect 946 109708 970 109710
rect 1026 109708 1050 109710
rect 1106 109708 1130 109710
rect 968 109656 970 109708
rect 1032 109656 1044 109708
rect 1106 109656 1108 109708
rect 946 109654 970 109656
rect 1026 109654 1050 109656
rect 1106 109654 1130 109656
rect 890 109634 1186 109654
rect 890 108622 1186 108642
rect 946 108620 970 108622
rect 1026 108620 1050 108622
rect 1106 108620 1130 108622
rect 968 108568 970 108620
rect 1032 108568 1044 108620
rect 1106 108568 1108 108620
rect 946 108566 970 108568
rect 1026 108566 1050 108568
rect 1106 108566 1130 108568
rect 890 108546 1186 108566
rect 890 107534 1186 107554
rect 946 107532 970 107534
rect 1026 107532 1050 107534
rect 1106 107532 1130 107534
rect 968 107480 970 107532
rect 1032 107480 1044 107532
rect 1106 107480 1108 107532
rect 946 107478 970 107480
rect 1026 107478 1050 107480
rect 1106 107478 1130 107480
rect 890 107458 1186 107478
rect 890 106446 1186 106466
rect 946 106444 970 106446
rect 1026 106444 1050 106446
rect 1106 106444 1130 106446
rect 968 106392 970 106444
rect 1032 106392 1044 106444
rect 1106 106392 1108 106444
rect 946 106390 970 106392
rect 1026 106390 1050 106392
rect 1106 106390 1130 106392
rect 890 106370 1186 106390
rect 890 105358 1186 105378
rect 946 105356 970 105358
rect 1026 105356 1050 105358
rect 1106 105356 1130 105358
rect 968 105304 970 105356
rect 1032 105304 1044 105356
rect 1106 105304 1108 105356
rect 946 105302 970 105304
rect 1026 105302 1050 105304
rect 1106 105302 1130 105304
rect 890 105282 1186 105302
rect 890 104270 1186 104290
rect 946 104268 970 104270
rect 1026 104268 1050 104270
rect 1106 104268 1130 104270
rect 968 104216 970 104268
rect 1032 104216 1044 104268
rect 1106 104216 1108 104268
rect 946 104214 970 104216
rect 1026 104214 1050 104216
rect 1106 104214 1130 104216
rect 890 104194 1186 104214
rect 890 103182 1186 103202
rect 946 103180 970 103182
rect 1026 103180 1050 103182
rect 1106 103180 1130 103182
rect 968 103128 970 103180
rect 1032 103128 1044 103180
rect 1106 103128 1108 103180
rect 946 103126 970 103128
rect 1026 103126 1050 103128
rect 1106 103126 1130 103128
rect 890 103106 1186 103126
rect 890 102094 1186 102114
rect 946 102092 970 102094
rect 1026 102092 1050 102094
rect 1106 102092 1130 102094
rect 968 102040 970 102092
rect 1032 102040 1044 102092
rect 1106 102040 1108 102092
rect 946 102038 970 102040
rect 1026 102038 1050 102040
rect 1106 102038 1130 102040
rect 890 102018 1186 102038
rect 890 101006 1186 101026
rect 946 101004 970 101006
rect 1026 101004 1050 101006
rect 1106 101004 1130 101006
rect 968 100952 970 101004
rect 1032 100952 1044 101004
rect 1106 100952 1108 101004
rect 946 100950 970 100952
rect 1026 100950 1050 100952
rect 1106 100950 1130 100952
rect 890 100930 1186 100950
rect 890 99918 1186 99938
rect 946 99916 970 99918
rect 1026 99916 1050 99918
rect 1106 99916 1130 99918
rect 968 99864 970 99916
rect 1032 99864 1044 99916
rect 1106 99864 1108 99916
rect 946 99862 970 99864
rect 1026 99862 1050 99864
rect 1106 99862 1130 99864
rect 890 99842 1186 99862
rect 890 98830 1186 98850
rect 946 98828 970 98830
rect 1026 98828 1050 98830
rect 1106 98828 1130 98830
rect 968 98776 970 98828
rect 1032 98776 1044 98828
rect 1106 98776 1108 98828
rect 946 98774 970 98776
rect 1026 98774 1050 98776
rect 1106 98774 1130 98776
rect 890 98754 1186 98774
rect 890 97742 1186 97762
rect 946 97740 970 97742
rect 1026 97740 1050 97742
rect 1106 97740 1130 97742
rect 968 97688 970 97740
rect 1032 97688 1044 97740
rect 1106 97688 1108 97740
rect 946 97686 970 97688
rect 1026 97686 1050 97688
rect 1106 97686 1130 97688
rect 890 97666 1186 97686
rect 890 96654 1186 96674
rect 946 96652 970 96654
rect 1026 96652 1050 96654
rect 1106 96652 1130 96654
rect 968 96600 970 96652
rect 1032 96600 1044 96652
rect 1106 96600 1108 96652
rect 946 96598 970 96600
rect 1026 96598 1050 96600
rect 1106 96598 1130 96600
rect 890 96578 1186 96598
rect 890 95566 1186 95586
rect 946 95564 970 95566
rect 1026 95564 1050 95566
rect 1106 95564 1130 95566
rect 968 95512 970 95564
rect 1032 95512 1044 95564
rect 1106 95512 1108 95564
rect 946 95510 970 95512
rect 1026 95510 1050 95512
rect 1106 95510 1130 95512
rect 890 95490 1186 95510
rect 890 94478 1186 94498
rect 946 94476 970 94478
rect 1026 94476 1050 94478
rect 1106 94476 1130 94478
rect 968 94424 970 94476
rect 1032 94424 1044 94476
rect 1106 94424 1108 94476
rect 946 94422 970 94424
rect 1026 94422 1050 94424
rect 1106 94422 1130 94424
rect 890 94402 1186 94422
rect 890 93390 1186 93410
rect 946 93388 970 93390
rect 1026 93388 1050 93390
rect 1106 93388 1130 93390
rect 968 93336 970 93388
rect 1032 93336 1044 93388
rect 1106 93336 1108 93388
rect 946 93334 970 93336
rect 1026 93334 1050 93336
rect 1106 93334 1130 93336
rect 890 93314 1186 93334
rect 890 92302 1186 92322
rect 946 92300 970 92302
rect 1026 92300 1050 92302
rect 1106 92300 1130 92302
rect 968 92248 970 92300
rect 1032 92248 1044 92300
rect 1106 92248 1108 92300
rect 946 92246 970 92248
rect 1026 92246 1050 92248
rect 1106 92246 1130 92248
rect 890 92226 1186 92246
rect 890 91214 1186 91234
rect 946 91212 970 91214
rect 1026 91212 1050 91214
rect 1106 91212 1130 91214
rect 968 91160 970 91212
rect 1032 91160 1044 91212
rect 1106 91160 1108 91212
rect 946 91158 970 91160
rect 1026 91158 1050 91160
rect 1106 91158 1130 91160
rect 890 91138 1186 91158
rect 890 90126 1186 90146
rect 946 90124 970 90126
rect 1026 90124 1050 90126
rect 1106 90124 1130 90126
rect 968 90072 970 90124
rect 1032 90072 1044 90124
rect 1106 90072 1108 90124
rect 946 90070 970 90072
rect 1026 90070 1050 90072
rect 1106 90070 1130 90072
rect 890 90050 1186 90070
rect 890 89038 1186 89058
rect 946 89036 970 89038
rect 1026 89036 1050 89038
rect 1106 89036 1130 89038
rect 968 88984 970 89036
rect 1032 88984 1044 89036
rect 1106 88984 1108 89036
rect 946 88982 970 88984
rect 1026 88982 1050 88984
rect 1106 88982 1130 88984
rect 890 88962 1186 88982
rect 890 87950 1186 87970
rect 946 87948 970 87950
rect 1026 87948 1050 87950
rect 1106 87948 1130 87950
rect 968 87896 970 87948
rect 1032 87896 1044 87948
rect 1106 87896 1108 87948
rect 946 87894 970 87896
rect 1026 87894 1050 87896
rect 1106 87894 1130 87896
rect 890 87874 1186 87894
rect 890 86862 1186 86882
rect 946 86860 970 86862
rect 1026 86860 1050 86862
rect 1106 86860 1130 86862
rect 968 86808 970 86860
rect 1032 86808 1044 86860
rect 1106 86808 1108 86860
rect 946 86806 970 86808
rect 1026 86806 1050 86808
rect 1106 86806 1130 86808
rect 890 86786 1186 86806
rect 890 85774 1186 85794
rect 946 85772 970 85774
rect 1026 85772 1050 85774
rect 1106 85772 1130 85774
rect 968 85720 970 85772
rect 1032 85720 1044 85772
rect 1106 85720 1108 85772
rect 946 85718 970 85720
rect 1026 85718 1050 85720
rect 1106 85718 1130 85720
rect 890 85698 1186 85718
rect 890 84686 1186 84706
rect 946 84684 970 84686
rect 1026 84684 1050 84686
rect 1106 84684 1130 84686
rect 968 84632 970 84684
rect 1032 84632 1044 84684
rect 1106 84632 1108 84684
rect 946 84630 970 84632
rect 1026 84630 1050 84632
rect 1106 84630 1130 84632
rect 890 84610 1186 84630
rect 890 83598 1186 83618
rect 946 83596 970 83598
rect 1026 83596 1050 83598
rect 1106 83596 1130 83598
rect 968 83544 970 83596
rect 1032 83544 1044 83596
rect 1106 83544 1108 83596
rect 946 83542 970 83544
rect 1026 83542 1050 83544
rect 1106 83542 1130 83544
rect 890 83522 1186 83542
rect 890 82510 1186 82530
rect 946 82508 970 82510
rect 1026 82508 1050 82510
rect 1106 82508 1130 82510
rect 968 82456 970 82508
rect 1032 82456 1044 82508
rect 1106 82456 1108 82508
rect 946 82454 970 82456
rect 1026 82454 1050 82456
rect 1106 82454 1130 82456
rect 890 82434 1186 82454
rect 890 81422 1186 81442
rect 946 81420 970 81422
rect 1026 81420 1050 81422
rect 1106 81420 1130 81422
rect 968 81368 970 81420
rect 1032 81368 1044 81420
rect 1106 81368 1108 81420
rect 946 81366 970 81368
rect 1026 81366 1050 81368
rect 1106 81366 1130 81368
rect 890 81346 1186 81366
rect 890 80334 1186 80354
rect 946 80332 970 80334
rect 1026 80332 1050 80334
rect 1106 80332 1130 80334
rect 968 80280 970 80332
rect 1032 80280 1044 80332
rect 1106 80280 1108 80332
rect 946 80278 970 80280
rect 1026 80278 1050 80280
rect 1106 80278 1130 80280
rect 890 80258 1186 80278
rect 890 79246 1186 79266
rect 946 79244 970 79246
rect 1026 79244 1050 79246
rect 1106 79244 1130 79246
rect 968 79192 970 79244
rect 1032 79192 1044 79244
rect 1106 79192 1108 79244
rect 946 79190 970 79192
rect 1026 79190 1050 79192
rect 1106 79190 1130 79192
rect 890 79170 1186 79190
rect 890 78158 1186 78178
rect 946 78156 970 78158
rect 1026 78156 1050 78158
rect 1106 78156 1130 78158
rect 968 78104 970 78156
rect 1032 78104 1044 78156
rect 1106 78104 1108 78156
rect 946 78102 970 78104
rect 1026 78102 1050 78104
rect 1106 78102 1130 78104
rect 890 78082 1186 78102
rect 890 77070 1186 77090
rect 946 77068 970 77070
rect 1026 77068 1050 77070
rect 1106 77068 1130 77070
rect 968 77016 970 77068
rect 1032 77016 1044 77068
rect 1106 77016 1108 77068
rect 946 77014 970 77016
rect 1026 77014 1050 77016
rect 1106 77014 1130 77016
rect 890 76994 1186 77014
rect 890 75982 1186 76002
rect 946 75980 970 75982
rect 1026 75980 1050 75982
rect 1106 75980 1130 75982
rect 968 75928 970 75980
rect 1032 75928 1044 75980
rect 1106 75928 1108 75980
rect 946 75926 970 75928
rect 1026 75926 1050 75928
rect 1106 75926 1130 75928
rect 890 75906 1186 75926
rect 890 74894 1186 74914
rect 946 74892 970 74894
rect 1026 74892 1050 74894
rect 1106 74892 1130 74894
rect 968 74840 970 74892
rect 1032 74840 1044 74892
rect 1106 74840 1108 74892
rect 946 74838 970 74840
rect 1026 74838 1050 74840
rect 1106 74838 1130 74840
rect 890 74818 1186 74838
rect 890 73806 1186 73826
rect 946 73804 970 73806
rect 1026 73804 1050 73806
rect 1106 73804 1130 73806
rect 968 73752 970 73804
rect 1032 73752 1044 73804
rect 1106 73752 1108 73804
rect 946 73750 970 73752
rect 1026 73750 1050 73752
rect 1106 73750 1130 73752
rect 890 73730 1186 73750
rect 890 72718 1186 72738
rect 946 72716 970 72718
rect 1026 72716 1050 72718
rect 1106 72716 1130 72718
rect 968 72664 970 72716
rect 1032 72664 1044 72716
rect 1106 72664 1108 72716
rect 946 72662 970 72664
rect 1026 72662 1050 72664
rect 1106 72662 1130 72664
rect 890 72642 1186 72662
rect 890 71630 1186 71650
rect 946 71628 970 71630
rect 1026 71628 1050 71630
rect 1106 71628 1130 71630
rect 968 71576 970 71628
rect 1032 71576 1044 71628
rect 1106 71576 1108 71628
rect 946 71574 970 71576
rect 1026 71574 1050 71576
rect 1106 71574 1130 71576
rect 890 71554 1186 71574
rect 890 70542 1186 70562
rect 946 70540 970 70542
rect 1026 70540 1050 70542
rect 1106 70540 1130 70542
rect 968 70488 970 70540
rect 1032 70488 1044 70540
rect 1106 70488 1108 70540
rect 946 70486 970 70488
rect 1026 70486 1050 70488
rect 1106 70486 1130 70488
rect 890 70466 1186 70486
rect 890 69454 1186 69474
rect 946 69452 970 69454
rect 1026 69452 1050 69454
rect 1106 69452 1130 69454
rect 968 69400 970 69452
rect 1032 69400 1044 69452
rect 1106 69400 1108 69452
rect 946 69398 970 69400
rect 1026 69398 1050 69400
rect 1106 69398 1130 69400
rect 890 69378 1186 69398
rect 890 68366 1186 68386
rect 946 68364 970 68366
rect 1026 68364 1050 68366
rect 1106 68364 1130 68366
rect 968 68312 970 68364
rect 1032 68312 1044 68364
rect 1106 68312 1108 68364
rect 946 68310 970 68312
rect 1026 68310 1050 68312
rect 1106 68310 1130 68312
rect 890 68290 1186 68310
rect 890 67278 1186 67298
rect 946 67276 970 67278
rect 1026 67276 1050 67278
rect 1106 67276 1130 67278
rect 968 67224 970 67276
rect 1032 67224 1044 67276
rect 1106 67224 1108 67276
rect 946 67222 970 67224
rect 1026 67222 1050 67224
rect 1106 67222 1130 67224
rect 890 67202 1186 67222
rect 890 66190 1186 66210
rect 946 66188 970 66190
rect 1026 66188 1050 66190
rect 1106 66188 1130 66190
rect 968 66136 970 66188
rect 1032 66136 1044 66188
rect 1106 66136 1108 66188
rect 946 66134 970 66136
rect 1026 66134 1050 66136
rect 1106 66134 1130 66136
rect 890 66114 1186 66134
rect 890 65102 1186 65122
rect 946 65100 970 65102
rect 1026 65100 1050 65102
rect 1106 65100 1130 65102
rect 968 65048 970 65100
rect 1032 65048 1044 65100
rect 1106 65048 1108 65100
rect 946 65046 970 65048
rect 1026 65046 1050 65048
rect 1106 65046 1130 65048
rect 890 65026 1186 65046
rect 890 64014 1186 64034
rect 946 64012 970 64014
rect 1026 64012 1050 64014
rect 1106 64012 1130 64014
rect 968 63960 970 64012
rect 1032 63960 1044 64012
rect 1106 63960 1108 64012
rect 946 63958 970 63960
rect 1026 63958 1050 63960
rect 1106 63958 1130 63960
rect 890 63938 1186 63958
rect 890 62926 1186 62946
rect 946 62924 970 62926
rect 1026 62924 1050 62926
rect 1106 62924 1130 62926
rect 968 62872 970 62924
rect 1032 62872 1044 62924
rect 1106 62872 1108 62924
rect 946 62870 970 62872
rect 1026 62870 1050 62872
rect 1106 62870 1130 62872
rect 890 62850 1186 62870
rect 890 61838 1186 61858
rect 946 61836 970 61838
rect 1026 61836 1050 61838
rect 1106 61836 1130 61838
rect 968 61784 970 61836
rect 1032 61784 1044 61836
rect 1106 61784 1108 61836
rect 946 61782 970 61784
rect 1026 61782 1050 61784
rect 1106 61782 1130 61784
rect 890 61762 1186 61782
rect 890 60750 1186 60770
rect 946 60748 970 60750
rect 1026 60748 1050 60750
rect 1106 60748 1130 60750
rect 968 60696 970 60748
rect 1032 60696 1044 60748
rect 1106 60696 1108 60748
rect 946 60694 970 60696
rect 1026 60694 1050 60696
rect 1106 60694 1130 60696
rect 890 60674 1186 60694
rect 890 59662 1186 59682
rect 946 59660 970 59662
rect 1026 59660 1050 59662
rect 1106 59660 1130 59662
rect 968 59608 970 59660
rect 1032 59608 1044 59660
rect 1106 59608 1108 59660
rect 946 59606 970 59608
rect 1026 59606 1050 59608
rect 1106 59606 1130 59608
rect 890 59586 1186 59606
rect 890 58574 1186 58594
rect 946 58572 970 58574
rect 1026 58572 1050 58574
rect 1106 58572 1130 58574
rect 968 58520 970 58572
rect 1032 58520 1044 58572
rect 1106 58520 1108 58572
rect 946 58518 970 58520
rect 1026 58518 1050 58520
rect 1106 58518 1130 58520
rect 890 58498 1186 58518
rect 890 57486 1186 57506
rect 946 57484 970 57486
rect 1026 57484 1050 57486
rect 1106 57484 1130 57486
rect 968 57432 970 57484
rect 1032 57432 1044 57484
rect 1106 57432 1108 57484
rect 946 57430 970 57432
rect 1026 57430 1050 57432
rect 1106 57430 1130 57432
rect 890 57410 1186 57430
rect 890 56398 1186 56418
rect 946 56396 970 56398
rect 1026 56396 1050 56398
rect 1106 56396 1130 56398
rect 968 56344 970 56396
rect 1032 56344 1044 56396
rect 1106 56344 1108 56396
rect 946 56342 970 56344
rect 1026 56342 1050 56344
rect 1106 56342 1130 56344
rect 890 56322 1186 56342
rect 890 55310 1186 55330
rect 946 55308 970 55310
rect 1026 55308 1050 55310
rect 1106 55308 1130 55310
rect 968 55256 970 55308
rect 1032 55256 1044 55308
rect 1106 55256 1108 55308
rect 946 55254 970 55256
rect 1026 55254 1050 55256
rect 1106 55254 1130 55256
rect 890 55234 1186 55254
rect 890 54222 1186 54242
rect 946 54220 970 54222
rect 1026 54220 1050 54222
rect 1106 54220 1130 54222
rect 968 54168 970 54220
rect 1032 54168 1044 54220
rect 1106 54168 1108 54220
rect 946 54166 970 54168
rect 1026 54166 1050 54168
rect 1106 54166 1130 54168
rect 890 54146 1186 54166
rect 890 53134 1186 53154
rect 946 53132 970 53134
rect 1026 53132 1050 53134
rect 1106 53132 1130 53134
rect 968 53080 970 53132
rect 1032 53080 1044 53132
rect 1106 53080 1108 53132
rect 946 53078 970 53080
rect 1026 53078 1050 53080
rect 1106 53078 1130 53080
rect 890 53058 1186 53078
rect 890 52046 1186 52066
rect 946 52044 970 52046
rect 1026 52044 1050 52046
rect 1106 52044 1130 52046
rect 968 51992 970 52044
rect 1032 51992 1044 52044
rect 1106 51992 1108 52044
rect 946 51990 970 51992
rect 1026 51990 1050 51992
rect 1106 51990 1130 51992
rect 890 51970 1186 51990
rect 890 50958 1186 50978
rect 946 50956 970 50958
rect 1026 50956 1050 50958
rect 1106 50956 1130 50958
rect 968 50904 970 50956
rect 1032 50904 1044 50956
rect 1106 50904 1108 50956
rect 946 50902 970 50904
rect 1026 50902 1050 50904
rect 1106 50902 1130 50904
rect 890 50882 1186 50902
rect 890 49870 1186 49890
rect 946 49868 970 49870
rect 1026 49868 1050 49870
rect 1106 49868 1130 49870
rect 968 49816 970 49868
rect 1032 49816 1044 49868
rect 1106 49816 1108 49868
rect 946 49814 970 49816
rect 1026 49814 1050 49816
rect 1106 49814 1130 49816
rect 890 49794 1186 49814
rect 890 48782 1186 48802
rect 946 48780 970 48782
rect 1026 48780 1050 48782
rect 1106 48780 1130 48782
rect 968 48728 970 48780
rect 1032 48728 1044 48780
rect 1106 48728 1108 48780
rect 946 48726 970 48728
rect 1026 48726 1050 48728
rect 1106 48726 1130 48728
rect 890 48706 1186 48726
rect 890 47694 1186 47714
rect 946 47692 970 47694
rect 1026 47692 1050 47694
rect 1106 47692 1130 47694
rect 968 47640 970 47692
rect 1032 47640 1044 47692
rect 1106 47640 1108 47692
rect 946 47638 970 47640
rect 1026 47638 1050 47640
rect 1106 47638 1130 47640
rect 890 47618 1186 47638
rect 890 46606 1186 46626
rect 946 46604 970 46606
rect 1026 46604 1050 46606
rect 1106 46604 1130 46606
rect 968 46552 970 46604
rect 1032 46552 1044 46604
rect 1106 46552 1108 46604
rect 946 46550 970 46552
rect 1026 46550 1050 46552
rect 1106 46550 1130 46552
rect 890 46530 1186 46550
rect 890 45518 1186 45538
rect 946 45516 970 45518
rect 1026 45516 1050 45518
rect 1106 45516 1130 45518
rect 968 45464 970 45516
rect 1032 45464 1044 45516
rect 1106 45464 1108 45516
rect 946 45462 970 45464
rect 1026 45462 1050 45464
rect 1106 45462 1130 45464
rect 890 45442 1186 45462
rect 890 44430 1186 44450
rect 946 44428 970 44430
rect 1026 44428 1050 44430
rect 1106 44428 1130 44430
rect 968 44376 970 44428
rect 1032 44376 1044 44428
rect 1106 44376 1108 44428
rect 946 44374 970 44376
rect 1026 44374 1050 44376
rect 1106 44374 1130 44376
rect 890 44354 1186 44374
rect 890 43342 1186 43362
rect 946 43340 970 43342
rect 1026 43340 1050 43342
rect 1106 43340 1130 43342
rect 968 43288 970 43340
rect 1032 43288 1044 43340
rect 1106 43288 1108 43340
rect 946 43286 970 43288
rect 1026 43286 1050 43288
rect 1106 43286 1130 43288
rect 890 43266 1186 43286
rect 890 42254 1186 42274
rect 946 42252 970 42254
rect 1026 42252 1050 42254
rect 1106 42252 1130 42254
rect 968 42200 970 42252
rect 1032 42200 1044 42252
rect 1106 42200 1108 42252
rect 946 42198 970 42200
rect 1026 42198 1050 42200
rect 1106 42198 1130 42200
rect 890 42178 1186 42198
rect 890 41166 1186 41186
rect 946 41164 970 41166
rect 1026 41164 1050 41166
rect 1106 41164 1130 41166
rect 968 41112 970 41164
rect 1032 41112 1044 41164
rect 1106 41112 1108 41164
rect 946 41110 970 41112
rect 1026 41110 1050 41112
rect 1106 41110 1130 41112
rect 890 41090 1186 41110
rect 890 40078 1186 40098
rect 946 40076 970 40078
rect 1026 40076 1050 40078
rect 1106 40076 1130 40078
rect 968 40024 970 40076
rect 1032 40024 1044 40076
rect 1106 40024 1108 40076
rect 946 40022 970 40024
rect 1026 40022 1050 40024
rect 1106 40022 1130 40024
rect 890 40002 1186 40022
rect 890 38990 1186 39010
rect 946 38988 970 38990
rect 1026 38988 1050 38990
rect 1106 38988 1130 38990
rect 968 38936 970 38988
rect 1032 38936 1044 38988
rect 1106 38936 1108 38988
rect 946 38934 970 38936
rect 1026 38934 1050 38936
rect 1106 38934 1130 38936
rect 890 38914 1186 38934
rect 890 37902 1186 37922
rect 946 37900 970 37902
rect 1026 37900 1050 37902
rect 1106 37900 1130 37902
rect 968 37848 970 37900
rect 1032 37848 1044 37900
rect 1106 37848 1108 37900
rect 946 37846 970 37848
rect 1026 37846 1050 37848
rect 1106 37846 1130 37848
rect 890 37826 1186 37846
rect 890 36814 1186 36834
rect 946 36812 970 36814
rect 1026 36812 1050 36814
rect 1106 36812 1130 36814
rect 968 36760 970 36812
rect 1032 36760 1044 36812
rect 1106 36760 1108 36812
rect 946 36758 970 36760
rect 1026 36758 1050 36760
rect 1106 36758 1130 36760
rect 890 36738 1186 36758
rect 890 35726 1186 35746
rect 946 35724 970 35726
rect 1026 35724 1050 35726
rect 1106 35724 1130 35726
rect 968 35672 970 35724
rect 1032 35672 1044 35724
rect 1106 35672 1108 35724
rect 946 35670 970 35672
rect 1026 35670 1050 35672
rect 1106 35670 1130 35672
rect 890 35650 1186 35670
rect 890 34638 1186 34658
rect 946 34636 970 34638
rect 1026 34636 1050 34638
rect 1106 34636 1130 34638
rect 968 34584 970 34636
rect 1032 34584 1044 34636
rect 1106 34584 1108 34636
rect 946 34582 970 34584
rect 1026 34582 1050 34584
rect 1106 34582 1130 34584
rect 890 34562 1186 34582
rect 890 33550 1186 33570
rect 946 33548 970 33550
rect 1026 33548 1050 33550
rect 1106 33548 1130 33550
rect 968 33496 970 33548
rect 1032 33496 1044 33548
rect 1106 33496 1108 33548
rect 946 33494 970 33496
rect 1026 33494 1050 33496
rect 1106 33494 1130 33496
rect 890 33474 1186 33494
rect 890 32462 1186 32482
rect 946 32460 970 32462
rect 1026 32460 1050 32462
rect 1106 32460 1130 32462
rect 968 32408 970 32460
rect 1032 32408 1044 32460
rect 1106 32408 1108 32460
rect 946 32406 970 32408
rect 1026 32406 1050 32408
rect 1106 32406 1130 32408
rect 890 32386 1186 32406
rect 890 31374 1186 31394
rect 946 31372 970 31374
rect 1026 31372 1050 31374
rect 1106 31372 1130 31374
rect 968 31320 970 31372
rect 1032 31320 1044 31372
rect 1106 31320 1108 31372
rect 946 31318 970 31320
rect 1026 31318 1050 31320
rect 1106 31318 1130 31320
rect 890 31298 1186 31318
rect 890 30286 1186 30306
rect 946 30284 970 30286
rect 1026 30284 1050 30286
rect 1106 30284 1130 30286
rect 968 30232 970 30284
rect 1032 30232 1044 30284
rect 1106 30232 1108 30284
rect 946 30230 970 30232
rect 1026 30230 1050 30232
rect 1106 30230 1130 30232
rect 890 30210 1186 30230
rect 890 29198 1186 29218
rect 946 29196 970 29198
rect 1026 29196 1050 29198
rect 1106 29196 1130 29198
rect 968 29144 970 29196
rect 1032 29144 1044 29196
rect 1106 29144 1108 29196
rect 946 29142 970 29144
rect 1026 29142 1050 29144
rect 1106 29142 1130 29144
rect 890 29122 1186 29142
rect 890 28110 1186 28130
rect 946 28108 970 28110
rect 1026 28108 1050 28110
rect 1106 28108 1130 28110
rect 968 28056 970 28108
rect 1032 28056 1044 28108
rect 1106 28056 1108 28108
rect 946 28054 970 28056
rect 1026 28054 1050 28056
rect 1106 28054 1130 28056
rect 890 28034 1186 28054
rect 890 27022 1186 27042
rect 946 27020 970 27022
rect 1026 27020 1050 27022
rect 1106 27020 1130 27022
rect 968 26968 970 27020
rect 1032 26968 1044 27020
rect 1106 26968 1108 27020
rect 946 26966 970 26968
rect 1026 26966 1050 26968
rect 1106 26966 1130 26968
rect 890 26946 1186 26966
rect 890 25934 1186 25954
rect 946 25932 970 25934
rect 1026 25932 1050 25934
rect 1106 25932 1130 25934
rect 968 25880 970 25932
rect 1032 25880 1044 25932
rect 1106 25880 1108 25932
rect 946 25878 970 25880
rect 1026 25878 1050 25880
rect 1106 25878 1130 25880
rect 890 25858 1186 25878
rect 890 24846 1186 24866
rect 946 24844 970 24846
rect 1026 24844 1050 24846
rect 1106 24844 1130 24846
rect 968 24792 970 24844
rect 1032 24792 1044 24844
rect 1106 24792 1108 24844
rect 946 24790 970 24792
rect 1026 24790 1050 24792
rect 1106 24790 1130 24792
rect 890 24770 1186 24790
rect 890 23758 1186 23778
rect 946 23756 970 23758
rect 1026 23756 1050 23758
rect 1106 23756 1130 23758
rect 968 23704 970 23756
rect 1032 23704 1044 23756
rect 1106 23704 1108 23756
rect 946 23702 970 23704
rect 1026 23702 1050 23704
rect 1106 23702 1130 23704
rect 890 23682 1186 23702
rect 890 22670 1186 22690
rect 946 22668 970 22670
rect 1026 22668 1050 22670
rect 1106 22668 1130 22670
rect 968 22616 970 22668
rect 1032 22616 1044 22668
rect 1106 22616 1108 22668
rect 946 22614 970 22616
rect 1026 22614 1050 22616
rect 1106 22614 1130 22616
rect 890 22594 1186 22614
rect 890 21582 1186 21602
rect 946 21580 970 21582
rect 1026 21580 1050 21582
rect 1106 21580 1130 21582
rect 968 21528 970 21580
rect 1032 21528 1044 21580
rect 1106 21528 1108 21580
rect 946 21526 970 21528
rect 1026 21526 1050 21528
rect 1106 21526 1130 21528
rect 890 21506 1186 21526
rect 890 20494 1186 20514
rect 946 20492 970 20494
rect 1026 20492 1050 20494
rect 1106 20492 1130 20494
rect 968 20440 970 20492
rect 1032 20440 1044 20492
rect 1106 20440 1108 20492
rect 946 20438 970 20440
rect 1026 20438 1050 20440
rect 1106 20438 1130 20440
rect 890 20418 1186 20438
rect 890 19406 1186 19426
rect 946 19404 970 19406
rect 1026 19404 1050 19406
rect 1106 19404 1130 19406
rect 968 19352 970 19404
rect 1032 19352 1044 19404
rect 1106 19352 1108 19404
rect 946 19350 970 19352
rect 1026 19350 1050 19352
rect 1106 19350 1130 19352
rect 890 19330 1186 19350
rect 890 18318 1186 18338
rect 946 18316 970 18318
rect 1026 18316 1050 18318
rect 1106 18316 1130 18318
rect 968 18264 970 18316
rect 1032 18264 1044 18316
rect 1106 18264 1108 18316
rect 946 18262 970 18264
rect 1026 18262 1050 18264
rect 1106 18262 1130 18264
rect 890 18242 1186 18262
rect 890 17230 1186 17250
rect 946 17228 970 17230
rect 1026 17228 1050 17230
rect 1106 17228 1130 17230
rect 968 17176 970 17228
rect 1032 17176 1044 17228
rect 1106 17176 1108 17228
rect 946 17174 970 17176
rect 1026 17174 1050 17176
rect 1106 17174 1130 17176
rect 890 17154 1186 17174
rect 890 16142 1186 16162
rect 946 16140 970 16142
rect 1026 16140 1050 16142
rect 1106 16140 1130 16142
rect 968 16088 970 16140
rect 1032 16088 1044 16140
rect 1106 16088 1108 16140
rect 946 16086 970 16088
rect 1026 16086 1050 16088
rect 1106 16086 1130 16088
rect 890 16066 1186 16086
rect 890 15054 1186 15074
rect 946 15052 970 15054
rect 1026 15052 1050 15054
rect 1106 15052 1130 15054
rect 968 15000 970 15052
rect 1032 15000 1044 15052
rect 1106 15000 1108 15052
rect 946 14998 970 15000
rect 1026 14998 1050 15000
rect 1106 14998 1130 15000
rect 890 14978 1186 14998
rect 890 13966 1186 13986
rect 946 13964 970 13966
rect 1026 13964 1050 13966
rect 1106 13964 1130 13966
rect 968 13912 970 13964
rect 1032 13912 1044 13964
rect 1106 13912 1108 13964
rect 946 13910 970 13912
rect 1026 13910 1050 13912
rect 1106 13910 1130 13912
rect 890 13890 1186 13910
rect 890 12878 1186 12898
rect 946 12876 970 12878
rect 1026 12876 1050 12878
rect 1106 12876 1130 12878
rect 968 12824 970 12876
rect 1032 12824 1044 12876
rect 1106 12824 1108 12876
rect 946 12822 970 12824
rect 1026 12822 1050 12824
rect 1106 12822 1130 12824
rect 890 12802 1186 12822
rect 890 11790 1186 11810
rect 946 11788 970 11790
rect 1026 11788 1050 11790
rect 1106 11788 1130 11790
rect 968 11736 970 11788
rect 1032 11736 1044 11788
rect 1106 11736 1108 11788
rect 946 11734 970 11736
rect 1026 11734 1050 11736
rect 1106 11734 1130 11736
rect 890 11714 1186 11734
rect 890 10702 1186 10722
rect 946 10700 970 10702
rect 1026 10700 1050 10702
rect 1106 10700 1130 10702
rect 968 10648 970 10700
rect 1032 10648 1044 10700
rect 1106 10648 1108 10700
rect 946 10646 970 10648
rect 1026 10646 1050 10648
rect 1106 10646 1130 10648
rect 890 10626 1186 10646
rect 890 9614 1186 9634
rect 946 9612 970 9614
rect 1026 9612 1050 9614
rect 1106 9612 1130 9614
rect 968 9560 970 9612
rect 1032 9560 1044 9612
rect 1106 9560 1108 9612
rect 946 9558 970 9560
rect 1026 9558 1050 9560
rect 1106 9558 1130 9560
rect 890 9538 1186 9558
rect 890 8526 1186 8546
rect 946 8524 970 8526
rect 1026 8524 1050 8526
rect 1106 8524 1130 8526
rect 968 8472 970 8524
rect 1032 8472 1044 8524
rect 1106 8472 1108 8524
rect 946 8470 970 8472
rect 1026 8470 1050 8472
rect 1106 8470 1130 8472
rect 890 8450 1186 8470
rect 890 7438 1186 7458
rect 946 7436 970 7438
rect 1026 7436 1050 7438
rect 1106 7436 1130 7438
rect 968 7384 970 7436
rect 1032 7384 1044 7436
rect 1106 7384 1108 7436
rect 946 7382 970 7384
rect 1026 7382 1050 7384
rect 1106 7382 1130 7384
rect 890 7362 1186 7382
rect 890 6350 1186 6370
rect 946 6348 970 6350
rect 1026 6348 1050 6350
rect 1106 6348 1130 6350
rect 968 6296 970 6348
rect 1032 6296 1044 6348
rect 1106 6296 1108 6348
rect 946 6294 970 6296
rect 1026 6294 1050 6296
rect 1106 6294 1130 6296
rect 890 6274 1186 6294
rect 890 5262 1186 5282
rect 946 5260 970 5262
rect 1026 5260 1050 5262
rect 1106 5260 1130 5262
rect 968 5208 970 5260
rect 1032 5208 1044 5260
rect 1106 5208 1108 5260
rect 946 5206 970 5208
rect 1026 5206 1050 5208
rect 1106 5206 1130 5208
rect 890 5186 1186 5206
rect 1266 4908 1294 187233
rect 1358 97372 1386 187816
rect 1436 186754 1492 186763
rect 1436 186689 1492 186698
rect 1346 97366 1398 97372
rect 1346 97308 1398 97314
rect 1358 97032 1386 97308
rect 1346 97026 1398 97032
rect 1346 96968 1398 96974
rect 1358 5044 1386 96968
rect 1450 5180 1478 186689
rect 1990 186582 2042 186588
rect 1990 186524 2042 186530
rect 1896 171114 1952 171123
rect 1896 171049 1952 171058
rect 1910 162176 1938 171049
rect 1898 162170 1950 162176
rect 1898 162112 1950 162118
rect 1898 162034 1950 162040
rect 1898 161976 1950 161982
rect 1910 153132 1938 161976
rect 1898 153126 1950 153132
rect 1898 153068 1950 153074
rect 1898 145986 1950 145992
rect 1898 145928 1950 145934
rect 1910 141572 1938 145928
rect 1898 141566 1950 141572
rect 1898 141508 1950 141514
rect 1898 133746 1950 133752
rect 1898 133688 1950 133694
rect 1910 124776 1938 133688
rect 1898 124770 1950 124776
rect 1898 124712 1950 124718
rect 1898 98386 1950 98392
rect 1898 98328 1950 98334
rect 1714 96754 1766 96760
rect 1714 96696 1766 96702
rect 1726 96556 1754 96696
rect 1714 96550 1766 96556
rect 1714 96492 1766 96498
rect 1714 95870 1766 95876
rect 1714 95812 1766 95818
rect 1622 94782 1674 94788
rect 1622 94724 1674 94730
rect 1450 5152 1570 5180
rect 1358 5016 1478 5044
rect 1266 4880 1386 4908
rect 890 4174 1186 4194
rect 946 4172 970 4174
rect 1026 4172 1050 4174
rect 1106 4172 1130 4174
rect 968 4120 970 4172
rect 1032 4120 1044 4172
rect 1106 4120 1108 4172
rect 946 4118 970 4120
rect 1026 4118 1050 4120
rect 1106 4118 1130 4120
rect 890 4098 1186 4118
rect 1358 3192 1386 4880
rect 1346 3186 1398 3192
rect 1346 3128 1398 3134
rect 890 3086 1186 3106
rect 946 3084 970 3086
rect 1026 3084 1050 3086
rect 1106 3084 1130 3086
rect 968 3032 970 3084
rect 1032 3032 1044 3084
rect 1106 3032 1108 3084
rect 946 3030 970 3032
rect 1026 3030 1050 3032
rect 1106 3030 1130 3032
rect 890 3010 1186 3030
rect 1358 2891 1386 3128
rect 1344 2882 1400 2891
rect 1344 2817 1400 2826
rect 978 2642 1030 2648
rect 978 2584 1030 2590
rect 990 2444 1018 2584
rect 1450 2444 1478 5016
rect 1542 4280 1570 5152
rect 1530 4274 1582 4280
rect 1530 4216 1582 4222
rect 978 2438 1030 2444
rect 978 2380 1030 2386
rect 1438 2438 1490 2444
rect 1438 2380 1490 2386
rect 1634 2188 1662 94724
rect 1726 3260 1754 95812
rect 1910 94788 1938 98328
rect 1898 94782 1950 94788
rect 1898 94724 1950 94730
rect 2002 4076 2030 186524
rect 2094 97576 2122 188088
rect 2174 180190 2226 180196
rect 2174 180132 2226 180138
rect 2186 173668 2214 180132
rect 2174 173662 2226 173668
rect 2174 173604 2226 173610
rect 2266 173594 2318 173600
rect 2266 173536 2318 173542
rect 2278 171123 2306 173536
rect 2264 171114 2320 171123
rect 2264 171049 2320 171058
rect 2266 162170 2318 162176
rect 2266 162112 2318 162118
rect 2278 162040 2306 162112
rect 2266 162034 2318 162040
rect 2266 161976 2318 161982
rect 2266 153126 2318 153132
rect 2266 153068 2318 153074
rect 2278 145992 2306 153068
rect 2266 145986 2318 145992
rect 2266 145928 2318 145934
rect 2174 141566 2226 141572
rect 2174 141508 2226 141514
rect 2186 138324 2214 141508
rect 2186 138296 2306 138324
rect 2278 133752 2306 138296
rect 2266 133746 2318 133752
rect 2266 133688 2318 133694
rect 2174 124770 2226 124776
rect 2172 124738 2174 124747
rect 2226 124738 2228 124747
rect 2172 124673 2228 124682
rect 2172 108146 2228 108155
rect 2172 108081 2228 108090
rect 2082 97570 2134 97576
rect 2082 97512 2134 97518
rect 2094 97304 2122 97512
rect 2082 97298 2134 97304
rect 2082 97240 2134 97246
rect 1990 4070 2042 4076
rect 1990 4012 2042 4018
rect 2094 3464 2122 97240
rect 2186 96420 2214 108081
rect 2266 97842 2318 97848
rect 2266 97784 2318 97790
rect 2174 96414 2226 96420
rect 2174 96356 2226 96362
rect 2174 96278 2226 96284
rect 2174 96220 2226 96226
rect 2082 3458 2134 3464
rect 2082 3400 2134 3406
rect 1804 3290 1860 3299
rect 1714 3254 1766 3260
rect 1804 3225 1860 3234
rect 1714 3196 1766 3202
rect 1818 2920 1846 3225
rect 1806 2914 1858 2920
rect 1806 2856 1858 2862
rect 1634 2160 1754 2188
rect 2186 2172 2214 96220
rect 2278 94652 2306 97784
rect 2370 97304 2398 188224
rect 2450 187942 2502 187948
rect 2450 187884 2502 187890
rect 2462 97848 2490 187884
rect 2450 97842 2502 97848
rect 2450 97784 2502 97790
rect 2358 97298 2410 97304
rect 2358 97240 2410 97246
rect 2542 97298 2594 97304
rect 2542 97240 2594 97246
rect 2554 97003 2582 97240
rect 2540 96994 2596 97003
rect 2540 96929 2596 96938
rect 2358 96210 2410 96216
rect 2358 96152 2410 96158
rect 2370 95876 2398 96152
rect 2554 96028 2582 96929
rect 2462 96000 2582 96028
rect 2646 96012 2674 188292
rect 2818 188214 2870 188220
rect 2818 188156 2870 188162
rect 2726 188078 2778 188084
rect 2726 188020 2778 188026
rect 2738 97660 2766 188020
rect 2830 98392 2858 188156
rect 4750 187602 4802 187608
rect 4750 187544 4802 187550
rect 2890 187502 3186 187522
rect 2946 187500 2970 187502
rect 3026 187500 3050 187502
rect 3106 187500 3130 187502
rect 2968 187448 2970 187500
rect 3032 187448 3044 187500
rect 3106 187448 3108 187500
rect 2946 187446 2970 187448
rect 3026 187446 3050 187448
rect 3106 187446 3130 187448
rect 2890 187426 3186 187446
rect 4566 187330 4618 187336
rect 4566 187272 4618 187278
rect 4474 187194 4526 187200
rect 4474 187136 4526 187142
rect 4198 187058 4250 187064
rect 4198 187000 4250 187006
rect 4106 186786 4158 186792
rect 4106 186728 4158 186734
rect 3370 186650 3422 186656
rect 3370 186592 3422 186598
rect 2890 186414 3186 186434
rect 2946 186412 2970 186414
rect 3026 186412 3050 186414
rect 3106 186412 3130 186414
rect 2968 186360 2970 186412
rect 3032 186360 3044 186412
rect 3106 186360 3108 186412
rect 2946 186358 2970 186360
rect 3026 186358 3050 186360
rect 3106 186358 3130 186360
rect 2890 186338 3186 186358
rect 2890 185326 3186 185346
rect 2946 185324 2970 185326
rect 3026 185324 3050 185326
rect 3106 185324 3130 185326
rect 2968 185272 2970 185324
rect 3032 185272 3044 185324
rect 3106 185272 3108 185324
rect 2946 185270 2970 185272
rect 3026 185270 3050 185272
rect 3106 185270 3130 185272
rect 2890 185250 3186 185270
rect 2890 184238 3186 184258
rect 2946 184236 2970 184238
rect 3026 184236 3050 184238
rect 3106 184236 3130 184238
rect 2968 184184 2970 184236
rect 3032 184184 3044 184236
rect 3106 184184 3108 184236
rect 2946 184182 2970 184184
rect 3026 184182 3050 184184
rect 3106 184182 3130 184184
rect 2890 184162 3186 184182
rect 2890 183150 3186 183170
rect 2946 183148 2970 183150
rect 3026 183148 3050 183150
rect 3106 183148 3130 183150
rect 2968 183096 2970 183148
rect 3032 183096 3044 183148
rect 3106 183096 3108 183148
rect 2946 183094 2970 183096
rect 3026 183094 3050 183096
rect 3106 183094 3130 183096
rect 2890 183074 3186 183094
rect 2890 182062 3186 182082
rect 2946 182060 2970 182062
rect 3026 182060 3050 182062
rect 3106 182060 3130 182062
rect 2968 182008 2970 182060
rect 3032 182008 3044 182060
rect 3106 182008 3108 182060
rect 2946 182006 2970 182008
rect 3026 182006 3050 182008
rect 3106 182006 3130 182008
rect 2890 181986 3186 182006
rect 2890 180974 3186 180994
rect 2946 180972 2970 180974
rect 3026 180972 3050 180974
rect 3106 180972 3130 180974
rect 2968 180920 2970 180972
rect 3032 180920 3044 180972
rect 3106 180920 3108 180972
rect 2946 180918 2970 180920
rect 3026 180918 3050 180920
rect 3106 180918 3130 180920
rect 2890 180898 3186 180918
rect 2890 179886 3186 179906
rect 2946 179884 2970 179886
rect 3026 179884 3050 179886
rect 3106 179884 3130 179886
rect 2968 179832 2970 179884
rect 3032 179832 3044 179884
rect 3106 179832 3108 179884
rect 2946 179830 2970 179832
rect 3026 179830 3050 179832
rect 3106 179830 3130 179832
rect 2890 179810 3186 179830
rect 2890 178798 3186 178818
rect 2946 178796 2970 178798
rect 3026 178796 3050 178798
rect 3106 178796 3130 178798
rect 2968 178744 2970 178796
rect 3032 178744 3044 178796
rect 3106 178744 3108 178796
rect 2946 178742 2970 178744
rect 3026 178742 3050 178744
rect 3106 178742 3130 178744
rect 2890 178722 3186 178742
rect 2890 177710 3186 177730
rect 2946 177708 2970 177710
rect 3026 177708 3050 177710
rect 3106 177708 3130 177710
rect 2968 177656 2970 177708
rect 3032 177656 3044 177708
rect 3106 177656 3108 177708
rect 2946 177654 2970 177656
rect 3026 177654 3050 177656
rect 3106 177654 3130 177656
rect 2890 177634 3186 177654
rect 2890 176622 3186 176642
rect 2946 176620 2970 176622
rect 3026 176620 3050 176622
rect 3106 176620 3130 176622
rect 2968 176568 2970 176620
rect 3032 176568 3044 176620
rect 3106 176568 3108 176620
rect 2946 176566 2970 176568
rect 3026 176566 3050 176568
rect 3106 176566 3130 176568
rect 2890 176546 3186 176566
rect 3276 175738 3332 175747
rect 3276 175673 3332 175682
rect 3290 175640 3318 175673
rect 3278 175634 3330 175640
rect 3278 175576 3330 175582
rect 2890 175534 3186 175554
rect 2946 175532 2970 175534
rect 3026 175532 3050 175534
rect 3106 175532 3130 175534
rect 2968 175480 2970 175532
rect 3032 175480 3044 175532
rect 3106 175480 3108 175532
rect 2946 175478 2970 175480
rect 3026 175478 3050 175480
rect 3106 175478 3130 175480
rect 2890 175458 3186 175478
rect 2890 174446 3186 174466
rect 2946 174444 2970 174446
rect 3026 174444 3050 174446
rect 3106 174444 3130 174446
rect 2968 174392 2970 174444
rect 3032 174392 3044 174444
rect 3106 174392 3108 174444
rect 2946 174390 2970 174392
rect 3026 174390 3050 174392
rect 3106 174390 3130 174392
rect 2890 174370 3186 174390
rect 2890 173358 3186 173378
rect 2946 173356 2970 173358
rect 3026 173356 3050 173358
rect 3106 173356 3130 173358
rect 2968 173304 2970 173356
rect 3032 173304 3044 173356
rect 3106 173304 3108 173356
rect 2946 173302 2970 173304
rect 3026 173302 3050 173304
rect 3106 173302 3130 173304
rect 2890 173282 3186 173302
rect 2890 172270 3186 172290
rect 2946 172268 2970 172270
rect 3026 172268 3050 172270
rect 3106 172268 3130 172270
rect 2968 172216 2970 172268
rect 3032 172216 3044 172268
rect 3106 172216 3108 172268
rect 2946 172214 2970 172216
rect 3026 172214 3050 172216
rect 3106 172214 3130 172216
rect 2890 172194 3186 172214
rect 2890 171182 3186 171202
rect 2946 171180 2970 171182
rect 3026 171180 3050 171182
rect 3106 171180 3130 171182
rect 2968 171128 2970 171180
rect 3032 171128 3044 171180
rect 3106 171128 3108 171180
rect 2946 171126 2970 171128
rect 3026 171126 3050 171128
rect 3106 171126 3130 171128
rect 2890 171106 3186 171126
rect 2890 170094 3186 170114
rect 2946 170092 2970 170094
rect 3026 170092 3050 170094
rect 3106 170092 3130 170094
rect 2968 170040 2970 170092
rect 3032 170040 3044 170092
rect 3106 170040 3108 170092
rect 2946 170038 2970 170040
rect 3026 170038 3050 170040
rect 3106 170038 3130 170040
rect 2890 170018 3186 170038
rect 2890 169006 3186 169026
rect 2946 169004 2970 169006
rect 3026 169004 3050 169006
rect 3106 169004 3130 169006
rect 2968 168952 2970 169004
rect 3032 168952 3044 169004
rect 3106 168952 3108 169004
rect 2946 168950 2970 168952
rect 3026 168950 3050 168952
rect 3106 168950 3130 168952
rect 2890 168930 3186 168950
rect 2890 167918 3186 167938
rect 2946 167916 2970 167918
rect 3026 167916 3050 167918
rect 3106 167916 3130 167918
rect 2968 167864 2970 167916
rect 3032 167864 3044 167916
rect 3106 167864 3108 167916
rect 2946 167862 2970 167864
rect 3026 167862 3050 167864
rect 3106 167862 3130 167864
rect 2890 167842 3186 167862
rect 2890 166830 3186 166850
rect 2946 166828 2970 166830
rect 3026 166828 3050 166830
rect 3106 166828 3130 166830
rect 2968 166776 2970 166828
rect 3032 166776 3044 166828
rect 3106 166776 3108 166828
rect 2946 166774 2970 166776
rect 3026 166774 3050 166776
rect 3106 166774 3130 166776
rect 2890 166754 3186 166774
rect 2890 165742 3186 165762
rect 2946 165740 2970 165742
rect 3026 165740 3050 165742
rect 3106 165740 3130 165742
rect 2968 165688 2970 165740
rect 3032 165688 3044 165740
rect 3106 165688 3108 165740
rect 2946 165686 2970 165688
rect 3026 165686 3050 165688
rect 3106 165686 3130 165688
rect 2890 165666 3186 165686
rect 2890 164654 3186 164674
rect 2946 164652 2970 164654
rect 3026 164652 3050 164654
rect 3106 164652 3130 164654
rect 2968 164600 2970 164652
rect 3032 164600 3044 164652
rect 3106 164600 3108 164652
rect 2946 164598 2970 164600
rect 3026 164598 3050 164600
rect 3106 164598 3130 164600
rect 2890 164578 3186 164598
rect 2890 163566 3186 163586
rect 2946 163564 2970 163566
rect 3026 163564 3050 163566
rect 3106 163564 3130 163566
rect 2968 163512 2970 163564
rect 3032 163512 3044 163564
rect 3106 163512 3108 163564
rect 2946 163510 2970 163512
rect 3026 163510 3050 163512
rect 3106 163510 3130 163512
rect 2890 163490 3186 163510
rect 2890 162478 3186 162498
rect 2946 162476 2970 162478
rect 3026 162476 3050 162478
rect 3106 162476 3130 162478
rect 2968 162424 2970 162476
rect 3032 162424 3044 162476
rect 3106 162424 3108 162476
rect 2946 162422 2970 162424
rect 3026 162422 3050 162424
rect 3106 162422 3130 162424
rect 2890 162402 3186 162422
rect 2890 161390 3186 161410
rect 2946 161388 2970 161390
rect 3026 161388 3050 161390
rect 3106 161388 3130 161390
rect 2968 161336 2970 161388
rect 3032 161336 3044 161388
rect 3106 161336 3108 161388
rect 2946 161334 2970 161336
rect 3026 161334 3050 161336
rect 3106 161334 3130 161336
rect 2890 161314 3186 161334
rect 2890 160302 3186 160322
rect 2946 160300 2970 160302
rect 3026 160300 3050 160302
rect 3106 160300 3130 160302
rect 2968 160248 2970 160300
rect 3032 160248 3044 160300
rect 3106 160248 3108 160300
rect 2946 160246 2970 160248
rect 3026 160246 3050 160248
rect 3106 160246 3130 160248
rect 2890 160226 3186 160246
rect 2890 159214 3186 159234
rect 2946 159212 2970 159214
rect 3026 159212 3050 159214
rect 3106 159212 3130 159214
rect 2968 159160 2970 159212
rect 3032 159160 3044 159212
rect 3106 159160 3108 159212
rect 2946 159158 2970 159160
rect 3026 159158 3050 159160
rect 3106 159158 3130 159160
rect 2890 159138 3186 159158
rect 2890 158126 3186 158146
rect 2946 158124 2970 158126
rect 3026 158124 3050 158126
rect 3106 158124 3130 158126
rect 2968 158072 2970 158124
rect 3032 158072 3044 158124
rect 3106 158072 3108 158124
rect 2946 158070 2970 158072
rect 3026 158070 3050 158072
rect 3106 158070 3130 158072
rect 2890 158050 3186 158070
rect 2890 157038 3186 157058
rect 2946 157036 2970 157038
rect 3026 157036 3050 157038
rect 3106 157036 3130 157038
rect 2968 156984 2970 157036
rect 3032 156984 3044 157036
rect 3106 156984 3108 157036
rect 2946 156982 2970 156984
rect 3026 156982 3050 156984
rect 3106 156982 3130 156984
rect 2890 156962 3186 156982
rect 2890 155950 3186 155970
rect 2946 155948 2970 155950
rect 3026 155948 3050 155950
rect 3106 155948 3130 155950
rect 2968 155896 2970 155948
rect 3032 155896 3044 155948
rect 3106 155896 3108 155948
rect 2946 155894 2970 155896
rect 3026 155894 3050 155896
rect 3106 155894 3130 155896
rect 2890 155874 3186 155894
rect 2890 154862 3186 154882
rect 2946 154860 2970 154862
rect 3026 154860 3050 154862
rect 3106 154860 3130 154862
rect 2968 154808 2970 154860
rect 3032 154808 3044 154860
rect 3106 154808 3108 154860
rect 2946 154806 2970 154808
rect 3026 154806 3050 154808
rect 3106 154806 3130 154808
rect 2890 154786 3186 154806
rect 2890 153774 3186 153794
rect 2946 153772 2970 153774
rect 3026 153772 3050 153774
rect 3106 153772 3130 153774
rect 2968 153720 2970 153772
rect 3032 153720 3044 153772
rect 3106 153720 3108 153772
rect 2946 153718 2970 153720
rect 3026 153718 3050 153720
rect 3106 153718 3130 153720
rect 2890 153698 3186 153718
rect 2890 152686 3186 152706
rect 2946 152684 2970 152686
rect 3026 152684 3050 152686
rect 3106 152684 3130 152686
rect 2968 152632 2970 152684
rect 3032 152632 3044 152684
rect 3106 152632 3108 152684
rect 2946 152630 2970 152632
rect 3026 152630 3050 152632
rect 3106 152630 3130 152632
rect 2890 152610 3186 152630
rect 2890 151598 3186 151618
rect 2946 151596 2970 151598
rect 3026 151596 3050 151598
rect 3106 151596 3130 151598
rect 2968 151544 2970 151596
rect 3032 151544 3044 151596
rect 3106 151544 3108 151596
rect 2946 151542 2970 151544
rect 3026 151542 3050 151544
rect 3106 151542 3130 151544
rect 2890 151522 3186 151542
rect 2890 150510 3186 150530
rect 2946 150508 2970 150510
rect 3026 150508 3050 150510
rect 3106 150508 3130 150510
rect 2968 150456 2970 150508
rect 3032 150456 3044 150508
rect 3106 150456 3108 150508
rect 2946 150454 2970 150456
rect 3026 150454 3050 150456
rect 3106 150454 3130 150456
rect 2890 150434 3186 150454
rect 2890 149422 3186 149442
rect 2946 149420 2970 149422
rect 3026 149420 3050 149422
rect 3106 149420 3130 149422
rect 2968 149368 2970 149420
rect 3032 149368 3044 149420
rect 3106 149368 3108 149420
rect 2946 149366 2970 149368
rect 3026 149366 3050 149368
rect 3106 149366 3130 149368
rect 2890 149346 3186 149366
rect 2890 148334 3186 148354
rect 2946 148332 2970 148334
rect 3026 148332 3050 148334
rect 3106 148332 3130 148334
rect 2968 148280 2970 148332
rect 3032 148280 3044 148332
rect 3106 148280 3108 148332
rect 2946 148278 2970 148280
rect 3026 148278 3050 148280
rect 3106 148278 3130 148280
rect 2890 148258 3186 148278
rect 2890 147246 3186 147266
rect 2946 147244 2970 147246
rect 3026 147244 3050 147246
rect 3106 147244 3130 147246
rect 2968 147192 2970 147244
rect 3032 147192 3044 147244
rect 3106 147192 3108 147244
rect 2946 147190 2970 147192
rect 3026 147190 3050 147192
rect 3106 147190 3130 147192
rect 2890 147170 3186 147190
rect 2890 146158 3186 146178
rect 2946 146156 2970 146158
rect 3026 146156 3050 146158
rect 3106 146156 3130 146158
rect 2968 146104 2970 146156
rect 3032 146104 3044 146156
rect 3106 146104 3108 146156
rect 2946 146102 2970 146104
rect 3026 146102 3050 146104
rect 3106 146102 3130 146104
rect 2890 146082 3186 146102
rect 2890 145070 3186 145090
rect 2946 145068 2970 145070
rect 3026 145068 3050 145070
rect 3106 145068 3130 145070
rect 2968 145016 2970 145068
rect 3032 145016 3044 145068
rect 3106 145016 3108 145068
rect 2946 145014 2970 145016
rect 3026 145014 3050 145016
rect 3106 145014 3130 145016
rect 2890 144994 3186 145014
rect 2890 143982 3186 144002
rect 2946 143980 2970 143982
rect 3026 143980 3050 143982
rect 3106 143980 3130 143982
rect 2968 143928 2970 143980
rect 3032 143928 3044 143980
rect 3106 143928 3108 143980
rect 2946 143926 2970 143928
rect 3026 143926 3050 143928
rect 3106 143926 3130 143928
rect 2890 143906 3186 143926
rect 2890 142894 3186 142914
rect 2946 142892 2970 142894
rect 3026 142892 3050 142894
rect 3106 142892 3130 142894
rect 2968 142840 2970 142892
rect 3032 142840 3044 142892
rect 3106 142840 3108 142892
rect 2946 142838 2970 142840
rect 3026 142838 3050 142840
rect 3106 142838 3130 142840
rect 2890 142818 3186 142838
rect 2890 141806 3186 141826
rect 2946 141804 2970 141806
rect 3026 141804 3050 141806
rect 3106 141804 3130 141806
rect 2968 141752 2970 141804
rect 3032 141752 3044 141804
rect 3106 141752 3108 141804
rect 2946 141750 2970 141752
rect 3026 141750 3050 141752
rect 3106 141750 3130 141752
rect 2890 141730 3186 141750
rect 2890 140718 3186 140738
rect 2946 140716 2970 140718
rect 3026 140716 3050 140718
rect 3106 140716 3130 140718
rect 2968 140664 2970 140716
rect 3032 140664 3044 140716
rect 3106 140664 3108 140716
rect 2946 140662 2970 140664
rect 3026 140662 3050 140664
rect 3106 140662 3130 140664
rect 2890 140642 3186 140662
rect 2890 139630 3186 139650
rect 2946 139628 2970 139630
rect 3026 139628 3050 139630
rect 3106 139628 3130 139630
rect 2968 139576 2970 139628
rect 3032 139576 3044 139628
rect 3106 139576 3108 139628
rect 2946 139574 2970 139576
rect 3026 139574 3050 139576
rect 3106 139574 3130 139576
rect 2890 139554 3186 139574
rect 2890 138542 3186 138562
rect 2946 138540 2970 138542
rect 3026 138540 3050 138542
rect 3106 138540 3130 138542
rect 2968 138488 2970 138540
rect 3032 138488 3044 138540
rect 3106 138488 3108 138540
rect 2946 138486 2970 138488
rect 3026 138486 3050 138488
rect 3106 138486 3130 138488
rect 2890 138466 3186 138486
rect 2890 137454 3186 137474
rect 2946 137452 2970 137454
rect 3026 137452 3050 137454
rect 3106 137452 3130 137454
rect 2968 137400 2970 137452
rect 3032 137400 3044 137452
rect 3106 137400 3108 137452
rect 2946 137398 2970 137400
rect 3026 137398 3050 137400
rect 3106 137398 3130 137400
rect 2890 137378 3186 137398
rect 2890 136366 3186 136386
rect 2946 136364 2970 136366
rect 3026 136364 3050 136366
rect 3106 136364 3130 136366
rect 2968 136312 2970 136364
rect 3032 136312 3044 136364
rect 3106 136312 3108 136364
rect 2946 136310 2970 136312
rect 3026 136310 3050 136312
rect 3106 136310 3130 136312
rect 2890 136290 3186 136310
rect 2890 135278 3186 135298
rect 2946 135276 2970 135278
rect 3026 135276 3050 135278
rect 3106 135276 3130 135278
rect 2968 135224 2970 135276
rect 3032 135224 3044 135276
rect 3106 135224 3108 135276
rect 2946 135222 2970 135224
rect 3026 135222 3050 135224
rect 3106 135222 3130 135224
rect 2890 135202 3186 135222
rect 2890 134190 3186 134210
rect 2946 134188 2970 134190
rect 3026 134188 3050 134190
rect 3106 134188 3130 134190
rect 2968 134136 2970 134188
rect 3032 134136 3044 134188
rect 3106 134136 3108 134188
rect 2946 134134 2970 134136
rect 3026 134134 3050 134136
rect 3106 134134 3130 134136
rect 2890 134114 3186 134134
rect 2890 133102 3186 133122
rect 2946 133100 2970 133102
rect 3026 133100 3050 133102
rect 3106 133100 3130 133102
rect 2968 133048 2970 133100
rect 3032 133048 3044 133100
rect 3106 133048 3108 133100
rect 2946 133046 2970 133048
rect 3026 133046 3050 133048
rect 3106 133046 3130 133048
rect 2890 133026 3186 133046
rect 2890 132014 3186 132034
rect 2946 132012 2970 132014
rect 3026 132012 3050 132014
rect 3106 132012 3130 132014
rect 2968 131960 2970 132012
rect 3032 131960 3044 132012
rect 3106 131960 3108 132012
rect 2946 131958 2970 131960
rect 3026 131958 3050 131960
rect 3106 131958 3130 131960
rect 2890 131938 3186 131958
rect 2890 130926 3186 130946
rect 2946 130924 2970 130926
rect 3026 130924 3050 130926
rect 3106 130924 3130 130926
rect 2968 130872 2970 130924
rect 3032 130872 3044 130924
rect 3106 130872 3108 130924
rect 2946 130870 2970 130872
rect 3026 130870 3050 130872
rect 3106 130870 3130 130872
rect 2890 130850 3186 130870
rect 2890 129838 3186 129858
rect 2946 129836 2970 129838
rect 3026 129836 3050 129838
rect 3106 129836 3130 129838
rect 2968 129784 2970 129836
rect 3032 129784 3044 129836
rect 3106 129784 3108 129836
rect 2946 129782 2970 129784
rect 3026 129782 3050 129784
rect 3106 129782 3130 129784
rect 2890 129762 3186 129782
rect 2890 128750 3186 128770
rect 2946 128748 2970 128750
rect 3026 128748 3050 128750
rect 3106 128748 3130 128750
rect 2968 128696 2970 128748
rect 3032 128696 3044 128748
rect 3106 128696 3108 128748
rect 2946 128694 2970 128696
rect 3026 128694 3050 128696
rect 3106 128694 3130 128696
rect 2890 128674 3186 128694
rect 2890 127662 3186 127682
rect 2946 127660 2970 127662
rect 3026 127660 3050 127662
rect 3106 127660 3130 127662
rect 2968 127608 2970 127660
rect 3032 127608 3044 127660
rect 3106 127608 3108 127660
rect 2946 127606 2970 127608
rect 3026 127606 3050 127608
rect 3106 127606 3130 127608
rect 2890 127586 3186 127606
rect 2890 126574 3186 126594
rect 2946 126572 2970 126574
rect 3026 126572 3050 126574
rect 3106 126572 3130 126574
rect 2968 126520 2970 126572
rect 3032 126520 3044 126572
rect 3106 126520 3108 126572
rect 2946 126518 2970 126520
rect 3026 126518 3050 126520
rect 3106 126518 3130 126520
rect 2890 126498 3186 126518
rect 2890 125486 3186 125506
rect 2946 125484 2970 125486
rect 3026 125484 3050 125486
rect 3106 125484 3130 125486
rect 2968 125432 2970 125484
rect 3032 125432 3044 125484
rect 3106 125432 3108 125484
rect 2946 125430 2970 125432
rect 3026 125430 3050 125432
rect 3106 125430 3130 125432
rect 2890 125410 3186 125430
rect 2890 124398 3186 124418
rect 2946 124396 2970 124398
rect 3026 124396 3050 124398
rect 3106 124396 3130 124398
rect 2968 124344 2970 124396
rect 3032 124344 3044 124396
rect 3106 124344 3108 124396
rect 2946 124342 2970 124344
rect 3026 124342 3050 124344
rect 3106 124342 3130 124344
rect 2890 124322 3186 124342
rect 2890 123310 3186 123330
rect 2946 123308 2970 123310
rect 3026 123308 3050 123310
rect 3106 123308 3130 123310
rect 2968 123256 2970 123308
rect 3032 123256 3044 123308
rect 3106 123256 3108 123308
rect 2946 123254 2970 123256
rect 3026 123254 3050 123256
rect 3106 123254 3130 123256
rect 2890 123234 3186 123254
rect 2890 122222 3186 122242
rect 2946 122220 2970 122222
rect 3026 122220 3050 122222
rect 3106 122220 3130 122222
rect 2968 122168 2970 122220
rect 3032 122168 3044 122220
rect 3106 122168 3108 122220
rect 2946 122166 2970 122168
rect 3026 122166 3050 122168
rect 3106 122166 3130 122168
rect 2890 122146 3186 122166
rect 2890 121134 3186 121154
rect 2946 121132 2970 121134
rect 3026 121132 3050 121134
rect 3106 121132 3130 121134
rect 2968 121080 2970 121132
rect 3032 121080 3044 121132
rect 3106 121080 3108 121132
rect 2946 121078 2970 121080
rect 3026 121078 3050 121080
rect 3106 121078 3130 121080
rect 2890 121058 3186 121078
rect 2890 120046 3186 120066
rect 2946 120044 2970 120046
rect 3026 120044 3050 120046
rect 3106 120044 3130 120046
rect 2968 119992 2970 120044
rect 3032 119992 3044 120044
rect 3106 119992 3108 120044
rect 2946 119990 2970 119992
rect 3026 119990 3050 119992
rect 3106 119990 3130 119992
rect 2890 119970 3186 119990
rect 2890 118958 3186 118978
rect 2946 118956 2970 118958
rect 3026 118956 3050 118958
rect 3106 118956 3130 118958
rect 2968 118904 2970 118956
rect 3032 118904 3044 118956
rect 3106 118904 3108 118956
rect 2946 118902 2970 118904
rect 3026 118902 3050 118904
rect 3106 118902 3130 118904
rect 2890 118882 3186 118902
rect 2890 117870 3186 117890
rect 2946 117868 2970 117870
rect 3026 117868 3050 117870
rect 3106 117868 3130 117870
rect 2968 117816 2970 117868
rect 3032 117816 3044 117868
rect 3106 117816 3108 117868
rect 2946 117814 2970 117816
rect 3026 117814 3050 117816
rect 3106 117814 3130 117816
rect 2890 117794 3186 117814
rect 2890 116782 3186 116802
rect 2946 116780 2970 116782
rect 3026 116780 3050 116782
rect 3106 116780 3130 116782
rect 2968 116728 2970 116780
rect 3032 116728 3044 116780
rect 3106 116728 3108 116780
rect 2946 116726 2970 116728
rect 3026 116726 3050 116728
rect 3106 116726 3130 116728
rect 2890 116706 3186 116726
rect 2890 115694 3186 115714
rect 2946 115692 2970 115694
rect 3026 115692 3050 115694
rect 3106 115692 3130 115694
rect 2968 115640 2970 115692
rect 3032 115640 3044 115692
rect 3106 115640 3108 115692
rect 2946 115638 2970 115640
rect 3026 115638 3050 115640
rect 3106 115638 3130 115640
rect 2890 115618 3186 115638
rect 2890 114606 3186 114626
rect 2946 114604 2970 114606
rect 3026 114604 3050 114606
rect 3106 114604 3130 114606
rect 2968 114552 2970 114604
rect 3032 114552 3044 114604
rect 3106 114552 3108 114604
rect 2946 114550 2970 114552
rect 3026 114550 3050 114552
rect 3106 114550 3130 114552
rect 2890 114530 3186 114550
rect 2890 113518 3186 113538
rect 2946 113516 2970 113518
rect 3026 113516 3050 113518
rect 3106 113516 3130 113518
rect 2968 113464 2970 113516
rect 3032 113464 3044 113516
rect 3106 113464 3108 113516
rect 2946 113462 2970 113464
rect 3026 113462 3050 113464
rect 3106 113462 3130 113464
rect 2890 113442 3186 113462
rect 2890 112430 3186 112450
rect 2946 112428 2970 112430
rect 3026 112428 3050 112430
rect 3106 112428 3130 112430
rect 2968 112376 2970 112428
rect 3032 112376 3044 112428
rect 3106 112376 3108 112428
rect 2946 112374 2970 112376
rect 3026 112374 3050 112376
rect 3106 112374 3130 112376
rect 2890 112354 3186 112374
rect 2890 111342 3186 111362
rect 2946 111340 2970 111342
rect 3026 111340 3050 111342
rect 3106 111340 3130 111342
rect 2968 111288 2970 111340
rect 3032 111288 3044 111340
rect 3106 111288 3108 111340
rect 2946 111286 2970 111288
rect 3026 111286 3050 111288
rect 3106 111286 3130 111288
rect 2890 111266 3186 111286
rect 2890 110254 3186 110274
rect 2946 110252 2970 110254
rect 3026 110252 3050 110254
rect 3106 110252 3130 110254
rect 2968 110200 2970 110252
rect 3032 110200 3044 110252
rect 3106 110200 3108 110252
rect 2946 110198 2970 110200
rect 3026 110198 3050 110200
rect 3106 110198 3130 110200
rect 2890 110178 3186 110198
rect 2890 109166 3186 109186
rect 2946 109164 2970 109166
rect 3026 109164 3050 109166
rect 3106 109164 3130 109166
rect 2968 109112 2970 109164
rect 3032 109112 3044 109164
rect 3106 109112 3108 109164
rect 2946 109110 2970 109112
rect 3026 109110 3050 109112
rect 3106 109110 3130 109112
rect 2890 109090 3186 109110
rect 2890 108078 3186 108098
rect 2946 108076 2970 108078
rect 3026 108076 3050 108078
rect 3106 108076 3130 108078
rect 2968 108024 2970 108076
rect 3032 108024 3044 108076
rect 3106 108024 3108 108076
rect 2946 108022 2970 108024
rect 3026 108022 3050 108024
rect 3106 108022 3130 108024
rect 2890 108002 3186 108022
rect 2890 106990 3186 107010
rect 2946 106988 2970 106990
rect 3026 106988 3050 106990
rect 3106 106988 3130 106990
rect 2968 106936 2970 106988
rect 3032 106936 3044 106988
rect 3106 106936 3108 106988
rect 2946 106934 2970 106936
rect 3026 106934 3050 106936
rect 3106 106934 3130 106936
rect 2890 106914 3186 106934
rect 2890 105902 3186 105922
rect 2946 105900 2970 105902
rect 3026 105900 3050 105902
rect 3106 105900 3130 105902
rect 2968 105848 2970 105900
rect 3032 105848 3044 105900
rect 3106 105848 3108 105900
rect 2946 105846 2970 105848
rect 3026 105846 3050 105848
rect 3106 105846 3130 105848
rect 2890 105826 3186 105846
rect 2890 104814 3186 104834
rect 2946 104812 2970 104814
rect 3026 104812 3050 104814
rect 3106 104812 3130 104814
rect 2968 104760 2970 104812
rect 3032 104760 3044 104812
rect 3106 104760 3108 104812
rect 2946 104758 2970 104760
rect 3026 104758 3050 104760
rect 3106 104758 3130 104760
rect 2890 104738 3186 104758
rect 2890 103726 3186 103746
rect 2946 103724 2970 103726
rect 3026 103724 3050 103726
rect 3106 103724 3130 103726
rect 2968 103672 2970 103724
rect 3032 103672 3044 103724
rect 3106 103672 3108 103724
rect 2946 103670 2970 103672
rect 3026 103670 3050 103672
rect 3106 103670 3130 103672
rect 2890 103650 3186 103670
rect 2890 102638 3186 102658
rect 2946 102636 2970 102638
rect 3026 102636 3050 102638
rect 3106 102636 3130 102638
rect 2968 102584 2970 102636
rect 3032 102584 3044 102636
rect 3106 102584 3108 102636
rect 2946 102582 2970 102584
rect 3026 102582 3050 102584
rect 3106 102582 3130 102584
rect 2890 102562 3186 102582
rect 2890 101550 3186 101570
rect 2946 101548 2970 101550
rect 3026 101548 3050 101550
rect 3106 101548 3130 101550
rect 2968 101496 2970 101548
rect 3032 101496 3044 101548
rect 3106 101496 3108 101548
rect 2946 101494 2970 101496
rect 3026 101494 3050 101496
rect 3106 101494 3130 101496
rect 2890 101474 3186 101494
rect 2890 100462 3186 100482
rect 2946 100460 2970 100462
rect 3026 100460 3050 100462
rect 3106 100460 3130 100462
rect 2968 100408 2970 100460
rect 3032 100408 3044 100460
rect 3106 100408 3108 100460
rect 2946 100406 2970 100408
rect 3026 100406 3050 100408
rect 3106 100406 3130 100408
rect 2890 100386 3186 100406
rect 2890 99374 3186 99394
rect 2946 99372 2970 99374
rect 3026 99372 3050 99374
rect 3106 99372 3130 99374
rect 2968 99320 2970 99372
rect 3032 99320 3044 99372
rect 3106 99320 3108 99372
rect 2946 99318 2970 99320
rect 3026 99318 3050 99320
rect 3106 99318 3130 99320
rect 2890 99298 3186 99318
rect 2818 98386 2870 98392
rect 2818 98328 2870 98334
rect 2890 98286 3186 98306
rect 2946 98284 2970 98286
rect 3026 98284 3050 98286
rect 3106 98284 3130 98286
rect 2968 98232 2970 98284
rect 3032 98232 3044 98284
rect 3106 98232 3108 98284
rect 2946 98230 2970 98232
rect 3026 98230 3050 98232
rect 3106 98230 3130 98232
rect 2890 98210 3186 98230
rect 2738 97644 2858 97660
rect 2738 97638 2870 97644
rect 2738 97632 2818 97638
rect 2738 96420 2766 97632
rect 2818 97580 2870 97586
rect 2818 97434 2870 97440
rect 2818 97376 2870 97382
rect 2726 96414 2778 96420
rect 2726 96356 2778 96362
rect 2634 96006 2686 96012
rect 2358 95870 2410 95876
rect 2358 95812 2410 95818
rect 2462 95756 2490 96000
rect 2634 95948 2686 95954
rect 2646 95892 2674 95948
rect 2370 95728 2490 95756
rect 2554 95864 2674 95892
rect 2266 94646 2318 94652
rect 2266 94588 2318 94594
rect 2370 5860 2398 95728
rect 2370 5832 2490 5860
rect 2266 4070 2318 4076
rect 2266 4012 2318 4018
rect 1726 2104 1754 2160
rect 2174 2166 2226 2172
rect 2174 2108 2226 2114
rect 1714 2098 1766 2104
rect 1714 2040 1766 2046
rect 890 1998 1186 2018
rect 946 1996 970 1998
rect 1026 1996 1050 1998
rect 1106 1996 1130 1998
rect 968 1944 970 1996
rect 1032 1944 1044 1996
rect 1106 1944 1108 1996
rect 946 1942 970 1944
rect 1026 1942 1050 1944
rect 1106 1942 1130 1944
rect 890 1922 1186 1942
rect 1726 1900 1754 2040
rect 1714 1894 1766 1900
rect 1714 1836 1766 1842
rect 2278 1084 2306 4012
rect 2358 3458 2410 3464
rect 2358 3400 2410 3406
rect 2370 2988 2398 3400
rect 2462 3192 2490 5832
rect 2554 4076 2582 95864
rect 2738 95196 2766 96356
rect 2726 95190 2778 95196
rect 2726 95132 2778 95138
rect 2634 94646 2686 94652
rect 2634 94588 2686 94594
rect 2646 88756 2674 94588
rect 2726 94306 2778 94312
rect 2726 94248 2778 94254
rect 2738 88820 2766 94248
rect 2830 88922 2858 97376
rect 2890 97198 3186 97218
rect 2946 97196 2970 97198
rect 3026 97196 3050 97198
rect 3106 97196 3130 97198
rect 2968 97144 2970 97196
rect 3032 97144 3044 97196
rect 3106 97144 3108 97196
rect 2946 97142 2970 97144
rect 3026 97142 3050 97144
rect 3106 97142 3130 97144
rect 2890 97122 3186 97142
rect 3002 96754 3054 96760
rect 3000 96722 3002 96731
rect 3054 96722 3056 96731
rect 3000 96657 3056 96666
rect 3186 96346 3238 96352
rect 3184 96314 3186 96323
rect 3238 96314 3240 96323
rect 3184 96249 3240 96258
rect 2890 96110 3186 96130
rect 2946 96108 2970 96110
rect 3026 96108 3050 96110
rect 3106 96108 3130 96110
rect 2968 96056 2970 96108
rect 3032 96056 3044 96108
rect 3106 96056 3108 96108
rect 2946 96054 2970 96056
rect 3026 96054 3050 96056
rect 3106 96054 3130 96056
rect 2890 96034 3186 96054
rect 2890 95022 3186 95042
rect 2946 95020 2970 95022
rect 3026 95020 3050 95022
rect 3106 95020 3130 95022
rect 2968 94968 2970 95020
rect 3032 94968 3044 95020
rect 3106 94968 3108 95020
rect 2946 94966 2970 94968
rect 3026 94966 3050 94968
rect 3106 94966 3130 94968
rect 2890 94946 3186 94966
rect 2890 93934 3186 93954
rect 2946 93932 2970 93934
rect 3026 93932 3050 93934
rect 3106 93932 3130 93934
rect 2968 93880 2970 93932
rect 3032 93880 3044 93932
rect 3106 93880 3108 93932
rect 2946 93878 2970 93880
rect 3026 93878 3050 93880
rect 3106 93878 3130 93880
rect 2890 93858 3186 93878
rect 2890 92846 3186 92866
rect 2946 92844 2970 92846
rect 3026 92844 3050 92846
rect 3106 92844 3130 92846
rect 2968 92792 2970 92844
rect 3032 92792 3044 92844
rect 3106 92792 3108 92844
rect 2946 92790 2970 92792
rect 3026 92790 3050 92792
rect 3106 92790 3130 92792
rect 2890 92770 3186 92790
rect 2890 91758 3186 91778
rect 2946 91756 2970 91758
rect 3026 91756 3050 91758
rect 3106 91756 3130 91758
rect 2968 91704 2970 91756
rect 3032 91704 3044 91756
rect 3106 91704 3108 91756
rect 2946 91702 2970 91704
rect 3026 91702 3050 91704
rect 3106 91702 3130 91704
rect 2890 91682 3186 91702
rect 2890 90670 3186 90690
rect 2946 90668 2970 90670
rect 3026 90668 3050 90670
rect 3106 90668 3130 90670
rect 2968 90616 2970 90668
rect 3032 90616 3044 90668
rect 3106 90616 3108 90668
rect 2946 90614 2970 90616
rect 3026 90614 3050 90616
rect 3106 90614 3130 90616
rect 2890 90594 3186 90614
rect 2890 89582 3186 89602
rect 2946 89580 2970 89582
rect 3026 89580 3050 89582
rect 3106 89580 3130 89582
rect 2968 89528 2970 89580
rect 3032 89528 3044 89580
rect 3106 89528 3108 89580
rect 2946 89526 2970 89528
rect 3026 89526 3050 89528
rect 3106 89526 3130 89528
rect 2890 89506 3186 89526
rect 2830 88894 2950 88922
rect 2738 88792 2858 88820
rect 2646 88728 2766 88756
rect 2634 82270 2686 82276
rect 2634 82212 2686 82218
rect 2542 4070 2594 4076
rect 2542 4012 2594 4018
rect 2450 3186 2502 3192
rect 2450 3128 2502 3134
rect 2462 3027 2490 3128
rect 2448 3018 2504 3027
rect 2358 2982 2410 2988
rect 2448 2953 2504 2962
rect 2358 2924 2410 2930
rect 2266 1078 2318 1084
rect 2266 1020 2318 1026
rect 2554 880 2582 4012
rect 2646 2240 2674 82212
rect 2738 2852 2766 88728
rect 2830 4076 2858 88792
rect 2922 88668 2950 88894
rect 2910 88662 2962 88668
rect 2910 88604 2962 88610
rect 2890 88494 3186 88514
rect 2946 88492 2970 88494
rect 3026 88492 3050 88494
rect 3106 88492 3130 88494
rect 2968 88440 2970 88492
rect 3032 88440 3044 88492
rect 3106 88440 3108 88492
rect 2946 88438 2970 88440
rect 3026 88438 3050 88440
rect 3106 88438 3130 88440
rect 2890 88418 3186 88438
rect 2890 87406 3186 87426
rect 2946 87404 2970 87406
rect 3026 87404 3050 87406
rect 3106 87404 3130 87406
rect 2968 87352 2970 87404
rect 3032 87352 3044 87404
rect 3106 87352 3108 87404
rect 2946 87350 2970 87352
rect 3026 87350 3050 87352
rect 3106 87350 3130 87352
rect 2890 87330 3186 87350
rect 2890 86318 3186 86338
rect 2946 86316 2970 86318
rect 3026 86316 3050 86318
rect 3106 86316 3130 86318
rect 2968 86264 2970 86316
rect 3032 86264 3044 86316
rect 3106 86264 3108 86316
rect 2946 86262 2970 86264
rect 3026 86262 3050 86264
rect 3106 86262 3130 86264
rect 2890 86242 3186 86262
rect 2890 85230 3186 85250
rect 2946 85228 2970 85230
rect 3026 85228 3050 85230
rect 3106 85228 3130 85230
rect 2968 85176 2970 85228
rect 3032 85176 3044 85228
rect 3106 85176 3108 85228
rect 2946 85174 2970 85176
rect 3026 85174 3050 85176
rect 3106 85174 3130 85176
rect 2890 85154 3186 85174
rect 2890 84142 3186 84162
rect 2946 84140 2970 84142
rect 3026 84140 3050 84142
rect 3106 84140 3130 84142
rect 2968 84088 2970 84140
rect 3032 84088 3044 84140
rect 3106 84088 3108 84140
rect 2946 84086 2970 84088
rect 3026 84086 3050 84088
rect 3106 84086 3130 84088
rect 2890 84066 3186 84086
rect 2890 83054 3186 83074
rect 2946 83052 2970 83054
rect 3026 83052 3050 83054
rect 3106 83052 3130 83054
rect 2968 83000 2970 83052
rect 3032 83000 3044 83052
rect 3106 83000 3108 83052
rect 2946 82998 2970 83000
rect 3026 82998 3050 83000
rect 3106 82998 3130 83000
rect 2890 82978 3186 82998
rect 3290 82276 3318 175576
rect 3382 97644 3410 186592
rect 3934 182819 3962 182845
rect 3920 182810 3976 182819
rect 3920 182745 3922 182754
rect 3974 182745 3976 182754
rect 3922 182716 3974 182722
rect 3552 181722 3608 181731
rect 3552 181657 3554 181666
rect 3606 181657 3608 181666
rect 3554 181628 3606 181634
rect 3566 180348 3594 181628
rect 3566 180320 3778 180348
rect 3554 180190 3606 180196
rect 3554 180132 3606 180138
rect 3566 179963 3594 180132
rect 3552 179954 3608 179963
rect 3552 179889 3608 179898
rect 3644 176826 3700 176835
rect 3644 176761 3700 176770
rect 3658 176728 3686 176761
rect 3646 176722 3698 176728
rect 3646 176664 3698 176670
rect 3658 174212 3686 176664
rect 3646 174206 3698 174212
rect 3646 174148 3698 174154
rect 3644 174106 3700 174115
rect 3644 174041 3700 174050
rect 3658 174008 3686 174041
rect 3646 174002 3698 174008
rect 3646 173944 3698 173950
rect 3462 173662 3514 173668
rect 3462 173604 3514 173610
rect 3474 155716 3502 173604
rect 3462 155710 3514 155716
rect 3462 155652 3514 155658
rect 3554 155642 3606 155648
rect 3554 155584 3606 155590
rect 3462 151834 3514 151840
rect 3462 151776 3514 151782
rect 3474 114916 3502 151776
rect 3566 146808 3594 155584
rect 3554 146802 3606 146808
rect 3554 146744 3606 146750
rect 3554 141566 3606 141572
rect 3554 141508 3606 141514
rect 3566 128856 3594 141508
rect 3554 128850 3606 128856
rect 3554 128792 3606 128798
rect 3554 123478 3606 123484
rect 3554 123420 3606 123426
rect 3462 114910 3514 114916
rect 3462 114852 3514 114858
rect 3460 114810 3516 114819
rect 3460 114745 3462 114754
rect 3514 114745 3516 114754
rect 3462 114716 3514 114722
rect 3370 97638 3422 97644
rect 3370 97580 3422 97586
rect 3370 97298 3422 97304
rect 3370 97240 3422 97246
rect 3382 94924 3410 97240
rect 3370 94918 3422 94924
rect 3370 94860 3422 94866
rect 3370 94374 3422 94380
rect 3370 94316 3422 94322
rect 3382 89960 3410 94316
rect 3370 89954 3422 89960
rect 3370 89896 3422 89902
rect 3278 82270 3330 82276
rect 3278 82212 3330 82218
rect 3290 82043 3318 82212
rect 3276 82034 3332 82043
rect 2890 81966 3186 81986
rect 3276 81969 3332 81978
rect 2946 81964 2970 81966
rect 3026 81964 3050 81966
rect 3106 81964 3130 81966
rect 2968 81912 2970 81964
rect 3032 81912 3044 81964
rect 3106 81912 3108 81964
rect 2946 81910 2970 81912
rect 3026 81910 3050 81912
rect 3106 81910 3130 81912
rect 2890 81890 3186 81910
rect 3370 80978 3422 80984
rect 3370 80920 3422 80926
rect 2890 80878 3186 80898
rect 2946 80876 2970 80878
rect 3026 80876 3050 80878
rect 3106 80876 3130 80878
rect 2968 80824 2970 80876
rect 3032 80824 3044 80876
rect 3106 80824 3108 80876
rect 2946 80822 2970 80824
rect 3026 80822 3050 80824
rect 3106 80822 3130 80824
rect 2890 80802 3186 80822
rect 2890 79790 3186 79810
rect 2946 79788 2970 79790
rect 3026 79788 3050 79790
rect 3106 79788 3130 79790
rect 2968 79736 2970 79788
rect 3032 79736 3044 79788
rect 3106 79736 3108 79788
rect 2946 79734 2970 79736
rect 3026 79734 3050 79736
rect 3106 79734 3130 79736
rect 2890 79714 3186 79734
rect 2890 78702 3186 78722
rect 2946 78700 2970 78702
rect 3026 78700 3050 78702
rect 3106 78700 3130 78702
rect 2968 78648 2970 78700
rect 3032 78648 3044 78700
rect 3106 78648 3108 78700
rect 2946 78646 2970 78648
rect 3026 78646 3050 78648
rect 3106 78646 3130 78648
rect 2890 78626 3186 78646
rect 2890 77614 3186 77634
rect 2946 77612 2970 77614
rect 3026 77612 3050 77614
rect 3106 77612 3130 77614
rect 2968 77560 2970 77612
rect 3032 77560 3044 77612
rect 3106 77560 3108 77612
rect 2946 77558 2970 77560
rect 3026 77558 3050 77560
rect 3106 77558 3130 77560
rect 2890 77538 3186 77558
rect 2890 76526 3186 76546
rect 2946 76524 2970 76526
rect 3026 76524 3050 76526
rect 3106 76524 3130 76526
rect 2968 76472 2970 76524
rect 3032 76472 3044 76524
rect 3106 76472 3108 76524
rect 2946 76470 2970 76472
rect 3026 76470 3050 76472
rect 3106 76470 3130 76472
rect 2890 76450 3186 76470
rect 2890 75438 3186 75458
rect 2946 75436 2970 75438
rect 3026 75436 3050 75438
rect 3106 75436 3130 75438
rect 2968 75384 2970 75436
rect 3032 75384 3044 75436
rect 3106 75384 3108 75436
rect 2946 75382 2970 75384
rect 3026 75382 3050 75384
rect 3106 75382 3130 75384
rect 2890 75362 3186 75382
rect 2890 74350 3186 74370
rect 2946 74348 2970 74350
rect 3026 74348 3050 74350
rect 3106 74348 3130 74350
rect 2968 74296 2970 74348
rect 3032 74296 3044 74348
rect 3106 74296 3108 74348
rect 2946 74294 2970 74296
rect 3026 74294 3050 74296
rect 3106 74294 3130 74296
rect 2890 74274 3186 74294
rect 2890 73262 3186 73282
rect 2946 73260 2970 73262
rect 3026 73260 3050 73262
rect 3106 73260 3130 73262
rect 2968 73208 2970 73260
rect 3032 73208 3044 73260
rect 3106 73208 3108 73260
rect 2946 73206 2970 73208
rect 3026 73206 3050 73208
rect 3106 73206 3130 73208
rect 2890 73186 3186 73206
rect 2890 72174 3186 72194
rect 2946 72172 2970 72174
rect 3026 72172 3050 72174
rect 3106 72172 3130 72174
rect 2968 72120 2970 72172
rect 3032 72120 3044 72172
rect 3106 72120 3108 72172
rect 2946 72118 2970 72120
rect 3026 72118 3050 72120
rect 3106 72118 3130 72120
rect 2890 72098 3186 72118
rect 2890 71086 3186 71106
rect 2946 71084 2970 71086
rect 3026 71084 3050 71086
rect 3106 71084 3130 71086
rect 2968 71032 2970 71084
rect 3032 71032 3044 71084
rect 3106 71032 3108 71084
rect 2946 71030 2970 71032
rect 3026 71030 3050 71032
rect 3106 71030 3130 71032
rect 2890 71010 3186 71030
rect 2890 69998 3186 70018
rect 2946 69996 2970 69998
rect 3026 69996 3050 69998
rect 3106 69996 3130 69998
rect 2968 69944 2970 69996
rect 3032 69944 3044 69996
rect 3106 69944 3108 69996
rect 2946 69942 2970 69944
rect 3026 69942 3050 69944
rect 3106 69942 3130 69944
rect 2890 69922 3186 69942
rect 2890 68910 3186 68930
rect 2946 68908 2970 68910
rect 3026 68908 3050 68910
rect 3106 68908 3130 68910
rect 2968 68856 2970 68908
rect 3032 68856 3044 68908
rect 3106 68856 3108 68908
rect 2946 68854 2970 68856
rect 3026 68854 3050 68856
rect 3106 68854 3130 68856
rect 2890 68834 3186 68854
rect 2890 67822 3186 67842
rect 2946 67820 2970 67822
rect 3026 67820 3050 67822
rect 3106 67820 3130 67822
rect 2968 67768 2970 67820
rect 3032 67768 3044 67820
rect 3106 67768 3108 67820
rect 2946 67766 2970 67768
rect 3026 67766 3050 67768
rect 3106 67766 3130 67768
rect 2890 67746 3186 67766
rect 2890 66734 3186 66754
rect 2946 66732 2970 66734
rect 3026 66732 3050 66734
rect 3106 66732 3130 66734
rect 2968 66680 2970 66732
rect 3032 66680 3044 66732
rect 3106 66680 3108 66732
rect 2946 66678 2970 66680
rect 3026 66678 3050 66680
rect 3106 66678 3130 66680
rect 2890 66658 3186 66678
rect 2890 65646 3186 65666
rect 2946 65644 2970 65646
rect 3026 65644 3050 65646
rect 3106 65644 3130 65646
rect 2968 65592 2970 65644
rect 3032 65592 3044 65644
rect 3106 65592 3108 65644
rect 2946 65590 2970 65592
rect 3026 65590 3050 65592
rect 3106 65590 3130 65592
rect 2890 65570 3186 65590
rect 2890 64558 3186 64578
rect 2946 64556 2970 64558
rect 3026 64556 3050 64558
rect 3106 64556 3130 64558
rect 2968 64504 2970 64556
rect 3032 64504 3044 64556
rect 3106 64504 3108 64556
rect 2946 64502 2970 64504
rect 3026 64502 3050 64504
rect 3106 64502 3130 64504
rect 2890 64482 3186 64502
rect 2890 63470 3186 63490
rect 2946 63468 2970 63470
rect 3026 63468 3050 63470
rect 3106 63468 3130 63470
rect 2968 63416 2970 63468
rect 3032 63416 3044 63468
rect 3106 63416 3108 63468
rect 2946 63414 2970 63416
rect 3026 63414 3050 63416
rect 3106 63414 3130 63416
rect 2890 63394 3186 63414
rect 2890 62382 3186 62402
rect 2946 62380 2970 62382
rect 3026 62380 3050 62382
rect 3106 62380 3130 62382
rect 2968 62328 2970 62380
rect 3032 62328 3044 62380
rect 3106 62328 3108 62380
rect 2946 62326 2970 62328
rect 3026 62326 3050 62328
rect 3106 62326 3130 62328
rect 2890 62306 3186 62326
rect 2890 61294 3186 61314
rect 2946 61292 2970 61294
rect 3026 61292 3050 61294
rect 3106 61292 3130 61294
rect 2968 61240 2970 61292
rect 3032 61240 3044 61292
rect 3106 61240 3108 61292
rect 2946 61238 2970 61240
rect 3026 61238 3050 61240
rect 3106 61238 3130 61240
rect 2890 61218 3186 61238
rect 2890 60206 3186 60226
rect 2946 60204 2970 60206
rect 3026 60204 3050 60206
rect 3106 60204 3130 60206
rect 2968 60152 2970 60204
rect 3032 60152 3044 60204
rect 3106 60152 3108 60204
rect 2946 60150 2970 60152
rect 3026 60150 3050 60152
rect 3106 60150 3130 60152
rect 2890 60130 3186 60150
rect 2890 59118 3186 59138
rect 2946 59116 2970 59118
rect 3026 59116 3050 59118
rect 3106 59116 3130 59118
rect 2968 59064 2970 59116
rect 3032 59064 3044 59116
rect 3106 59064 3108 59116
rect 2946 59062 2970 59064
rect 3026 59062 3050 59064
rect 3106 59062 3130 59064
rect 2890 59042 3186 59062
rect 2890 58030 3186 58050
rect 2946 58028 2970 58030
rect 3026 58028 3050 58030
rect 3106 58028 3130 58030
rect 2968 57976 2970 58028
rect 3032 57976 3044 58028
rect 3106 57976 3108 58028
rect 2946 57974 2970 57976
rect 3026 57974 3050 57976
rect 3106 57974 3130 57976
rect 2890 57954 3186 57974
rect 2890 56942 3186 56962
rect 2946 56940 2970 56942
rect 3026 56940 3050 56942
rect 3106 56940 3130 56942
rect 2968 56888 2970 56940
rect 3032 56888 3044 56940
rect 3106 56888 3108 56940
rect 2946 56886 2970 56888
rect 3026 56886 3050 56888
rect 3106 56886 3130 56888
rect 2890 56866 3186 56886
rect 2890 55854 3186 55874
rect 2946 55852 2970 55854
rect 3026 55852 3050 55854
rect 3106 55852 3130 55854
rect 2968 55800 2970 55852
rect 3032 55800 3044 55852
rect 3106 55800 3108 55852
rect 2946 55798 2970 55800
rect 3026 55798 3050 55800
rect 3106 55798 3130 55800
rect 2890 55778 3186 55798
rect 2890 54766 3186 54786
rect 2946 54764 2970 54766
rect 3026 54764 3050 54766
rect 3106 54764 3130 54766
rect 2968 54712 2970 54764
rect 3032 54712 3044 54764
rect 3106 54712 3108 54764
rect 2946 54710 2970 54712
rect 3026 54710 3050 54712
rect 3106 54710 3130 54712
rect 2890 54690 3186 54710
rect 2890 53678 3186 53698
rect 2946 53676 2970 53678
rect 3026 53676 3050 53678
rect 3106 53676 3130 53678
rect 2968 53624 2970 53676
rect 3032 53624 3044 53676
rect 3106 53624 3108 53676
rect 2946 53622 2970 53624
rect 3026 53622 3050 53624
rect 3106 53622 3130 53624
rect 2890 53602 3186 53622
rect 2890 52590 3186 52610
rect 2946 52588 2970 52590
rect 3026 52588 3050 52590
rect 3106 52588 3130 52590
rect 2968 52536 2970 52588
rect 3032 52536 3044 52588
rect 3106 52536 3108 52588
rect 2946 52534 2970 52536
rect 3026 52534 3050 52536
rect 3106 52534 3130 52536
rect 2890 52514 3186 52534
rect 2890 51502 3186 51522
rect 2946 51500 2970 51502
rect 3026 51500 3050 51502
rect 3106 51500 3130 51502
rect 2968 51448 2970 51500
rect 3032 51448 3044 51500
rect 3106 51448 3108 51500
rect 2946 51446 2970 51448
rect 3026 51446 3050 51448
rect 3106 51446 3130 51448
rect 2890 51426 3186 51446
rect 2890 50414 3186 50434
rect 2946 50412 2970 50414
rect 3026 50412 3050 50414
rect 3106 50412 3130 50414
rect 2968 50360 2970 50412
rect 3032 50360 3044 50412
rect 3106 50360 3108 50412
rect 2946 50358 2970 50360
rect 3026 50358 3050 50360
rect 3106 50358 3130 50360
rect 2890 50338 3186 50358
rect 2890 49326 3186 49346
rect 2946 49324 2970 49326
rect 3026 49324 3050 49326
rect 3106 49324 3130 49326
rect 2968 49272 2970 49324
rect 3032 49272 3044 49324
rect 3106 49272 3108 49324
rect 2946 49270 2970 49272
rect 3026 49270 3050 49272
rect 3106 49270 3130 49272
rect 2890 49250 3186 49270
rect 2890 48238 3186 48258
rect 2946 48236 2970 48238
rect 3026 48236 3050 48238
rect 3106 48236 3130 48238
rect 2968 48184 2970 48236
rect 3032 48184 3044 48236
rect 3106 48184 3108 48236
rect 2946 48182 2970 48184
rect 3026 48182 3050 48184
rect 3106 48182 3130 48184
rect 2890 48162 3186 48182
rect 2890 47150 3186 47170
rect 2946 47148 2970 47150
rect 3026 47148 3050 47150
rect 3106 47148 3130 47150
rect 2968 47096 2970 47148
rect 3032 47096 3044 47148
rect 3106 47096 3108 47148
rect 2946 47094 2970 47096
rect 3026 47094 3050 47096
rect 3106 47094 3130 47096
rect 2890 47074 3186 47094
rect 2890 46062 3186 46082
rect 2946 46060 2970 46062
rect 3026 46060 3050 46062
rect 3106 46060 3130 46062
rect 2968 46008 2970 46060
rect 3032 46008 3044 46060
rect 3106 46008 3108 46060
rect 2946 46006 2970 46008
rect 3026 46006 3050 46008
rect 3106 46006 3130 46008
rect 2890 45986 3186 46006
rect 2890 44974 3186 44994
rect 2946 44972 2970 44974
rect 3026 44972 3050 44974
rect 3106 44972 3130 44974
rect 2968 44920 2970 44972
rect 3032 44920 3044 44972
rect 3106 44920 3108 44972
rect 2946 44918 2970 44920
rect 3026 44918 3050 44920
rect 3106 44918 3130 44920
rect 2890 44898 3186 44918
rect 3382 44876 3410 80920
rect 3370 44870 3422 44876
rect 3370 44812 3422 44818
rect 2890 43886 3186 43906
rect 2946 43884 2970 43886
rect 3026 43884 3050 43886
rect 3106 43884 3130 43886
rect 2968 43832 2970 43884
rect 3032 43832 3044 43884
rect 3106 43832 3108 43884
rect 2946 43830 2970 43832
rect 3026 43830 3050 43832
rect 3106 43830 3130 43832
rect 2890 43810 3186 43830
rect 2890 42798 3186 42818
rect 2946 42796 2970 42798
rect 3026 42796 3050 42798
rect 3106 42796 3130 42798
rect 2968 42744 2970 42796
rect 3032 42744 3044 42796
rect 3106 42744 3108 42796
rect 2946 42742 2970 42744
rect 3026 42742 3050 42744
rect 3106 42742 3130 42744
rect 2890 42722 3186 42742
rect 2890 41710 3186 41730
rect 2946 41708 2970 41710
rect 3026 41708 3050 41710
rect 3106 41708 3130 41710
rect 2968 41656 2970 41708
rect 3032 41656 3044 41708
rect 3106 41656 3108 41708
rect 2946 41654 2970 41656
rect 3026 41654 3050 41656
rect 3106 41654 3130 41656
rect 2890 41634 3186 41654
rect 2890 40622 3186 40642
rect 2946 40620 2970 40622
rect 3026 40620 3050 40622
rect 3106 40620 3130 40622
rect 2968 40568 2970 40620
rect 3032 40568 3044 40620
rect 3106 40568 3108 40620
rect 2946 40566 2970 40568
rect 3026 40566 3050 40568
rect 3106 40566 3130 40568
rect 2890 40546 3186 40566
rect 2890 39534 3186 39554
rect 2946 39532 2970 39534
rect 3026 39532 3050 39534
rect 3106 39532 3130 39534
rect 2968 39480 2970 39532
rect 3032 39480 3044 39532
rect 3106 39480 3108 39532
rect 2946 39478 2970 39480
rect 3026 39478 3050 39480
rect 3106 39478 3130 39480
rect 2890 39458 3186 39478
rect 2890 38446 3186 38466
rect 2946 38444 2970 38446
rect 3026 38444 3050 38446
rect 3106 38444 3130 38446
rect 2968 38392 2970 38444
rect 3032 38392 3044 38444
rect 3106 38392 3108 38444
rect 2946 38390 2970 38392
rect 3026 38390 3050 38392
rect 3106 38390 3130 38392
rect 2890 38370 3186 38390
rect 2890 37358 3186 37378
rect 2946 37356 2970 37358
rect 3026 37356 3050 37358
rect 3106 37356 3130 37358
rect 2968 37304 2970 37356
rect 3032 37304 3044 37356
rect 3106 37304 3108 37356
rect 2946 37302 2970 37304
rect 3026 37302 3050 37304
rect 3106 37302 3130 37304
rect 2890 37282 3186 37302
rect 2890 36270 3186 36290
rect 2946 36268 2970 36270
rect 3026 36268 3050 36270
rect 3106 36268 3130 36270
rect 2968 36216 2970 36268
rect 3032 36216 3044 36268
rect 3106 36216 3108 36268
rect 2946 36214 2970 36216
rect 3026 36214 3050 36216
rect 3106 36214 3130 36216
rect 2890 36194 3186 36214
rect 3278 35894 3330 35900
rect 3278 35836 3330 35842
rect 2890 35182 3186 35202
rect 2946 35180 2970 35182
rect 3026 35180 3050 35182
rect 3106 35180 3130 35182
rect 2968 35128 2970 35180
rect 3032 35128 3044 35180
rect 3106 35128 3108 35180
rect 2946 35126 2970 35128
rect 3026 35126 3050 35128
rect 3106 35126 3130 35128
rect 2890 35106 3186 35126
rect 3290 34579 3318 35836
rect 3276 34570 3332 34579
rect 3276 34505 3332 34514
rect 2890 34094 3186 34114
rect 2946 34092 2970 34094
rect 3026 34092 3050 34094
rect 3106 34092 3130 34094
rect 2968 34040 2970 34092
rect 3032 34040 3044 34092
rect 3106 34040 3108 34092
rect 2946 34038 2970 34040
rect 3026 34038 3050 34040
rect 3106 34038 3130 34040
rect 2890 34018 3186 34038
rect 2890 33006 3186 33026
rect 2946 33004 2970 33006
rect 3026 33004 3050 33006
rect 3106 33004 3130 33006
rect 2968 32952 2970 33004
rect 3032 32952 3044 33004
rect 3106 32952 3108 33004
rect 2946 32950 2970 32952
rect 3026 32950 3050 32952
rect 3106 32950 3130 32952
rect 2890 32930 3186 32950
rect 2890 31918 3186 31938
rect 2946 31916 2970 31918
rect 3026 31916 3050 31918
rect 3106 31916 3130 31918
rect 2968 31864 2970 31916
rect 3032 31864 3044 31916
rect 3106 31864 3108 31916
rect 2946 31862 2970 31864
rect 3026 31862 3050 31864
rect 3106 31862 3130 31864
rect 2890 31842 3186 31862
rect 2890 30830 3186 30850
rect 2946 30828 2970 30830
rect 3026 30828 3050 30830
rect 3106 30828 3130 30830
rect 2968 30776 2970 30828
rect 3032 30776 3044 30828
rect 3106 30776 3108 30828
rect 2946 30774 2970 30776
rect 3026 30774 3050 30776
rect 3106 30774 3130 30776
rect 2890 30754 3186 30774
rect 2890 29742 3186 29762
rect 2946 29740 2970 29742
rect 3026 29740 3050 29742
rect 3106 29740 3130 29742
rect 2968 29688 2970 29740
rect 3032 29688 3044 29740
rect 3106 29688 3108 29740
rect 2946 29686 2970 29688
rect 3026 29686 3050 29688
rect 3106 29686 3130 29688
rect 2890 29666 3186 29686
rect 2890 28654 3186 28674
rect 2946 28652 2970 28654
rect 3026 28652 3050 28654
rect 3106 28652 3130 28654
rect 2968 28600 2970 28652
rect 3032 28600 3044 28652
rect 3106 28600 3108 28652
rect 2946 28598 2970 28600
rect 3026 28598 3050 28600
rect 3106 28598 3130 28600
rect 2890 28578 3186 28598
rect 2890 27566 3186 27586
rect 2946 27564 2970 27566
rect 3026 27564 3050 27566
rect 3106 27564 3130 27566
rect 2968 27512 2970 27564
rect 3032 27512 3044 27564
rect 3106 27512 3108 27564
rect 2946 27510 2970 27512
rect 3026 27510 3050 27512
rect 3106 27510 3130 27512
rect 2890 27490 3186 27510
rect 2890 26478 3186 26498
rect 2946 26476 2970 26478
rect 3026 26476 3050 26478
rect 3106 26476 3130 26478
rect 2968 26424 2970 26476
rect 3032 26424 3044 26476
rect 3106 26424 3108 26476
rect 2946 26422 2970 26424
rect 3026 26422 3050 26424
rect 3106 26422 3130 26424
rect 2890 26402 3186 26422
rect 3368 25594 3424 25603
rect 3278 25558 3330 25564
rect 3368 25529 3370 25538
rect 3278 25500 3330 25506
rect 3422 25529 3424 25538
rect 3370 25500 3422 25506
rect 2890 25390 3186 25410
rect 2946 25388 2970 25390
rect 3026 25388 3050 25390
rect 3106 25388 3130 25390
rect 2968 25336 2970 25388
rect 3032 25336 3044 25388
rect 3106 25336 3108 25388
rect 2946 25334 2970 25336
rect 3026 25334 3050 25336
rect 3106 25334 3130 25336
rect 2890 25314 3186 25334
rect 2890 24302 3186 24322
rect 2946 24300 2970 24302
rect 3026 24300 3050 24302
rect 3106 24300 3130 24302
rect 2968 24248 2970 24300
rect 3032 24248 3044 24300
rect 3106 24248 3108 24300
rect 2946 24246 2970 24248
rect 3026 24246 3050 24248
rect 3106 24246 3130 24248
rect 2890 24226 3186 24246
rect 3290 24204 3318 25500
rect 3278 24198 3330 24204
rect 3278 24140 3330 24146
rect 2890 23214 3186 23234
rect 2946 23212 2970 23214
rect 3026 23212 3050 23214
rect 3106 23212 3130 23214
rect 2968 23160 2970 23212
rect 3032 23160 3044 23212
rect 3106 23160 3108 23212
rect 2946 23158 2970 23160
rect 3026 23158 3050 23160
rect 3106 23158 3130 23160
rect 2890 23138 3186 23158
rect 2890 22126 3186 22146
rect 2946 22124 2970 22126
rect 3026 22124 3050 22126
rect 3106 22124 3130 22126
rect 2968 22072 2970 22124
rect 3032 22072 3044 22124
rect 3106 22072 3108 22124
rect 2946 22070 2970 22072
rect 3026 22070 3050 22072
rect 3106 22070 3130 22072
rect 2890 22050 3186 22070
rect 2890 21038 3186 21058
rect 2946 21036 2970 21038
rect 3026 21036 3050 21038
rect 3106 21036 3130 21038
rect 2968 20984 2970 21036
rect 3032 20984 3044 21036
rect 3106 20984 3108 21036
rect 2946 20982 2970 20984
rect 3026 20982 3050 20984
rect 3106 20982 3130 20984
rect 2890 20962 3186 20982
rect 2890 19950 3186 19970
rect 2946 19948 2970 19950
rect 3026 19948 3050 19950
rect 3106 19948 3130 19950
rect 2968 19896 2970 19948
rect 3032 19896 3044 19948
rect 3106 19896 3108 19948
rect 2946 19894 2970 19896
rect 3026 19894 3050 19896
rect 3106 19894 3130 19896
rect 2890 19874 3186 19894
rect 2890 18862 3186 18882
rect 2946 18860 2970 18862
rect 3026 18860 3050 18862
rect 3106 18860 3130 18862
rect 2968 18808 2970 18860
rect 3032 18808 3044 18860
rect 3106 18808 3108 18860
rect 2946 18806 2970 18808
rect 3026 18806 3050 18808
rect 3106 18806 3130 18808
rect 2890 18786 3186 18806
rect 2890 17774 3186 17794
rect 2946 17772 2970 17774
rect 3026 17772 3050 17774
rect 3106 17772 3130 17774
rect 2968 17720 2970 17772
rect 3032 17720 3044 17772
rect 3106 17720 3108 17772
rect 2946 17718 2970 17720
rect 3026 17718 3050 17720
rect 3106 17718 3130 17720
rect 2890 17698 3186 17718
rect 3474 17035 3502 114716
rect 3566 110700 3594 123420
rect 3554 110694 3606 110700
rect 3554 110636 3606 110642
rect 3554 105458 3606 105464
rect 3554 105400 3606 105406
rect 3566 83160 3594 105400
rect 3554 83154 3606 83160
rect 3552 83122 3554 83131
rect 3606 83122 3608 83131
rect 3552 83057 3608 83066
rect 3460 17026 3516 17035
rect 3460 16961 3516 16970
rect 2890 16686 3186 16706
rect 2946 16684 2970 16686
rect 3026 16684 3050 16686
rect 3106 16684 3130 16686
rect 2968 16632 2970 16684
rect 3032 16632 3044 16684
rect 3106 16632 3108 16684
rect 2946 16630 2970 16632
rect 3026 16630 3050 16632
rect 3106 16630 3130 16632
rect 2890 16610 3186 16630
rect 3460 16618 3516 16627
rect 3460 16553 3516 16562
rect 2890 15598 3186 15618
rect 2946 15596 2970 15598
rect 3026 15596 3050 15598
rect 3106 15596 3130 15598
rect 2968 15544 2970 15596
rect 3032 15544 3044 15596
rect 3106 15544 3108 15596
rect 2946 15542 2970 15544
rect 3026 15542 3050 15544
rect 3106 15542 3130 15544
rect 2890 15522 3186 15542
rect 3278 15290 3330 15296
rect 3278 15232 3330 15238
rect 2890 14510 3186 14530
rect 2946 14508 2970 14510
rect 3026 14508 3050 14510
rect 3106 14508 3130 14510
rect 2968 14456 2970 14508
rect 3032 14456 3044 14508
rect 3106 14456 3108 14508
rect 2946 14454 2970 14456
rect 3026 14454 3050 14456
rect 3106 14454 3130 14456
rect 2890 14434 3186 14454
rect 3290 13664 3318 15232
rect 3278 13658 3330 13664
rect 3278 13600 3330 13606
rect 2890 13422 3186 13442
rect 2946 13420 2970 13422
rect 3026 13420 3050 13422
rect 3106 13420 3130 13422
rect 2968 13368 2970 13420
rect 3032 13368 3044 13420
rect 3106 13368 3108 13420
rect 2946 13366 2970 13368
rect 3026 13366 3050 13368
rect 3106 13366 3130 13368
rect 2890 13346 3186 13366
rect 2890 12334 3186 12354
rect 2946 12332 2970 12334
rect 3026 12332 3050 12334
rect 3106 12332 3130 12334
rect 2968 12280 2970 12332
rect 3032 12280 3044 12332
rect 3106 12280 3108 12332
rect 2946 12278 2970 12280
rect 3026 12278 3050 12280
rect 3106 12278 3130 12280
rect 2890 12258 3186 12278
rect 2890 11246 3186 11266
rect 2946 11244 2970 11246
rect 3026 11244 3050 11246
rect 3106 11244 3130 11246
rect 2968 11192 2970 11244
rect 3032 11192 3044 11244
rect 3106 11192 3108 11244
rect 2946 11190 2970 11192
rect 3026 11190 3050 11192
rect 3106 11190 3130 11192
rect 2890 11170 3186 11190
rect 2890 10158 3186 10178
rect 2946 10156 2970 10158
rect 3026 10156 3050 10158
rect 3106 10156 3130 10158
rect 2968 10104 2970 10156
rect 3032 10104 3044 10156
rect 3106 10104 3108 10156
rect 2946 10102 2970 10104
rect 3026 10102 3050 10104
rect 3106 10102 3130 10104
rect 2890 10082 3186 10102
rect 2890 9070 3186 9090
rect 2946 9068 2970 9070
rect 3026 9068 3050 9070
rect 3106 9068 3130 9070
rect 2968 9016 2970 9068
rect 3032 9016 3044 9068
rect 3106 9016 3108 9068
rect 2946 9014 2970 9016
rect 3026 9014 3050 9016
rect 3106 9014 3130 9016
rect 2890 8994 3186 9014
rect 2890 7982 3186 8002
rect 2946 7980 2970 7982
rect 3026 7980 3050 7982
rect 3106 7980 3130 7982
rect 2968 7928 2970 7980
rect 3032 7928 3044 7980
rect 3106 7928 3108 7980
rect 2946 7926 2970 7928
rect 3026 7926 3050 7928
rect 3106 7926 3130 7928
rect 2890 7906 3186 7926
rect 2890 6894 3186 6914
rect 2946 6892 2970 6894
rect 3026 6892 3050 6894
rect 3106 6892 3130 6894
rect 2968 6840 2970 6892
rect 3032 6840 3044 6892
rect 3106 6840 3108 6892
rect 2946 6838 2970 6840
rect 3026 6838 3050 6840
rect 3106 6838 3130 6840
rect 2890 6818 3186 6838
rect 2890 5806 3186 5826
rect 2946 5804 2970 5806
rect 3026 5804 3050 5806
rect 3106 5804 3130 5806
rect 2968 5752 2970 5804
rect 3032 5752 3044 5804
rect 3106 5752 3108 5804
rect 2946 5750 2970 5752
rect 3026 5750 3050 5752
rect 3106 5750 3130 5752
rect 2890 5730 3186 5750
rect 2890 4718 3186 4738
rect 2946 4716 2970 4718
rect 3026 4716 3050 4718
rect 3106 4716 3130 4718
rect 2968 4664 2970 4716
rect 3032 4664 3044 4716
rect 3106 4664 3108 4716
rect 2946 4662 2970 4664
rect 3026 4662 3050 4664
rect 3106 4662 3130 4664
rect 2890 4642 3186 4662
rect 2910 4274 2962 4280
rect 2908 4242 2910 4251
rect 2962 4242 2964 4251
rect 2908 4177 2964 4186
rect 2818 4070 2870 4076
rect 2818 4012 2870 4018
rect 3370 4002 3422 4008
rect 3370 3944 3422 3950
rect 2890 3630 3186 3650
rect 2946 3628 2970 3630
rect 3026 3628 3050 3630
rect 3106 3628 3130 3630
rect 2968 3576 2970 3628
rect 3032 3576 3044 3628
rect 3106 3576 3108 3628
rect 2946 3574 2970 3576
rect 3026 3574 3050 3576
rect 3106 3574 3130 3576
rect 2890 3554 3186 3574
rect 3276 3562 3332 3571
rect 3276 3497 3278 3506
rect 3330 3497 3332 3506
rect 3278 3468 3330 3474
rect 2818 3390 2870 3396
rect 2818 3332 2870 3338
rect 2830 2988 2858 3332
rect 3000 3154 3056 3163
rect 3000 3089 3056 3098
rect 2818 2982 2870 2988
rect 2818 2924 2870 2930
rect 2726 2846 2778 2852
rect 2726 2788 2778 2794
rect 2724 2746 2780 2755
rect 2724 2681 2726 2690
rect 2778 2681 2780 2690
rect 2726 2652 2778 2658
rect 2634 2234 2686 2240
rect 2634 2176 2686 2182
rect 2830 2188 2858 2924
rect 3014 2920 3042 3089
rect 3290 2988 3318 3468
rect 3278 2982 3330 2988
rect 3278 2924 3330 2930
rect 3002 2914 3054 2920
rect 3382 2868 3410 3944
rect 3002 2856 3054 2862
rect 3290 2840 3410 2868
rect 2890 2542 3186 2562
rect 2946 2540 2970 2542
rect 3026 2540 3050 2542
rect 3106 2540 3130 2542
rect 2968 2488 2970 2540
rect 3032 2488 3044 2540
rect 3106 2488 3108 2540
rect 2946 2486 2970 2488
rect 3026 2486 3050 2488
rect 3106 2486 3130 2488
rect 2890 2466 3186 2486
rect 2830 2160 2950 2188
rect 2818 2098 2870 2104
rect 2818 2040 2870 2046
rect 2830 1832 2858 2040
rect 2818 1826 2870 1832
rect 2818 1768 2870 1774
rect 2542 874 2594 880
rect 2542 816 2594 822
rect 2922 676 2950 2160
rect 2910 670 2962 676
rect 2910 612 2962 618
rect 3290 540 3318 2840
rect 3474 1531 3502 16553
rect 3566 2376 3594 83057
rect 3658 80003 3686 173944
rect 3750 164760 3778 180320
rect 3828 179954 3884 179963
rect 3828 179889 3884 179898
rect 3738 164754 3790 164760
rect 3738 164696 3790 164702
rect 3738 164550 3790 164556
rect 3738 164492 3790 164498
rect 3750 155648 3778 164492
rect 3738 155642 3790 155648
rect 3738 155584 3790 155590
rect 3738 155506 3790 155512
rect 3738 155448 3790 155454
rect 3750 146779 3778 155448
rect 3736 146770 3792 146779
rect 3736 146705 3792 146714
rect 3738 141634 3790 141640
rect 3738 141576 3790 141582
rect 3750 128652 3778 141576
rect 3738 128646 3790 128652
rect 3738 128588 3790 128594
rect 3738 123546 3790 123552
rect 3738 123488 3790 123494
rect 3750 110632 3778 123488
rect 3738 110626 3790 110632
rect 3738 110568 3790 110574
rect 3738 105526 3790 105532
rect 3738 105468 3790 105474
rect 3750 97100 3778 105468
rect 3738 97094 3790 97100
rect 3738 97036 3790 97042
rect 3738 95394 3790 95400
rect 3738 95336 3790 95342
rect 3750 94380 3778 95336
rect 3738 94374 3790 94380
rect 3738 94316 3790 94322
rect 3738 94238 3790 94244
rect 3738 94180 3790 94186
rect 3750 88843 3778 94180
rect 3736 88834 3792 88843
rect 3736 88769 3792 88778
rect 3738 88662 3790 88668
rect 3738 88604 3790 88610
rect 3750 87852 3778 88604
rect 3738 87846 3790 87852
rect 3738 87788 3790 87794
rect 3750 87619 3778 87788
rect 3736 87610 3792 87619
rect 3736 87545 3792 87554
rect 3644 79994 3700 80003
rect 3644 79929 3700 79938
rect 3658 79896 3686 79929
rect 3646 79890 3698 79896
rect 3646 79832 3698 79838
rect 3658 63372 3686 79832
rect 3750 63388 3778 87545
rect 3842 85880 3870 179889
rect 3934 97440 3962 182716
rect 4014 178898 4066 178904
rect 4012 178866 4014 178875
rect 4066 178866 4068 178875
rect 4012 178801 4068 178810
rect 4026 155580 4054 178801
rect 4014 155574 4066 155580
rect 4014 155516 4066 155522
rect 4014 155370 4066 155376
rect 4014 155312 4066 155318
rect 4026 146876 4054 155312
rect 4014 146870 4066 146876
rect 4014 146812 4066 146818
rect 4012 146770 4068 146779
rect 4012 146705 4068 146714
rect 3922 97434 3974 97440
rect 3922 97376 3974 97382
rect 3922 97094 3974 97100
rect 3922 97036 3974 97042
rect 3934 88668 3962 97036
rect 3922 88662 3974 88668
rect 3922 88604 3974 88610
rect 3920 88562 3976 88571
rect 3920 88497 3976 88506
rect 3830 85874 3882 85880
rect 3830 85816 3882 85822
rect 3646 63366 3698 63372
rect 3750 63360 3870 63388
rect 3646 63308 3698 63314
rect 3842 63139 3870 63360
rect 3828 63130 3884 63139
rect 3828 63065 3884 63074
rect 3934 63032 3962 88497
rect 4026 84860 4054 146705
rect 4118 116480 4146 186728
rect 4106 116474 4158 116480
rect 4106 116416 4158 116422
rect 4106 98386 4158 98392
rect 4104 98354 4106 98363
rect 4158 98354 4160 98363
rect 4104 98289 4160 98298
rect 4104 98218 4160 98227
rect 4104 98153 4106 98162
rect 4158 98153 4160 98162
rect 4106 98124 4158 98130
rect 4106 97502 4158 97508
rect 4106 97444 4158 97450
rect 4118 97032 4146 97444
rect 4106 97026 4158 97032
rect 4106 96968 4158 96974
rect 4106 96550 4158 96556
rect 4106 96492 4158 96498
rect 4118 96459 4146 96492
rect 4104 96450 4160 96459
rect 4104 96385 4160 96394
rect 4210 96323 4238 187000
rect 4290 116474 4342 116480
rect 4288 116442 4290 116451
rect 4342 116442 4344 116451
rect 4288 116377 4344 116386
rect 4290 114910 4342 114916
rect 4290 114852 4342 114858
rect 4302 96352 4330 114852
rect 4382 98998 4434 99004
rect 4382 98940 4434 98946
rect 4394 97796 4422 98940
rect 4486 98363 4514 187136
rect 4578 99140 4606 187272
rect 4658 186854 4710 186860
rect 4658 186796 4710 186802
rect 4566 99134 4618 99140
rect 4566 99076 4618 99082
rect 4670 99020 4698 186796
rect 4578 98992 4698 99020
rect 4762 99004 4790 187544
rect 5118 187398 5170 187404
rect 5118 187340 5170 187346
rect 4934 187126 4986 187132
rect 4934 187068 4986 187074
rect 4842 186718 4894 186724
rect 4842 186660 4894 186666
rect 4750 98998 4802 99004
rect 4472 98354 4528 98363
rect 4472 98289 4528 98298
rect 4394 97768 4514 97796
rect 4382 97638 4434 97644
rect 4382 97580 4434 97586
rect 4394 96624 4422 97580
rect 4486 97100 4514 97768
rect 4474 97094 4526 97100
rect 4474 97036 4526 97042
rect 4382 96618 4434 96624
rect 4382 96560 4434 96566
rect 4290 96346 4342 96352
rect 4196 96314 4252 96323
rect 4290 96288 4342 96294
rect 4196 96249 4252 96258
rect 4210 95332 4238 96249
rect 4290 96210 4342 96216
rect 4290 96152 4342 96158
rect 4198 95326 4250 95332
rect 4198 95268 4250 95274
rect 4302 95264 4330 96152
rect 4290 95258 4342 95264
rect 4290 95200 4342 95206
rect 4288 95090 4344 95099
rect 4288 95025 4344 95034
rect 4302 94516 4330 95025
rect 4290 94510 4342 94516
rect 4290 94452 4342 94458
rect 4106 88594 4158 88600
rect 4104 88562 4106 88571
rect 4158 88562 4160 88571
rect 4104 88497 4160 88506
rect 4014 84854 4066 84860
rect 4014 84796 4066 84802
rect 4026 84763 4054 84796
rect 4012 84754 4068 84763
rect 4012 84689 4068 84698
rect 3646 63026 3698 63032
rect 3830 63026 3882 63032
rect 3646 62968 3698 62974
rect 3736 62994 3792 63003
rect 3658 44876 3686 62968
rect 3830 62968 3882 62974
rect 3922 63026 3974 63032
rect 3922 62968 3974 62974
rect 3736 62929 3792 62938
rect 3750 44876 3778 62929
rect 3842 61604 3870 62968
rect 3830 61598 3882 61604
rect 3830 61540 3882 61546
rect 3830 56294 3882 56300
rect 3830 56236 3882 56242
rect 3646 44870 3698 44876
rect 3646 44812 3698 44818
rect 3738 44870 3790 44876
rect 3738 44812 3790 44818
rect 3842 44808 3870 56236
rect 3830 44802 3882 44808
rect 3830 44744 3882 44750
rect 3646 44598 3698 44604
rect 3646 44540 3698 44546
rect 3738 44598 3790 44604
rect 3738 44540 3790 44546
rect 3658 6252 3686 44540
rect 3646 6246 3698 6252
rect 3646 6188 3698 6194
rect 3644 5194 3700 5203
rect 3644 5129 3646 5138
rect 3698 5129 3700 5138
rect 3646 5100 3698 5106
rect 3554 2370 3606 2376
rect 3554 2312 3606 2318
rect 3460 1522 3516 1531
rect 3460 1457 3516 1466
rect 3658 1016 3686 5100
rect 3750 1803 3778 44540
rect 3830 44530 3882 44536
rect 3830 44472 3882 44478
rect 3842 35900 3870 44472
rect 3922 38342 3974 38348
rect 3922 38284 3974 38290
rect 3830 35894 3882 35900
rect 3830 35836 3882 35842
rect 3934 35780 3962 38284
rect 3842 35752 3962 35780
rect 3842 29508 3870 35752
rect 3920 34570 3976 34579
rect 3920 34505 3976 34514
rect 3830 29502 3882 29508
rect 3830 29444 3882 29450
rect 3830 29366 3882 29372
rect 3830 29308 3882 29314
rect 3842 22980 3870 29308
rect 3934 25603 3962 34505
rect 3920 25594 3976 25603
rect 3920 25529 3976 25538
rect 3830 22974 3882 22980
rect 3830 22916 3882 22922
rect 3828 22874 3884 22883
rect 3828 22809 3884 22818
rect 3842 22572 3870 22809
rect 3830 22566 3882 22572
rect 3830 22508 3882 22514
rect 3922 16582 3974 16588
rect 3922 16524 3974 16530
rect 3934 11488 3962 16524
rect 3922 11482 3974 11488
rect 3922 11424 3974 11430
rect 3830 11414 3882 11420
rect 3830 11356 3882 11362
rect 3842 1832 3870 11356
rect 3922 4070 3974 4076
rect 3922 4012 3974 4018
rect 3830 1826 3882 1832
rect 3736 1794 3792 1803
rect 3830 1768 3882 1774
rect 3736 1729 3792 1738
rect 3842 1220 3870 1768
rect 3934 1560 3962 4012
rect 4026 2075 4054 84689
rect 4118 2512 4146 88497
rect 4196 85978 4252 85987
rect 4196 85913 4252 85922
rect 4210 85880 4238 85913
rect 4198 85874 4250 85880
rect 4198 85816 4250 85822
rect 4106 2506 4158 2512
rect 4106 2448 4158 2454
rect 4012 2066 4068 2075
rect 4012 2001 4068 2010
rect 4210 1939 4238 85816
rect 4302 20600 4330 20631
rect 4290 20594 4342 20600
rect 4288 20562 4290 20571
rect 4342 20562 4344 20571
rect 4288 20497 4344 20506
rect 4196 1930 4252 1939
rect 4196 1865 4252 1874
rect 3922 1554 3974 1560
rect 3922 1496 3974 1502
rect 3830 1214 3882 1220
rect 3830 1156 3882 1162
rect 3646 1010 3698 1016
rect 3646 952 3698 958
rect 3278 534 3330 540
rect 3278 476 3330 482
rect 4302 132 4330 20497
rect 4394 4772 4422 96560
rect 4486 96556 4514 97036
rect 4578 96896 4606 98992
rect 4750 98940 4802 98946
rect 4854 98748 4882 186660
rect 4658 98726 4710 98732
rect 4658 98668 4710 98674
rect 4762 98720 4882 98748
rect 4946 98732 4974 187068
rect 4934 98726 4986 98732
rect 4566 96890 4618 96896
rect 4566 96832 4618 96838
rect 4578 96692 4606 96832
rect 4566 96686 4618 96692
rect 4566 96628 4618 96634
rect 4474 96550 4526 96556
rect 4474 96492 4526 96498
rect 4578 96300 4606 96628
rect 4486 96272 4606 96300
rect 4486 95212 4514 96272
rect 4670 96012 4698 98668
rect 4658 96006 4710 96012
rect 4658 95948 4710 95954
rect 4670 95348 4698 95948
rect 4762 95740 4790 98720
rect 4934 98668 4986 98674
rect 5130 98612 5158 187340
rect 4854 98584 5158 98612
rect 4750 95734 4802 95740
rect 4750 95676 4802 95682
rect 4854 95468 4882 98584
rect 5118 98182 5170 98188
rect 5118 98124 5170 98130
rect 4934 96754 4986 96760
rect 4934 96696 4986 96702
rect 4842 95462 4894 95468
rect 4842 95404 4894 95410
rect 4670 95320 4882 95348
rect 4854 95264 4882 95320
rect 4842 95258 4894 95264
rect 4486 95184 4698 95212
rect 4842 95200 4894 95206
rect 4474 95122 4526 95128
rect 4474 95064 4526 95070
rect 4566 95122 4618 95128
rect 4566 95064 4618 95070
rect 4486 4892 4514 95064
rect 4474 4886 4526 4892
rect 4474 4828 4526 4834
rect 4394 4744 4514 4772
rect 4380 4650 4436 4659
rect 4380 4585 4382 4594
rect 4434 4585 4436 4594
rect 4382 4556 4434 4562
rect 4382 4478 4434 4484
rect 4382 4420 4434 4426
rect 4394 3299 4422 4420
rect 4486 3396 4514 4744
rect 4474 3390 4526 3396
rect 4474 3332 4526 3338
rect 4380 3290 4436 3299
rect 4380 3225 4436 3234
rect 4394 2755 4422 3225
rect 4578 2920 4606 95064
rect 4566 2914 4618 2920
rect 4566 2856 4618 2862
rect 4380 2746 4436 2755
rect 4380 2681 4436 2690
rect 4578 812 4606 2856
rect 4670 2104 4698 95184
rect 4750 95122 4802 95128
rect 4750 95064 4802 95070
rect 4762 2619 4790 95064
rect 4748 2610 4804 2619
rect 4748 2545 4804 2554
rect 4854 2308 4882 95200
rect 4946 94856 4974 96696
rect 5026 96550 5078 96556
rect 5026 96492 5078 96498
rect 5038 95128 5066 96492
rect 5026 95122 5078 95128
rect 5026 95064 5078 95070
rect 5130 94940 5158 98124
rect 5222 96964 5250 188428
rect 5302 188418 5354 188424
rect 5302 188360 5354 188366
rect 5314 97032 5342 188360
rect 5762 187262 5814 187268
rect 5762 187204 5814 187210
rect 5578 151834 5630 151840
rect 5576 151802 5578 151811
rect 5630 151802 5632 151811
rect 5576 151737 5632 151746
rect 5302 97026 5354 97032
rect 5302 96968 5354 96974
rect 5210 96958 5262 96964
rect 5210 96900 5262 96906
rect 5222 96731 5250 96900
rect 5208 96722 5264 96731
rect 5208 96657 5264 96666
rect 5774 96148 5802 187204
rect 5866 96760 5894 188496
rect 82122 188350 82174 188356
rect 82122 188292 82174 188298
rect 81846 188282 81898 188288
rect 81846 188224 81898 188230
rect 81752 187978 81808 187987
rect 81752 187913 81808 187922
rect 81766 163944 81794 187913
rect 81754 163938 81806 163944
rect 81754 163880 81806 163886
rect 81858 162856 81886 188224
rect 81938 188146 81990 188152
rect 81938 188088 81990 188094
rect 81846 162850 81898 162856
rect 81846 162792 81898 162798
rect 81950 145312 81978 188088
rect 82030 187330 82082 187336
rect 82030 187272 82082 187278
rect 81938 145306 81990 145312
rect 81938 145248 81990 145254
rect 82042 143884 82070 187272
rect 82134 146604 82162 188292
rect 82398 188214 82450 188220
rect 82398 188156 82450 188162
rect 82214 188010 82266 188016
rect 82214 187952 82266 187958
rect 82226 147896 82254 187952
rect 82306 187874 82358 187880
rect 82306 187816 82358 187822
rect 82318 149188 82346 187816
rect 82410 150140 82438 188156
rect 82502 156940 82530 188496
rect 84342 188492 84370 189137
rect 84330 188486 84382 188492
rect 84330 188428 84382 188434
rect 85158 188418 85210 188424
rect 85158 188360 85210 188366
rect 82582 188078 82634 188084
rect 82582 188020 82634 188026
rect 82594 160748 82622 188020
rect 85170 187987 85198 188360
rect 85156 187978 85212 187987
rect 83226 187942 83278 187948
rect 85156 187913 85212 187922
rect 83226 187884 83278 187890
rect 82582 160742 82634 160748
rect 82582 160684 82634 160690
rect 82490 156934 82542 156940
rect 82490 156876 82542 156882
rect 82488 151802 82544 151811
rect 82488 151737 82544 151746
rect 82398 150134 82450 150140
rect 82398 150076 82450 150082
rect 82306 149182 82358 149188
rect 82306 149124 82358 149130
rect 82214 147890 82266 147896
rect 82214 147832 82266 147838
rect 82122 146598 82174 146604
rect 82122 146540 82174 146546
rect 82030 143878 82082 143884
rect 82030 143820 82082 143826
rect 81938 137690 81990 137696
rect 81938 137632 81990 137638
rect 81846 109334 81898 109340
rect 81846 109276 81898 109282
rect 81662 108178 81714 108184
rect 81662 108120 81714 108126
rect 81478 97502 81530 97508
rect 81478 97444 81530 97450
rect 81294 97298 81346 97304
rect 81294 97240 81346 97246
rect 81306 97116 81334 97240
rect 22138 97094 22190 97100
rect 22138 97036 22190 97042
rect 45322 97094 45374 97100
rect 45322 97036 45374 97042
rect 81214 97088 81334 97116
rect 81386 97094 81438 97100
rect 14594 97026 14646 97032
rect 14594 96968 14646 96974
rect 14606 96867 14634 96968
rect 14592 96858 14648 96867
rect 14592 96793 14648 96802
rect 5854 96754 5906 96760
rect 22150 96731 22178 97036
rect 28486 97026 28538 97032
rect 28486 96968 28538 96974
rect 28498 96867 28526 96968
rect 28484 96858 28540 96867
rect 25266 96822 25318 96828
rect 28484 96793 28540 96802
rect 25266 96764 25318 96770
rect 25278 96731 25306 96764
rect 5854 96696 5906 96702
rect 22136 96722 22192 96731
rect 22136 96657 22192 96666
rect 25264 96722 25320 96731
rect 25264 96657 25320 96666
rect 28944 96722 29000 96731
rect 28944 96657 28946 96666
rect 28998 96657 29000 96666
rect 29956 96722 30012 96731
rect 35016 96722 35072 96731
rect 29956 96657 30012 96666
rect 34926 96686 34978 96692
rect 28946 96628 28998 96634
rect 29970 96624 29998 96657
rect 35016 96657 35072 96666
rect 36856 96722 36912 96731
rect 36856 96657 36912 96666
rect 37040 96722 37096 96731
rect 37040 96657 37042 96666
rect 34926 96628 34978 96634
rect 29958 96618 30010 96624
rect 15696 96586 15752 96595
rect 24712 96586 24768 96595
rect 15696 96521 15752 96530
rect 24634 96544 24712 96572
rect 15710 96420 15738 96521
rect 15698 96414 15750 96420
rect 15698 96356 15750 96362
rect 24438 96414 24490 96420
rect 24438 96356 24490 96362
rect 24450 96300 24478 96356
rect 24634 96300 24662 96544
rect 29958 96560 30010 96566
rect 24712 96521 24768 96530
rect 33636 96450 33692 96459
rect 33558 96408 33636 96436
rect 24450 96272 24662 96300
rect 24988 96314 25044 96323
rect 33558 96284 33586 96408
rect 33636 96385 33692 96394
rect 24988 96249 24990 96258
rect 25042 96249 25044 96258
rect 33546 96278 33598 96284
rect 24990 96220 25042 96226
rect 33546 96220 33598 96226
rect 34466 96278 34518 96284
rect 34466 96220 34518 96226
rect 5486 96142 5538 96148
rect 5486 96084 5538 96090
rect 5762 96142 5814 96148
rect 5762 96084 5814 96090
rect 5498 95604 5526 96084
rect 18364 96042 18420 96051
rect 18364 95977 18366 95986
rect 18418 95977 18420 95986
rect 23424 96042 23480 96051
rect 23424 95977 23480 95986
rect 18366 95948 18418 95954
rect 14040 95906 14096 95915
rect 14040 95841 14096 95850
rect 16984 95906 17040 95915
rect 16984 95841 17040 95850
rect 14054 95740 14082 95841
rect 14042 95734 14094 95740
rect 14042 95676 14094 95682
rect 5486 95598 5538 95604
rect 5486 95540 5538 95546
rect 5038 94912 5158 94940
rect 4934 94850 4986 94856
rect 4934 94792 4986 94798
rect 4946 2852 4974 94792
rect 5038 94584 5066 94912
rect 5026 94578 5078 94584
rect 5026 94520 5078 94526
rect 5038 4008 5066 94520
rect 5394 93898 5446 93904
rect 5394 93840 5446 93846
rect 5406 91948 5434 93840
rect 5314 91920 5434 91948
rect 5314 28051 5342 91920
rect 5498 91812 5526 95540
rect 16998 95507 17026 95841
rect 18378 95536 18406 95948
rect 23438 95944 23466 95977
rect 23426 95938 23478 95944
rect 23426 95880 23478 95886
rect 23976 95906 24032 95915
rect 23976 95841 23978 95850
rect 24030 95841 24032 95850
rect 23978 95812 24030 95818
rect 25726 95802 25778 95808
rect 19836 95770 19892 95779
rect 25726 95744 25778 95750
rect 19836 95705 19892 95714
rect 18366 95530 18418 95536
rect 16984 95498 17040 95507
rect 11834 95462 11886 95468
rect 18366 95472 18418 95478
rect 16984 95433 17040 95442
rect 11834 95404 11886 95410
rect 8166 95128 8194 95159
rect 8154 95122 8206 95128
rect 8152 95090 8154 95099
rect 11846 95099 11874 95404
rect 16998 95196 17026 95433
rect 19850 95400 19878 95705
rect 19838 95394 19890 95400
rect 20758 95394 20810 95400
rect 19838 95336 19890 95342
rect 20756 95362 20758 95371
rect 20810 95362 20812 95371
rect 20756 95297 20812 95306
rect 25738 95235 25766 95744
rect 27196 95634 27252 95643
rect 27196 95569 27252 95578
rect 26646 95530 26698 95536
rect 26646 95472 26698 95478
rect 26658 95235 26686 95472
rect 24436 95226 24492 95235
rect 16986 95190 17038 95196
rect 24436 95161 24438 95170
rect 16986 95132 17038 95138
rect 24490 95161 24492 95170
rect 25724 95226 25780 95235
rect 25724 95161 25780 95170
rect 26644 95226 26700 95235
rect 26644 95161 26700 95170
rect 24438 95132 24490 95138
rect 8206 95090 8208 95099
rect 8152 95025 8208 95034
rect 11832 95090 11888 95099
rect 11832 95025 11888 95034
rect 8166 94924 8194 95025
rect 11096 94954 11152 94963
rect 8154 94918 8206 94924
rect 11096 94889 11152 94898
rect 23332 94954 23388 94963
rect 23332 94889 23388 94898
rect 25908 94954 25964 94963
rect 25908 94889 25910 94898
rect 8154 94860 8206 94866
rect 11110 94856 11138 94889
rect 11098 94850 11150 94856
rect 11098 94792 11150 94798
rect 18180 94818 18236 94827
rect 18180 94753 18236 94762
rect 19836 94818 19892 94827
rect 19836 94753 19892 94762
rect 20848 94818 20904 94827
rect 20848 94753 20904 94762
rect 5854 94034 5906 94040
rect 5854 93976 5906 93982
rect 5406 91784 5526 91812
rect 5406 89960 5434 91784
rect 5394 89954 5446 89960
rect 5394 89896 5446 89902
rect 5578 83426 5630 83432
rect 5578 83368 5630 83374
rect 5300 28042 5356 28051
rect 5300 27977 5356 27986
rect 5590 11488 5618 83368
rect 5866 38364 5894 93976
rect 18194 93972 18222 94753
rect 18272 94410 18328 94419
rect 18272 94345 18328 94354
rect 18286 94040 18314 94345
rect 18274 94034 18326 94040
rect 18274 93976 18326 93982
rect 18182 93966 18234 93972
rect 18182 93908 18234 93914
rect 19850 93904 19878 94753
rect 20862 94720 20890 94753
rect 20850 94714 20902 94720
rect 20850 94656 20902 94662
rect 23346 94244 23374 94889
rect 25962 94889 25964 94898
rect 25910 94860 25962 94866
rect 26000 94818 26056 94827
rect 26000 94753 26002 94762
rect 26054 94753 26056 94762
rect 26002 94724 26054 94730
rect 23334 94238 23386 94244
rect 23334 94180 23386 94186
rect 24620 94138 24676 94147
rect 24620 94073 24676 94082
rect 24634 94040 24662 94073
rect 24622 94034 24674 94040
rect 24622 93976 24674 93982
rect 19838 93898 19890 93904
rect 19838 93840 19890 93846
rect 27210 93331 27238 95569
rect 31154 95326 31206 95332
rect 31154 95268 31206 95274
rect 29774 95190 29826 95196
rect 29774 95132 29826 95138
rect 29682 94918 29734 94924
rect 29682 94860 29734 94866
rect 27288 94682 27344 94691
rect 27288 94617 27290 94626
rect 27342 94617 27344 94626
rect 27290 94588 27342 94594
rect 28392 94138 28448 94147
rect 28392 94073 28394 94082
rect 28446 94073 28448 94082
rect 28394 94044 28446 94050
rect 29694 93467 29722 94860
rect 29786 94652 29814 95132
rect 31166 95099 31194 95268
rect 34478 95235 34506 96220
rect 34938 95672 34966 96628
rect 35030 96556 35058 96657
rect 35018 96550 35070 96556
rect 35018 96492 35070 96498
rect 36870 96488 36898 96657
rect 37094 96657 37096 96666
rect 37042 96628 37094 96634
rect 38606 96550 38658 96556
rect 38606 96492 38658 96498
rect 36858 96482 36910 96488
rect 36858 96424 36910 96430
rect 38144 96178 38200 96187
rect 38144 96113 38200 96122
rect 37502 96074 37554 96080
rect 37502 96016 37554 96022
rect 34926 95666 34978 95672
rect 34926 95608 34978 95614
rect 35018 95530 35070 95536
rect 35018 95472 35070 95478
rect 34464 95226 34520 95235
rect 34464 95161 34520 95170
rect 31152 95090 31208 95099
rect 31152 95025 31208 95034
rect 35030 94963 35058 95472
rect 36214 95462 36266 95468
rect 36214 95404 36266 95410
rect 35662 95326 35714 95332
rect 35662 95268 35714 95274
rect 35674 95235 35702 95268
rect 36226 95235 36254 95404
rect 36306 95258 36358 95264
rect 35660 95226 35716 95235
rect 35660 95161 35716 95170
rect 36212 95226 36268 95235
rect 37514 95235 37542 96016
rect 38158 95604 38186 96113
rect 38146 95598 38198 95604
rect 38146 95540 38198 95546
rect 38618 95235 38646 96492
rect 41826 96346 41878 96352
rect 41826 96288 41878 96294
rect 44494 96346 44546 96352
rect 44494 96288 44546 96294
rect 41838 95235 41866 96288
rect 43758 95870 43810 95876
rect 43758 95812 43810 95818
rect 43770 95235 43798 95812
rect 44506 95235 44534 96288
rect 45334 96284 45362 97036
rect 56638 97026 56690 97032
rect 48724 96994 48780 97003
rect 48724 96929 48780 96938
rect 55532 96994 55588 97003
rect 56638 96968 56690 96974
rect 60870 97026 60922 97032
rect 60870 96968 60922 96974
rect 77980 96994 78036 97003
rect 55532 96929 55588 96938
rect 46608 96858 46664 96867
rect 46608 96793 46664 96802
rect 46622 96595 46650 96793
rect 48738 96731 48766 96929
rect 50198 96890 50250 96896
rect 50198 96832 50250 96838
rect 51024 96858 51080 96867
rect 50210 96731 50238 96832
rect 51024 96793 51080 96802
rect 51670 96822 51722 96828
rect 48724 96722 48780 96731
rect 48724 96657 48780 96666
rect 48908 96722 48964 96731
rect 48908 96657 48910 96666
rect 48962 96657 48964 96666
rect 50196 96722 50252 96731
rect 50196 96657 50252 96666
rect 48910 96628 48962 96634
rect 46608 96586 46664 96595
rect 46608 96521 46664 96530
rect 46518 96414 46570 96420
rect 46518 96356 46570 96362
rect 45322 96278 45374 96284
rect 45322 96220 45374 96226
rect 45322 95462 45374 95468
rect 45322 95404 45374 95410
rect 36306 95200 36358 95206
rect 37500 95226 37556 95235
rect 36212 95161 36268 95170
rect 36318 95099 36346 95200
rect 37500 95161 37556 95170
rect 38604 95226 38660 95235
rect 38604 95161 38660 95170
rect 41824 95226 41880 95235
rect 41824 95161 41880 95170
rect 43756 95226 43812 95235
rect 43756 95161 43812 95170
rect 44492 95226 44548 95235
rect 44492 95161 44548 95170
rect 36304 95090 36360 95099
rect 36304 95025 36360 95034
rect 37316 95090 37372 95099
rect 37316 95025 37318 95034
rect 37370 95025 37372 95034
rect 38788 95090 38844 95099
rect 38788 95025 38844 95034
rect 43940 95090 43996 95099
rect 43940 95025 43996 95034
rect 37318 94996 37370 95002
rect 38802 94992 38830 95025
rect 38790 94986 38842 94992
rect 35016 94954 35072 94963
rect 38790 94928 38842 94934
rect 43954 94924 43982 95025
rect 35016 94889 35072 94898
rect 43942 94918 43994 94924
rect 43942 94860 43994 94866
rect 30694 94714 30746 94720
rect 38790 94714 38842 94720
rect 30694 94656 30746 94662
rect 32440 94682 32496 94691
rect 29774 94646 29826 94652
rect 29774 94588 29826 94594
rect 29772 94410 29828 94419
rect 29772 94345 29774 94354
rect 29826 94345 29828 94354
rect 29774 94316 29826 94322
rect 30706 93875 30734 94656
rect 38790 94656 38842 94662
rect 41734 94714 41786 94720
rect 41734 94656 41786 94662
rect 32440 94617 32496 94626
rect 32454 94584 32482 94617
rect 32442 94578 32494 94584
rect 32442 94520 32494 94526
rect 33454 94374 33506 94380
rect 33454 94316 33506 94322
rect 31060 94002 31116 94011
rect 31060 93937 31116 93946
rect 30692 93866 30748 93875
rect 30692 93801 30748 93810
rect 29680 93458 29736 93467
rect 29680 93393 29736 93402
rect 27196 93322 27252 93331
rect 27196 93257 27252 93266
rect 31074 93224 31102 93937
rect 32348 93866 32404 93875
rect 32348 93801 32404 93810
rect 32362 93292 32390 93801
rect 33466 93360 33494 94316
rect 38054 94306 38106 94312
rect 38054 94248 38106 94254
rect 36306 94102 36358 94108
rect 36306 94044 36358 94050
rect 33636 93866 33692 93875
rect 33636 93801 33692 93810
rect 34924 93866 34980 93875
rect 34924 93801 34980 93810
rect 36212 93866 36268 93875
rect 36212 93801 36268 93810
rect 33650 93564 33678 93801
rect 34938 93632 34966 93801
rect 34926 93626 34978 93632
rect 34926 93568 34978 93574
rect 33638 93558 33690 93564
rect 33638 93500 33690 93506
rect 33454 93354 33506 93360
rect 33454 93296 33506 93302
rect 32350 93286 32402 93292
rect 32350 93228 32402 93234
rect 31062 93218 31114 93224
rect 31062 93160 31114 93166
rect 36226 93020 36254 93801
rect 36318 93739 36346 94044
rect 36304 93730 36360 93739
rect 36304 93665 36360 93674
rect 38066 93603 38094 94248
rect 38238 94034 38290 94040
rect 38238 93976 38290 93982
rect 38250 93603 38278 93976
rect 38052 93594 38108 93603
rect 38052 93529 38108 93538
rect 38236 93594 38292 93603
rect 38236 93529 38292 93538
rect 36214 93014 36266 93020
rect 36214 92956 36266 92962
rect 38802 92952 38830 94656
rect 40170 94646 40222 94652
rect 40170 94588 40222 94594
rect 40076 94546 40132 94555
rect 40076 94481 40132 94490
rect 40090 94448 40118 94481
rect 40078 94442 40130 94448
rect 40078 94384 40130 94390
rect 38880 93866 38936 93875
rect 38880 93801 38936 93810
rect 38894 93768 38922 93801
rect 38882 93762 38934 93768
rect 38882 93704 38934 93710
rect 38790 92946 38842 92952
rect 38790 92888 38842 92894
rect 40182 92544 40210 94588
rect 41456 94546 41512 94555
rect 41456 94481 41458 94490
rect 41510 94481 41512 94490
rect 41458 94452 41510 94458
rect 41746 94419 41774 94656
rect 42652 94546 42708 94555
rect 42652 94481 42654 94490
rect 42706 94481 42708 94490
rect 42654 94452 42706 94458
rect 41272 94410 41328 94419
rect 41272 94345 41328 94354
rect 41732 94410 41788 94419
rect 41732 94345 41788 94354
rect 43940 94410 43996 94419
rect 43940 94345 43996 94354
rect 45228 94410 45284 94419
rect 45228 94345 45284 94354
rect 41286 94176 41314 94345
rect 42654 94306 42706 94312
rect 42654 94248 42706 94254
rect 41274 94170 41326 94176
rect 42666 94147 42694 94248
rect 41274 94112 41326 94118
rect 42652 94138 42708 94147
rect 42652 94073 42708 94082
rect 43954 94040 43982 94345
rect 45242 94108 45270 94345
rect 45230 94102 45282 94108
rect 45230 94044 45282 94050
rect 43942 94034 43994 94040
rect 43942 93976 43994 93982
rect 42744 93866 42800 93875
rect 42744 93801 42800 93810
rect 42758 93496 42786 93801
rect 45334 93700 45362 95404
rect 45414 95394 45466 95400
rect 45414 95336 45466 95342
rect 45322 93694 45374 93700
rect 45322 93636 45374 93642
rect 42746 93490 42798 93496
rect 42746 93432 42798 93438
rect 45426 93088 45454 95336
rect 46530 95235 46558 96356
rect 50198 96278 50250 96284
rect 50198 96220 50250 96226
rect 47806 96210 47858 96216
rect 47620 96178 47676 96187
rect 47806 96152 47858 96158
rect 47620 96113 47676 96122
rect 47634 95672 47662 96113
rect 47622 95666 47674 95672
rect 47622 95608 47674 95614
rect 47818 95235 47846 96152
rect 50210 95235 50238 96220
rect 46516 95226 46572 95235
rect 46516 95161 46572 95170
rect 47804 95226 47860 95235
rect 47804 95161 47860 95170
rect 48724 95226 48780 95235
rect 48724 95161 48726 95170
rect 48778 95161 48780 95170
rect 50196 95226 50252 95235
rect 50196 95161 50252 95170
rect 48726 95132 48778 95138
rect 49094 95122 49146 95128
rect 49092 95090 49094 95099
rect 49146 95090 49148 95099
rect 49092 95025 49148 95034
rect 50380 95090 50436 95099
rect 50380 95025 50436 95034
rect 50394 94856 50422 95025
rect 51038 94924 51066 96793
rect 51670 96764 51722 96770
rect 51578 96142 51630 96148
rect 51578 96084 51630 96090
rect 51484 95634 51540 95643
rect 51484 95569 51540 95578
rect 51498 95536 51526 95569
rect 51486 95530 51538 95536
rect 51486 95472 51538 95478
rect 51590 95235 51618 96084
rect 51576 95226 51632 95235
rect 51576 95161 51632 95170
rect 51682 95128 51710 96764
rect 53050 96482 53102 96488
rect 55546 96459 55574 96929
rect 53050 96424 53102 96430
rect 55532 96450 55588 96459
rect 53062 96080 53090 96424
rect 55532 96385 55588 96394
rect 53050 96074 53102 96080
rect 53050 96016 53102 96022
rect 53142 95462 53194 95468
rect 53142 95404 53194 95410
rect 51762 95326 51814 95332
rect 51762 95268 51814 95274
rect 53050 95326 53102 95332
rect 53050 95268 53102 95274
rect 51670 95122 51722 95128
rect 51670 95064 51722 95070
rect 51026 94918 51078 94924
rect 51026 94860 51078 94866
rect 50382 94850 50434 94856
rect 50288 94818 50344 94827
rect 50382 94792 50434 94798
rect 50288 94753 50290 94762
rect 50342 94753 50344 94762
rect 50290 94724 50342 94730
rect 49092 94682 49148 94691
rect 49092 94617 49148 94626
rect 49106 94584 49134 94617
rect 49094 94578 49146 94584
rect 49094 94520 49146 94526
rect 51668 94410 51724 94419
rect 51668 94345 51670 94354
rect 51722 94345 51724 94354
rect 51670 94316 51722 94322
rect 48818 94238 48870 94244
rect 48818 94180 48870 94186
rect 46148 94002 46204 94011
rect 46148 93937 46204 93946
rect 48450 93966 48502 93972
rect 46162 93904 46190 93937
rect 48450 93908 48502 93914
rect 46150 93898 46202 93904
rect 46150 93840 46202 93846
rect 48462 93156 48490 93908
rect 48450 93150 48502 93156
rect 48450 93092 48502 93098
rect 45414 93082 45466 93088
rect 48830 93059 48858 94180
rect 45414 93024 45466 93030
rect 48816 93050 48872 93059
rect 48816 92985 48872 92994
rect 51774 92884 51802 95268
rect 53062 95060 53090 95268
rect 53050 95054 53102 95060
rect 53050 94996 53102 95002
rect 52956 94682 53012 94691
rect 52956 94617 52958 94626
rect 53010 94617 53012 94626
rect 52958 94588 53010 94594
rect 53154 94448 53182 95404
rect 53234 95394 53286 95400
rect 53234 95336 53286 95342
rect 53142 94442 53194 94448
rect 53142 94384 53194 94390
rect 53246 93768 53274 95336
rect 56650 95235 56678 96968
rect 56822 96482 56874 96488
rect 56822 96424 56874 96430
rect 56636 95226 56692 95235
rect 54154 95190 54206 95196
rect 56636 95161 56692 95170
rect 54154 95132 54206 95138
rect 54166 94924 54194 95132
rect 54244 95090 54300 95099
rect 54244 95025 54300 95034
rect 54154 94918 54206 94924
rect 54154 94860 54206 94866
rect 54152 94818 54208 94827
rect 54152 94753 54208 94762
rect 54166 94011 54194 94753
rect 54258 94448 54286 95025
rect 56834 94788 56862 96424
rect 57926 96006 57978 96012
rect 57926 95948 57978 95954
rect 57938 95235 57966 95948
rect 58018 95394 58070 95400
rect 58018 95336 58070 95342
rect 57924 95226 57980 95235
rect 57924 95161 57980 95170
rect 58030 95128 58058 95336
rect 58110 95258 58162 95264
rect 59398 95258 59450 95264
rect 58110 95200 58162 95206
rect 59396 95226 59398 95235
rect 59450 95226 59452 95235
rect 58018 95122 58070 95128
rect 58122 95099 58150 95200
rect 59396 95161 59452 95170
rect 58018 95064 58070 95070
rect 58108 95090 58164 95099
rect 58108 95025 58164 95034
rect 56822 94782 56874 94788
rect 56822 94724 56874 94730
rect 54246 94442 54298 94448
rect 54246 94384 54298 94390
rect 56360 94410 56416 94419
rect 56360 94345 56416 94354
rect 54152 94002 54208 94011
rect 54152 93937 54208 93946
rect 53692 93866 53748 93875
rect 53692 93801 53748 93810
rect 53706 93768 53734 93801
rect 53234 93762 53286 93768
rect 53234 93704 53286 93710
rect 53694 93762 53746 93768
rect 53694 93704 53746 93710
rect 56374 93700 56402 94345
rect 60778 94306 60830 94312
rect 56912 94274 56968 94283
rect 60778 94248 60830 94254
rect 56912 94209 56968 94218
rect 56362 93694 56414 93700
rect 56362 93636 56414 93642
rect 51762 92878 51814 92884
rect 51762 92820 51814 92826
rect 56926 92787 56954 94209
rect 60042 93762 60094 93768
rect 60042 93704 60094 93710
rect 60054 92952 60082 93704
rect 60790 93700 60818 94248
rect 60778 93694 60830 93700
rect 60778 93636 60830 93642
rect 60502 93490 60554 93496
rect 60502 93432 60554 93438
rect 60042 92946 60094 92952
rect 60042 92888 60094 92894
rect 56912 92778 56968 92787
rect 56912 92713 56968 92722
rect 60514 92651 60542 93432
rect 60882 92816 60910 96968
rect 77980 96929 78036 96938
rect 80282 96958 80334 96964
rect 64548 96722 64604 96731
rect 66572 96722 66628 96731
rect 64604 96680 64958 96708
rect 64548 96657 64604 96666
rect 64930 96595 64958 96680
rect 66572 96657 66628 96666
rect 73472 96722 73528 96731
rect 73472 96657 73528 96666
rect 64916 96586 64972 96595
rect 61974 96550 62026 96556
rect 61974 96492 62026 96498
rect 62526 96550 62578 96556
rect 64916 96521 64972 96530
rect 62526 96492 62578 96498
rect 61986 96300 62014 96492
rect 62066 96482 62118 96488
rect 62064 96450 62066 96459
rect 62118 96450 62120 96459
rect 62064 96385 62120 96394
rect 61986 96272 62198 96300
rect 61790 95938 61842 95944
rect 61790 95880 61842 95886
rect 61802 95235 61830 95880
rect 61974 95530 62026 95536
rect 61974 95472 62026 95478
rect 61788 95226 61844 95235
rect 61788 95161 61844 95170
rect 61986 94283 62014 95472
rect 62170 94856 62198 96272
rect 62432 96178 62488 96187
rect 62432 96113 62488 96122
rect 62342 95598 62394 95604
rect 62342 95540 62394 95546
rect 62250 95462 62302 95468
rect 62250 95404 62302 95410
rect 62158 94850 62210 94856
rect 62158 94792 62210 94798
rect 61972 94274 62028 94283
rect 61972 94209 62028 94218
rect 62262 93768 62290 95404
rect 62250 93762 62302 93768
rect 62250 93704 62302 93710
rect 60870 92810 60922 92816
rect 60870 92752 60922 92758
rect 62354 92748 62382 95540
rect 62446 92884 62474 96113
rect 62538 93156 62566 96492
rect 66586 96488 66614 96657
rect 66574 96482 66626 96488
rect 66574 96424 66626 96430
rect 73486 96436 73514 96657
rect 77994 96595 78022 96929
rect 80282 96900 80334 96906
rect 80190 96890 80242 96896
rect 80190 96832 80242 96838
rect 80098 96754 80150 96760
rect 80098 96696 80150 96702
rect 77980 96586 78036 96595
rect 74394 96550 74446 96556
rect 74394 96492 74446 96498
rect 77430 96550 77482 96556
rect 77980 96521 78036 96530
rect 77430 96492 77482 96498
rect 73564 96450 73620 96459
rect 73486 96408 73564 96436
rect 73564 96385 73620 96394
rect 62802 95870 62854 95876
rect 62802 95812 62854 95818
rect 62814 95235 62842 95812
rect 63446 95802 63498 95808
rect 63446 95744 63498 95750
rect 63354 95258 63406 95264
rect 62800 95226 62856 95235
rect 63354 95200 63406 95206
rect 62800 95161 62856 95170
rect 63262 94442 63314 94448
rect 63262 94384 63314 94390
rect 62526 93150 62578 93156
rect 62526 93092 62578 93098
rect 63274 93088 63302 94384
rect 63366 93836 63394 95200
rect 63354 93830 63406 93836
rect 63354 93772 63406 93778
rect 63458 93428 63486 95744
rect 68966 95734 69018 95740
rect 68966 95676 69018 95682
rect 68874 95462 68926 95468
rect 68874 95404 68926 95410
rect 68414 95258 68466 95264
rect 68414 95200 68466 95206
rect 66482 95122 66534 95128
rect 66480 95090 66482 95099
rect 66534 95090 66536 95099
rect 66480 95025 66536 95034
rect 68426 94720 68454 95200
rect 68414 94714 68466 94720
rect 68414 94656 68466 94662
rect 68506 94714 68558 94720
rect 68506 94656 68558 94662
rect 68518 94555 68546 94656
rect 68504 94546 68560 94555
rect 68504 94481 68560 94490
rect 66482 94442 66534 94448
rect 66480 94410 66482 94419
rect 66534 94410 66536 94419
rect 66480 94345 66536 94354
rect 63446 93422 63498 93428
rect 63446 93364 63498 93370
rect 63262 93082 63314 93088
rect 63262 93024 63314 93030
rect 62434 92878 62486 92884
rect 62434 92820 62486 92826
rect 62342 92742 62394 92748
rect 62342 92684 62394 92690
rect 68886 92680 68914 95404
rect 68978 93700 69006 95676
rect 71174 95666 71226 95672
rect 71174 95608 71226 95614
rect 69058 95598 69110 95604
rect 69058 95540 69110 95546
rect 69070 94788 69098 95540
rect 69242 95394 69294 95400
rect 69242 95336 69294 95342
rect 69150 94850 69202 94856
rect 69150 94792 69202 94798
rect 69058 94782 69110 94788
rect 69058 94724 69110 94730
rect 69058 94306 69110 94312
rect 69058 94248 69110 94254
rect 68966 93694 69018 93700
rect 68966 93636 69018 93642
rect 68874 92674 68926 92680
rect 55348 92642 55404 92651
rect 55348 92577 55350 92586
rect 55402 92577 55404 92586
rect 60500 92642 60556 92651
rect 68874 92616 68926 92622
rect 69070 92612 69098 94248
rect 69162 94244 69190 94792
rect 69150 94238 69202 94244
rect 69150 94180 69202 94186
rect 69254 93156 69282 95336
rect 69886 95326 69938 95332
rect 69886 95268 69938 95274
rect 69794 94170 69846 94176
rect 69794 94112 69846 94118
rect 69242 93150 69294 93156
rect 69242 93092 69294 93098
rect 69806 93088 69834 94112
rect 69898 93428 69926 95268
rect 71082 95122 71134 95128
rect 71082 95064 71134 95070
rect 70990 94714 71042 94720
rect 70990 94656 71042 94662
rect 71002 94555 71030 94656
rect 70988 94546 71044 94555
rect 70988 94481 71044 94490
rect 70990 94442 71042 94448
rect 70988 94410 70990 94419
rect 71042 94410 71044 94419
rect 70988 94345 71044 94354
rect 71094 93700 71122 95064
rect 71082 93694 71134 93700
rect 71082 93636 71134 93642
rect 69886 93422 69938 93428
rect 69886 93364 69938 93370
rect 69794 93082 69846 93088
rect 69794 93024 69846 93030
rect 71186 92952 71214 95608
rect 72462 94714 72514 94720
rect 72462 94656 72514 94662
rect 72370 94510 72422 94516
rect 72370 94452 72422 94458
rect 72382 94176 72410 94452
rect 72370 94170 72422 94176
rect 72370 94112 72422 94118
rect 72474 93836 72502 94656
rect 72554 94510 72606 94516
rect 72554 94452 72606 94458
rect 72566 93972 72594 94452
rect 74406 94448 74434 96492
rect 77442 95604 77470 96492
rect 80110 95779 80138 96696
rect 80096 95770 80152 95779
rect 80096 95705 80152 95714
rect 80202 95672 80230 96832
rect 80294 95944 80322 96900
rect 81214 96012 81242 97088
rect 81386 97036 81438 97042
rect 81398 96980 81426 97036
rect 81306 96952 81426 96980
rect 81202 96006 81254 96012
rect 81202 95948 81254 95954
rect 80282 95938 80334 95944
rect 80282 95880 80334 95886
rect 81306 95740 81334 96952
rect 81490 96731 81518 97444
rect 81476 96722 81532 96731
rect 81476 96657 81532 96666
rect 81490 96488 81518 96657
rect 81478 96482 81530 96488
rect 81478 96424 81530 96430
rect 81674 95915 81702 108120
rect 81754 101650 81806 101656
rect 81754 101592 81806 101598
rect 81660 95906 81716 95915
rect 81660 95841 81716 95850
rect 81294 95734 81346 95740
rect 81294 95676 81346 95682
rect 80190 95666 80242 95672
rect 80190 95608 80242 95614
rect 77430 95598 77482 95604
rect 77430 95540 77482 95546
rect 77430 95462 77482 95468
rect 77430 95404 77482 95410
rect 77442 95060 77470 95404
rect 80098 95394 80150 95400
rect 80098 95336 80150 95342
rect 77430 95054 77482 95060
rect 77430 94996 77482 95002
rect 80110 94963 80138 95336
rect 80190 95190 80242 95196
rect 80190 95132 80242 95138
rect 80096 94954 80152 94963
rect 80096 94889 80152 94898
rect 80202 94516 80230 95132
rect 80190 94510 80242 94516
rect 80190 94452 80242 94458
rect 74394 94442 74446 94448
rect 74394 94384 74446 94390
rect 81202 94442 81254 94448
rect 81766 94419 81794 101592
rect 81858 96051 81886 109276
rect 81844 96042 81900 96051
rect 81844 95977 81900 95986
rect 81950 95876 81978 137632
rect 82030 124770 82082 124776
rect 82030 124712 82082 124718
rect 81938 95870 81990 95876
rect 81938 95812 81990 95818
rect 82042 94992 82070 124712
rect 82122 123954 82174 123960
rect 82122 123896 82174 123902
rect 82134 96216 82162 123896
rect 82214 119670 82266 119676
rect 82214 119612 82266 119618
rect 82122 96210 82174 96216
rect 82122 96152 82174 96158
rect 82226 96080 82254 119612
rect 82502 119404 82530 151737
rect 83238 150723 83266 187884
rect 86890 187502 87186 187522
rect 86946 187500 86970 187502
rect 87026 187500 87050 187502
rect 87106 187500 87130 187502
rect 86968 187448 86970 187500
rect 87032 187448 87044 187500
rect 87106 187448 87108 187500
rect 86946 187446 86970 187448
rect 87026 187446 87050 187448
rect 87106 187446 87130 187448
rect 84236 187434 84292 187443
rect 86890 187426 87186 187446
rect 84236 187369 84292 187378
rect 84790 187398 84842 187404
rect 84054 187262 84106 187268
rect 84054 187204 84106 187210
rect 83318 187194 83370 187200
rect 83318 187136 83370 187142
rect 83330 165411 83358 187136
rect 83962 186582 84014 186588
rect 83962 186524 84014 186530
rect 83974 180779 84002 186524
rect 83960 180770 84016 180779
rect 83960 180705 84016 180714
rect 84066 180620 84094 187204
rect 84146 186786 84198 186792
rect 84146 186728 84198 186734
rect 83974 180592 84094 180620
rect 83776 176826 83832 176835
rect 83776 176761 83832 176770
rect 83316 165402 83372 165411
rect 83316 165337 83372 165346
rect 83224 150714 83280 150723
rect 83224 150649 83280 150658
rect 83316 136162 83372 136171
rect 83316 136097 83372 136106
rect 83226 129938 83278 129944
rect 83226 129880 83278 129886
rect 83134 128646 83186 128652
rect 83134 128588 83186 128594
rect 83042 120894 83094 120900
rect 83042 120836 83094 120842
rect 82490 119398 82542 119404
rect 82490 119340 82542 119346
rect 82398 116678 82450 116684
rect 82398 116620 82450 116626
rect 82306 114706 82358 114712
rect 82306 114648 82358 114654
rect 82214 96074 82266 96080
rect 82214 96016 82266 96022
rect 82030 94986 82082 94992
rect 82030 94928 82082 94934
rect 82318 94788 82346 114648
rect 82410 96352 82438 116620
rect 82950 115590 83002 115596
rect 82950 115532 83002 115538
rect 82490 112054 82542 112060
rect 82490 111996 82542 112002
rect 82398 96346 82450 96352
rect 82398 96288 82450 96294
rect 82502 96187 82530 111996
rect 82858 111986 82910 111992
rect 82858 111928 82910 111934
rect 82582 106614 82634 106620
rect 82582 106556 82634 106562
rect 82488 96178 82544 96187
rect 82488 96113 82544 96122
rect 82594 95808 82622 106556
rect 82766 102874 82818 102880
rect 82766 102816 82818 102822
rect 82674 98182 82726 98188
rect 82674 98124 82726 98130
rect 82582 95802 82634 95808
rect 82582 95744 82634 95750
rect 82306 94782 82358 94788
rect 82306 94724 82358 94730
rect 82686 94691 82714 98124
rect 82778 96148 82806 102816
rect 82870 96964 82898 111928
rect 82962 97100 82990 115532
rect 83054 97168 83082 120836
rect 83146 97372 83174 128588
rect 83134 97366 83186 97372
rect 83134 97308 83186 97314
rect 83042 97162 83094 97168
rect 83042 97104 83094 97110
rect 82950 97094 83002 97100
rect 82950 97036 83002 97042
rect 82858 96958 82910 96964
rect 82858 96900 82910 96906
rect 82766 96142 82818 96148
rect 82766 96084 82818 96090
rect 83238 95371 83266 129880
rect 83224 95362 83280 95371
rect 83224 95297 83280 95306
rect 83330 94856 83358 136097
rect 83592 130178 83648 130187
rect 83592 130113 83648 130122
rect 83410 127422 83462 127428
rect 83410 127364 83462 127370
rect 83318 94850 83370 94856
rect 83318 94792 83370 94798
rect 82766 94782 82818 94788
rect 82766 94724 82818 94730
rect 82672 94682 82728 94691
rect 82672 94617 82728 94626
rect 81202 94384 81254 94390
rect 81752 94410 81808 94419
rect 72554 93966 72606 93972
rect 72554 93908 72606 93914
rect 78440 93866 78496 93875
rect 72462 93830 72514 93836
rect 78440 93801 78496 93810
rect 72462 93772 72514 93778
rect 78454 93700 78482 93801
rect 78442 93694 78494 93700
rect 78442 93636 78494 93642
rect 78454 93496 78482 93636
rect 78442 93490 78494 93496
rect 78442 93432 78494 93438
rect 80190 93422 80242 93428
rect 80190 93364 80242 93370
rect 71174 92946 71226 92952
rect 71174 92888 71226 92894
rect 73750 92946 73802 92952
rect 73750 92888 73802 92894
rect 73762 92651 73790 92888
rect 80096 92778 80152 92787
rect 80096 92713 80152 92722
rect 73748 92642 73804 92651
rect 60500 92577 60556 92586
rect 69058 92606 69110 92612
rect 55350 92548 55402 92554
rect 73748 92577 73804 92586
rect 69058 92548 69110 92554
rect 80110 92544 80138 92713
rect 80202 92612 80230 93364
rect 81214 92816 81242 94384
rect 81752 94345 81808 94354
rect 81294 93898 81346 93904
rect 81294 93840 81346 93846
rect 81202 92810 81254 92816
rect 81202 92752 81254 92758
rect 80190 92606 80242 92612
rect 80190 92548 80242 92554
rect 40170 92538 40222 92544
rect 40170 92480 40222 92486
rect 80098 92538 80150 92544
rect 80098 92480 80150 92486
rect 81306 92068 81334 93840
rect 81844 93730 81900 93739
rect 81844 93665 81900 93674
rect 81660 93594 81716 93603
rect 81660 93529 81716 93538
rect 81384 93186 81440 93195
rect 81384 93121 81440 93130
rect 81294 92062 81346 92068
rect 81294 92004 81346 92010
rect 81398 89960 81426 93121
rect 81386 89954 81438 89960
rect 81386 89896 81438 89902
rect 81674 77380 81702 93529
rect 81662 77374 81714 77380
rect 81662 77316 81714 77322
rect 81858 74524 81886 93665
rect 82674 93558 82726 93564
rect 82674 93500 82726 93506
rect 82582 93490 82634 93496
rect 82488 93458 82544 93467
rect 82582 93432 82634 93438
rect 82488 93393 82544 93402
rect 82214 93354 82266 93360
rect 82120 93322 82176 93331
rect 82214 93296 82266 93302
rect 82120 93257 82176 93266
rect 81938 92810 81990 92816
rect 81938 92752 81990 92758
rect 81846 74518 81898 74524
rect 81846 74460 81898 74466
rect 81950 62828 81978 92752
rect 82030 92538 82082 92544
rect 82030 92480 82082 92486
rect 82042 66636 82070 92480
rect 82134 73164 82162 93257
rect 82226 83772 82254 93296
rect 82304 93050 82360 93059
rect 82304 92985 82360 92994
rect 82214 83766 82266 83772
rect 82214 83708 82266 83714
rect 82122 73158 82174 73164
rect 82122 73100 82174 73106
rect 82318 73096 82346 92985
rect 82502 74456 82530 93393
rect 82490 74450 82542 74456
rect 82490 74392 82542 74398
rect 82306 73090 82358 73096
rect 82306 73032 82358 73038
rect 82030 66630 82082 66636
rect 82030 66572 82082 66578
rect 81938 62822 81990 62828
rect 81938 62764 81990 62770
rect 81938 56498 81990 56504
rect 81938 56440 81990 56446
rect 5774 38336 5894 38364
rect 5774 29547 5802 38336
rect 5760 29538 5816 29547
rect 5760 29473 5816 29482
rect 81846 29502 81898 29508
rect 81846 29444 81898 29450
rect 81754 28550 81806 28556
rect 81754 28492 81806 28498
rect 81662 25626 81714 25632
rect 81662 25568 81714 25574
rect 5578 11482 5630 11488
rect 5578 11424 5630 11430
rect 5486 11414 5538 11420
rect 5486 11356 5538 11362
rect 5498 4092 5526 11356
rect 81570 7062 81622 7068
rect 81570 7004 81622 7010
rect 5762 6246 5814 6252
rect 5762 6188 5814 6194
rect 5314 4064 5526 4092
rect 5026 4002 5078 4008
rect 5026 3944 5078 3950
rect 5314 3940 5342 4064
rect 5302 3934 5354 3940
rect 5302 3876 5354 3882
rect 4934 2846 4986 2852
rect 4934 2788 4986 2794
rect 4842 2302 4894 2308
rect 4842 2244 4894 2250
rect 4658 2098 4710 2104
rect 4658 2040 4710 2046
rect 4670 1492 4698 2040
rect 4658 1486 4710 1492
rect 4658 1428 4710 1434
rect 4854 1424 4882 2244
rect 4842 1418 4894 1424
rect 4842 1360 4894 1366
rect 4946 948 4974 2788
rect 4934 942 4986 948
rect 4934 884 4986 890
rect 4566 806 4618 812
rect 4566 748 4618 754
rect 5314 336 5342 3876
rect 5774 2308 5802 6188
rect 81476 3290 81532 3299
rect 81476 3225 81532 3234
rect 81384 3154 81440 3163
rect 81306 3112 81384 3140
rect 8706 3050 8758 3056
rect 8706 2992 8758 2998
rect 36950 3050 37002 3056
rect 36950 2992 37002 2998
rect 7878 2506 7930 2512
rect 7876 2474 7878 2483
rect 7930 2474 7932 2483
rect 7876 2409 7932 2418
rect 5762 2302 5814 2308
rect 5762 2244 5814 2250
rect 8718 1667 8746 2992
rect 33730 2982 33782 2988
rect 33730 2924 33782 2930
rect 23978 2914 24030 2920
rect 19744 2882 19800 2891
rect 19744 2817 19800 2826
rect 22136 2882 22192 2891
rect 22136 2817 22192 2826
rect 23976 2882 23978 2891
rect 33742 2891 33770 2924
rect 34834 2914 34886 2920
rect 24030 2882 24032 2891
rect 23976 2817 24032 2826
rect 25080 2882 25136 2891
rect 25080 2817 25136 2826
rect 27472 2882 27528 2891
rect 27472 2817 27474 2826
rect 19758 2716 19786 2817
rect 22150 2784 22178 2817
rect 22138 2778 22190 2784
rect 22138 2720 22190 2726
rect 19746 2710 19798 2716
rect 19746 2652 19798 2658
rect 19470 2642 19522 2648
rect 19468 2610 19470 2619
rect 24622 2642 24674 2648
rect 19522 2610 19524 2619
rect 19468 2545 19524 2554
rect 24620 2610 24622 2619
rect 24674 2610 24676 2619
rect 25094 2580 25122 2817
rect 27526 2817 27528 2826
rect 31060 2882 31116 2891
rect 31060 2817 31116 2826
rect 33728 2882 33784 2891
rect 36962 2891 36990 2992
rect 53694 2982 53746 2988
rect 53694 2924 53746 2930
rect 34834 2856 34886 2862
rect 36948 2882 37004 2891
rect 33728 2817 33784 2826
rect 27474 2788 27526 2794
rect 24620 2545 24676 2554
rect 25082 2574 25134 2580
rect 25082 2516 25134 2522
rect 26002 2506 26054 2512
rect 26000 2474 26002 2483
rect 28394 2506 28446 2512
rect 26054 2474 26056 2483
rect 28394 2448 28446 2454
rect 26000 2409 26056 2418
rect 28406 2347 28434 2448
rect 31074 2444 31102 2817
rect 31062 2438 31114 2444
rect 31062 2380 31114 2386
rect 18272 2338 18328 2347
rect 18272 2273 18328 2282
rect 28392 2338 28448 2347
rect 28392 2273 28448 2282
rect 18286 2172 18314 2273
rect 19376 2202 19432 2211
rect 18274 2166 18326 2172
rect 19560 2202 19616 2211
rect 19432 2160 19560 2188
rect 19376 2137 19432 2146
rect 19560 2137 19616 2146
rect 26368 2202 26424 2211
rect 26368 2137 26424 2146
rect 18274 2108 18326 2114
rect 26382 1900 26410 2137
rect 26370 1894 26422 1900
rect 26370 1836 26422 1842
rect 8704 1658 8760 1667
rect 8704 1593 8760 1602
rect 22412 1658 22468 1667
rect 22412 1593 22468 1602
rect 24712 1658 24768 1667
rect 24712 1593 24768 1602
rect 29220 1658 29276 1667
rect 29220 1593 29276 1602
rect 5302 330 5354 336
rect 5302 272 5354 278
rect 4290 126 4342 132
rect 4290 68 4342 74
rect 8718 64 8746 1593
rect 22426 1220 22454 1593
rect 24726 1288 24754 1593
rect 29234 1492 29262 1593
rect 29222 1486 29274 1492
rect 29222 1428 29274 1434
rect 33084 1386 33140 1395
rect 33084 1321 33140 1330
rect 24714 1282 24766 1288
rect 24714 1224 24766 1230
rect 20850 1214 20902 1220
rect 20850 1156 20902 1162
rect 22414 1214 22466 1220
rect 22414 1156 22466 1162
rect 18918 1146 18970 1152
rect 18918 1088 18970 1094
rect 11834 1078 11886 1084
rect 11834 1020 11886 1026
rect 11846 987 11874 1020
rect 14410 1010 14462 1016
rect 11648 978 11704 987
rect 11832 978 11888 987
rect 11704 948 11782 964
rect 11704 942 11794 948
rect 11704 936 11742 942
rect 11648 913 11704 922
rect 11832 913 11888 922
rect 14408 978 14410 987
rect 18930 987 18958 1088
rect 20862 987 20890 1156
rect 33098 1084 33126 1321
rect 28302 1078 28354 1084
rect 28302 1020 28354 1026
rect 33086 1078 33138 1084
rect 33086 1020 33138 1026
rect 28314 987 28342 1020
rect 29406 1010 29458 1016
rect 14462 978 14464 987
rect 14408 913 14464 922
rect 16984 978 17040 987
rect 16984 913 17040 922
rect 18088 978 18144 987
rect 18088 913 18144 922
rect 18916 978 18972 987
rect 18916 913 18972 922
rect 20848 978 20904 987
rect 20848 913 20904 922
rect 21308 978 21364 987
rect 21308 913 21310 922
rect 11742 884 11794 890
rect 11754 472 11782 884
rect 16998 812 17026 913
rect 16986 806 17038 812
rect 16986 748 17038 754
rect 18102 608 18130 913
rect 21362 913 21364 922
rect 23424 978 23480 987
rect 23424 913 23480 922
rect 24252 978 24308 987
rect 24252 913 24308 922
rect 28300 978 28356 987
rect 28300 913 28356 922
rect 29404 978 29406 987
rect 29458 978 29460 987
rect 29404 913 29460 922
rect 31060 978 31116 987
rect 31060 913 31116 922
rect 31888 978 31944 987
rect 31888 913 31944 922
rect 32900 978 32956 987
rect 32900 913 32956 922
rect 34740 978 34796 987
rect 34740 913 34796 922
rect 21310 884 21362 890
rect 23438 880 23466 913
rect 24266 880 24294 913
rect 23426 874 23478 880
rect 23426 816 23478 822
rect 24254 874 24306 880
rect 24254 816 24306 822
rect 31074 812 31102 913
rect 31062 806 31114 812
rect 31062 748 31114 754
rect 31902 744 31930 913
rect 31890 738 31942 744
rect 20756 706 20812 715
rect 20756 641 20812 650
rect 29864 706 29920 715
rect 31890 680 31942 686
rect 32914 676 32942 913
rect 29864 641 29866 650
rect 18090 602 18142 608
rect 18090 544 18142 550
rect 11742 466 11794 472
rect 11742 408 11794 414
rect 20770 404 20798 641
rect 29918 641 29920 650
rect 32902 670 32954 676
rect 29866 612 29918 618
rect 32902 612 32954 618
rect 34754 608 34782 913
rect 34742 602 34794 608
rect 32440 570 32496 579
rect 34742 544 34794 550
rect 34846 540 34874 2856
rect 36948 2817 37004 2826
rect 38788 2882 38844 2891
rect 38788 2817 38790 2826
rect 38842 2817 38844 2826
rect 41364 2882 41420 2891
rect 41364 2817 41420 2826
rect 38790 2788 38842 2794
rect 37594 2778 37646 2784
rect 37594 2720 37646 2726
rect 35016 2202 35072 2211
rect 35016 2137 35018 2146
rect 35070 2137 35072 2146
rect 35018 2108 35070 2114
rect 36304 1658 36360 1667
rect 36304 1593 36360 1602
rect 36488 1658 36544 1667
rect 36488 1593 36544 1602
rect 36318 1424 36346 1593
rect 36306 1418 36358 1424
rect 36502 1395 36530 1593
rect 36306 1360 36358 1366
rect 36488 1386 36544 1395
rect 36488 1321 36544 1330
rect 37606 1016 37634 2720
rect 41378 2716 41406 2817
rect 41366 2710 41418 2716
rect 41366 2652 41418 2658
rect 53706 2619 53734 2924
rect 81306 2868 81334 3112
rect 81384 3089 81440 3098
rect 61974 2846 62026 2852
rect 61974 2788 62026 2794
rect 81214 2840 81334 2868
rect 50196 2610 50252 2619
rect 53692 2610 53748 2619
rect 50196 2545 50252 2554
rect 50474 2574 50526 2580
rect 50210 2444 50238 2545
rect 61986 2580 62014 2788
rect 78072 2746 78128 2755
rect 78072 2681 78128 2690
rect 53692 2545 53748 2554
rect 61974 2574 62026 2580
rect 50474 2516 50526 2522
rect 61974 2516 62026 2522
rect 50198 2438 50250 2444
rect 50198 2380 50250 2386
rect 41824 2202 41880 2211
rect 45228 2202 45284 2211
rect 41824 2137 41880 2146
rect 42470 2166 42522 2172
rect 39986 1758 40038 1764
rect 39986 1700 40038 1706
rect 37594 1010 37646 1016
rect 35292 978 35348 987
rect 37594 952 37646 958
rect 38328 978 38384 987
rect 35292 913 35348 922
rect 38328 913 38384 922
rect 35306 540 35334 913
rect 32440 505 32442 514
rect 32494 505 32496 514
rect 34834 534 34886 540
rect 32442 476 32494 482
rect 34834 476 34886 482
rect 35294 534 35346 540
rect 35294 476 35346 482
rect 38052 434 38108 443
rect 20758 398 20810 404
rect 38052 369 38108 378
rect 20758 340 20810 346
rect 38066 336 38094 369
rect 38342 336 38370 913
rect 39998 404 40026 1700
rect 41838 1560 41866 2137
rect 45228 2137 45284 2146
rect 46700 2202 46756 2211
rect 46700 2137 46756 2146
rect 47896 2202 47952 2211
rect 47896 2137 47952 2146
rect 49828 2202 49884 2211
rect 49828 2137 49884 2146
rect 50012 2202 50068 2211
rect 50012 2137 50068 2146
rect 42470 2108 42522 2114
rect 41826 1554 41878 1560
rect 41826 1496 41878 1502
rect 42482 1395 42510 2108
rect 45242 1424 45270 2137
rect 46714 2104 46742 2137
rect 46702 2098 46754 2104
rect 46702 2040 46754 2046
rect 47910 1832 47938 2137
rect 47898 1826 47950 1832
rect 47898 1768 47950 1774
rect 49842 1560 49870 2137
rect 49830 1554 49882 1560
rect 49830 1496 49882 1502
rect 45230 1418 45282 1424
rect 42284 1386 42340 1395
rect 42284 1321 42286 1330
rect 42338 1321 42340 1330
rect 42468 1386 42524 1395
rect 50026 1395 50054 2137
rect 45230 1360 45282 1366
rect 50012 1386 50068 1395
rect 42468 1321 42524 1330
rect 50012 1321 50068 1330
rect 42286 1292 42338 1298
rect 50486 987 50514 2516
rect 78086 2483 78114 2681
rect 78072 2474 78128 2483
rect 78072 2409 78128 2418
rect 54244 2338 54300 2347
rect 54244 2273 54300 2282
rect 54258 1628 54286 2273
rect 80740 1658 80796 1667
rect 54246 1622 54298 1628
rect 80740 1593 80796 1602
rect 54246 1564 54298 1570
rect 51486 1486 51538 1492
rect 51486 1428 51538 1434
rect 51498 1395 51526 1428
rect 80754 1395 80782 1593
rect 51484 1386 51540 1395
rect 51484 1321 51540 1330
rect 80740 1386 80796 1395
rect 80740 1321 80796 1330
rect 40076 978 40132 987
rect 40076 913 40132 922
rect 43940 978 43996 987
rect 43940 913 43996 922
rect 46148 978 46204 987
rect 46148 913 46204 922
rect 50472 978 50528 987
rect 50472 913 50528 922
rect 40090 404 40118 913
rect 39986 398 40038 404
rect 39986 340 40038 346
rect 40078 398 40130 404
rect 40078 340 40130 346
rect 38054 330 38106 336
rect 38054 272 38106 278
rect 38330 330 38382 336
rect 38330 272 38382 278
rect 43954 268 43982 913
rect 43942 262 43994 268
rect 43942 204 43994 210
rect 46162 200 46190 913
rect 46150 194 46202 200
rect 81214 171 81242 2840
rect 81292 2746 81348 2755
rect 81292 2681 81348 2690
rect 81386 2710 81438 2716
rect 81306 2240 81334 2681
rect 81386 2652 81438 2658
rect 81398 2444 81426 2652
rect 81386 2438 81438 2444
rect 81386 2380 81438 2386
rect 81294 2234 81346 2240
rect 81294 2176 81346 2182
rect 81490 2052 81518 3225
rect 81306 2024 81518 2052
rect 81306 307 81334 2024
rect 81292 298 81348 307
rect 81582 268 81610 7004
rect 81674 1152 81702 25568
rect 81662 1146 81714 1152
rect 81662 1088 81714 1094
rect 81766 851 81794 28492
rect 81752 842 81808 851
rect 81752 777 81808 786
rect 81858 336 81886 29444
rect 81950 1560 81978 56440
rect 82030 50106 82082 50112
rect 82030 50048 82082 50054
rect 82042 7068 82070 50048
rect 82122 48882 82174 48888
rect 82122 48824 82174 48830
rect 82030 7062 82082 7068
rect 82030 7004 82082 7010
rect 82030 6926 82082 6932
rect 82030 6868 82082 6874
rect 81938 1554 81990 1560
rect 81938 1496 81990 1502
rect 82042 540 82070 6868
rect 82134 1356 82162 48824
rect 82214 43646 82266 43652
rect 82214 43588 82266 43594
rect 82226 3056 82254 43588
rect 82306 39974 82358 39980
rect 82306 39916 82358 39922
rect 82214 3050 82266 3056
rect 82214 2992 82266 2998
rect 82122 1350 82174 1356
rect 82122 1292 82174 1298
rect 82318 676 82346 39916
rect 82398 35486 82450 35492
rect 82398 35428 82450 35434
rect 82410 6932 82438 35428
rect 82490 32086 82542 32092
rect 82490 32028 82542 32034
rect 82502 17851 82530 32028
rect 82594 19648 82622 93432
rect 82686 87852 82714 93500
rect 82778 92476 82806 94724
rect 83422 94720 83450 127364
rect 83606 96896 83634 130113
rect 83790 97796 83818 176761
rect 83868 175874 83924 175883
rect 83868 175809 83924 175818
rect 83882 98188 83910 175809
rect 83974 164896 84002 180592
rect 84158 179555 84186 186728
rect 84250 182411 84278 187369
rect 84790 187340 84842 187346
rect 84422 187126 84474 187132
rect 84422 187068 84474 187074
rect 84330 187058 84382 187064
rect 84330 187000 84382 187006
rect 84342 185432 84370 187000
rect 84330 185426 84382 185432
rect 84330 185368 84382 185374
rect 84236 182402 84292 182411
rect 84236 182337 84292 182346
rect 84434 182304 84462 187068
rect 84604 187026 84660 187035
rect 84604 186961 84660 186970
rect 84514 186650 84566 186656
rect 84514 186592 84566 186598
rect 84238 182298 84290 182304
rect 84238 182240 84290 182246
rect 84422 182298 84474 182304
rect 84422 182240 84474 182246
rect 84144 179546 84200 179555
rect 84144 179481 84200 179490
rect 84144 174786 84200 174795
rect 84144 174721 84200 174730
rect 84052 173562 84108 173571
rect 84052 173497 84108 173506
rect 83962 164890 84014 164896
rect 83962 164832 84014 164838
rect 83962 164550 84014 164556
rect 83962 164492 84014 164498
rect 83974 157931 84002 164492
rect 83960 157922 84016 157931
rect 83960 157857 84016 157866
rect 83962 150134 84014 150140
rect 83962 150076 84014 150082
rect 83974 149635 84002 150076
rect 83960 149626 84016 149635
rect 83960 149561 84016 149570
rect 83962 149182 84014 149188
rect 83962 149124 84014 149130
rect 83974 148547 84002 149124
rect 83960 148538 84016 148547
rect 83960 148473 84016 148482
rect 83962 147890 84014 147896
rect 83962 147832 84014 147838
rect 83974 147051 84002 147832
rect 83960 147042 84016 147051
rect 83960 146977 84016 146986
rect 83962 146598 84014 146604
rect 83962 146540 84014 146546
rect 83974 145827 84002 146540
rect 83960 145818 84016 145827
rect 83960 145753 84016 145762
rect 83962 145306 84014 145312
rect 83962 145248 84014 145254
rect 83974 144739 84002 145248
rect 83960 144730 84016 144739
rect 83960 144665 84016 144674
rect 83960 121882 84016 121891
rect 83960 121817 84016 121826
rect 83974 116684 84002 121817
rect 83962 116678 84014 116684
rect 83962 116620 84014 116626
rect 83960 115898 84016 115907
rect 83960 115833 84016 115842
rect 83974 111992 84002 115833
rect 83962 111986 84014 111992
rect 83962 111928 84014 111934
rect 83960 109370 84016 109379
rect 83960 109305 83962 109314
rect 84014 109305 84016 109314
rect 83962 109276 84014 109282
rect 83960 108282 84016 108291
rect 83960 108217 84016 108226
rect 83974 108184 84002 108217
rect 83962 108178 84014 108184
rect 83962 108120 84014 108126
rect 83960 107330 84016 107339
rect 83960 107265 84016 107274
rect 83870 98182 83922 98188
rect 83870 98124 83922 98130
rect 83790 97768 83910 97796
rect 83776 97674 83832 97683
rect 83776 97609 83832 97618
rect 83790 97576 83818 97609
rect 83778 97570 83830 97576
rect 83778 97512 83830 97518
rect 83790 97139 83818 97512
rect 83776 97130 83832 97139
rect 83698 97088 83776 97116
rect 83594 96890 83646 96896
rect 83500 96858 83556 96867
rect 83594 96832 83646 96838
rect 83500 96793 83556 96802
rect 83410 94714 83462 94720
rect 83410 94656 83462 94662
rect 83224 94546 83280 94555
rect 83224 94481 83280 94490
rect 82766 92470 82818 92476
rect 82766 92412 82818 92418
rect 82674 87846 82726 87852
rect 82674 87788 82726 87794
rect 83238 80984 83266 94481
rect 83410 93286 83462 93292
rect 83410 93228 83462 93234
rect 83318 93218 83370 93224
rect 83318 93160 83370 93166
rect 83042 80978 83094 80984
rect 83042 80920 83094 80926
rect 83226 80978 83278 80984
rect 83226 80920 83278 80926
rect 83054 71956 83082 80920
rect 83330 76195 83358 93160
rect 83422 84792 83450 93228
rect 83410 84786 83462 84792
rect 83410 84728 83462 84734
rect 83316 76186 83372 76195
rect 83316 76121 83372 76130
rect 83054 71928 83174 71956
rect 83146 63139 83174 71928
rect 83132 63130 83188 63139
rect 83132 63065 83188 63074
rect 83132 62994 83188 63003
rect 83132 62929 83188 62938
rect 83146 56572 83174 62929
rect 83316 61634 83372 61643
rect 83316 61569 83372 61578
rect 83134 56566 83186 56572
rect 83134 56508 83186 56514
rect 83134 56430 83186 56436
rect 83134 56372 83186 56378
rect 83146 52628 83174 56372
rect 82858 52622 82910 52628
rect 82858 52564 82910 52570
rect 83134 52622 83186 52628
rect 83134 52564 83186 52570
rect 82870 43691 82898 52564
rect 82856 43682 82912 43691
rect 82856 43617 82912 43626
rect 83040 43682 83096 43691
rect 83040 43617 83096 43626
rect 83054 43532 83082 43617
rect 83054 43504 83266 43532
rect 83132 38786 83188 38795
rect 83132 38721 83188 38730
rect 83040 37698 83096 37707
rect 83040 37633 83096 37642
rect 82950 30930 83002 30936
rect 82950 30872 83002 30878
rect 82858 28210 82910 28216
rect 82672 28178 82728 28187
rect 82858 28152 82910 28158
rect 82672 28113 82728 28122
rect 82686 24379 82714 28113
rect 82672 24370 82728 24379
rect 82672 24305 82728 24314
rect 82672 24234 82728 24243
rect 82672 24169 82728 24178
rect 82582 19642 82634 19648
rect 82582 19584 82634 19590
rect 82488 17842 82544 17851
rect 82488 17777 82544 17786
rect 82686 15403 82714 24169
rect 82764 17842 82820 17851
rect 82764 17777 82820 17786
rect 82672 15394 82728 15403
rect 82672 15329 82728 15338
rect 82778 8875 82806 17777
rect 82580 8866 82636 8875
rect 82580 8801 82582 8810
rect 82634 8801 82636 8810
rect 82764 8866 82820 8875
rect 82764 8801 82820 8810
rect 82582 8772 82634 8778
rect 82488 8594 82544 8603
rect 82488 8529 82544 8538
rect 82398 6926 82450 6932
rect 82398 6868 82450 6874
rect 82398 3662 82450 3668
rect 82398 3604 82450 3610
rect 82410 3260 82438 3604
rect 82398 3254 82450 3260
rect 82398 3196 82450 3202
rect 82410 2716 82438 3196
rect 82398 2710 82450 2716
rect 82398 2652 82450 2658
rect 82306 670 82358 676
rect 82306 612 82358 618
rect 82030 534 82082 540
rect 82030 476 82082 482
rect 82502 404 82530 8529
rect 82582 7606 82634 7612
rect 82582 7548 82634 7554
rect 82594 1803 82622 7548
rect 82672 6146 82728 6155
rect 82672 6081 82728 6090
rect 82686 3027 82714 6081
rect 82764 3834 82820 3843
rect 82764 3769 82820 3778
rect 82778 3668 82806 3769
rect 82766 3662 82818 3668
rect 82766 3604 82818 3610
rect 82766 3526 82818 3532
rect 82766 3468 82818 3474
rect 82672 3018 82728 3027
rect 82672 2953 82674 2962
rect 82726 2953 82728 2962
rect 82674 2924 82726 2930
rect 82686 2893 82714 2924
rect 82580 1794 82636 1803
rect 82580 1729 82636 1738
rect 82778 579 82806 3468
rect 82870 1220 82898 28152
rect 82962 1288 82990 30872
rect 82950 1282 83002 1288
rect 82950 1224 83002 1230
rect 82858 1214 82910 1220
rect 82858 1156 82910 1162
rect 83054 812 83082 37633
rect 83042 806 83094 812
rect 83042 748 83094 754
rect 83146 744 83174 38721
rect 83238 28284 83266 43504
rect 83226 28278 83278 28284
rect 83226 28220 83278 28226
rect 83224 27906 83280 27915
rect 83224 27841 83280 27850
rect 83238 948 83266 27841
rect 83330 1628 83358 61569
rect 83408 53338 83464 53347
rect 83408 53273 83464 53282
rect 83318 1622 83370 1628
rect 83318 1564 83370 1570
rect 83226 942 83278 948
rect 83226 884 83278 890
rect 83134 738 83186 744
rect 83134 680 83186 686
rect 82764 570 82820 579
rect 82764 505 82820 514
rect 82490 398 82542 404
rect 82490 340 82542 346
rect 81846 330 81898 336
rect 81846 272 81898 278
rect 81292 233 81348 242
rect 81570 262 81622 268
rect 81570 204 81622 210
rect 83422 200 83450 53273
rect 83514 28187 83542 96793
rect 83592 96314 83648 96323
rect 83592 96249 83648 96258
rect 83606 88056 83634 96249
rect 83594 88050 83646 88056
rect 83594 87992 83646 87998
rect 83592 51842 83648 51851
rect 83592 51777 83648 51786
rect 83500 28178 83556 28187
rect 83500 28113 83556 28122
rect 83502 26034 83554 26040
rect 83502 25976 83554 25982
rect 83514 25739 83542 25976
rect 83500 25730 83556 25739
rect 83500 25665 83556 25674
rect 83514 20260 83542 25665
rect 83502 20254 83554 20260
rect 83502 20196 83554 20202
rect 83502 20050 83554 20056
rect 83502 19992 83554 19998
rect 83514 18424 83542 19992
rect 83502 18418 83554 18424
rect 83502 18360 83554 18366
rect 83500 17842 83556 17851
rect 83500 17777 83556 17786
rect 83514 8875 83542 17777
rect 83500 8866 83556 8875
rect 83500 8801 83556 8810
rect 83606 3736 83634 51777
rect 83698 32024 83726 97088
rect 83776 97065 83832 97074
rect 83778 96890 83830 96896
rect 83776 96858 83778 96867
rect 83830 96858 83832 96867
rect 83776 96793 83832 96802
rect 83882 96556 83910 97768
rect 83974 97644 84002 107265
rect 84066 102744 84094 173497
rect 84054 102738 84106 102744
rect 84054 102680 84106 102686
rect 84158 102556 84186 174721
rect 84250 164828 84278 182240
rect 84422 182162 84474 182168
rect 84422 182104 84474 182110
rect 84330 180190 84382 180196
rect 84330 180132 84382 180138
rect 84342 173668 84370 180132
rect 84330 173662 84382 173668
rect 84330 173604 84382 173610
rect 84330 171078 84382 171084
rect 84330 171020 84382 171026
rect 84238 164822 84290 164828
rect 84238 164764 84290 164770
rect 84342 164708 84370 171020
rect 84434 165003 84462 182104
rect 84420 164994 84476 165003
rect 84420 164929 84476 164938
rect 84422 164890 84474 164896
rect 84422 164832 84474 164838
rect 84250 164680 84370 164708
rect 84250 164556 84278 164680
rect 84434 164572 84462 164832
rect 84342 164556 84462 164572
rect 84238 164550 84290 164556
rect 84238 164492 84290 164498
rect 84330 164550 84462 164556
rect 84382 164544 84462 164550
rect 84330 164492 84382 164498
rect 84236 164450 84292 164459
rect 84236 164385 84292 164394
rect 84250 159268 84278 164385
rect 84420 164314 84476 164323
rect 84420 164249 84476 164258
rect 84330 162850 84382 162856
rect 84330 162792 84382 162798
rect 84342 162691 84370 162792
rect 84328 162682 84384 162691
rect 84328 162617 84384 162626
rect 84330 161830 84382 161836
rect 84330 161772 84382 161778
rect 84342 159427 84370 161772
rect 84434 160680 84462 164249
rect 84422 160674 84474 160680
rect 84422 160616 84474 160622
rect 84526 160204 84554 186592
rect 84618 182168 84646 186961
rect 84698 186854 84750 186860
rect 84698 186796 84750 186802
rect 84606 182162 84658 182168
rect 84606 182104 84658 182110
rect 84604 181994 84660 182003
rect 84604 181929 84660 181938
rect 84618 178603 84646 181929
rect 84604 178594 84660 178603
rect 84710 178564 84738 186796
rect 84802 185539 84830 187340
rect 84890 186958 85186 186978
rect 84946 186956 84970 186958
rect 85026 186956 85050 186958
rect 85106 186956 85130 186958
rect 84968 186904 84970 186956
rect 85032 186904 85044 186956
rect 85106 186904 85108 186956
rect 84946 186902 84970 186904
rect 85026 186902 85050 186904
rect 85106 186902 85130 186904
rect 84890 186882 85186 186902
rect 85156 186754 85212 186763
rect 85156 186689 85158 186698
rect 85210 186689 85212 186698
rect 85158 186660 85210 186666
rect 86890 186414 87186 186434
rect 86946 186412 86970 186414
rect 87026 186412 87050 186414
rect 87106 186412 87130 186414
rect 86968 186360 86970 186412
rect 87032 186360 87044 186412
rect 87106 186360 87108 186412
rect 86946 186358 86970 186360
rect 87026 186358 87050 186360
rect 87106 186358 87130 186360
rect 86890 186338 87186 186358
rect 84890 185870 85186 185890
rect 84946 185868 84970 185870
rect 85026 185868 85050 185870
rect 85106 185868 85130 185870
rect 84968 185816 84970 185868
rect 85032 185816 85044 185868
rect 85106 185816 85108 185868
rect 84946 185814 84970 185816
rect 85026 185814 85050 185816
rect 85106 185814 85130 185816
rect 84890 185794 85186 185814
rect 84788 185530 84844 185539
rect 84788 185465 84844 185474
rect 84790 185426 84842 185432
rect 84790 185368 84842 185374
rect 84604 178529 84660 178538
rect 84698 178558 84750 178564
rect 84698 178500 84750 178506
rect 84698 178354 84750 178360
rect 84698 178296 84750 178302
rect 84606 175634 84658 175640
rect 84606 175576 84658 175582
rect 84618 164867 84646 175576
rect 84604 164858 84660 164867
rect 84604 164793 84660 164802
rect 84606 164754 84658 164760
rect 84606 164696 84658 164702
rect 84618 161836 84646 164696
rect 84606 161830 84658 161836
rect 84606 161772 84658 161778
rect 84606 160742 84658 160748
rect 84606 160684 84658 160690
rect 84618 160515 84646 160684
rect 84604 160506 84660 160515
rect 84604 160441 84660 160450
rect 84514 160198 84566 160204
rect 84514 160140 84566 160146
rect 84514 159994 84566 160000
rect 84514 159936 84566 159942
rect 84328 159418 84384 159427
rect 84328 159353 84384 159362
rect 84250 159240 84462 159268
rect 84434 155619 84462 159240
rect 84420 155610 84476 155619
rect 84420 155545 84476 155554
rect 84526 153035 84554 159936
rect 84512 153026 84568 153035
rect 84512 152961 84568 152970
rect 84710 151947 84738 178296
rect 84802 175640 84830 185368
rect 86890 185326 87186 185346
rect 86946 185324 86970 185326
rect 87026 185324 87050 185326
rect 87106 185324 87130 185326
rect 86968 185272 86970 185324
rect 87032 185272 87044 185324
rect 87106 185272 87108 185324
rect 86946 185270 86970 185272
rect 87026 185270 87050 185272
rect 87106 185270 87130 185272
rect 86890 185250 87186 185270
rect 84890 184782 85186 184802
rect 84946 184780 84970 184782
rect 85026 184780 85050 184782
rect 85106 184780 85130 184782
rect 84968 184728 84970 184780
rect 85032 184728 85044 184780
rect 85106 184728 85108 184780
rect 84946 184726 84970 184728
rect 85026 184726 85050 184728
rect 85106 184726 85130 184728
rect 84890 184706 85186 184726
rect 86890 184238 87186 184258
rect 86946 184236 86970 184238
rect 87026 184236 87050 184238
rect 87106 184236 87130 184238
rect 86968 184184 86970 184236
rect 87032 184184 87044 184236
rect 87106 184184 87108 184236
rect 86946 184182 86970 184184
rect 87026 184182 87050 184184
rect 87106 184182 87130 184184
rect 86890 184162 87186 184182
rect 84890 183694 85186 183714
rect 84946 183692 84970 183694
rect 85026 183692 85050 183694
rect 85106 183692 85130 183694
rect 84968 183640 84970 183692
rect 85032 183640 85044 183692
rect 85106 183640 85108 183692
rect 84946 183638 84970 183640
rect 85026 183638 85050 183640
rect 85106 183638 85130 183640
rect 84890 183618 85186 183638
rect 86890 183150 87186 183170
rect 86946 183148 86970 183150
rect 87026 183148 87050 183150
rect 87106 183148 87130 183150
rect 86968 183096 86970 183148
rect 87032 183096 87044 183148
rect 87106 183096 87108 183148
rect 86946 183094 86970 183096
rect 87026 183094 87050 183096
rect 87106 183094 87130 183096
rect 86890 183074 87186 183094
rect 84890 182606 85186 182626
rect 84946 182604 84970 182606
rect 85026 182604 85050 182606
rect 85106 182604 85130 182606
rect 84968 182552 84970 182604
rect 85032 182552 85044 182604
rect 85106 182552 85108 182604
rect 84946 182550 84970 182552
rect 85026 182550 85050 182552
rect 85106 182550 85130 182552
rect 84890 182530 85186 182550
rect 86890 182062 87186 182082
rect 86946 182060 86970 182062
rect 87026 182060 87050 182062
rect 87106 182060 87130 182062
rect 86968 182008 86970 182060
rect 87032 182008 87044 182060
rect 87106 182008 87108 182060
rect 86946 182006 86970 182008
rect 87026 182006 87050 182008
rect 87106 182006 87130 182008
rect 86890 181986 87186 182006
rect 84890 181518 85186 181538
rect 84946 181516 84970 181518
rect 85026 181516 85050 181518
rect 85106 181516 85130 181518
rect 84968 181464 84970 181516
rect 85032 181464 85044 181516
rect 85106 181464 85108 181516
rect 84946 181462 84970 181464
rect 85026 181462 85050 181464
rect 85106 181462 85130 181464
rect 84890 181442 85186 181462
rect 86890 180974 87186 180994
rect 86946 180972 86970 180974
rect 87026 180972 87050 180974
rect 87106 180972 87130 180974
rect 86968 180920 86970 180972
rect 87032 180920 87044 180972
rect 87106 180920 87108 180972
rect 86946 180918 86970 180920
rect 87026 180918 87050 180920
rect 87106 180918 87130 180920
rect 86890 180898 87186 180918
rect 84890 180430 85186 180450
rect 84946 180428 84970 180430
rect 85026 180428 85050 180430
rect 85106 180428 85130 180430
rect 84968 180376 84970 180428
rect 85032 180376 85044 180428
rect 85106 180376 85108 180428
rect 84946 180374 84970 180376
rect 85026 180374 85050 180376
rect 85106 180374 85130 180376
rect 84890 180354 85186 180374
rect 86890 179886 87186 179906
rect 86946 179884 86970 179886
rect 87026 179884 87050 179886
rect 87106 179884 87130 179886
rect 86968 179832 86970 179884
rect 87032 179832 87044 179884
rect 87106 179832 87108 179884
rect 86946 179830 86970 179832
rect 87026 179830 87050 179832
rect 87106 179830 87130 179832
rect 86890 179810 87186 179830
rect 84890 179342 85186 179362
rect 84946 179340 84970 179342
rect 85026 179340 85050 179342
rect 85106 179340 85130 179342
rect 84968 179288 84970 179340
rect 85032 179288 85044 179340
rect 85106 179288 85108 179340
rect 84946 179286 84970 179288
rect 85026 179286 85050 179288
rect 85106 179286 85130 179288
rect 84890 179266 85186 179286
rect 86890 178798 87186 178818
rect 86946 178796 86970 178798
rect 87026 178796 87050 178798
rect 87106 178796 87130 178798
rect 86968 178744 86970 178796
rect 87032 178744 87044 178796
rect 87106 178744 87108 178796
rect 86946 178742 86970 178744
rect 87026 178742 87050 178744
rect 87106 178742 87130 178744
rect 86890 178722 87186 178742
rect 84890 178254 85186 178274
rect 84946 178252 84970 178254
rect 85026 178252 85050 178254
rect 85106 178252 85130 178254
rect 84968 178200 84970 178252
rect 85032 178200 85044 178252
rect 85106 178200 85108 178252
rect 84946 178198 84970 178200
rect 85026 178198 85050 178200
rect 85106 178198 85130 178200
rect 84890 178178 85186 178198
rect 86890 177710 87186 177730
rect 86946 177708 86970 177710
rect 87026 177708 87050 177710
rect 87106 177708 87130 177710
rect 86968 177656 86970 177708
rect 87032 177656 87044 177708
rect 87106 177656 87108 177708
rect 86946 177654 86970 177656
rect 87026 177654 87050 177656
rect 87106 177654 87130 177656
rect 86890 177634 87186 177654
rect 84890 177166 85186 177186
rect 84946 177164 84970 177166
rect 85026 177164 85050 177166
rect 85106 177164 85130 177166
rect 84968 177112 84970 177164
rect 85032 177112 85044 177164
rect 85106 177112 85108 177164
rect 84946 177110 84970 177112
rect 85026 177110 85050 177112
rect 85106 177110 85130 177112
rect 84890 177090 85186 177110
rect 86890 176622 87186 176642
rect 86946 176620 86970 176622
rect 87026 176620 87050 176622
rect 87106 176620 87130 176622
rect 86968 176568 86970 176620
rect 87032 176568 87044 176620
rect 87106 176568 87108 176620
rect 86946 176566 86970 176568
rect 87026 176566 87050 176568
rect 87106 176566 87130 176568
rect 86890 176546 87186 176566
rect 84890 176078 85186 176098
rect 84946 176076 84970 176078
rect 85026 176076 85050 176078
rect 85106 176076 85130 176078
rect 84968 176024 84970 176076
rect 85032 176024 85044 176076
rect 85106 176024 85108 176076
rect 84946 176022 84970 176024
rect 85026 176022 85050 176024
rect 85106 176022 85130 176024
rect 84890 176002 85186 176022
rect 84790 175634 84842 175640
rect 84790 175576 84842 175582
rect 86890 175534 87186 175554
rect 86946 175532 86970 175534
rect 87026 175532 87050 175534
rect 87106 175532 87130 175534
rect 86968 175480 86970 175532
rect 87032 175480 87044 175532
rect 87106 175480 87108 175532
rect 86946 175478 86970 175480
rect 87026 175478 87050 175480
rect 87106 175478 87130 175480
rect 86890 175458 87186 175478
rect 84890 174990 85186 175010
rect 84946 174988 84970 174990
rect 85026 174988 85050 174990
rect 85106 174988 85130 174990
rect 84968 174936 84970 174988
rect 85032 174936 85044 174988
rect 85106 174936 85108 174988
rect 84946 174934 84970 174936
rect 85026 174934 85050 174936
rect 85106 174934 85130 174936
rect 84890 174914 85186 174934
rect 86890 174446 87186 174466
rect 86946 174444 86970 174446
rect 87026 174444 87050 174446
rect 87106 174444 87130 174446
rect 86968 174392 86970 174444
rect 87032 174392 87044 174444
rect 87106 174392 87108 174444
rect 86946 174390 86970 174392
rect 87026 174390 87050 174392
rect 87106 174390 87130 174392
rect 86890 174370 87186 174390
rect 84890 173902 85186 173922
rect 84946 173900 84970 173902
rect 85026 173900 85050 173902
rect 85106 173900 85130 173902
rect 84968 173848 84970 173900
rect 85032 173848 85044 173900
rect 85106 173848 85108 173900
rect 84946 173846 84970 173848
rect 85026 173846 85050 173848
rect 85106 173846 85130 173848
rect 84890 173826 85186 173846
rect 84790 173662 84842 173668
rect 84790 173604 84842 173610
rect 84802 171084 84830 173604
rect 86890 173358 87186 173378
rect 86946 173356 86970 173358
rect 87026 173356 87050 173358
rect 87106 173356 87130 173358
rect 86968 173304 86970 173356
rect 87032 173304 87044 173356
rect 87106 173304 87108 173356
rect 86946 173302 86970 173304
rect 87026 173302 87050 173304
rect 87106 173302 87130 173304
rect 86890 173282 87186 173302
rect 84890 172814 85186 172834
rect 84946 172812 84970 172814
rect 85026 172812 85050 172814
rect 85106 172812 85130 172814
rect 84968 172760 84970 172812
rect 85032 172760 85044 172812
rect 85106 172760 85108 172812
rect 84946 172758 84970 172760
rect 85026 172758 85050 172760
rect 85106 172758 85130 172760
rect 84890 172738 85186 172758
rect 86890 172270 87186 172290
rect 86946 172268 86970 172270
rect 87026 172268 87050 172270
rect 87106 172268 87130 172270
rect 86968 172216 86970 172268
rect 87032 172216 87044 172268
rect 87106 172216 87108 172268
rect 86946 172214 86970 172216
rect 87026 172214 87050 172216
rect 87106 172214 87130 172216
rect 86890 172194 87186 172214
rect 84890 171726 85186 171746
rect 84946 171724 84970 171726
rect 85026 171724 85050 171726
rect 85106 171724 85130 171726
rect 84968 171672 84970 171724
rect 85032 171672 85044 171724
rect 85106 171672 85108 171724
rect 84946 171670 84970 171672
rect 85026 171670 85050 171672
rect 85106 171670 85130 171672
rect 84890 171650 85186 171670
rect 86890 171182 87186 171202
rect 86946 171180 86970 171182
rect 87026 171180 87050 171182
rect 87106 171180 87130 171182
rect 86968 171128 86970 171180
rect 87032 171128 87044 171180
rect 87106 171128 87108 171180
rect 86946 171126 86970 171128
rect 87026 171126 87050 171128
rect 87106 171126 87130 171128
rect 86890 171106 87186 171126
rect 84790 171078 84842 171084
rect 84790 171020 84842 171026
rect 84788 170978 84844 170987
rect 84788 170913 84844 170922
rect 84696 151938 84752 151947
rect 84696 151873 84752 151882
rect 84238 143878 84290 143884
rect 84238 143820 84290 143826
rect 84250 143787 84278 143820
rect 84236 143778 84292 143787
rect 84236 143713 84292 143722
rect 84512 142146 84568 142155
rect 84512 142081 84568 142090
rect 84236 138338 84292 138347
rect 84236 138273 84292 138282
rect 84250 137696 84278 138273
rect 84238 137690 84290 137696
rect 84238 137632 84290 137638
rect 84420 133850 84476 133859
rect 84420 133785 84476 133794
rect 84328 132898 84384 132907
rect 84328 132833 84384 132842
rect 84236 131810 84292 131819
rect 84236 131745 84292 131754
rect 84250 127428 84278 131745
rect 84238 127422 84290 127428
rect 84238 127364 84290 127370
rect 84236 125282 84292 125291
rect 84236 125217 84292 125226
rect 84250 124776 84278 125217
rect 84238 124770 84290 124776
rect 84238 124712 84290 124718
rect 84342 120900 84370 132833
rect 84434 128652 84462 133785
rect 84526 129944 84554 142081
rect 84604 139834 84660 139843
rect 84604 139769 84660 139778
rect 84514 129938 84566 129944
rect 84514 129880 84566 129886
rect 84422 128646 84474 128652
rect 84422 128588 84474 128594
rect 84512 127866 84568 127875
rect 84512 127801 84568 127810
rect 84420 124194 84476 124203
rect 84420 124129 84476 124138
rect 84434 123960 84462 124129
rect 84422 123954 84474 123960
rect 84422 123896 84474 123902
rect 84420 122970 84476 122979
rect 84420 122905 84476 122914
rect 84330 120894 84382 120900
rect 84330 120836 84382 120842
rect 84236 120250 84292 120259
rect 84236 120185 84292 120194
rect 84250 119676 84278 120185
rect 84238 119670 84290 119676
rect 84238 119612 84290 119618
rect 84328 118210 84384 118219
rect 84328 118145 84384 118154
rect 84236 116986 84292 116995
rect 84236 116921 84292 116930
rect 84250 106620 84278 116921
rect 84342 115596 84370 118145
rect 84330 115590 84382 115596
rect 84330 115532 84382 115538
rect 84328 114810 84384 114819
rect 84328 114745 84384 114754
rect 84342 114712 84370 114745
rect 84330 114706 84382 114712
rect 84330 114648 84382 114654
rect 84328 113314 84384 113323
rect 84328 113249 84384 113258
rect 84238 106614 84290 106620
rect 84238 106556 84290 106562
rect 84236 106242 84292 106251
rect 84236 106177 84292 106186
rect 84066 102528 84186 102556
rect 84066 100568 84094 102528
rect 84144 102434 84200 102443
rect 84144 102369 84200 102378
rect 84054 100562 84106 100568
rect 84054 100504 84106 100510
rect 84054 100358 84106 100364
rect 84054 100300 84106 100306
rect 83962 97638 84014 97644
rect 83962 97580 84014 97586
rect 84066 97388 84094 100300
rect 83974 97360 84094 97388
rect 83870 96550 83922 96556
rect 83870 96492 83922 96498
rect 83778 96346 83830 96352
rect 83776 96314 83778 96323
rect 83870 96346 83922 96352
rect 83830 96314 83832 96323
rect 83870 96288 83922 96294
rect 83776 96249 83832 96258
rect 83882 94011 83910 96288
rect 83974 94652 84002 97360
rect 84158 97252 84186 102369
rect 84066 97224 84186 97252
rect 84066 95196 84094 97224
rect 84144 97130 84200 97139
rect 84144 97065 84146 97074
rect 84198 97065 84200 97074
rect 84146 97036 84198 97042
rect 84158 96731 84186 97036
rect 84250 96828 84278 106177
rect 84342 101656 84370 113249
rect 84330 101650 84382 101656
rect 84330 101592 84382 101598
rect 84330 100562 84382 100568
rect 84330 100504 84382 100510
rect 84342 98052 84370 100504
rect 84330 98046 84382 98052
rect 84330 97988 84382 97994
rect 84328 97946 84384 97955
rect 84328 97881 84384 97890
rect 84238 96822 84290 96828
rect 84238 96764 84290 96770
rect 84144 96722 84200 96731
rect 84144 96657 84200 96666
rect 84146 96550 84198 96556
rect 84146 96492 84198 96498
rect 84158 96012 84186 96492
rect 84146 96006 84198 96012
rect 84146 95948 84198 95954
rect 84054 95190 84106 95196
rect 84054 95132 84106 95138
rect 83962 94646 84014 94652
rect 83962 94588 84014 94594
rect 84158 94555 84186 95948
rect 84144 94546 84200 94555
rect 84144 94481 84200 94490
rect 84342 94380 84370 97881
rect 84434 96420 84462 122905
rect 84526 102880 84554 127801
rect 84514 102874 84566 102880
rect 84514 102816 84566 102822
rect 84514 102738 84566 102744
rect 84514 102680 84566 102686
rect 84526 97644 84554 102680
rect 84618 100244 84646 139769
rect 84696 135074 84752 135083
rect 84696 135009 84752 135018
rect 84710 100364 84738 135009
rect 84802 103492 84830 170913
rect 84890 170638 85186 170658
rect 84946 170636 84970 170638
rect 85026 170636 85050 170638
rect 85106 170636 85130 170638
rect 84968 170584 84970 170636
rect 85032 170584 85044 170636
rect 85106 170584 85108 170636
rect 84946 170582 84970 170584
rect 85026 170582 85050 170584
rect 85106 170582 85130 170584
rect 84890 170562 85186 170582
rect 86890 170094 87186 170114
rect 86946 170092 86970 170094
rect 87026 170092 87050 170094
rect 87106 170092 87130 170094
rect 86968 170040 86970 170092
rect 87032 170040 87044 170092
rect 87106 170040 87108 170092
rect 86946 170038 86970 170040
rect 87026 170038 87050 170040
rect 87106 170038 87130 170040
rect 86890 170018 87186 170038
rect 84890 169550 85186 169570
rect 84946 169548 84970 169550
rect 85026 169548 85050 169550
rect 85106 169548 85130 169550
rect 84968 169496 84970 169548
rect 85032 169496 85044 169548
rect 85106 169496 85108 169548
rect 84946 169494 84970 169496
rect 85026 169494 85050 169496
rect 85106 169494 85130 169496
rect 84890 169474 85186 169494
rect 86890 169006 87186 169026
rect 86946 169004 86970 169006
rect 87026 169004 87050 169006
rect 87106 169004 87130 169006
rect 86968 168952 86970 169004
rect 87032 168952 87044 169004
rect 87106 168952 87108 169004
rect 86946 168950 86970 168952
rect 87026 168950 87050 168952
rect 87106 168950 87130 168952
rect 86890 168930 87186 168950
rect 84890 168462 85186 168482
rect 84946 168460 84970 168462
rect 85026 168460 85050 168462
rect 85106 168460 85130 168462
rect 84968 168408 84970 168460
rect 85032 168408 85044 168460
rect 85106 168408 85108 168460
rect 84946 168406 84970 168408
rect 85026 168406 85050 168408
rect 85106 168406 85130 168408
rect 84890 168386 85186 168406
rect 86890 167918 87186 167938
rect 86946 167916 86970 167918
rect 87026 167916 87050 167918
rect 87106 167916 87130 167918
rect 86968 167864 86970 167916
rect 87032 167864 87044 167916
rect 87106 167864 87108 167916
rect 86946 167862 86970 167864
rect 87026 167862 87050 167864
rect 87106 167862 87130 167864
rect 86890 167842 87186 167862
rect 84890 167374 85186 167394
rect 84946 167372 84970 167374
rect 85026 167372 85050 167374
rect 85106 167372 85130 167374
rect 84968 167320 84970 167372
rect 85032 167320 85044 167372
rect 85106 167320 85108 167372
rect 84946 167318 84970 167320
rect 85026 167318 85050 167320
rect 85106 167318 85130 167320
rect 84890 167298 85186 167318
rect 86890 166830 87186 166850
rect 86946 166828 86970 166830
rect 87026 166828 87050 166830
rect 87106 166828 87130 166830
rect 86968 166776 86970 166828
rect 87032 166776 87044 166828
rect 87106 166776 87108 166828
rect 86946 166774 86970 166776
rect 87026 166774 87050 166776
rect 87106 166774 87130 166776
rect 86890 166754 87186 166774
rect 84890 166286 85186 166306
rect 84946 166284 84970 166286
rect 85026 166284 85050 166286
rect 85106 166284 85130 166286
rect 84968 166232 84970 166284
rect 85032 166232 85044 166284
rect 85106 166232 85108 166284
rect 84946 166230 84970 166232
rect 85026 166230 85050 166232
rect 85106 166230 85130 166232
rect 84890 166210 85186 166230
rect 86890 165742 87186 165762
rect 86946 165740 86970 165742
rect 87026 165740 87050 165742
rect 87106 165740 87130 165742
rect 86968 165688 86970 165740
rect 87032 165688 87044 165740
rect 87106 165688 87108 165740
rect 86946 165686 86970 165688
rect 87026 165686 87050 165688
rect 87106 165686 87130 165688
rect 86890 165666 87186 165686
rect 84890 165198 85186 165218
rect 84946 165196 84970 165198
rect 85026 165196 85050 165198
rect 85106 165196 85130 165198
rect 84968 165144 84970 165196
rect 85032 165144 85044 165196
rect 85106 165144 85108 165196
rect 84946 165142 84970 165144
rect 85026 165142 85050 165144
rect 85106 165142 85130 165144
rect 84890 165122 85186 165142
rect 86890 164654 87186 164674
rect 86946 164652 86970 164654
rect 87026 164652 87050 164654
rect 87106 164652 87130 164654
rect 86968 164600 86970 164652
rect 87032 164600 87044 164652
rect 87106 164600 87108 164652
rect 86946 164598 86970 164600
rect 87026 164598 87050 164600
rect 87106 164598 87130 164600
rect 86890 164578 87186 164598
rect 85158 164550 85210 164556
rect 85158 164492 85210 164498
rect 85170 164300 85198 164492
rect 85170 164272 85290 164300
rect 84890 164110 85186 164130
rect 84946 164108 84970 164110
rect 85026 164108 85050 164110
rect 85106 164108 85130 164110
rect 84968 164056 84970 164108
rect 85032 164056 85044 164108
rect 85106 164056 85108 164108
rect 84946 164054 84970 164056
rect 85026 164054 85050 164056
rect 85106 164054 85130 164056
rect 84890 164034 85186 164054
rect 85158 163938 85210 163944
rect 85156 163906 85158 163915
rect 85210 163906 85212 163915
rect 85156 163841 85212 163850
rect 84890 163022 85186 163042
rect 84946 163020 84970 163022
rect 85026 163020 85050 163022
rect 85106 163020 85130 163022
rect 84968 162968 84970 163020
rect 85032 162968 85044 163020
rect 85106 162968 85108 163020
rect 84946 162966 84970 162968
rect 85026 162966 85050 162968
rect 85106 162966 85130 162968
rect 84890 162946 85186 162966
rect 85262 162804 85290 164272
rect 86890 163566 87186 163586
rect 86946 163564 86970 163566
rect 87026 163564 87050 163566
rect 87106 163564 87130 163566
rect 86968 163512 86970 163564
rect 87032 163512 87044 163564
rect 87106 163512 87108 163564
rect 86946 163510 86970 163512
rect 87026 163510 87050 163512
rect 87106 163510 87130 163512
rect 86890 163490 87186 163510
rect 85170 162776 85290 162804
rect 85170 162124 85198 162776
rect 86890 162478 87186 162498
rect 86946 162476 86970 162478
rect 87026 162476 87050 162478
rect 87106 162476 87130 162478
rect 86968 162424 86970 162476
rect 87032 162424 87044 162476
rect 87106 162424 87108 162476
rect 86946 162422 86970 162424
rect 87026 162422 87050 162424
rect 87106 162422 87130 162424
rect 86890 162402 87186 162422
rect 85170 162096 85290 162124
rect 84890 161934 85186 161954
rect 84946 161932 84970 161934
rect 85026 161932 85050 161934
rect 85106 161932 85130 161934
rect 84968 161880 84970 161932
rect 85032 161880 85044 161932
rect 85106 161880 85108 161932
rect 84946 161878 84970 161880
rect 85026 161878 85050 161880
rect 85106 161878 85130 161880
rect 84890 161858 85186 161878
rect 85262 161716 85290 162096
rect 85170 161688 85290 161716
rect 85170 161603 85198 161688
rect 85156 161594 85212 161603
rect 85156 161529 85212 161538
rect 86890 161390 87186 161410
rect 86946 161388 86970 161390
rect 87026 161388 87050 161390
rect 87106 161388 87130 161390
rect 86968 161336 86970 161388
rect 87032 161336 87044 161388
rect 87106 161336 87108 161388
rect 86946 161334 86970 161336
rect 87026 161334 87050 161336
rect 87106 161334 87130 161336
rect 86890 161314 87186 161334
rect 84890 160846 85186 160866
rect 84946 160844 84970 160846
rect 85026 160844 85050 160846
rect 85106 160844 85130 160846
rect 84968 160792 84970 160844
rect 85032 160792 85044 160844
rect 85106 160792 85108 160844
rect 84946 160790 84970 160792
rect 85026 160790 85050 160792
rect 85106 160790 85130 160792
rect 84890 160770 85186 160790
rect 85342 160674 85394 160680
rect 85342 160616 85394 160622
rect 84890 159758 85186 159778
rect 84946 159756 84970 159758
rect 85026 159756 85050 159758
rect 85106 159756 85130 159758
rect 84968 159704 84970 159756
rect 85032 159704 85044 159756
rect 85106 159704 85108 159756
rect 84946 159702 84970 159704
rect 85026 159702 85050 159704
rect 85106 159702 85130 159704
rect 84890 159682 85186 159702
rect 84890 158670 85186 158690
rect 84946 158668 84970 158670
rect 85026 158668 85050 158670
rect 85106 158668 85130 158670
rect 84968 158616 84970 158668
rect 85032 158616 85044 158668
rect 85106 158616 85108 158668
rect 84946 158614 84970 158616
rect 85026 158614 85050 158616
rect 85106 158614 85130 158616
rect 84890 158594 85186 158614
rect 84890 157582 85186 157602
rect 84946 157580 84970 157582
rect 85026 157580 85050 157582
rect 85106 157580 85130 157582
rect 84968 157528 84970 157580
rect 85032 157528 85044 157580
rect 85106 157528 85108 157580
rect 84946 157526 84970 157528
rect 85026 157526 85050 157528
rect 85106 157526 85130 157528
rect 84890 157506 85186 157526
rect 85066 156934 85118 156940
rect 85066 156876 85118 156882
rect 85078 156707 85106 156876
rect 85064 156698 85120 156707
rect 85064 156633 85120 156642
rect 84890 156494 85186 156514
rect 84946 156492 84970 156494
rect 85026 156492 85050 156494
rect 85106 156492 85130 156494
rect 84968 156440 84970 156492
rect 85032 156440 85044 156492
rect 85106 156440 85108 156492
rect 84946 156438 84970 156440
rect 85026 156438 85050 156440
rect 85106 156438 85130 156440
rect 84890 156418 85186 156438
rect 84890 155406 85186 155426
rect 84946 155404 84970 155406
rect 85026 155404 85050 155406
rect 85106 155404 85130 155406
rect 84968 155352 84970 155404
rect 85032 155352 85044 155404
rect 85106 155352 85108 155404
rect 84946 155350 84970 155352
rect 85026 155350 85050 155352
rect 85106 155350 85130 155352
rect 84890 155330 85186 155350
rect 84890 154318 85186 154338
rect 84946 154316 84970 154318
rect 85026 154316 85050 154318
rect 85106 154316 85130 154318
rect 84968 154264 84970 154316
rect 85032 154264 85044 154316
rect 85106 154264 85108 154316
rect 84946 154262 84970 154264
rect 85026 154262 85050 154264
rect 85106 154262 85130 154264
rect 84890 154242 85186 154262
rect 85354 154259 85382 160616
rect 86890 160302 87186 160322
rect 86946 160300 86970 160302
rect 87026 160300 87050 160302
rect 87106 160300 87130 160302
rect 86968 160248 86970 160300
rect 87032 160248 87044 160300
rect 87106 160248 87108 160300
rect 86946 160246 86970 160248
rect 87026 160246 87050 160248
rect 87106 160246 87130 160248
rect 86890 160226 87186 160246
rect 86890 159214 87186 159234
rect 86946 159212 86970 159214
rect 87026 159212 87050 159214
rect 87106 159212 87130 159214
rect 86968 159160 86970 159212
rect 87032 159160 87044 159212
rect 87106 159160 87108 159212
rect 86946 159158 86970 159160
rect 87026 159158 87050 159160
rect 87106 159158 87130 159160
rect 86890 159138 87186 159158
rect 86890 158126 87186 158146
rect 86946 158124 86970 158126
rect 87026 158124 87050 158126
rect 87106 158124 87130 158126
rect 86968 158072 86970 158124
rect 87032 158072 87044 158124
rect 87106 158072 87108 158124
rect 86946 158070 86970 158072
rect 87026 158070 87050 158072
rect 87106 158070 87130 158072
rect 86890 158050 87186 158070
rect 86890 157038 87186 157058
rect 86946 157036 86970 157038
rect 87026 157036 87050 157038
rect 87106 157036 87130 157038
rect 86968 156984 86970 157036
rect 87032 156984 87044 157036
rect 87106 156984 87108 157036
rect 86946 156982 86970 156984
rect 87026 156982 87050 156984
rect 87106 156982 87130 156984
rect 86890 156962 87186 156982
rect 86890 155950 87186 155970
rect 86946 155948 86970 155950
rect 87026 155948 87050 155950
rect 87106 155948 87130 155950
rect 86968 155896 86970 155948
rect 87032 155896 87044 155948
rect 87106 155896 87108 155948
rect 86946 155894 86970 155896
rect 87026 155894 87050 155896
rect 87106 155894 87130 155896
rect 86890 155874 87186 155894
rect 86890 154862 87186 154882
rect 86946 154860 86970 154862
rect 87026 154860 87050 154862
rect 87106 154860 87130 154862
rect 86968 154808 86970 154860
rect 87032 154808 87044 154860
rect 87106 154808 87108 154860
rect 86946 154806 86970 154808
rect 87026 154806 87050 154808
rect 87106 154806 87130 154808
rect 86890 154786 87186 154806
rect 85340 154250 85396 154259
rect 85340 154185 85396 154194
rect 86890 153774 87186 153794
rect 86946 153772 86970 153774
rect 87026 153772 87050 153774
rect 87106 153772 87130 153774
rect 86968 153720 86970 153772
rect 87032 153720 87044 153772
rect 87106 153720 87108 153772
rect 86946 153718 86970 153720
rect 87026 153718 87050 153720
rect 87106 153718 87130 153720
rect 86890 153698 87186 153718
rect 84890 153230 85186 153250
rect 84946 153228 84970 153230
rect 85026 153228 85050 153230
rect 85106 153228 85130 153230
rect 84968 153176 84970 153228
rect 85032 153176 85044 153228
rect 85106 153176 85108 153228
rect 84946 153174 84970 153176
rect 85026 153174 85050 153176
rect 85106 153174 85130 153176
rect 84890 153154 85186 153174
rect 86890 152686 87186 152706
rect 86946 152684 86970 152686
rect 87026 152684 87050 152686
rect 87106 152684 87130 152686
rect 86968 152632 86970 152684
rect 87032 152632 87044 152684
rect 87106 152632 87108 152684
rect 86946 152630 86970 152632
rect 87026 152630 87050 152632
rect 87106 152630 87130 152632
rect 86890 152610 87186 152630
rect 84890 152142 85186 152162
rect 84946 152140 84970 152142
rect 85026 152140 85050 152142
rect 85106 152140 85130 152142
rect 84968 152088 84970 152140
rect 85032 152088 85044 152140
rect 85106 152088 85108 152140
rect 84946 152086 84970 152088
rect 85026 152086 85050 152088
rect 85106 152086 85130 152088
rect 84890 152066 85186 152086
rect 86890 151598 87186 151618
rect 86946 151596 86970 151598
rect 87026 151596 87050 151598
rect 87106 151596 87130 151598
rect 86968 151544 86970 151596
rect 87032 151544 87044 151596
rect 87106 151544 87108 151596
rect 86946 151542 86970 151544
rect 87026 151542 87050 151544
rect 87106 151542 87130 151544
rect 86890 151522 87186 151542
rect 84890 151054 85186 151074
rect 84946 151052 84970 151054
rect 85026 151052 85050 151054
rect 85106 151052 85130 151054
rect 84968 151000 84970 151052
rect 85032 151000 85044 151052
rect 85106 151000 85108 151052
rect 84946 150998 84970 151000
rect 85026 150998 85050 151000
rect 85106 150998 85130 151000
rect 84890 150978 85186 150998
rect 86890 150510 87186 150530
rect 86946 150508 86970 150510
rect 87026 150508 87050 150510
rect 87106 150508 87130 150510
rect 86968 150456 86970 150508
rect 87032 150456 87044 150508
rect 87106 150456 87108 150508
rect 86946 150454 86970 150456
rect 87026 150454 87050 150456
rect 87106 150454 87130 150456
rect 86890 150434 87186 150454
rect 84890 149966 85186 149986
rect 84946 149964 84970 149966
rect 85026 149964 85050 149966
rect 85106 149964 85130 149966
rect 84968 149912 84970 149964
rect 85032 149912 85044 149964
rect 85106 149912 85108 149964
rect 84946 149910 84970 149912
rect 85026 149910 85050 149912
rect 85106 149910 85130 149912
rect 84890 149890 85186 149910
rect 86890 149422 87186 149442
rect 86946 149420 86970 149422
rect 87026 149420 87050 149422
rect 87106 149420 87130 149422
rect 86968 149368 86970 149420
rect 87032 149368 87044 149420
rect 87106 149368 87108 149420
rect 86946 149366 86970 149368
rect 87026 149366 87050 149368
rect 87106 149366 87130 149368
rect 86890 149346 87186 149366
rect 84890 148878 85186 148898
rect 84946 148876 84970 148878
rect 85026 148876 85050 148878
rect 85106 148876 85130 148878
rect 84968 148824 84970 148876
rect 85032 148824 85044 148876
rect 85106 148824 85108 148876
rect 84946 148822 84970 148824
rect 85026 148822 85050 148824
rect 85106 148822 85130 148824
rect 84890 148802 85186 148822
rect 86890 148334 87186 148354
rect 86946 148332 86970 148334
rect 87026 148332 87050 148334
rect 87106 148332 87130 148334
rect 86968 148280 86970 148332
rect 87032 148280 87044 148332
rect 87106 148280 87108 148332
rect 86946 148278 86970 148280
rect 87026 148278 87050 148280
rect 87106 148278 87130 148280
rect 86890 148258 87186 148278
rect 84890 147790 85186 147810
rect 84946 147788 84970 147790
rect 85026 147788 85050 147790
rect 85106 147788 85130 147790
rect 84968 147736 84970 147788
rect 85032 147736 85044 147788
rect 85106 147736 85108 147788
rect 84946 147734 84970 147736
rect 85026 147734 85050 147736
rect 85106 147734 85130 147736
rect 84890 147714 85186 147734
rect 86890 147246 87186 147266
rect 86946 147244 86970 147246
rect 87026 147244 87050 147246
rect 87106 147244 87130 147246
rect 86968 147192 86970 147244
rect 87032 147192 87044 147244
rect 87106 147192 87108 147244
rect 86946 147190 86970 147192
rect 87026 147190 87050 147192
rect 87106 147190 87130 147192
rect 86890 147170 87186 147190
rect 84890 146702 85186 146722
rect 84946 146700 84970 146702
rect 85026 146700 85050 146702
rect 85106 146700 85130 146702
rect 84968 146648 84970 146700
rect 85032 146648 85044 146700
rect 85106 146648 85108 146700
rect 84946 146646 84970 146648
rect 85026 146646 85050 146648
rect 85106 146646 85130 146648
rect 84890 146626 85186 146646
rect 86890 146158 87186 146178
rect 86946 146156 86970 146158
rect 87026 146156 87050 146158
rect 87106 146156 87130 146158
rect 86968 146104 86970 146156
rect 87032 146104 87044 146156
rect 87106 146104 87108 146156
rect 86946 146102 86970 146104
rect 87026 146102 87050 146104
rect 87106 146102 87130 146104
rect 86890 146082 87186 146102
rect 84890 145614 85186 145634
rect 84946 145612 84970 145614
rect 85026 145612 85050 145614
rect 85106 145612 85130 145614
rect 84968 145560 84970 145612
rect 85032 145560 85044 145612
rect 85106 145560 85108 145612
rect 84946 145558 84970 145560
rect 85026 145558 85050 145560
rect 85106 145558 85130 145560
rect 84890 145538 85186 145558
rect 86890 145070 87186 145090
rect 86946 145068 86970 145070
rect 87026 145068 87050 145070
rect 87106 145068 87130 145070
rect 86968 145016 86970 145068
rect 87032 145016 87044 145068
rect 87106 145016 87108 145068
rect 86946 145014 86970 145016
rect 87026 145014 87050 145016
rect 87106 145014 87130 145016
rect 86890 144994 87186 145014
rect 84890 144526 85186 144546
rect 84946 144524 84970 144526
rect 85026 144524 85050 144526
rect 85106 144524 85130 144526
rect 84968 144472 84970 144524
rect 85032 144472 85044 144524
rect 85106 144472 85108 144524
rect 84946 144470 84970 144472
rect 85026 144470 85050 144472
rect 85106 144470 85130 144472
rect 84890 144450 85186 144470
rect 86890 143982 87186 144002
rect 86946 143980 86970 143982
rect 87026 143980 87050 143982
rect 87106 143980 87130 143982
rect 86968 143928 86970 143980
rect 87032 143928 87044 143980
rect 87106 143928 87108 143980
rect 86946 143926 86970 143928
rect 87026 143926 87050 143928
rect 87106 143926 87130 143928
rect 86890 143906 87186 143926
rect 84890 143438 85186 143458
rect 84946 143436 84970 143438
rect 85026 143436 85050 143438
rect 85106 143436 85130 143438
rect 84968 143384 84970 143436
rect 85032 143384 85044 143436
rect 85106 143384 85108 143436
rect 84946 143382 84970 143384
rect 85026 143382 85050 143384
rect 85106 143382 85130 143384
rect 84890 143362 85186 143382
rect 86890 142894 87186 142914
rect 86946 142892 86970 142894
rect 87026 142892 87050 142894
rect 87106 142892 87130 142894
rect 86968 142840 86970 142892
rect 87032 142840 87044 142892
rect 87106 142840 87108 142892
rect 86946 142838 86970 142840
rect 87026 142838 87050 142840
rect 87106 142838 87130 142840
rect 86890 142818 87186 142838
rect 84890 142350 85186 142370
rect 84946 142348 84970 142350
rect 85026 142348 85050 142350
rect 85106 142348 85130 142350
rect 84968 142296 84970 142348
rect 85032 142296 85044 142348
rect 85106 142296 85108 142348
rect 84946 142294 84970 142296
rect 85026 142294 85050 142296
rect 85106 142294 85130 142296
rect 84890 142274 85186 142294
rect 86890 141806 87186 141826
rect 86946 141804 86970 141806
rect 87026 141804 87050 141806
rect 87106 141804 87130 141806
rect 86968 141752 86970 141804
rect 87032 141752 87044 141804
rect 87106 141752 87108 141804
rect 86946 141750 86970 141752
rect 87026 141750 87050 141752
rect 87106 141750 87130 141752
rect 86890 141730 87186 141750
rect 84890 141262 85186 141282
rect 84946 141260 84970 141262
rect 85026 141260 85050 141262
rect 85106 141260 85130 141262
rect 84968 141208 84970 141260
rect 85032 141208 85044 141260
rect 85106 141208 85108 141260
rect 84946 141206 84970 141208
rect 85026 141206 85050 141208
rect 85106 141206 85130 141208
rect 84890 141186 85186 141206
rect 86890 140718 87186 140738
rect 86946 140716 86970 140718
rect 87026 140716 87050 140718
rect 87106 140716 87130 140718
rect 86968 140664 86970 140716
rect 87032 140664 87044 140716
rect 87106 140664 87108 140716
rect 86946 140662 86970 140664
rect 87026 140662 87050 140664
rect 87106 140662 87130 140664
rect 86890 140642 87186 140662
rect 84890 140174 85186 140194
rect 84946 140172 84970 140174
rect 85026 140172 85050 140174
rect 85106 140172 85130 140174
rect 84968 140120 84970 140172
rect 85032 140120 85044 140172
rect 85106 140120 85108 140172
rect 84946 140118 84970 140120
rect 85026 140118 85050 140120
rect 85106 140118 85130 140120
rect 84890 140098 85186 140118
rect 86890 139630 87186 139650
rect 86946 139628 86970 139630
rect 87026 139628 87050 139630
rect 87106 139628 87130 139630
rect 86968 139576 86970 139628
rect 87032 139576 87044 139628
rect 87106 139576 87108 139628
rect 86946 139574 86970 139576
rect 87026 139574 87050 139576
rect 87106 139574 87130 139576
rect 86890 139554 87186 139574
rect 84890 139086 85186 139106
rect 84946 139084 84970 139086
rect 85026 139084 85050 139086
rect 85106 139084 85130 139086
rect 84968 139032 84970 139084
rect 85032 139032 85044 139084
rect 85106 139032 85108 139084
rect 84946 139030 84970 139032
rect 85026 139030 85050 139032
rect 85106 139030 85130 139032
rect 84890 139010 85186 139030
rect 86890 138542 87186 138562
rect 86946 138540 86970 138542
rect 87026 138540 87050 138542
rect 87106 138540 87130 138542
rect 86968 138488 86970 138540
rect 87032 138488 87044 138540
rect 87106 138488 87108 138540
rect 86946 138486 86970 138488
rect 87026 138486 87050 138488
rect 87106 138486 87130 138488
rect 86890 138466 87186 138486
rect 84890 137998 85186 138018
rect 84946 137996 84970 137998
rect 85026 137996 85050 137998
rect 85106 137996 85130 137998
rect 84968 137944 84970 137996
rect 85032 137944 85044 137996
rect 85106 137944 85108 137996
rect 84946 137942 84970 137944
rect 85026 137942 85050 137944
rect 85106 137942 85130 137944
rect 84890 137922 85186 137942
rect 86890 137454 87186 137474
rect 86946 137452 86970 137454
rect 87026 137452 87050 137454
rect 87106 137452 87130 137454
rect 86968 137400 86970 137452
rect 87032 137400 87044 137452
rect 87106 137400 87108 137452
rect 86946 137398 86970 137400
rect 87026 137398 87050 137400
rect 87106 137398 87130 137400
rect 86890 137378 87186 137398
rect 85800 137250 85856 137259
rect 85800 137185 85856 137194
rect 84890 136910 85186 136930
rect 84946 136908 84970 136910
rect 85026 136908 85050 136910
rect 85106 136908 85130 136910
rect 84968 136856 84970 136908
rect 85032 136856 85044 136908
rect 85106 136856 85108 136908
rect 84946 136854 84970 136856
rect 85026 136854 85050 136856
rect 85106 136854 85130 136856
rect 84890 136834 85186 136854
rect 84890 135822 85186 135842
rect 84946 135820 84970 135822
rect 85026 135820 85050 135822
rect 85106 135820 85130 135822
rect 84968 135768 84970 135820
rect 85032 135768 85044 135820
rect 85106 135768 85108 135820
rect 84946 135766 84970 135768
rect 85026 135766 85050 135768
rect 85106 135766 85130 135768
rect 84890 135746 85186 135766
rect 84890 134734 85186 134754
rect 84946 134732 84970 134734
rect 85026 134732 85050 134734
rect 85106 134732 85130 134734
rect 84968 134680 84970 134732
rect 85032 134680 85044 134732
rect 85106 134680 85108 134732
rect 84946 134678 84970 134680
rect 85026 134678 85050 134680
rect 85106 134678 85130 134680
rect 84890 134658 85186 134678
rect 84890 133646 85186 133666
rect 84946 133644 84970 133646
rect 85026 133644 85050 133646
rect 85106 133644 85130 133646
rect 84968 133592 84970 133644
rect 85032 133592 85044 133644
rect 85106 133592 85108 133644
rect 84946 133590 84970 133592
rect 85026 133590 85050 133592
rect 85106 133590 85130 133592
rect 84890 133570 85186 133590
rect 84890 132558 85186 132578
rect 84946 132556 84970 132558
rect 85026 132556 85050 132558
rect 85106 132556 85130 132558
rect 84968 132504 84970 132556
rect 85032 132504 85044 132556
rect 85106 132504 85108 132556
rect 84946 132502 84970 132504
rect 85026 132502 85050 132504
rect 85106 132502 85130 132504
rect 84890 132482 85186 132502
rect 84890 131470 85186 131490
rect 84946 131468 84970 131470
rect 85026 131468 85050 131470
rect 85106 131468 85130 131470
rect 84968 131416 84970 131468
rect 85032 131416 85044 131468
rect 85106 131416 85108 131468
rect 84946 131414 84970 131416
rect 85026 131414 85050 131416
rect 85106 131414 85130 131416
rect 84890 131394 85186 131414
rect 84890 130382 85186 130402
rect 84946 130380 84970 130382
rect 85026 130380 85050 130382
rect 85106 130380 85130 130382
rect 84968 130328 84970 130380
rect 85032 130328 85044 130380
rect 85106 130328 85108 130380
rect 84946 130326 84970 130328
rect 85026 130326 85050 130328
rect 85106 130326 85130 130328
rect 84890 130306 85186 130326
rect 84890 129294 85186 129314
rect 84946 129292 84970 129294
rect 85026 129292 85050 129294
rect 85106 129292 85130 129294
rect 84968 129240 84970 129292
rect 85032 129240 85044 129292
rect 85106 129240 85108 129292
rect 84946 129238 84970 129240
rect 85026 129238 85050 129240
rect 85106 129238 85130 129240
rect 84890 129218 85186 129238
rect 84890 128206 85186 128226
rect 84946 128204 84970 128206
rect 85026 128204 85050 128206
rect 85106 128204 85130 128206
rect 84968 128152 84970 128204
rect 85032 128152 85044 128204
rect 85106 128152 85108 128204
rect 84946 128150 84970 128152
rect 85026 128150 85050 128152
rect 85106 128150 85130 128152
rect 84890 128130 85186 128150
rect 84890 127118 85186 127138
rect 84946 127116 84970 127118
rect 85026 127116 85050 127118
rect 85106 127116 85130 127118
rect 84968 127064 84970 127116
rect 85032 127064 85044 127116
rect 85106 127064 85108 127116
rect 84946 127062 84970 127064
rect 85026 127062 85050 127064
rect 85106 127062 85130 127064
rect 84890 127042 85186 127062
rect 84890 126030 85186 126050
rect 84946 126028 84970 126030
rect 85026 126028 85050 126030
rect 85106 126028 85130 126030
rect 84968 125976 84970 126028
rect 85032 125976 85044 126028
rect 85106 125976 85108 126028
rect 84946 125974 84970 125976
rect 85026 125974 85050 125976
rect 85106 125974 85130 125976
rect 84890 125954 85186 125974
rect 84890 124942 85186 124962
rect 84946 124940 84970 124942
rect 85026 124940 85050 124942
rect 85106 124940 85130 124942
rect 84968 124888 84970 124940
rect 85032 124888 85044 124940
rect 85106 124888 85108 124940
rect 84946 124886 84970 124888
rect 85026 124886 85050 124888
rect 85106 124886 85130 124888
rect 84890 124866 85186 124886
rect 84890 123854 85186 123874
rect 84946 123852 84970 123854
rect 85026 123852 85050 123854
rect 85106 123852 85130 123854
rect 84968 123800 84970 123852
rect 85032 123800 85044 123852
rect 85106 123800 85108 123852
rect 84946 123798 84970 123800
rect 85026 123798 85050 123800
rect 85106 123798 85130 123800
rect 84890 123778 85186 123798
rect 84890 122766 85186 122786
rect 84946 122764 84970 122766
rect 85026 122764 85050 122766
rect 85106 122764 85130 122766
rect 84968 122712 84970 122764
rect 85032 122712 85044 122764
rect 85106 122712 85108 122764
rect 84946 122710 84970 122712
rect 85026 122710 85050 122712
rect 85106 122710 85130 122712
rect 84890 122690 85186 122710
rect 84890 121678 85186 121698
rect 84946 121676 84970 121678
rect 85026 121676 85050 121678
rect 85106 121676 85130 121678
rect 84968 121624 84970 121676
rect 85032 121624 85044 121676
rect 85106 121624 85108 121676
rect 84946 121622 84970 121624
rect 85026 121622 85050 121624
rect 85106 121622 85130 121624
rect 84890 121602 85186 121622
rect 84890 120590 85186 120610
rect 84946 120588 84970 120590
rect 85026 120588 85050 120590
rect 85106 120588 85130 120590
rect 84968 120536 84970 120588
rect 85032 120536 85044 120588
rect 85106 120536 85108 120588
rect 84946 120534 84970 120536
rect 85026 120534 85050 120536
rect 85106 120534 85130 120536
rect 84890 120514 85186 120534
rect 84890 119502 85186 119522
rect 84946 119500 84970 119502
rect 85026 119500 85050 119502
rect 85106 119500 85130 119502
rect 84968 119448 84970 119500
rect 85032 119448 85044 119500
rect 85106 119448 85108 119500
rect 84946 119446 84970 119448
rect 85026 119446 85050 119448
rect 85106 119446 85130 119448
rect 84890 119426 85186 119446
rect 85340 119434 85396 119443
rect 85340 119369 85342 119378
rect 85394 119369 85396 119378
rect 85342 119340 85394 119346
rect 84890 118414 85186 118434
rect 84946 118412 84970 118414
rect 85026 118412 85050 118414
rect 85106 118412 85130 118414
rect 84968 118360 84970 118412
rect 85032 118360 85044 118412
rect 85106 118360 85108 118412
rect 84946 118358 84970 118360
rect 85026 118358 85050 118360
rect 85106 118358 85130 118360
rect 84890 118338 85186 118358
rect 84890 117326 85186 117346
rect 84946 117324 84970 117326
rect 85026 117324 85050 117326
rect 85106 117324 85130 117326
rect 84968 117272 84970 117324
rect 85032 117272 85044 117324
rect 85106 117272 85108 117324
rect 84946 117270 84970 117272
rect 85026 117270 85050 117272
rect 85106 117270 85130 117272
rect 84890 117250 85186 117270
rect 84890 116238 85186 116258
rect 84946 116236 84970 116238
rect 85026 116236 85050 116238
rect 85106 116236 85130 116238
rect 84968 116184 84970 116236
rect 85032 116184 85044 116236
rect 85106 116184 85108 116236
rect 84946 116182 84970 116184
rect 85026 116182 85050 116184
rect 85106 116182 85130 116184
rect 84890 116162 85186 116182
rect 84890 115150 85186 115170
rect 84946 115148 84970 115150
rect 85026 115148 85050 115150
rect 85106 115148 85130 115150
rect 84968 115096 84970 115148
rect 85032 115096 85044 115148
rect 85106 115096 85108 115148
rect 84946 115094 84970 115096
rect 85026 115094 85050 115096
rect 85106 115094 85130 115096
rect 84890 115074 85186 115094
rect 84890 114062 85186 114082
rect 84946 114060 84970 114062
rect 85026 114060 85050 114062
rect 85106 114060 85130 114062
rect 84968 114008 84970 114060
rect 85032 114008 85044 114060
rect 85106 114008 85108 114060
rect 84946 114006 84970 114008
rect 85026 114006 85050 114008
rect 85106 114006 85130 114008
rect 84890 113986 85186 114006
rect 84890 112974 85186 112994
rect 84946 112972 84970 112974
rect 85026 112972 85050 112974
rect 85106 112972 85130 112974
rect 84968 112920 84970 112972
rect 85032 112920 85044 112972
rect 85106 112920 85108 112972
rect 84946 112918 84970 112920
rect 85026 112918 85050 112920
rect 85106 112918 85130 112920
rect 84890 112898 85186 112918
rect 84880 112226 84936 112235
rect 84880 112161 84936 112170
rect 84894 112060 84922 112161
rect 84882 112054 84934 112060
rect 84882 111996 84934 112002
rect 84890 111886 85186 111906
rect 84946 111884 84970 111886
rect 85026 111884 85050 111886
rect 85106 111884 85130 111886
rect 84968 111832 84970 111884
rect 85032 111832 85044 111884
rect 85106 111832 85108 111884
rect 84946 111830 84970 111832
rect 85026 111830 85050 111832
rect 85106 111830 85130 111832
rect 84890 111810 85186 111830
rect 84890 110798 85186 110818
rect 84946 110796 84970 110798
rect 85026 110796 85050 110798
rect 85106 110796 85130 110798
rect 84968 110744 84970 110796
rect 85032 110744 85044 110796
rect 85106 110744 85108 110796
rect 84946 110742 84970 110744
rect 85026 110742 85050 110744
rect 85106 110742 85130 110744
rect 84890 110722 85186 110742
rect 84890 109710 85186 109730
rect 84946 109708 84970 109710
rect 85026 109708 85050 109710
rect 85106 109708 85130 109710
rect 84968 109656 84970 109708
rect 85032 109656 85044 109708
rect 85106 109656 85108 109708
rect 84946 109654 84970 109656
rect 85026 109654 85050 109656
rect 85106 109654 85130 109656
rect 84890 109634 85186 109654
rect 84890 108622 85186 108642
rect 84946 108620 84970 108622
rect 85026 108620 85050 108622
rect 85106 108620 85130 108622
rect 84968 108568 84970 108620
rect 85032 108568 85044 108620
rect 85106 108568 85108 108620
rect 84946 108566 84970 108568
rect 85026 108566 85050 108568
rect 85106 108566 85130 108568
rect 84890 108546 85186 108566
rect 84890 107534 85186 107554
rect 84946 107532 84970 107534
rect 85026 107532 85050 107534
rect 85106 107532 85130 107534
rect 84968 107480 84970 107532
rect 85032 107480 85044 107532
rect 85106 107480 85108 107532
rect 84946 107478 84970 107480
rect 85026 107478 85050 107480
rect 85106 107478 85130 107480
rect 84890 107458 85186 107478
rect 84890 106446 85186 106466
rect 84946 106444 84970 106446
rect 85026 106444 85050 106446
rect 85106 106444 85130 106446
rect 84968 106392 84970 106444
rect 85032 106392 85044 106444
rect 85106 106392 85108 106444
rect 84946 106390 84970 106392
rect 85026 106390 85050 106392
rect 85106 106390 85130 106392
rect 84890 106370 85186 106390
rect 84890 105358 85186 105378
rect 84946 105356 84970 105358
rect 85026 105356 85050 105358
rect 85106 105356 85130 105358
rect 84968 105304 84970 105356
rect 85032 105304 85044 105356
rect 85106 105304 85108 105356
rect 84946 105302 84970 105304
rect 85026 105302 85050 105304
rect 85106 105302 85130 105304
rect 84890 105282 85186 105302
rect 84890 104270 85186 104290
rect 84946 104268 84970 104270
rect 85026 104268 85050 104270
rect 85106 104268 85130 104270
rect 84968 104216 84970 104268
rect 85032 104216 85044 104268
rect 85106 104216 85108 104268
rect 84946 104214 84970 104216
rect 85026 104214 85050 104216
rect 85106 104214 85130 104216
rect 84890 104194 85186 104214
rect 84790 103486 84842 103492
rect 84790 103428 84842 103434
rect 85250 103486 85302 103492
rect 85250 103428 85302 103434
rect 84890 103182 85186 103202
rect 84946 103180 84970 103182
rect 85026 103180 85050 103182
rect 85106 103180 85130 103182
rect 84968 103128 84970 103180
rect 85032 103128 85044 103180
rect 85106 103128 85108 103180
rect 84946 103126 84970 103128
rect 85026 103126 85050 103128
rect 85106 103126 85130 103128
rect 84890 103106 85186 103126
rect 84890 102094 85186 102114
rect 84946 102092 84970 102094
rect 85026 102092 85050 102094
rect 85106 102092 85130 102094
rect 84968 102040 84970 102092
rect 85032 102040 85044 102092
rect 85106 102040 85108 102092
rect 84946 102038 84970 102040
rect 85026 102038 85050 102040
rect 85106 102038 85130 102040
rect 84890 102018 85186 102038
rect 84890 101006 85186 101026
rect 84946 101004 84970 101006
rect 85026 101004 85050 101006
rect 85106 101004 85130 101006
rect 84968 100952 84970 101004
rect 85032 100952 85044 101004
rect 85106 100952 85108 101004
rect 84946 100950 84970 100952
rect 85026 100950 85050 100952
rect 85106 100950 85130 100952
rect 84890 100930 85186 100950
rect 84698 100358 84750 100364
rect 84698 100300 84750 100306
rect 84618 100216 84830 100244
rect 84696 100122 84752 100131
rect 84696 100057 84752 100066
rect 84604 99034 84660 99043
rect 84604 98969 84660 98978
rect 84514 97638 84566 97644
rect 84514 97580 84566 97586
rect 84514 96890 84566 96896
rect 84514 96832 84566 96838
rect 84422 96414 84474 96420
rect 84422 96356 84474 96362
rect 84526 95507 84554 96832
rect 84512 95498 84568 95507
rect 84512 95433 84568 95442
rect 84618 94924 84646 98969
rect 84710 95468 84738 100057
rect 84802 96896 84830 100216
rect 84890 99918 85186 99938
rect 84946 99916 84970 99918
rect 85026 99916 85050 99918
rect 85106 99916 85130 99918
rect 84968 99864 84970 99916
rect 85032 99864 85044 99916
rect 85106 99864 85108 99916
rect 84946 99862 84970 99864
rect 85026 99862 85050 99864
rect 85106 99862 85130 99864
rect 84890 99842 85186 99862
rect 85262 99004 85290 103428
rect 85708 101346 85764 101355
rect 85708 101281 85764 101290
rect 85250 98998 85302 99004
rect 85250 98940 85302 98946
rect 84890 98830 85186 98850
rect 84946 98828 84970 98830
rect 85026 98828 85050 98830
rect 85106 98828 85130 98830
rect 84968 98776 84970 98828
rect 85032 98776 85044 98828
rect 85106 98776 85108 98828
rect 84946 98774 84970 98776
rect 85026 98774 85050 98776
rect 85106 98774 85130 98776
rect 84890 98754 85186 98774
rect 85158 98046 85210 98052
rect 85158 97988 85210 97994
rect 85170 97932 85198 97988
rect 85170 97904 85290 97932
rect 84890 97742 85186 97762
rect 84946 97740 84970 97742
rect 85026 97740 85050 97742
rect 85106 97740 85130 97742
rect 84968 97688 84970 97740
rect 85032 97688 85044 97740
rect 85106 97688 85108 97740
rect 84946 97686 84970 97688
rect 85026 97686 85050 97688
rect 85106 97686 85130 97688
rect 84890 97666 85186 97686
rect 85262 97524 85290 97904
rect 85170 97496 85290 97524
rect 84790 96890 84842 96896
rect 84790 96832 84842 96838
rect 85170 96844 85198 97496
rect 85340 96858 85396 96867
rect 85170 96816 85290 96844
rect 84890 96654 85186 96674
rect 84946 96652 84970 96654
rect 85026 96652 85050 96654
rect 85106 96652 85130 96654
rect 84968 96600 84970 96652
rect 85032 96600 85044 96652
rect 85106 96600 85108 96652
rect 84946 96598 84970 96600
rect 85026 96598 85050 96600
rect 85106 96598 85130 96600
rect 84890 96578 85186 96598
rect 85262 96436 85290 96816
rect 85340 96793 85396 96802
rect 85354 96760 85382 96793
rect 85342 96754 85394 96760
rect 85342 96696 85394 96702
rect 85354 96488 85382 96696
rect 85432 96586 85488 96595
rect 85432 96521 85488 96530
rect 85170 96408 85290 96436
rect 85342 96482 85394 96488
rect 85342 96424 85394 96430
rect 85170 96352 85198 96408
rect 85158 96346 85210 96352
rect 85158 96288 85210 96294
rect 85446 96216 85474 96521
rect 85434 96210 85486 96216
rect 85434 96152 85486 96158
rect 84890 95566 85186 95586
rect 84946 95564 84970 95566
rect 85026 95564 85050 95566
rect 85106 95564 85130 95566
rect 84968 95512 84970 95564
rect 85032 95512 85044 95564
rect 85106 95512 85108 95564
rect 84946 95510 84970 95512
rect 85026 95510 85050 95512
rect 85106 95510 85130 95512
rect 84890 95490 85186 95510
rect 84698 95462 84750 95468
rect 84698 95404 84750 95410
rect 85156 95362 85212 95371
rect 85156 95297 85212 95306
rect 85170 95264 85198 95297
rect 85158 95258 85210 95264
rect 85158 95200 85210 95206
rect 84606 94918 84658 94924
rect 84606 94860 84658 94866
rect 85722 94788 85750 101281
rect 85814 97372 85842 137185
rect 86890 136366 87186 136386
rect 86946 136364 86970 136366
rect 87026 136364 87050 136366
rect 87106 136364 87130 136366
rect 86968 136312 86970 136364
rect 87032 136312 87044 136364
rect 87106 136312 87108 136364
rect 86946 136310 86970 136312
rect 87026 136310 87050 136312
rect 87106 136310 87130 136312
rect 86890 136290 87186 136310
rect 86890 135278 87186 135298
rect 86946 135276 86970 135278
rect 87026 135276 87050 135278
rect 87106 135276 87130 135278
rect 86968 135224 86970 135276
rect 87032 135224 87044 135276
rect 87106 135224 87108 135276
rect 86946 135222 86970 135224
rect 87026 135222 87050 135224
rect 87106 135222 87130 135224
rect 86890 135202 87186 135222
rect 86890 134190 87186 134210
rect 86946 134188 86970 134190
rect 87026 134188 87050 134190
rect 87106 134188 87130 134190
rect 86968 134136 86970 134188
rect 87032 134136 87044 134188
rect 87106 134136 87108 134188
rect 86946 134134 86970 134136
rect 87026 134134 87050 134136
rect 87106 134134 87130 134136
rect 86890 134114 87186 134134
rect 86890 133102 87186 133122
rect 86946 133100 86970 133102
rect 87026 133100 87050 133102
rect 87106 133100 87130 133102
rect 86968 133048 86970 133100
rect 87032 133048 87044 133100
rect 87106 133048 87108 133100
rect 86946 133046 86970 133048
rect 87026 133046 87050 133048
rect 87106 133046 87130 133048
rect 86890 133026 87186 133046
rect 86890 132014 87186 132034
rect 86946 132012 86970 132014
rect 87026 132012 87050 132014
rect 87106 132012 87130 132014
rect 86968 131960 86970 132012
rect 87032 131960 87044 132012
rect 87106 131960 87108 132012
rect 86946 131958 86970 131960
rect 87026 131958 87050 131960
rect 87106 131958 87130 131960
rect 86890 131938 87186 131958
rect 86890 130926 87186 130946
rect 86946 130924 86970 130926
rect 87026 130924 87050 130926
rect 87106 130924 87130 130926
rect 86968 130872 86970 130924
rect 87032 130872 87044 130924
rect 87106 130872 87108 130924
rect 86946 130870 86970 130872
rect 87026 130870 87050 130872
rect 87106 130870 87130 130872
rect 86890 130850 87186 130870
rect 86890 129838 87186 129858
rect 86946 129836 86970 129838
rect 87026 129836 87050 129838
rect 87106 129836 87130 129838
rect 86968 129784 86970 129836
rect 87032 129784 87044 129836
rect 87106 129784 87108 129836
rect 86946 129782 86970 129784
rect 87026 129782 87050 129784
rect 87106 129782 87130 129784
rect 86890 129762 87186 129782
rect 85892 129090 85948 129099
rect 85892 129025 85948 129034
rect 85802 97366 85854 97372
rect 85802 97308 85854 97314
rect 85906 94827 85934 129025
rect 86890 128750 87186 128770
rect 86946 128748 86970 128750
rect 87026 128748 87050 128750
rect 87106 128748 87130 128750
rect 86968 128696 86970 128748
rect 87032 128696 87044 128748
rect 87106 128696 87108 128748
rect 86946 128694 86970 128696
rect 87026 128694 87050 128696
rect 87106 128694 87130 128696
rect 86890 128674 87186 128694
rect 86890 127662 87186 127682
rect 86946 127660 86970 127662
rect 87026 127660 87050 127662
rect 87106 127660 87130 127662
rect 86968 127608 86970 127660
rect 87032 127608 87044 127660
rect 87106 127608 87108 127660
rect 86946 127606 86970 127608
rect 87026 127606 87050 127608
rect 87106 127606 87130 127608
rect 86890 127586 87186 127606
rect 86890 126574 87186 126594
rect 86946 126572 86970 126574
rect 87026 126572 87050 126574
rect 87106 126572 87130 126574
rect 86968 126520 86970 126572
rect 87032 126520 87044 126572
rect 87106 126520 87108 126572
rect 86946 126518 86970 126520
rect 87026 126518 87050 126520
rect 87106 126518 87130 126520
rect 86890 126498 87186 126518
rect 85984 126370 86040 126379
rect 85984 126305 86040 126314
rect 85998 96284 86026 126305
rect 86890 125486 87186 125506
rect 86946 125484 86970 125486
rect 87026 125484 87050 125486
rect 87106 125484 87130 125486
rect 86968 125432 86970 125484
rect 87032 125432 87044 125484
rect 87106 125432 87108 125484
rect 86946 125430 86970 125432
rect 87026 125430 87050 125432
rect 87106 125430 87130 125432
rect 86890 125410 87186 125430
rect 86890 124398 87186 124418
rect 86946 124396 86970 124398
rect 87026 124396 87050 124398
rect 87106 124396 87130 124398
rect 86968 124344 86970 124396
rect 87032 124344 87044 124396
rect 87106 124344 87108 124396
rect 86946 124342 86970 124344
rect 87026 124342 87050 124344
rect 87106 124342 87130 124344
rect 86890 124322 87186 124342
rect 86890 123310 87186 123330
rect 86946 123308 86970 123310
rect 87026 123308 87050 123310
rect 87106 123308 87130 123310
rect 86968 123256 86970 123308
rect 87032 123256 87044 123308
rect 87106 123256 87108 123308
rect 86946 123254 86970 123256
rect 87026 123254 87050 123256
rect 87106 123254 87130 123256
rect 86890 123234 87186 123254
rect 86890 122222 87186 122242
rect 86946 122220 86970 122222
rect 87026 122220 87050 122222
rect 87106 122220 87130 122222
rect 86968 122168 86970 122220
rect 87032 122168 87044 122220
rect 87106 122168 87108 122220
rect 86946 122166 86970 122168
rect 87026 122166 87050 122168
rect 87106 122166 87130 122168
rect 86890 122146 87186 122166
rect 86890 121134 87186 121154
rect 86946 121132 86970 121134
rect 87026 121132 87050 121134
rect 87106 121132 87130 121134
rect 86968 121080 86970 121132
rect 87032 121080 87044 121132
rect 87106 121080 87108 121132
rect 86946 121078 86970 121080
rect 87026 121078 87050 121080
rect 87106 121078 87130 121080
rect 86890 121058 87186 121078
rect 86890 120046 87186 120066
rect 86946 120044 86970 120046
rect 87026 120044 87050 120046
rect 87106 120044 87130 120046
rect 86968 119992 86970 120044
rect 87032 119992 87044 120044
rect 87106 119992 87108 120044
rect 86946 119990 86970 119992
rect 87026 119990 87050 119992
rect 87106 119990 87130 119992
rect 86890 119970 87186 119990
rect 86890 118958 87186 118978
rect 86946 118956 86970 118958
rect 87026 118956 87050 118958
rect 87106 118956 87130 118958
rect 86968 118904 86970 118956
rect 87032 118904 87044 118956
rect 87106 118904 87108 118956
rect 86946 118902 86970 118904
rect 87026 118902 87050 118904
rect 87106 118902 87130 118904
rect 86890 118882 87186 118902
rect 86890 117870 87186 117890
rect 86946 117868 86970 117870
rect 87026 117868 87050 117870
rect 87106 117868 87130 117870
rect 86968 117816 86970 117868
rect 87032 117816 87044 117868
rect 87106 117816 87108 117868
rect 86946 117814 86970 117816
rect 87026 117814 87050 117816
rect 87106 117814 87130 117816
rect 86890 117794 87186 117814
rect 86890 116782 87186 116802
rect 86946 116780 86970 116782
rect 87026 116780 87050 116782
rect 87106 116780 87130 116782
rect 86968 116728 86970 116780
rect 87032 116728 87044 116780
rect 87106 116728 87108 116780
rect 86946 116726 86970 116728
rect 87026 116726 87050 116728
rect 87106 116726 87130 116728
rect 86890 116706 87186 116726
rect 86890 115694 87186 115714
rect 86946 115692 86970 115694
rect 87026 115692 87050 115694
rect 87106 115692 87130 115694
rect 86968 115640 86970 115692
rect 87032 115640 87044 115692
rect 87106 115640 87108 115692
rect 86946 115638 86970 115640
rect 87026 115638 87050 115640
rect 87106 115638 87130 115640
rect 86890 115618 87186 115638
rect 86890 114606 87186 114626
rect 86946 114604 86970 114606
rect 87026 114604 87050 114606
rect 87106 114604 87130 114606
rect 86968 114552 86970 114604
rect 87032 114552 87044 114604
rect 87106 114552 87108 114604
rect 86946 114550 86970 114552
rect 87026 114550 87050 114552
rect 87106 114550 87130 114552
rect 86890 114530 87186 114550
rect 86890 113518 87186 113538
rect 86946 113516 86970 113518
rect 87026 113516 87050 113518
rect 87106 113516 87130 113518
rect 86968 113464 86970 113516
rect 87032 113464 87044 113516
rect 87106 113464 87108 113516
rect 86946 113462 86970 113464
rect 87026 113462 87050 113464
rect 87106 113462 87130 113464
rect 86890 113442 87186 113462
rect 86890 112430 87186 112450
rect 86946 112428 86970 112430
rect 87026 112428 87050 112430
rect 87106 112428 87130 112430
rect 86968 112376 86970 112428
rect 87032 112376 87044 112428
rect 87106 112376 87108 112428
rect 86946 112374 86970 112376
rect 87026 112374 87050 112376
rect 87106 112374 87130 112376
rect 86890 112354 87186 112374
rect 86890 111342 87186 111362
rect 86946 111340 86970 111342
rect 87026 111340 87050 111342
rect 87106 111340 87130 111342
rect 86968 111288 86970 111340
rect 87032 111288 87044 111340
rect 87106 111288 87108 111340
rect 86946 111286 86970 111288
rect 87026 111286 87050 111288
rect 87106 111286 87130 111288
rect 86890 111266 87186 111286
rect 86076 111002 86132 111011
rect 86076 110937 86132 110946
rect 86090 97440 86118 110937
rect 86890 110254 87186 110274
rect 86946 110252 86970 110254
rect 87026 110252 87050 110254
rect 87106 110252 87130 110254
rect 86968 110200 86970 110252
rect 87032 110200 87044 110252
rect 87106 110200 87108 110252
rect 86946 110198 86970 110200
rect 87026 110198 87050 110200
rect 87106 110198 87130 110200
rect 86890 110178 87186 110198
rect 86890 109166 87186 109186
rect 86946 109164 86970 109166
rect 87026 109164 87050 109166
rect 87106 109164 87130 109166
rect 86968 109112 86970 109164
rect 87032 109112 87044 109164
rect 87106 109112 87108 109164
rect 86946 109110 86970 109112
rect 87026 109110 87050 109112
rect 87106 109110 87130 109112
rect 86890 109090 87186 109110
rect 86890 108078 87186 108098
rect 86946 108076 86970 108078
rect 87026 108076 87050 108078
rect 87106 108076 87130 108078
rect 86968 108024 86970 108076
rect 87032 108024 87044 108076
rect 87106 108024 87108 108076
rect 86946 108022 86970 108024
rect 87026 108022 87050 108024
rect 87106 108022 87130 108024
rect 86890 108002 87186 108022
rect 86890 106990 87186 107010
rect 86946 106988 86970 106990
rect 87026 106988 87050 106990
rect 87106 106988 87130 106990
rect 86968 106936 86970 106988
rect 87032 106936 87044 106988
rect 87106 106936 87108 106988
rect 86946 106934 86970 106936
rect 87026 106934 87050 106936
rect 87106 106934 87130 106936
rect 86890 106914 87186 106934
rect 86890 105902 87186 105922
rect 86946 105900 86970 105902
rect 87026 105900 87050 105902
rect 87106 105900 87130 105902
rect 86968 105848 86970 105900
rect 87032 105848 87044 105900
rect 87106 105848 87108 105900
rect 86946 105846 86970 105848
rect 87026 105846 87050 105848
rect 87106 105846 87130 105848
rect 86890 105826 87186 105846
rect 86168 105018 86224 105027
rect 86168 104953 86224 104962
rect 86078 97434 86130 97440
rect 86078 97376 86130 97382
rect 85986 96278 86038 96284
rect 85986 96220 86038 96226
rect 85892 94818 85948 94827
rect 85710 94782 85762 94788
rect 85892 94753 85948 94762
rect 85710 94724 85762 94730
rect 84790 94578 84842 94584
rect 84790 94520 84842 94526
rect 84330 94374 84382 94380
rect 84330 94316 84382 94322
rect 84422 94170 84474 94176
rect 84802 94147 84830 94520
rect 84890 94478 85186 94498
rect 84946 94476 84970 94478
rect 85026 94476 85050 94478
rect 85106 94476 85130 94478
rect 84968 94424 84970 94476
rect 85032 94424 85044 94476
rect 85106 94424 85108 94476
rect 84946 94422 84970 94424
rect 85026 94422 85050 94424
rect 85106 94422 85130 94424
rect 84890 94402 85186 94422
rect 84422 94112 84474 94118
rect 84788 94138 84844 94147
rect 84054 94102 84106 94108
rect 84054 94044 84106 94050
rect 83868 94002 83924 94011
rect 83868 93937 83924 93946
rect 83962 93762 84014 93768
rect 83962 93704 84014 93710
rect 83778 92946 83830 92952
rect 83778 92888 83830 92894
rect 83686 32018 83738 32024
rect 83686 31960 83738 31966
rect 83684 30490 83740 30499
rect 83684 30425 83740 30434
rect 83594 3730 83646 3736
rect 83594 3672 83646 3678
rect 83502 2642 83554 2648
rect 83500 2610 83502 2619
rect 83554 2610 83556 2619
rect 83500 2545 83556 2554
rect 83500 2338 83556 2347
rect 83500 2273 83556 2282
rect 83514 2172 83542 2273
rect 83502 2166 83554 2172
rect 83502 2108 83554 2114
rect 83514 1492 83542 2108
rect 83502 1486 83554 1492
rect 83502 1428 83554 1434
rect 83698 880 83726 30425
rect 83790 13868 83818 92888
rect 83974 92628 84002 93704
rect 83882 92600 84002 92628
rect 83882 92492 83910 92600
rect 83882 92464 84002 92492
rect 83870 92402 83922 92408
rect 83870 92344 83922 92350
rect 83882 89280 83910 92344
rect 83974 92000 84002 92464
rect 83962 91994 84014 92000
rect 83962 91936 84014 91942
rect 83962 91858 84014 91864
rect 83960 91826 83962 91835
rect 84014 91826 84016 91835
rect 83960 91761 84016 91770
rect 83870 89274 83922 89280
rect 83870 89216 83922 89222
rect 83870 88050 83922 88056
rect 83870 87992 83922 87998
rect 83882 80984 83910 87992
rect 83870 80978 83922 80984
rect 83870 80920 83922 80926
rect 83868 46946 83924 46955
rect 83868 46881 83924 46890
rect 83882 17851 83910 46881
rect 83974 23427 84002 91761
rect 84066 90883 84094 94044
rect 84146 94034 84198 94040
rect 84146 93976 84198 93982
rect 84052 90874 84108 90883
rect 84052 90809 84108 90818
rect 84054 89954 84106 89960
rect 84054 89896 84106 89902
rect 84066 75000 84094 89896
rect 84158 89387 84186 93976
rect 84238 93150 84290 93156
rect 84238 93092 84290 93098
rect 84144 89378 84200 89387
rect 84144 89313 84200 89322
rect 84146 89274 84198 89280
rect 84146 89216 84198 89222
rect 84158 88056 84186 89216
rect 84146 88050 84198 88056
rect 84146 87992 84198 87998
rect 84146 87846 84198 87852
rect 84146 87788 84198 87794
rect 84158 85880 84186 87788
rect 84146 85874 84198 85880
rect 84146 85816 84198 85822
rect 84146 84786 84198 84792
rect 84146 84728 84198 84734
rect 84158 77283 84186 84728
rect 84250 84491 84278 93092
rect 84330 92742 84382 92748
rect 84330 92684 84382 92690
rect 84342 85987 84370 92684
rect 84434 88163 84462 94112
rect 84788 94073 84844 94082
rect 86182 94011 86210 104953
rect 86890 104814 87186 104834
rect 86946 104812 86970 104814
rect 87026 104812 87050 104814
rect 87106 104812 87130 104814
rect 86968 104760 86970 104812
rect 87032 104760 87044 104812
rect 87106 104760 87108 104812
rect 86946 104758 86970 104760
rect 87026 104758 87050 104760
rect 87106 104758 87130 104760
rect 86890 104738 87186 104758
rect 86890 103726 87186 103746
rect 86946 103724 86970 103726
rect 87026 103724 87050 103726
rect 87106 103724 87130 103726
rect 86968 103672 86970 103724
rect 87032 103672 87044 103724
rect 87106 103672 87108 103724
rect 86946 103670 86970 103672
rect 87026 103670 87050 103672
rect 87106 103670 87130 103672
rect 86890 103650 87186 103670
rect 86260 103522 86316 103531
rect 86260 103457 86316 103466
rect 86274 95400 86302 103457
rect 86890 102638 87186 102658
rect 86946 102636 86970 102638
rect 87026 102636 87050 102638
rect 87106 102636 87130 102638
rect 86968 102584 86970 102636
rect 87032 102584 87044 102636
rect 87106 102584 87108 102636
rect 86946 102582 86970 102584
rect 87026 102582 87050 102584
rect 87106 102582 87130 102584
rect 86890 102562 87186 102582
rect 86890 101550 87186 101570
rect 86946 101548 86970 101550
rect 87026 101548 87050 101550
rect 87106 101548 87130 101550
rect 86968 101496 86970 101548
rect 87032 101496 87044 101548
rect 87106 101496 87108 101548
rect 86946 101494 86970 101496
rect 87026 101494 87050 101496
rect 87106 101494 87130 101496
rect 86890 101474 87186 101494
rect 86890 100462 87186 100482
rect 86946 100460 86970 100462
rect 87026 100460 87050 100462
rect 87106 100460 87130 100462
rect 86968 100408 86970 100460
rect 87032 100408 87044 100460
rect 87106 100408 87108 100460
rect 86946 100406 86970 100408
rect 87026 100406 87050 100408
rect 87106 100406 87130 100408
rect 86890 100386 87186 100406
rect 86890 99374 87186 99394
rect 86946 99372 86970 99374
rect 87026 99372 87050 99374
rect 87106 99372 87130 99374
rect 86968 99320 86970 99372
rect 87032 99320 87044 99372
rect 87106 99320 87108 99372
rect 86946 99318 86970 99320
rect 87026 99318 87050 99320
rect 87106 99318 87130 99320
rect 86890 99298 87186 99318
rect 86538 98930 86590 98936
rect 86538 98872 86590 98878
rect 86550 96828 86578 98872
rect 86890 98286 87186 98306
rect 86946 98284 86970 98286
rect 87026 98284 87050 98286
rect 87106 98284 87130 98286
rect 86968 98232 86970 98284
rect 87032 98232 87044 98284
rect 87106 98232 87108 98284
rect 86946 98230 86970 98232
rect 87026 98230 87050 98232
rect 87106 98230 87130 98232
rect 86890 98210 87186 98230
rect 86890 97198 87186 97218
rect 86946 97196 86970 97198
rect 87026 97196 87050 97198
rect 87106 97196 87130 97198
rect 86968 97144 86970 97196
rect 87032 97144 87044 97196
rect 87106 97144 87108 97196
rect 86946 97142 86970 97144
rect 87026 97142 87050 97144
rect 87106 97142 87130 97144
rect 86890 97122 87186 97142
rect 86538 96822 86590 96828
rect 86538 96764 86590 96770
rect 86262 95394 86314 95400
rect 86262 95336 86314 95342
rect 86168 94002 86224 94011
rect 86168 93937 86224 93946
rect 84606 93626 84658 93632
rect 84606 93568 84658 93574
rect 84514 91994 84566 92000
rect 84514 91936 84566 91942
rect 84420 88154 84476 88163
rect 84420 88089 84476 88098
rect 84422 88050 84474 88056
rect 84422 87992 84474 87998
rect 84328 85978 84384 85987
rect 84328 85913 84384 85922
rect 84330 85874 84382 85880
rect 84330 85816 84382 85822
rect 84236 84482 84292 84491
rect 84236 84417 84292 84426
rect 84342 84332 84370 85816
rect 84250 84304 84370 84332
rect 84250 78507 84278 84304
rect 84330 83766 84382 83772
rect 84330 83708 84382 83714
rect 84342 79164 84370 83708
rect 84434 82179 84462 87992
rect 84526 83403 84554 91936
rect 84512 83394 84568 83403
rect 84512 83329 84568 83338
rect 84420 82170 84476 82179
rect 84420 82105 84476 82114
rect 84618 80003 84646 93568
rect 84890 93390 85186 93410
rect 84946 93388 84970 93390
rect 85026 93388 85050 93390
rect 85106 93388 85130 93390
rect 84968 93336 84970 93388
rect 85032 93336 85044 93388
rect 85106 93336 85108 93388
rect 84946 93334 84970 93336
rect 85026 93334 85050 93336
rect 85106 93334 85130 93336
rect 84890 93314 85186 93334
rect 85156 93050 85212 93059
rect 84790 93014 84842 93020
rect 85156 92985 85212 92994
rect 84790 92956 84842 92962
rect 84698 92198 84750 92204
rect 84698 92140 84750 92146
rect 84710 87075 84738 92140
rect 84696 87066 84752 87075
rect 84696 87001 84752 87010
rect 84802 80683 84830 92956
rect 85170 92680 85198 92985
rect 85158 92674 85210 92680
rect 85158 92616 85210 92622
rect 84890 92302 85186 92322
rect 84946 92300 84970 92302
rect 85026 92300 85050 92302
rect 85106 92300 85130 92302
rect 84968 92248 84970 92300
rect 85032 92248 85044 92300
rect 85106 92248 85108 92300
rect 84946 92246 84970 92248
rect 85026 92246 85050 92248
rect 85106 92246 85130 92248
rect 84890 92226 85186 92246
rect 85158 92062 85210 92068
rect 85158 92004 85210 92010
rect 85170 91971 85198 92004
rect 85156 91962 85212 91971
rect 85156 91897 85212 91906
rect 84890 91214 85186 91234
rect 84946 91212 84970 91214
rect 85026 91212 85050 91214
rect 85106 91212 85130 91214
rect 84968 91160 84970 91212
rect 85032 91160 85044 91212
rect 85106 91160 85108 91212
rect 84946 91158 84970 91160
rect 85026 91158 85050 91160
rect 85106 91158 85130 91160
rect 84890 91138 85186 91158
rect 84890 90126 85186 90146
rect 84946 90124 84970 90126
rect 85026 90124 85050 90126
rect 85106 90124 85130 90126
rect 84968 90072 84970 90124
rect 85032 90072 85044 90124
rect 85106 90072 85108 90124
rect 84946 90070 84970 90072
rect 85026 90070 85050 90072
rect 85106 90070 85130 90072
rect 84890 90050 85186 90070
rect 84890 89038 85186 89058
rect 84946 89036 84970 89038
rect 85026 89036 85050 89038
rect 85106 89036 85130 89038
rect 84968 88984 84970 89036
rect 85032 88984 85044 89036
rect 85106 88984 85108 89036
rect 84946 88982 84970 88984
rect 85026 88982 85050 88984
rect 85106 88982 85130 88984
rect 84890 88962 85186 88982
rect 84890 87950 85186 87970
rect 84946 87948 84970 87950
rect 85026 87948 85050 87950
rect 85106 87948 85130 87950
rect 84968 87896 84970 87948
rect 85032 87896 85044 87948
rect 85106 87896 85108 87948
rect 84946 87894 84970 87896
rect 85026 87894 85050 87896
rect 85106 87894 85130 87896
rect 84890 87874 85186 87894
rect 84890 86862 85186 86882
rect 84946 86860 84970 86862
rect 85026 86860 85050 86862
rect 85106 86860 85130 86862
rect 84968 86808 84970 86860
rect 85032 86808 85044 86860
rect 85106 86808 85108 86860
rect 84946 86806 84970 86808
rect 85026 86806 85050 86808
rect 85106 86806 85130 86808
rect 84890 86786 85186 86806
rect 84890 85774 85186 85794
rect 84946 85772 84970 85774
rect 85026 85772 85050 85774
rect 85106 85772 85130 85774
rect 84968 85720 84970 85772
rect 85032 85720 85044 85772
rect 85106 85720 85108 85772
rect 84946 85718 84970 85720
rect 85026 85718 85050 85720
rect 85106 85718 85130 85720
rect 84890 85698 85186 85718
rect 84890 84686 85186 84706
rect 84946 84684 84970 84686
rect 85026 84684 85050 84686
rect 85106 84684 85130 84686
rect 84968 84632 84970 84684
rect 85032 84632 85044 84684
rect 85106 84632 85108 84684
rect 84946 84630 84970 84632
rect 85026 84630 85050 84632
rect 85106 84630 85130 84632
rect 84890 84610 85186 84630
rect 84890 83598 85186 83618
rect 84946 83596 84970 83598
rect 85026 83596 85050 83598
rect 85106 83596 85130 83598
rect 84968 83544 84970 83596
rect 85032 83544 85044 83596
rect 85106 83544 85108 83596
rect 84946 83542 84970 83544
rect 85026 83542 85050 83544
rect 85106 83542 85130 83544
rect 84890 83522 85186 83542
rect 84890 82510 85186 82530
rect 84946 82508 84970 82510
rect 85026 82508 85050 82510
rect 85106 82508 85130 82510
rect 84968 82456 84970 82508
rect 85032 82456 85044 82508
rect 85106 82456 85108 82508
rect 84946 82454 84970 82456
rect 85026 82454 85050 82456
rect 85106 82454 85130 82456
rect 84890 82434 85186 82454
rect 84890 81422 85186 81442
rect 84946 81420 84970 81422
rect 85026 81420 85050 81422
rect 85106 81420 85130 81422
rect 84968 81368 84970 81420
rect 85032 81368 85044 81420
rect 85106 81368 85108 81420
rect 84946 81366 84970 81368
rect 85026 81366 85050 81368
rect 85106 81366 85130 81368
rect 84890 81346 85186 81366
rect 85250 80978 85302 80984
rect 85250 80920 85302 80926
rect 84788 80674 84844 80683
rect 84788 80609 84844 80618
rect 84890 80334 85186 80354
rect 84946 80332 84970 80334
rect 85026 80332 85050 80334
rect 85106 80332 85130 80334
rect 84968 80280 84970 80332
rect 85032 80280 85044 80332
rect 85106 80280 85108 80332
rect 84946 80278 84970 80280
rect 85026 80278 85050 80280
rect 85106 80278 85130 80280
rect 84890 80258 85186 80278
rect 84604 79994 84660 80003
rect 84604 79929 84660 79938
rect 84890 79246 85186 79266
rect 84946 79244 84970 79246
rect 85026 79244 85050 79246
rect 85106 79244 85130 79246
rect 84968 79192 84970 79244
rect 85032 79192 85044 79244
rect 85106 79192 85108 79244
rect 84946 79190 84970 79192
rect 85026 79190 85050 79192
rect 85106 79190 85130 79192
rect 84890 79170 85186 79190
rect 84342 79136 84830 79164
rect 84236 78498 84292 78507
rect 84236 78433 84292 78442
rect 84606 77374 84658 77380
rect 84606 77316 84658 77322
rect 84144 77274 84200 77283
rect 84144 77209 84200 77218
rect 84054 74994 84106 75000
rect 84054 74936 84106 74942
rect 84330 74450 84382 74456
rect 84330 74392 84382 74398
rect 84342 70211 84370 74392
rect 84618 73452 84646 77316
rect 84802 75107 84830 79136
rect 84890 78158 85186 78178
rect 84946 78156 84970 78158
rect 85026 78156 85050 78158
rect 85106 78156 85130 78158
rect 84968 78104 84970 78156
rect 85032 78104 85044 78156
rect 85106 78104 85108 78156
rect 84946 78102 84970 78104
rect 85026 78102 85050 78104
rect 85106 78102 85130 78104
rect 84890 78082 85186 78102
rect 84890 77070 85186 77090
rect 84946 77068 84970 77070
rect 85026 77068 85050 77070
rect 85106 77068 85130 77070
rect 84968 77016 84970 77068
rect 85032 77016 85044 77068
rect 85106 77016 85108 77068
rect 84946 77014 84970 77016
rect 85026 77014 85050 77016
rect 85106 77014 85130 77016
rect 84890 76994 85186 77014
rect 84890 75982 85186 76002
rect 84946 75980 84970 75982
rect 85026 75980 85050 75982
rect 85106 75980 85130 75982
rect 84968 75928 84970 75980
rect 85032 75928 85044 75980
rect 85106 75928 85108 75980
rect 84946 75926 84970 75928
rect 85026 75926 85050 75928
rect 85106 75926 85130 75928
rect 84890 75906 85186 75926
rect 84788 75098 84844 75107
rect 84788 75033 84844 75042
rect 84790 74994 84842 75000
rect 84790 74936 84842 74942
rect 84434 73424 84646 73452
rect 84328 70202 84384 70211
rect 84328 70137 84384 70146
rect 84434 69123 84462 73424
rect 84802 73316 84830 74936
rect 84890 74894 85186 74914
rect 84946 74892 84970 74894
rect 85026 74892 85050 74894
rect 85106 74892 85130 74894
rect 84968 74840 84970 74892
rect 85032 74840 85044 74892
rect 85106 74840 85108 74892
rect 84946 74838 84970 74840
rect 85026 74838 85050 74840
rect 85106 74838 85130 74840
rect 84890 74818 85186 74838
rect 84882 74518 84934 74524
rect 84882 74460 84934 74466
rect 84894 74019 84922 74460
rect 84880 74010 84936 74019
rect 84880 73945 84936 73954
rect 84890 73806 85186 73826
rect 84946 73804 84970 73806
rect 85026 73804 85050 73806
rect 85106 73804 85130 73806
rect 84968 73752 84970 73804
rect 85032 73752 85044 73804
rect 85106 73752 85108 73804
rect 84946 73750 84970 73752
rect 85026 73750 85050 73752
rect 85106 73750 85130 73752
rect 84890 73730 85186 73750
rect 84618 73288 84830 73316
rect 84618 71299 84646 73288
rect 84698 73158 84750 73164
rect 84698 73100 84750 73106
rect 84710 72523 84738 73100
rect 84790 73090 84842 73096
rect 84790 73032 84842 73038
rect 84696 72514 84752 72523
rect 84696 72449 84752 72458
rect 84604 71290 84660 71299
rect 84604 71225 84660 71234
rect 84420 69114 84476 69123
rect 84420 69049 84476 69058
rect 84802 68035 84830 73032
rect 84890 72718 85186 72738
rect 84946 72716 84970 72718
rect 85026 72716 85050 72718
rect 85106 72716 85130 72718
rect 84968 72664 84970 72716
rect 85032 72664 85044 72716
rect 85106 72664 85108 72716
rect 84946 72662 84970 72664
rect 85026 72662 85050 72664
rect 85106 72662 85130 72664
rect 84890 72642 85186 72662
rect 84890 71630 85186 71650
rect 84946 71628 84970 71630
rect 85026 71628 85050 71630
rect 85106 71628 85130 71630
rect 84968 71576 84970 71628
rect 85032 71576 85044 71628
rect 85106 71576 85108 71628
rect 84946 71574 84970 71576
rect 85026 71574 85050 71576
rect 85106 71574 85130 71576
rect 84890 71554 85186 71574
rect 84890 70542 85186 70562
rect 84946 70540 84970 70542
rect 85026 70540 85050 70542
rect 85106 70540 85130 70542
rect 84968 70488 84970 70540
rect 85032 70488 85044 70540
rect 85106 70488 85108 70540
rect 84946 70486 84970 70488
rect 85026 70486 85050 70488
rect 85106 70486 85130 70488
rect 84890 70466 85186 70486
rect 84890 69454 85186 69474
rect 84946 69452 84970 69454
rect 85026 69452 85050 69454
rect 85106 69452 85130 69454
rect 84968 69400 84970 69452
rect 85032 69400 85044 69452
rect 85106 69400 85108 69452
rect 84946 69398 84970 69400
rect 85026 69398 85050 69400
rect 85106 69398 85130 69400
rect 84890 69378 85186 69398
rect 84890 68366 85186 68386
rect 84946 68364 84970 68366
rect 85026 68364 85050 68366
rect 85106 68364 85130 68366
rect 84968 68312 84970 68364
rect 85032 68312 85044 68364
rect 85106 68312 85108 68364
rect 84946 68310 84970 68312
rect 85026 68310 85050 68312
rect 85106 68310 85130 68312
rect 84890 68290 85186 68310
rect 84788 68026 84844 68035
rect 84788 67961 84844 67970
rect 84890 67278 85186 67298
rect 84946 67276 84970 67278
rect 85026 67276 85050 67278
rect 85106 67276 85130 67278
rect 84968 67224 84970 67276
rect 85032 67224 85044 67276
rect 85106 67224 85108 67276
rect 84946 67222 84970 67224
rect 85026 67222 85050 67224
rect 85106 67222 85130 67224
rect 84890 67202 85186 67222
rect 85158 66630 85210 66636
rect 85158 66572 85210 66578
rect 85170 66539 85198 66572
rect 85156 66530 85212 66539
rect 85156 66465 85212 66474
rect 84890 66190 85186 66210
rect 84946 66188 84970 66190
rect 85026 66188 85050 66190
rect 85106 66188 85130 66190
rect 84968 66136 84970 66188
rect 85032 66136 85044 66188
rect 85106 66136 85108 66188
rect 84946 66134 84970 66136
rect 85026 66134 85050 66136
rect 85106 66134 85130 66136
rect 84890 66114 85186 66134
rect 84604 65306 84660 65315
rect 84604 65241 84660 65250
rect 84052 60546 84108 60555
rect 84052 60481 84108 60490
rect 84066 55251 84094 60481
rect 84420 55650 84476 55659
rect 84420 55585 84476 55594
rect 84052 55242 84108 55251
rect 84052 55177 84108 55186
rect 84328 45178 84384 45187
rect 84328 45113 84384 45122
rect 84144 42458 84200 42467
rect 84144 42393 84200 42402
rect 84158 35492 84186 42393
rect 84236 41370 84292 41379
rect 84236 41305 84292 41314
rect 84146 35486 84198 35492
rect 84146 35428 84198 35434
rect 84250 32092 84278 41305
rect 84238 32086 84290 32092
rect 84238 32028 84290 32034
rect 84144 31578 84200 31587
rect 84144 31513 84200 31522
rect 84054 31474 84106 31480
rect 84052 31442 84054 31451
rect 84106 31442 84108 31451
rect 84052 31377 84108 31386
rect 84158 30936 84186 31513
rect 84146 30930 84198 30936
rect 84146 30872 84198 30878
rect 84052 29946 84108 29955
rect 84052 29881 84054 29890
rect 84106 29881 84108 29890
rect 84054 29852 84106 29858
rect 83960 23418 84016 23427
rect 83960 23353 84016 23362
rect 83960 23146 84016 23155
rect 83960 23081 84016 23090
rect 83974 22980 84002 23081
rect 83962 22974 84014 22980
rect 83962 22916 84014 22922
rect 83974 18531 84002 22916
rect 84066 20056 84094 29852
rect 84342 29508 84370 45113
rect 84330 29502 84382 29508
rect 84330 29444 84382 29450
rect 84330 29366 84382 29372
rect 84330 29308 84382 29314
rect 84146 28754 84198 28760
rect 84144 28722 84146 28731
rect 84198 28722 84200 28731
rect 84144 28657 84200 28666
rect 84054 20050 84106 20056
rect 84054 19992 84106 19998
rect 84158 19868 84186 28657
rect 84238 27122 84290 27128
rect 84236 27090 84238 27099
rect 84290 27090 84292 27099
rect 84236 27025 84292 27034
rect 84342 26940 84370 29308
rect 84434 28556 84462 55585
rect 84512 54426 84568 54435
rect 84512 54361 84568 54370
rect 84422 28550 84474 28556
rect 84422 28492 84474 28498
rect 84250 26912 84370 26940
rect 84250 24068 84278 26912
rect 84328 26818 84384 26827
rect 84328 26753 84384 26762
rect 84238 24062 84290 24068
rect 84238 24004 84290 24010
rect 84236 23962 84292 23971
rect 84236 23897 84292 23906
rect 84250 23864 84278 23897
rect 84238 23858 84290 23864
rect 84238 23800 84290 23806
rect 84066 19840 84186 19868
rect 83960 18522 84016 18531
rect 83960 18457 84016 18466
rect 83962 18418 84014 18424
rect 83962 18360 84014 18366
rect 83868 17842 83924 17851
rect 83868 17777 83924 17786
rect 83778 13862 83830 13868
rect 83778 13804 83830 13810
rect 83974 12547 84002 18360
rect 84066 13635 84094 19840
rect 84250 19732 84278 23800
rect 84158 19704 84278 19732
rect 84158 17443 84186 19704
rect 84236 19610 84292 19619
rect 84236 19545 84292 19554
rect 84144 17434 84200 17443
rect 84144 17369 84200 17378
rect 84250 14859 84278 19545
rect 84342 15908 84370 26753
rect 84420 20834 84476 20843
rect 84420 20769 84476 20778
rect 84330 15902 84382 15908
rect 84330 15844 84382 15850
rect 84236 14850 84292 14859
rect 84236 14785 84292 14794
rect 84146 13862 84198 13868
rect 84146 13804 84198 13810
rect 84052 13626 84108 13635
rect 84052 13561 84108 13570
rect 83960 12538 84016 12547
rect 83960 12473 84016 12482
rect 84158 9963 84186 13804
rect 84144 9954 84200 9963
rect 84144 9889 84200 9898
rect 83960 8730 84016 8739
rect 83960 8665 84016 8674
rect 83776 4106 83832 4115
rect 83776 4041 83778 4050
rect 83830 4041 83832 4050
rect 83778 4012 83830 4018
rect 83778 3186 83830 3192
rect 83778 3128 83830 3134
rect 83790 2891 83818 3128
rect 83776 2882 83832 2891
rect 83776 2817 83832 2826
rect 83974 2483 84002 8665
rect 84330 7198 84382 7204
rect 84330 7140 84382 7146
rect 84144 5058 84200 5067
rect 84144 4993 84200 5002
rect 84052 3970 84108 3979
rect 84052 3905 84108 3914
rect 83960 2474 84016 2483
rect 83960 2409 84016 2418
rect 84066 2376 84094 3905
rect 84054 2370 84106 2376
rect 84054 2312 84106 2318
rect 83962 2302 84014 2308
rect 83962 2244 84014 2250
rect 83974 1531 84002 2244
rect 84158 2075 84186 4993
rect 84238 2982 84290 2988
rect 84238 2924 84290 2930
rect 84250 2619 84278 2924
rect 84342 2784 84370 7140
rect 84330 2778 84382 2784
rect 84330 2720 84382 2726
rect 84236 2610 84292 2619
rect 84236 2545 84292 2554
rect 84144 2066 84200 2075
rect 84144 2001 84200 2010
rect 83960 1522 84016 1531
rect 83960 1457 84016 1466
rect 83686 874 83738 880
rect 83686 816 83738 822
rect 83962 466 84014 472
rect 83960 434 83962 443
rect 84014 434 84016 443
rect 83960 369 84016 378
rect 83410 194 83462 200
rect 46150 136 46202 142
rect 81200 162 81256 171
rect 83410 136 83462 142
rect 84434 132 84462 20769
rect 84526 6812 84554 54361
rect 84618 28323 84646 65241
rect 84890 65102 85186 65122
rect 84946 65100 84970 65102
rect 85026 65100 85050 65102
rect 85106 65100 85130 65102
rect 84968 65048 84970 65100
rect 85032 65048 85044 65100
rect 85106 65048 85108 65100
rect 84946 65046 84970 65048
rect 85026 65046 85050 65048
rect 85106 65046 85130 65048
rect 84890 65026 85186 65046
rect 84890 64014 85186 64034
rect 84946 64012 84970 64014
rect 85026 64012 85050 64014
rect 85106 64012 85130 64014
rect 84968 63960 84970 64012
rect 85032 63960 85044 64012
rect 85106 63960 85108 64012
rect 84946 63958 84970 63960
rect 85026 63958 85050 63960
rect 85106 63958 85130 63960
rect 84890 63938 85186 63958
rect 84696 63810 84752 63819
rect 84696 63745 84752 63754
rect 84710 29411 84738 63745
rect 84890 62926 85186 62946
rect 84946 62924 84970 62926
rect 85026 62924 85050 62926
rect 85106 62924 85130 62926
rect 84968 62872 84970 62924
rect 85032 62872 85044 62924
rect 85106 62872 85108 62924
rect 84946 62870 84970 62872
rect 85026 62870 85050 62872
rect 85106 62870 85130 62872
rect 84890 62850 85186 62870
rect 84790 62822 84842 62828
rect 84790 62764 84842 62770
rect 84802 62731 84830 62764
rect 84788 62722 84844 62731
rect 84788 62657 84844 62666
rect 84890 61838 85186 61858
rect 84946 61836 84970 61838
rect 85026 61836 85050 61838
rect 85106 61836 85130 61838
rect 84968 61784 84970 61836
rect 85032 61784 85044 61836
rect 85106 61784 85108 61836
rect 84946 61782 84970 61784
rect 85026 61782 85050 61784
rect 85106 61782 85130 61784
rect 84890 61762 85186 61782
rect 84890 60750 85186 60770
rect 84946 60748 84970 60750
rect 85026 60748 85050 60750
rect 85106 60748 85130 60750
rect 84968 60696 84970 60748
rect 85032 60696 85044 60748
rect 85106 60696 85108 60748
rect 84946 60694 84970 60696
rect 85026 60694 85050 60696
rect 85106 60694 85130 60696
rect 84890 60674 85186 60694
rect 84890 59662 85186 59682
rect 84946 59660 84970 59662
rect 85026 59660 85050 59662
rect 85106 59660 85130 59662
rect 84968 59608 84970 59660
rect 85032 59608 85044 59660
rect 85106 59608 85108 59660
rect 84946 59606 84970 59608
rect 85026 59606 85050 59608
rect 85106 59606 85130 59608
rect 84890 59586 85186 59606
rect 84890 58574 85186 58594
rect 84946 58572 84970 58574
rect 85026 58572 85050 58574
rect 85106 58572 85130 58574
rect 84968 58520 84970 58572
rect 85032 58520 85044 58572
rect 85106 58520 85108 58572
rect 84946 58518 84970 58520
rect 85026 58518 85050 58520
rect 85106 58518 85130 58520
rect 84890 58498 85186 58518
rect 84890 57486 85186 57506
rect 84946 57484 84970 57486
rect 85026 57484 85050 57486
rect 85106 57484 85130 57486
rect 84968 57432 84970 57484
rect 85032 57432 85044 57484
rect 85106 57432 85108 57484
rect 84946 57430 84970 57432
rect 85026 57430 85050 57432
rect 85106 57430 85130 57432
rect 84890 57410 85186 57430
rect 84788 56738 84844 56747
rect 84788 56673 84844 56682
rect 84802 56504 84830 56673
rect 84790 56498 84842 56504
rect 84790 56440 84842 56446
rect 84890 56398 85186 56418
rect 84946 56396 84970 56398
rect 85026 56396 85050 56398
rect 85106 56396 85130 56398
rect 84968 56344 84970 56396
rect 85032 56344 85044 56396
rect 85106 56344 85108 56396
rect 84946 56342 84970 56344
rect 85026 56342 85050 56344
rect 85106 56342 85130 56344
rect 84890 56322 85186 56342
rect 84890 55310 85186 55330
rect 84946 55308 84970 55310
rect 85026 55308 85050 55310
rect 85106 55308 85130 55310
rect 84968 55256 84970 55308
rect 85032 55256 85044 55308
rect 85106 55256 85108 55308
rect 84946 55254 84970 55256
rect 85026 55254 85050 55256
rect 85106 55254 85130 55256
rect 84890 55234 85186 55254
rect 84890 54222 85186 54242
rect 84946 54220 84970 54222
rect 85026 54220 85050 54222
rect 85106 54220 85130 54222
rect 84968 54168 84970 54220
rect 85032 54168 85044 54220
rect 85106 54168 85108 54220
rect 84946 54166 84970 54168
rect 85026 54166 85050 54168
rect 85106 54166 85130 54168
rect 84890 54146 85186 54166
rect 84890 53134 85186 53154
rect 84946 53132 84970 53134
rect 85026 53132 85050 53134
rect 85106 53132 85130 53134
rect 84968 53080 84970 53132
rect 85032 53080 85044 53132
rect 85106 53080 85108 53132
rect 84946 53078 84970 53080
rect 85026 53078 85050 53080
rect 85106 53078 85130 53080
rect 84890 53058 85186 53078
rect 84890 52046 85186 52066
rect 84946 52044 84970 52046
rect 85026 52044 85050 52046
rect 85106 52044 85130 52046
rect 84968 51992 84970 52044
rect 85032 51992 85044 52044
rect 85106 51992 85108 52044
rect 84946 51990 84970 51992
rect 85026 51990 85050 51992
rect 85106 51990 85130 51992
rect 84890 51970 85186 51990
rect 84890 50958 85186 50978
rect 84946 50956 84970 50958
rect 85026 50956 85050 50958
rect 85106 50956 85130 50958
rect 84968 50904 84970 50956
rect 85032 50904 85044 50956
rect 85106 50904 85108 50956
rect 84946 50902 84970 50904
rect 85026 50902 85050 50904
rect 85106 50902 85130 50904
rect 84890 50882 85186 50902
rect 85156 50754 85212 50763
rect 85156 50689 85212 50698
rect 85170 50112 85198 50689
rect 85158 50106 85210 50112
rect 85158 50048 85210 50054
rect 84890 49870 85186 49890
rect 84946 49868 84970 49870
rect 85026 49868 85050 49870
rect 85106 49868 85130 49870
rect 84968 49816 84970 49868
rect 85032 49816 85044 49868
rect 85106 49816 85108 49868
rect 84946 49814 84970 49816
rect 85026 49814 85050 49816
rect 85106 49814 85130 49816
rect 84890 49794 85186 49814
rect 84788 49666 84844 49675
rect 84788 49601 84844 49610
rect 84802 48888 84830 49601
rect 84790 48882 84842 48888
rect 84790 48824 84842 48830
rect 84890 48782 85186 48802
rect 84946 48780 84970 48782
rect 85026 48780 85050 48782
rect 85106 48780 85130 48782
rect 84968 48728 84970 48780
rect 85032 48728 85044 48780
rect 85106 48728 85108 48780
rect 84946 48726 84970 48728
rect 85026 48726 85050 48728
rect 85106 48726 85130 48728
rect 84890 48706 85186 48726
rect 84890 47694 85186 47714
rect 84946 47692 84970 47694
rect 85026 47692 85050 47694
rect 85106 47692 85130 47694
rect 84968 47640 84970 47692
rect 85032 47640 85044 47692
rect 85106 47640 85108 47692
rect 84946 47638 84970 47640
rect 85026 47638 85050 47640
rect 85106 47638 85130 47640
rect 84890 47618 85186 47638
rect 84890 46606 85186 46626
rect 84946 46604 84970 46606
rect 85026 46604 85050 46606
rect 85106 46604 85130 46606
rect 84968 46552 84970 46604
rect 85032 46552 85044 46604
rect 85106 46552 85108 46604
rect 84946 46550 84970 46552
rect 85026 46550 85050 46552
rect 85106 46550 85130 46552
rect 84890 46530 85186 46550
rect 84890 45518 85186 45538
rect 84946 45516 84970 45518
rect 85026 45516 85050 45518
rect 85106 45516 85130 45518
rect 84968 45464 84970 45516
rect 85032 45464 85044 45516
rect 85106 45464 85108 45516
rect 84946 45462 84970 45464
rect 85026 45462 85050 45464
rect 85106 45462 85130 45464
rect 84890 45442 85186 45462
rect 84890 44430 85186 44450
rect 84946 44428 84970 44430
rect 85026 44428 85050 44430
rect 85106 44428 85130 44430
rect 84968 44376 84970 44428
rect 85032 44376 85044 44428
rect 85106 44376 85108 44428
rect 84946 44374 84970 44376
rect 85026 44374 85050 44376
rect 85106 44374 85130 44376
rect 84890 44354 85186 44374
rect 85156 43682 85212 43691
rect 85156 43617 85158 43626
rect 85210 43617 85212 43626
rect 85158 43588 85210 43594
rect 84890 43342 85186 43362
rect 84946 43340 84970 43342
rect 85026 43340 85050 43342
rect 85106 43340 85130 43342
rect 84968 43288 84970 43340
rect 85032 43288 85044 43340
rect 85106 43288 85108 43340
rect 84946 43286 84970 43288
rect 85026 43286 85050 43288
rect 85106 43286 85130 43288
rect 84890 43266 85186 43286
rect 84890 42254 85186 42274
rect 84946 42252 84970 42254
rect 85026 42252 85050 42254
rect 85106 42252 85130 42254
rect 84968 42200 84970 42252
rect 85032 42200 85044 42252
rect 85106 42200 85108 42252
rect 84946 42198 84970 42200
rect 85026 42198 85050 42200
rect 85106 42198 85130 42200
rect 84890 42178 85186 42198
rect 84890 41166 85186 41186
rect 84946 41164 84970 41166
rect 85026 41164 85050 41166
rect 85106 41164 85130 41166
rect 84968 41112 84970 41164
rect 85032 41112 85044 41164
rect 85106 41112 85108 41164
rect 84946 41110 84970 41112
rect 85026 41110 85050 41112
rect 85106 41110 85130 41112
rect 84890 41090 85186 41110
rect 84890 40078 85186 40098
rect 84946 40076 84970 40078
rect 85026 40076 85050 40078
rect 85106 40076 85130 40078
rect 84968 40024 84970 40076
rect 85032 40024 85044 40076
rect 85106 40024 85108 40076
rect 84946 40022 84970 40024
rect 85026 40022 85050 40024
rect 85106 40022 85130 40024
rect 84890 40002 85186 40022
rect 84790 39974 84842 39980
rect 84790 39916 84842 39922
rect 84802 39883 84830 39916
rect 84788 39874 84844 39883
rect 84788 39809 84844 39818
rect 84890 38990 85186 39010
rect 84946 38988 84970 38990
rect 85026 38988 85050 38990
rect 85106 38988 85130 38990
rect 84968 38936 84970 38988
rect 85032 38936 85044 38988
rect 85106 38936 85108 38988
rect 84946 38934 84970 38936
rect 85026 38934 85050 38936
rect 85106 38934 85130 38936
rect 84890 38914 85186 38934
rect 84890 37902 85186 37922
rect 84946 37900 84970 37902
rect 85026 37900 85050 37902
rect 85106 37900 85130 37902
rect 84968 37848 84970 37900
rect 85032 37848 85044 37900
rect 85106 37848 85108 37900
rect 84946 37846 84970 37848
rect 85026 37846 85050 37848
rect 85106 37846 85130 37848
rect 84890 37826 85186 37846
rect 84890 36814 85186 36834
rect 84946 36812 84970 36814
rect 85026 36812 85050 36814
rect 85106 36812 85130 36814
rect 84968 36760 84970 36812
rect 85032 36760 85044 36812
rect 85106 36760 85108 36812
rect 84946 36758 84970 36760
rect 85026 36758 85050 36760
rect 85106 36758 85130 36760
rect 84890 36738 85186 36758
rect 84788 36474 84844 36483
rect 84788 36409 84844 36418
rect 84802 29440 84830 36409
rect 84890 35726 85186 35746
rect 84946 35724 84970 35726
rect 85026 35724 85050 35726
rect 85106 35724 85130 35726
rect 84968 35672 84970 35724
rect 85032 35672 85044 35724
rect 85106 35672 85108 35724
rect 84946 35670 84970 35672
rect 85026 35670 85050 35672
rect 85106 35670 85130 35672
rect 84890 35650 85186 35670
rect 84890 34638 85186 34658
rect 84946 34636 84970 34638
rect 85026 34636 85050 34638
rect 85106 34636 85130 34638
rect 84968 34584 84970 34636
rect 85032 34584 85044 34636
rect 85106 34584 85108 34636
rect 84946 34582 84970 34584
rect 85026 34582 85050 34584
rect 85106 34582 85130 34584
rect 84890 34562 85186 34582
rect 84890 33550 85186 33570
rect 84946 33548 84970 33550
rect 85026 33548 85050 33550
rect 85106 33548 85130 33550
rect 84968 33496 84970 33548
rect 85032 33496 85044 33548
rect 85106 33496 85108 33548
rect 84946 33494 84970 33496
rect 85026 33494 85050 33496
rect 85106 33494 85130 33496
rect 84890 33474 85186 33494
rect 84890 32462 85186 32482
rect 84946 32460 84970 32462
rect 85026 32460 85050 32462
rect 85106 32460 85130 32462
rect 84968 32408 84970 32460
rect 85032 32408 85044 32460
rect 85106 32408 85108 32460
rect 84946 32406 84970 32408
rect 85026 32406 85050 32408
rect 85106 32406 85130 32408
rect 84890 32386 85186 32406
rect 84890 31374 85186 31394
rect 84946 31372 84970 31374
rect 85026 31372 85050 31374
rect 85106 31372 85130 31374
rect 84968 31320 84970 31372
rect 85032 31320 85044 31372
rect 85106 31320 85108 31372
rect 84946 31318 84970 31320
rect 85026 31318 85050 31320
rect 85106 31318 85130 31320
rect 84890 31298 85186 31318
rect 84890 30286 85186 30306
rect 84946 30284 84970 30286
rect 85026 30284 85050 30286
rect 85106 30284 85130 30286
rect 84968 30232 84970 30284
rect 85032 30232 85044 30284
rect 85106 30232 85108 30284
rect 84946 30230 84970 30232
rect 85026 30230 85050 30232
rect 85106 30230 85130 30232
rect 84890 30210 85186 30230
rect 84790 29434 84842 29440
rect 84696 29402 84752 29411
rect 84790 29376 84842 29382
rect 84696 29337 84752 29346
rect 84890 29198 85186 29218
rect 84946 29196 84970 29198
rect 85026 29196 85050 29198
rect 85106 29196 85130 29198
rect 84968 29144 84970 29196
rect 85032 29144 85044 29196
rect 85106 29144 85108 29196
rect 84946 29142 84970 29144
rect 85026 29142 85050 29144
rect 85106 29142 85130 29144
rect 84890 29122 85186 29142
rect 84696 28994 84752 29003
rect 84696 28929 84752 28938
rect 84604 28314 84660 28323
rect 84604 28249 84660 28258
rect 84710 28216 84738 28929
rect 84698 28210 84750 28216
rect 84698 28152 84750 28158
rect 84890 28110 85186 28130
rect 84946 28108 84970 28110
rect 85026 28108 85050 28110
rect 85106 28108 85130 28110
rect 84968 28056 84970 28108
rect 85032 28056 85044 28108
rect 85106 28056 85108 28108
rect 84946 28054 84970 28056
rect 85026 28054 85050 28056
rect 85106 28054 85130 28056
rect 84890 28034 85186 28054
rect 84698 27122 84750 27128
rect 84698 27064 84750 27070
rect 84604 24506 84660 24515
rect 84604 24441 84660 24450
rect 84618 16604 84646 24441
rect 84710 24243 84738 27064
rect 84890 27022 85186 27042
rect 84946 27020 84970 27022
rect 85026 27020 85050 27022
rect 85106 27020 85130 27022
rect 84968 26968 84970 27020
rect 85032 26968 85044 27020
rect 85106 26968 85108 27020
rect 84946 26966 84970 26968
rect 85026 26966 85050 26968
rect 85106 26966 85130 26968
rect 84890 26946 85186 26966
rect 84890 25934 85186 25954
rect 84946 25932 84970 25934
rect 85026 25932 85050 25934
rect 85106 25932 85130 25934
rect 84968 25880 84970 25932
rect 85032 25880 85044 25932
rect 85106 25880 85108 25932
rect 84946 25878 84970 25880
rect 85026 25878 85050 25880
rect 85106 25878 85130 25880
rect 84890 25858 85186 25878
rect 84882 25626 84934 25632
rect 84880 25594 84882 25603
rect 84934 25594 84936 25603
rect 84880 25529 84936 25538
rect 84890 24846 85186 24866
rect 84946 24844 84970 24846
rect 85026 24844 85050 24846
rect 85106 24844 85130 24846
rect 84968 24792 84970 24844
rect 85032 24792 85044 24844
rect 85106 24792 85108 24844
rect 84946 24790 84970 24792
rect 85026 24790 85050 24792
rect 85106 24790 85130 24792
rect 84890 24770 85186 24790
rect 84696 24234 84752 24243
rect 84696 24169 84752 24178
rect 84698 24062 84750 24068
rect 84698 24004 84750 24010
rect 84710 16740 84738 24004
rect 84890 23758 85186 23778
rect 84946 23756 84970 23758
rect 85026 23756 85050 23758
rect 85106 23756 85130 23758
rect 84968 23704 84970 23756
rect 85032 23704 85044 23756
rect 85106 23704 85108 23756
rect 84946 23702 84970 23704
rect 85026 23702 85050 23704
rect 85106 23702 85130 23704
rect 84890 23682 85186 23702
rect 84890 22670 85186 22690
rect 84946 22668 84970 22670
rect 85026 22668 85050 22670
rect 85106 22668 85130 22670
rect 84968 22616 84970 22668
rect 85032 22616 85044 22668
rect 85106 22616 85108 22668
rect 84946 22614 84970 22616
rect 85026 22614 85050 22616
rect 85106 22614 85130 22616
rect 84890 22594 85186 22614
rect 84890 21582 85186 21602
rect 84946 21580 84970 21582
rect 85026 21580 85050 21582
rect 85106 21580 85130 21582
rect 84968 21528 84970 21580
rect 85032 21528 85044 21580
rect 85106 21528 85108 21580
rect 84946 21526 84970 21528
rect 85026 21526 85050 21528
rect 85106 21526 85130 21528
rect 84890 21506 85186 21526
rect 84890 20494 85186 20514
rect 84946 20492 84970 20494
rect 85026 20492 85050 20494
rect 85106 20492 85130 20494
rect 84968 20440 84970 20492
rect 85032 20440 85044 20492
rect 85106 20440 85108 20492
rect 84946 20438 84970 20440
rect 85026 20438 85050 20440
rect 85106 20438 85130 20440
rect 84890 20418 85186 20438
rect 84790 20254 84842 20260
rect 84790 20196 84842 20202
rect 84802 17012 84830 20196
rect 84890 19406 85186 19426
rect 84946 19404 84970 19406
rect 85026 19404 85050 19406
rect 85106 19404 85130 19406
rect 84968 19352 84970 19404
rect 85032 19352 85044 19404
rect 85106 19352 85108 19404
rect 84946 19350 84970 19352
rect 85026 19350 85050 19352
rect 85106 19350 85130 19352
rect 84890 19330 85186 19350
rect 84890 18318 85186 18338
rect 84946 18316 84970 18318
rect 85026 18316 85050 18318
rect 85106 18316 85130 18318
rect 84968 18264 84970 18316
rect 85032 18264 85044 18316
rect 85106 18264 85108 18316
rect 84946 18262 84970 18264
rect 85026 18262 85050 18264
rect 85106 18262 85130 18264
rect 84890 18242 85186 18262
rect 84890 17230 85186 17250
rect 84946 17228 84970 17230
rect 85026 17228 85050 17230
rect 85106 17228 85130 17230
rect 84968 17176 84970 17228
rect 85032 17176 85044 17228
rect 85106 17176 85108 17228
rect 84946 17174 84970 17176
rect 85026 17174 85050 17176
rect 85106 17174 85130 17176
rect 84890 17154 85186 17174
rect 84802 16984 84922 17012
rect 84710 16712 84830 16740
rect 84618 16576 84738 16604
rect 84606 15902 84658 15908
rect 84606 15844 84658 15850
rect 84618 6948 84646 15844
rect 84710 7084 84738 16576
rect 84802 7204 84830 16712
rect 84894 16355 84922 16984
rect 84880 16346 84936 16355
rect 84880 16281 84936 16290
rect 84890 16142 85186 16162
rect 84946 16140 84970 16142
rect 85026 16140 85050 16142
rect 85106 16140 85130 16142
rect 84968 16088 84970 16140
rect 85032 16088 85044 16140
rect 85106 16088 85108 16140
rect 84946 16086 84970 16088
rect 85026 16086 85050 16088
rect 85106 16086 85130 16088
rect 84890 16066 85186 16086
rect 84890 15054 85186 15074
rect 84946 15052 84970 15054
rect 85026 15052 85050 15054
rect 85106 15052 85130 15054
rect 84968 15000 84970 15052
rect 85032 15000 85044 15052
rect 85106 15000 85108 15052
rect 84946 14998 84970 15000
rect 85026 14998 85050 15000
rect 85106 14998 85130 15000
rect 84890 14978 85186 14998
rect 84890 13966 85186 13986
rect 84946 13964 84970 13966
rect 85026 13964 85050 13966
rect 85106 13964 85130 13966
rect 84968 13912 84970 13964
rect 85032 13912 85044 13964
rect 85106 13912 85108 13964
rect 84946 13910 84970 13912
rect 85026 13910 85050 13912
rect 85106 13910 85130 13912
rect 84890 13890 85186 13910
rect 84890 12878 85186 12898
rect 84946 12876 84970 12878
rect 85026 12876 85050 12878
rect 85106 12876 85130 12878
rect 84968 12824 84970 12876
rect 85032 12824 85044 12876
rect 85106 12824 85108 12876
rect 84946 12822 84970 12824
rect 85026 12822 85050 12824
rect 85106 12822 85130 12824
rect 84890 12802 85186 12822
rect 84890 11790 85186 11810
rect 84946 11788 84970 11790
rect 85026 11788 85050 11790
rect 85106 11788 85130 11790
rect 84968 11736 84970 11788
rect 85032 11736 85044 11788
rect 85106 11736 85108 11788
rect 84946 11734 84970 11736
rect 85026 11734 85050 11736
rect 85106 11734 85130 11736
rect 84890 11714 85186 11734
rect 84890 10702 85186 10722
rect 84946 10700 84970 10702
rect 85026 10700 85050 10702
rect 85106 10700 85130 10702
rect 84968 10648 84970 10700
rect 85032 10648 85044 10700
rect 85106 10648 85108 10700
rect 84946 10646 84970 10648
rect 85026 10646 85050 10648
rect 85106 10646 85130 10648
rect 84890 10626 85186 10646
rect 84890 9614 85186 9634
rect 84946 9612 84970 9614
rect 85026 9612 85050 9614
rect 85106 9612 85130 9614
rect 84968 9560 84970 9612
rect 85032 9560 85044 9612
rect 85106 9560 85108 9612
rect 84946 9558 84970 9560
rect 85026 9558 85050 9560
rect 85106 9558 85130 9560
rect 84890 9538 85186 9558
rect 84890 8526 85186 8546
rect 84946 8524 84970 8526
rect 85026 8524 85050 8526
rect 85106 8524 85130 8526
rect 84968 8472 84970 8524
rect 85032 8472 85044 8524
rect 85106 8472 85108 8524
rect 84946 8470 84970 8472
rect 85026 8470 85050 8472
rect 85106 8470 85130 8472
rect 84890 8450 85186 8470
rect 85064 7642 85120 7651
rect 85064 7577 85066 7586
rect 85118 7577 85120 7586
rect 85066 7548 85118 7554
rect 84890 7438 85186 7458
rect 84946 7436 84970 7438
rect 85026 7436 85050 7438
rect 85106 7436 85130 7438
rect 84968 7384 84970 7436
rect 85032 7384 85044 7436
rect 85106 7384 85108 7436
rect 84946 7382 84970 7384
rect 85026 7382 85050 7384
rect 85106 7382 85130 7384
rect 84890 7362 85186 7382
rect 84790 7198 84842 7204
rect 84790 7140 84842 7146
rect 84710 7056 84830 7084
rect 84618 6920 84738 6948
rect 84526 6784 84646 6812
rect 84512 6554 84568 6563
rect 84512 6489 84568 6498
rect 84526 1939 84554 6489
rect 84512 1930 84568 1939
rect 84512 1865 84568 1874
rect 84618 1832 84646 6784
rect 84606 1826 84658 1832
rect 84606 1768 84658 1774
rect 84710 1764 84738 6920
rect 84802 2920 84830 7056
rect 84890 6350 85186 6370
rect 84946 6348 84970 6350
rect 85026 6348 85050 6350
rect 85106 6348 85130 6350
rect 84968 6296 84970 6348
rect 85032 6296 85044 6348
rect 85106 6296 85108 6348
rect 84946 6294 84970 6296
rect 85026 6294 85050 6296
rect 85106 6294 85130 6296
rect 84890 6274 85186 6294
rect 84890 5262 85186 5282
rect 84946 5260 84970 5262
rect 85026 5260 85050 5262
rect 85106 5260 85130 5262
rect 84968 5208 84970 5260
rect 85032 5208 85044 5260
rect 85106 5208 85108 5260
rect 84946 5206 84970 5208
rect 85026 5206 85050 5208
rect 85106 5206 85130 5208
rect 84890 5186 85186 5206
rect 84890 4174 85186 4194
rect 84946 4172 84970 4174
rect 85026 4172 85050 4174
rect 85106 4172 85130 4174
rect 84968 4120 84970 4172
rect 85032 4120 85044 4172
rect 85106 4120 85108 4172
rect 84946 4118 84970 4120
rect 85026 4118 85050 4120
rect 85106 4118 85130 4120
rect 84890 4098 85186 4118
rect 84890 3086 85186 3106
rect 84946 3084 84970 3086
rect 85026 3084 85050 3086
rect 85106 3084 85130 3086
rect 84968 3032 84970 3084
rect 85032 3032 85044 3084
rect 85106 3032 85108 3084
rect 84946 3030 84970 3032
rect 85026 3030 85050 3032
rect 85106 3030 85130 3032
rect 84890 3010 85186 3030
rect 84790 2914 84842 2920
rect 84790 2856 84842 2862
rect 84974 2914 85026 2920
rect 84974 2856 85026 2862
rect 84986 2648 85014 2856
rect 84974 2642 85026 2648
rect 84974 2584 85026 2590
rect 85262 2240 85290 80920
rect 85800 48442 85856 48451
rect 85800 48377 85856 48386
rect 85342 32018 85394 32024
rect 85342 31960 85394 31966
rect 85354 2988 85382 31960
rect 85434 28278 85486 28284
rect 85434 28220 85486 28226
rect 85446 3532 85474 28220
rect 85526 19642 85578 19648
rect 85524 19610 85526 19619
rect 85578 19610 85580 19619
rect 85524 19545 85580 19554
rect 85434 3526 85486 3532
rect 85434 3468 85486 3474
rect 85342 2982 85394 2988
rect 85342 2924 85394 2930
rect 85250 2234 85302 2240
rect 85250 2176 85302 2182
rect 84890 1998 85186 2018
rect 84946 1996 84970 1998
rect 85026 1996 85050 1998
rect 85106 1996 85130 1998
rect 84968 1944 84970 1996
rect 85032 1944 85044 1996
rect 85106 1944 85108 1996
rect 84946 1942 84970 1944
rect 85026 1942 85050 1944
rect 85106 1942 85130 1944
rect 84890 1922 85186 1942
rect 84698 1758 84750 1764
rect 84698 1700 84750 1706
rect 81200 97 81256 106
rect 84422 126 84474 132
rect 84422 68 84474 74
rect 85538 64 85566 19545
rect 85814 3396 85842 48377
rect 85892 45858 85948 45867
rect 85892 45793 85948 45802
rect 85802 3390 85854 3396
rect 85802 3332 85854 3338
rect 85906 2852 85934 45793
rect 85986 31474 86038 31480
rect 85986 31416 86038 31422
rect 85998 11051 86026 31416
rect 85984 11042 86040 11051
rect 85984 10977 86040 10986
rect 85894 2846 85946 2852
rect 85894 2788 85946 2794
rect 86550 2784 86578 96764
rect 86630 96754 86682 96760
rect 86630 96696 86682 96702
rect 86642 2920 86670 96696
rect 86890 96110 87186 96130
rect 86946 96108 86970 96110
rect 87026 96108 87050 96110
rect 87106 96108 87130 96110
rect 86968 96056 86970 96108
rect 87032 96056 87044 96108
rect 87106 96056 87108 96108
rect 86946 96054 86970 96056
rect 87026 96054 87050 96056
rect 87106 96054 87130 96056
rect 86890 96034 87186 96054
rect 86890 95022 87186 95042
rect 86946 95020 86970 95022
rect 87026 95020 87050 95022
rect 87106 95020 87130 95022
rect 86968 94968 86970 95020
rect 87032 94968 87044 95020
rect 87106 94968 87108 95020
rect 86946 94966 86970 94968
rect 87026 94966 87050 94968
rect 87106 94966 87130 94968
rect 86890 94946 87186 94966
rect 86890 93934 87186 93954
rect 86946 93932 86970 93934
rect 87026 93932 87050 93934
rect 87106 93932 87130 93934
rect 86968 93880 86970 93932
rect 87032 93880 87044 93932
rect 87106 93880 87108 93932
rect 86946 93878 86970 93880
rect 87026 93878 87050 93880
rect 87106 93878 87130 93880
rect 86890 93858 87186 93878
rect 86890 92846 87186 92866
rect 86946 92844 86970 92846
rect 87026 92844 87050 92846
rect 87106 92844 87130 92846
rect 86968 92792 86970 92844
rect 87032 92792 87044 92844
rect 87106 92792 87108 92844
rect 86946 92790 86970 92792
rect 87026 92790 87050 92792
rect 87106 92790 87130 92792
rect 86890 92770 87186 92790
rect 86890 91758 87186 91778
rect 86946 91756 86970 91758
rect 87026 91756 87050 91758
rect 87106 91756 87130 91758
rect 86968 91704 86970 91756
rect 87032 91704 87044 91756
rect 87106 91704 87108 91756
rect 86946 91702 86970 91704
rect 87026 91702 87050 91704
rect 87106 91702 87130 91704
rect 86890 91682 87186 91702
rect 86890 90670 87186 90690
rect 86946 90668 86970 90670
rect 87026 90668 87050 90670
rect 87106 90668 87130 90670
rect 86968 90616 86970 90668
rect 87032 90616 87044 90668
rect 87106 90616 87108 90668
rect 86946 90614 86970 90616
rect 87026 90614 87050 90616
rect 87106 90614 87130 90616
rect 86890 90594 87186 90614
rect 86890 89582 87186 89602
rect 86946 89580 86970 89582
rect 87026 89580 87050 89582
rect 87106 89580 87130 89582
rect 86968 89528 86970 89580
rect 87032 89528 87044 89580
rect 87106 89528 87108 89580
rect 86946 89526 86970 89528
rect 87026 89526 87050 89528
rect 87106 89526 87130 89528
rect 86890 89506 87186 89526
rect 86890 88494 87186 88514
rect 86946 88492 86970 88494
rect 87026 88492 87050 88494
rect 87106 88492 87130 88494
rect 86968 88440 86970 88492
rect 87032 88440 87044 88492
rect 87106 88440 87108 88492
rect 86946 88438 86970 88440
rect 87026 88438 87050 88440
rect 87106 88438 87130 88440
rect 86890 88418 87186 88438
rect 86890 87406 87186 87426
rect 86946 87404 86970 87406
rect 87026 87404 87050 87406
rect 87106 87404 87130 87406
rect 86968 87352 86970 87404
rect 87032 87352 87044 87404
rect 87106 87352 87108 87404
rect 86946 87350 86970 87352
rect 87026 87350 87050 87352
rect 87106 87350 87130 87352
rect 86890 87330 87186 87350
rect 86890 86318 87186 86338
rect 86946 86316 86970 86318
rect 87026 86316 87050 86318
rect 87106 86316 87130 86318
rect 86968 86264 86970 86316
rect 87032 86264 87044 86316
rect 87106 86264 87108 86316
rect 86946 86262 86970 86264
rect 87026 86262 87050 86264
rect 87106 86262 87130 86264
rect 86890 86242 87186 86262
rect 86890 85230 87186 85250
rect 86946 85228 86970 85230
rect 87026 85228 87050 85230
rect 87106 85228 87130 85230
rect 86968 85176 86970 85228
rect 87032 85176 87044 85228
rect 87106 85176 87108 85228
rect 86946 85174 86970 85176
rect 87026 85174 87050 85176
rect 87106 85174 87130 85176
rect 86890 85154 87186 85174
rect 86890 84142 87186 84162
rect 86946 84140 86970 84142
rect 87026 84140 87050 84142
rect 87106 84140 87130 84142
rect 86968 84088 86970 84140
rect 87032 84088 87044 84140
rect 87106 84088 87108 84140
rect 86946 84086 86970 84088
rect 87026 84086 87050 84088
rect 87106 84086 87130 84088
rect 86890 84066 87186 84086
rect 86890 83054 87186 83074
rect 86946 83052 86970 83054
rect 87026 83052 87050 83054
rect 87106 83052 87130 83054
rect 86968 83000 86970 83052
rect 87032 83000 87044 83052
rect 87106 83000 87108 83052
rect 86946 82998 86970 83000
rect 87026 82998 87050 83000
rect 87106 82998 87130 83000
rect 86890 82978 87186 82998
rect 86890 81966 87186 81986
rect 86946 81964 86970 81966
rect 87026 81964 87050 81966
rect 87106 81964 87130 81966
rect 86968 81912 86970 81964
rect 87032 81912 87044 81964
rect 87106 81912 87108 81964
rect 86946 81910 86970 81912
rect 87026 81910 87050 81912
rect 87106 81910 87130 81912
rect 86890 81890 87186 81910
rect 86890 80878 87186 80898
rect 86946 80876 86970 80878
rect 87026 80876 87050 80878
rect 87106 80876 87130 80878
rect 86968 80824 86970 80876
rect 87032 80824 87044 80876
rect 87106 80824 87108 80876
rect 86946 80822 86970 80824
rect 87026 80822 87050 80824
rect 87106 80822 87130 80824
rect 86890 80802 87186 80822
rect 86890 79790 87186 79810
rect 86946 79788 86970 79790
rect 87026 79788 87050 79790
rect 87106 79788 87130 79790
rect 86968 79736 86970 79788
rect 87032 79736 87044 79788
rect 87106 79736 87108 79788
rect 86946 79734 86970 79736
rect 87026 79734 87050 79736
rect 87106 79734 87130 79736
rect 86890 79714 87186 79734
rect 86890 78702 87186 78722
rect 86946 78700 86970 78702
rect 87026 78700 87050 78702
rect 87106 78700 87130 78702
rect 86968 78648 86970 78700
rect 87032 78648 87044 78700
rect 87106 78648 87108 78700
rect 86946 78646 86970 78648
rect 87026 78646 87050 78648
rect 87106 78646 87130 78648
rect 86890 78626 87186 78646
rect 86890 77614 87186 77634
rect 86946 77612 86970 77614
rect 87026 77612 87050 77614
rect 87106 77612 87130 77614
rect 86968 77560 86970 77612
rect 87032 77560 87044 77612
rect 87106 77560 87108 77612
rect 86946 77558 86970 77560
rect 87026 77558 87050 77560
rect 87106 77558 87130 77560
rect 86890 77538 87186 77558
rect 86890 76526 87186 76546
rect 86946 76524 86970 76526
rect 87026 76524 87050 76526
rect 87106 76524 87130 76526
rect 86968 76472 86970 76524
rect 87032 76472 87044 76524
rect 87106 76472 87108 76524
rect 86946 76470 86970 76472
rect 87026 76470 87050 76472
rect 87106 76470 87130 76472
rect 86890 76450 87186 76470
rect 86890 75438 87186 75458
rect 86946 75436 86970 75438
rect 87026 75436 87050 75438
rect 87106 75436 87130 75438
rect 86968 75384 86970 75436
rect 87032 75384 87044 75436
rect 87106 75384 87108 75436
rect 86946 75382 86970 75384
rect 87026 75382 87050 75384
rect 87106 75382 87130 75384
rect 86890 75362 87186 75382
rect 86890 74350 87186 74370
rect 86946 74348 86970 74350
rect 87026 74348 87050 74350
rect 87106 74348 87130 74350
rect 86968 74296 86970 74348
rect 87032 74296 87044 74348
rect 87106 74296 87108 74348
rect 86946 74294 86970 74296
rect 87026 74294 87050 74296
rect 87106 74294 87130 74296
rect 86890 74274 87186 74294
rect 86890 73262 87186 73282
rect 86946 73260 86970 73262
rect 87026 73260 87050 73262
rect 87106 73260 87130 73262
rect 86968 73208 86970 73260
rect 87032 73208 87044 73260
rect 87106 73208 87108 73260
rect 86946 73206 86970 73208
rect 87026 73206 87050 73208
rect 87106 73206 87130 73208
rect 86890 73186 87186 73206
rect 86890 72174 87186 72194
rect 86946 72172 86970 72174
rect 87026 72172 87050 72174
rect 87106 72172 87130 72174
rect 86968 72120 86970 72172
rect 87032 72120 87044 72172
rect 87106 72120 87108 72172
rect 86946 72118 86970 72120
rect 87026 72118 87050 72120
rect 87106 72118 87130 72120
rect 86890 72098 87186 72118
rect 86890 71086 87186 71106
rect 86946 71084 86970 71086
rect 87026 71084 87050 71086
rect 87106 71084 87130 71086
rect 86968 71032 86970 71084
rect 87032 71032 87044 71084
rect 87106 71032 87108 71084
rect 86946 71030 86970 71032
rect 87026 71030 87050 71032
rect 87106 71030 87130 71032
rect 86890 71010 87186 71030
rect 86890 69998 87186 70018
rect 86946 69996 86970 69998
rect 87026 69996 87050 69998
rect 87106 69996 87130 69998
rect 86968 69944 86970 69996
rect 87032 69944 87044 69996
rect 87106 69944 87108 69996
rect 86946 69942 86970 69944
rect 87026 69942 87050 69944
rect 87106 69942 87130 69944
rect 86890 69922 87186 69942
rect 86890 68910 87186 68930
rect 86946 68908 86970 68910
rect 87026 68908 87050 68910
rect 87106 68908 87130 68910
rect 86968 68856 86970 68908
rect 87032 68856 87044 68908
rect 87106 68856 87108 68908
rect 86946 68854 86970 68856
rect 87026 68854 87050 68856
rect 87106 68854 87130 68856
rect 86890 68834 87186 68854
rect 86890 67822 87186 67842
rect 86946 67820 86970 67822
rect 87026 67820 87050 67822
rect 87106 67820 87130 67822
rect 86968 67768 86970 67820
rect 87032 67768 87044 67820
rect 87106 67768 87108 67820
rect 86946 67766 86970 67768
rect 87026 67766 87050 67768
rect 87106 67766 87130 67768
rect 86890 67746 87186 67766
rect 86890 66734 87186 66754
rect 86946 66732 86970 66734
rect 87026 66732 87050 66734
rect 87106 66732 87130 66734
rect 86968 66680 86970 66732
rect 87032 66680 87044 66732
rect 87106 66680 87108 66732
rect 86946 66678 86970 66680
rect 87026 66678 87050 66680
rect 87106 66678 87130 66680
rect 86890 66658 87186 66678
rect 86890 65646 87186 65666
rect 86946 65644 86970 65646
rect 87026 65644 87050 65646
rect 87106 65644 87130 65646
rect 86968 65592 86970 65644
rect 87032 65592 87044 65644
rect 87106 65592 87108 65644
rect 86946 65590 86970 65592
rect 87026 65590 87050 65592
rect 87106 65590 87130 65592
rect 86890 65570 87186 65590
rect 86890 64558 87186 64578
rect 86946 64556 86970 64558
rect 87026 64556 87050 64558
rect 87106 64556 87130 64558
rect 86968 64504 86970 64556
rect 87032 64504 87044 64556
rect 87106 64504 87108 64556
rect 86946 64502 86970 64504
rect 87026 64502 87050 64504
rect 87106 64502 87130 64504
rect 86890 64482 87186 64502
rect 86890 63470 87186 63490
rect 86946 63468 86970 63470
rect 87026 63468 87050 63470
rect 87106 63468 87130 63470
rect 86968 63416 86970 63468
rect 87032 63416 87044 63468
rect 87106 63416 87108 63468
rect 86946 63414 86970 63416
rect 87026 63414 87050 63416
rect 87106 63414 87130 63416
rect 86890 63394 87186 63414
rect 86890 62382 87186 62402
rect 86946 62380 86970 62382
rect 87026 62380 87050 62382
rect 87106 62380 87130 62382
rect 86968 62328 86970 62380
rect 87032 62328 87044 62380
rect 87106 62328 87108 62380
rect 86946 62326 86970 62328
rect 87026 62326 87050 62328
rect 87106 62326 87130 62328
rect 86890 62306 87186 62326
rect 86890 61294 87186 61314
rect 86946 61292 86970 61294
rect 87026 61292 87050 61294
rect 87106 61292 87130 61294
rect 86968 61240 86970 61292
rect 87032 61240 87044 61292
rect 87106 61240 87108 61292
rect 86946 61238 86970 61240
rect 87026 61238 87050 61240
rect 87106 61238 87130 61240
rect 86890 61218 87186 61238
rect 86890 60206 87186 60226
rect 86946 60204 86970 60206
rect 87026 60204 87050 60206
rect 87106 60204 87130 60206
rect 86968 60152 86970 60204
rect 87032 60152 87044 60204
rect 87106 60152 87108 60204
rect 86946 60150 86970 60152
rect 87026 60150 87050 60152
rect 87106 60150 87130 60152
rect 86890 60130 87186 60150
rect 86890 59118 87186 59138
rect 86946 59116 86970 59118
rect 87026 59116 87050 59118
rect 87106 59116 87130 59118
rect 86968 59064 86970 59116
rect 87032 59064 87044 59116
rect 87106 59064 87108 59116
rect 86946 59062 86970 59064
rect 87026 59062 87050 59064
rect 87106 59062 87130 59064
rect 86890 59042 87186 59062
rect 86890 58030 87186 58050
rect 86946 58028 86970 58030
rect 87026 58028 87050 58030
rect 87106 58028 87130 58030
rect 86968 57976 86970 58028
rect 87032 57976 87044 58028
rect 87106 57976 87108 58028
rect 86946 57974 86970 57976
rect 87026 57974 87050 57976
rect 87106 57974 87130 57976
rect 86890 57954 87186 57974
rect 86890 56942 87186 56962
rect 86946 56940 86970 56942
rect 87026 56940 87050 56942
rect 87106 56940 87130 56942
rect 86968 56888 86970 56940
rect 87032 56888 87044 56940
rect 87106 56888 87108 56940
rect 86946 56886 86970 56888
rect 87026 56886 87050 56888
rect 87106 56886 87130 56888
rect 86890 56866 87186 56886
rect 86890 55854 87186 55874
rect 86946 55852 86970 55854
rect 87026 55852 87050 55854
rect 87106 55852 87130 55854
rect 86968 55800 86970 55852
rect 87032 55800 87044 55852
rect 87106 55800 87108 55852
rect 86946 55798 86970 55800
rect 87026 55798 87050 55800
rect 87106 55798 87130 55800
rect 86890 55778 87186 55798
rect 86890 54766 87186 54786
rect 86946 54764 86970 54766
rect 87026 54764 87050 54766
rect 87106 54764 87130 54766
rect 86968 54712 86970 54764
rect 87032 54712 87044 54764
rect 87106 54712 87108 54764
rect 86946 54710 86970 54712
rect 87026 54710 87050 54712
rect 87106 54710 87130 54712
rect 86890 54690 87186 54710
rect 86890 53678 87186 53698
rect 86946 53676 86970 53678
rect 87026 53676 87050 53678
rect 87106 53676 87130 53678
rect 86968 53624 86970 53676
rect 87032 53624 87044 53676
rect 87106 53624 87108 53676
rect 86946 53622 86970 53624
rect 87026 53622 87050 53624
rect 87106 53622 87130 53624
rect 86890 53602 87186 53622
rect 86890 52590 87186 52610
rect 86946 52588 86970 52590
rect 87026 52588 87050 52590
rect 87106 52588 87130 52590
rect 86968 52536 86970 52588
rect 87032 52536 87044 52588
rect 87106 52536 87108 52588
rect 86946 52534 86970 52536
rect 87026 52534 87050 52536
rect 87106 52534 87130 52536
rect 86890 52514 87186 52534
rect 86890 51502 87186 51522
rect 86946 51500 86970 51502
rect 87026 51500 87050 51502
rect 87106 51500 87130 51502
rect 86968 51448 86970 51500
rect 87032 51448 87044 51500
rect 87106 51448 87108 51500
rect 86946 51446 86970 51448
rect 87026 51446 87050 51448
rect 87106 51446 87130 51448
rect 86890 51426 87186 51446
rect 86890 50414 87186 50434
rect 86946 50412 86970 50414
rect 87026 50412 87050 50414
rect 87106 50412 87130 50414
rect 86968 50360 86970 50412
rect 87032 50360 87044 50412
rect 87106 50360 87108 50412
rect 86946 50358 86970 50360
rect 87026 50358 87050 50360
rect 87106 50358 87130 50360
rect 86890 50338 87186 50358
rect 86890 49326 87186 49346
rect 86946 49324 86970 49326
rect 87026 49324 87050 49326
rect 87106 49324 87130 49326
rect 86968 49272 86970 49324
rect 87032 49272 87044 49324
rect 87106 49272 87108 49324
rect 86946 49270 86970 49272
rect 87026 49270 87050 49272
rect 87106 49270 87130 49272
rect 86890 49250 87186 49270
rect 86890 48238 87186 48258
rect 86946 48236 86970 48238
rect 87026 48236 87050 48238
rect 87106 48236 87130 48238
rect 86968 48184 86970 48236
rect 87032 48184 87044 48236
rect 87106 48184 87108 48236
rect 86946 48182 86970 48184
rect 87026 48182 87050 48184
rect 87106 48182 87130 48184
rect 86890 48162 87186 48182
rect 86890 47150 87186 47170
rect 86946 47148 86970 47150
rect 87026 47148 87050 47150
rect 87106 47148 87130 47150
rect 86968 47096 86970 47148
rect 87032 47096 87044 47148
rect 87106 47096 87108 47148
rect 86946 47094 86970 47096
rect 87026 47094 87050 47096
rect 87106 47094 87130 47096
rect 86890 47074 87186 47094
rect 86890 46062 87186 46082
rect 86946 46060 86970 46062
rect 87026 46060 87050 46062
rect 87106 46060 87130 46062
rect 86968 46008 86970 46060
rect 87032 46008 87044 46060
rect 87106 46008 87108 46060
rect 86946 46006 86970 46008
rect 87026 46006 87050 46008
rect 87106 46006 87130 46008
rect 86890 45986 87186 46006
rect 86890 44974 87186 44994
rect 86946 44972 86970 44974
rect 87026 44972 87050 44974
rect 87106 44972 87130 44974
rect 86968 44920 86970 44972
rect 87032 44920 87044 44972
rect 87106 44920 87108 44972
rect 86946 44918 86970 44920
rect 87026 44918 87050 44920
rect 87106 44918 87130 44920
rect 86890 44898 87186 44918
rect 86890 43886 87186 43906
rect 86946 43884 86970 43886
rect 87026 43884 87050 43886
rect 87106 43884 87130 43886
rect 86968 43832 86970 43884
rect 87032 43832 87044 43884
rect 87106 43832 87108 43884
rect 86946 43830 86970 43832
rect 87026 43830 87050 43832
rect 87106 43830 87130 43832
rect 86890 43810 87186 43830
rect 86890 42798 87186 42818
rect 86946 42796 86970 42798
rect 87026 42796 87050 42798
rect 87106 42796 87130 42798
rect 86968 42744 86970 42796
rect 87032 42744 87044 42796
rect 87106 42744 87108 42796
rect 86946 42742 86970 42744
rect 87026 42742 87050 42744
rect 87106 42742 87130 42744
rect 86890 42722 87186 42742
rect 86890 41710 87186 41730
rect 86946 41708 86970 41710
rect 87026 41708 87050 41710
rect 87106 41708 87130 41710
rect 86968 41656 86970 41708
rect 87032 41656 87044 41708
rect 87106 41656 87108 41708
rect 86946 41654 86970 41656
rect 87026 41654 87050 41656
rect 87106 41654 87130 41656
rect 86890 41634 87186 41654
rect 86890 40622 87186 40642
rect 86946 40620 86970 40622
rect 87026 40620 87050 40622
rect 87106 40620 87130 40622
rect 86968 40568 86970 40620
rect 87032 40568 87044 40620
rect 87106 40568 87108 40620
rect 86946 40566 86970 40568
rect 87026 40566 87050 40568
rect 87106 40566 87130 40568
rect 86890 40546 87186 40566
rect 86890 39534 87186 39554
rect 86946 39532 86970 39534
rect 87026 39532 87050 39534
rect 87106 39532 87130 39534
rect 86968 39480 86970 39532
rect 87032 39480 87044 39532
rect 87106 39480 87108 39532
rect 86946 39478 86970 39480
rect 87026 39478 87050 39480
rect 87106 39478 87130 39480
rect 86890 39458 87186 39478
rect 86890 38446 87186 38466
rect 86946 38444 86970 38446
rect 87026 38444 87050 38446
rect 87106 38444 87130 38446
rect 86968 38392 86970 38444
rect 87032 38392 87044 38444
rect 87106 38392 87108 38444
rect 86946 38390 86970 38392
rect 87026 38390 87050 38392
rect 87106 38390 87130 38392
rect 86890 38370 87186 38390
rect 86890 37358 87186 37378
rect 86946 37356 86970 37358
rect 87026 37356 87050 37358
rect 87106 37356 87130 37358
rect 86968 37304 86970 37356
rect 87032 37304 87044 37356
rect 87106 37304 87108 37356
rect 86946 37302 86970 37304
rect 87026 37302 87050 37304
rect 87106 37302 87130 37304
rect 86890 37282 87186 37302
rect 86890 36270 87186 36290
rect 86946 36268 86970 36270
rect 87026 36268 87050 36270
rect 87106 36268 87130 36270
rect 86968 36216 86970 36268
rect 87032 36216 87044 36268
rect 87106 36216 87108 36268
rect 86946 36214 86970 36216
rect 87026 36214 87050 36216
rect 87106 36214 87130 36216
rect 86890 36194 87186 36214
rect 86890 35182 87186 35202
rect 86946 35180 86970 35182
rect 87026 35180 87050 35182
rect 87106 35180 87130 35182
rect 86968 35128 86970 35180
rect 87032 35128 87044 35180
rect 87106 35128 87108 35180
rect 86946 35126 86970 35128
rect 87026 35126 87050 35128
rect 87106 35126 87130 35128
rect 86890 35106 87186 35126
rect 86890 34094 87186 34114
rect 86946 34092 86970 34094
rect 87026 34092 87050 34094
rect 87106 34092 87130 34094
rect 86968 34040 86970 34092
rect 87032 34040 87044 34092
rect 87106 34040 87108 34092
rect 86946 34038 86970 34040
rect 87026 34038 87050 34040
rect 87106 34038 87130 34040
rect 86890 34018 87186 34038
rect 86890 33006 87186 33026
rect 86946 33004 86970 33006
rect 87026 33004 87050 33006
rect 87106 33004 87130 33006
rect 86968 32952 86970 33004
rect 87032 32952 87044 33004
rect 87106 32952 87108 33004
rect 86946 32950 86970 32952
rect 87026 32950 87050 32952
rect 87106 32950 87130 32952
rect 86890 32930 87186 32950
rect 86890 31918 87186 31938
rect 86946 31916 86970 31918
rect 87026 31916 87050 31918
rect 87106 31916 87130 31918
rect 86968 31864 86970 31916
rect 87032 31864 87044 31916
rect 87106 31864 87108 31916
rect 86946 31862 86970 31864
rect 87026 31862 87050 31864
rect 87106 31862 87130 31864
rect 86890 31842 87186 31862
rect 86890 30830 87186 30850
rect 86946 30828 86970 30830
rect 87026 30828 87050 30830
rect 87106 30828 87130 30830
rect 86968 30776 86970 30828
rect 87032 30776 87044 30828
rect 87106 30776 87108 30828
rect 86946 30774 86970 30776
rect 87026 30774 87050 30776
rect 87106 30774 87130 30776
rect 86890 30754 87186 30774
rect 86890 29742 87186 29762
rect 86946 29740 86970 29742
rect 87026 29740 87050 29742
rect 87106 29740 87130 29742
rect 86968 29688 86970 29740
rect 87032 29688 87044 29740
rect 87106 29688 87108 29740
rect 86946 29686 86970 29688
rect 87026 29686 87050 29688
rect 87106 29686 87130 29688
rect 86890 29666 87186 29686
rect 86890 28654 87186 28674
rect 86946 28652 86970 28654
rect 87026 28652 87050 28654
rect 87106 28652 87130 28654
rect 86968 28600 86970 28652
rect 87032 28600 87044 28652
rect 87106 28600 87108 28652
rect 86946 28598 86970 28600
rect 87026 28598 87050 28600
rect 87106 28598 87130 28600
rect 86890 28578 87186 28598
rect 86890 27566 87186 27586
rect 86946 27564 86970 27566
rect 87026 27564 87050 27566
rect 87106 27564 87130 27566
rect 86968 27512 86970 27564
rect 87032 27512 87044 27564
rect 87106 27512 87108 27564
rect 86946 27510 86970 27512
rect 87026 27510 87050 27512
rect 87106 27510 87130 27512
rect 86890 27490 87186 27510
rect 86890 26478 87186 26498
rect 86946 26476 86970 26478
rect 87026 26476 87050 26478
rect 87106 26476 87130 26478
rect 86968 26424 86970 26476
rect 87032 26424 87044 26476
rect 87106 26424 87108 26476
rect 86946 26422 86970 26424
rect 87026 26422 87050 26424
rect 87106 26422 87130 26424
rect 86890 26402 87186 26422
rect 86890 25390 87186 25410
rect 86946 25388 86970 25390
rect 87026 25388 87050 25390
rect 87106 25388 87130 25390
rect 86968 25336 86970 25388
rect 87032 25336 87044 25388
rect 87106 25336 87108 25388
rect 86946 25334 86970 25336
rect 87026 25334 87050 25336
rect 87106 25334 87130 25336
rect 86890 25314 87186 25334
rect 86890 24302 87186 24322
rect 86946 24300 86970 24302
rect 87026 24300 87050 24302
rect 87106 24300 87130 24302
rect 86968 24248 86970 24300
rect 87032 24248 87044 24300
rect 87106 24248 87108 24300
rect 86946 24246 86970 24248
rect 87026 24246 87050 24248
rect 87106 24246 87130 24248
rect 86890 24226 87186 24246
rect 86890 23214 87186 23234
rect 86946 23212 86970 23214
rect 87026 23212 87050 23214
rect 87106 23212 87130 23214
rect 86968 23160 86970 23212
rect 87032 23160 87044 23212
rect 87106 23160 87108 23212
rect 86946 23158 86970 23160
rect 87026 23158 87050 23160
rect 87106 23158 87130 23160
rect 86890 23138 87186 23158
rect 86890 22126 87186 22146
rect 86946 22124 86970 22126
rect 87026 22124 87050 22126
rect 87106 22124 87130 22126
rect 86968 22072 86970 22124
rect 87032 22072 87044 22124
rect 87106 22072 87108 22124
rect 86946 22070 86970 22072
rect 87026 22070 87050 22072
rect 87106 22070 87130 22072
rect 86890 22050 87186 22070
rect 86890 21038 87186 21058
rect 86946 21036 86970 21038
rect 87026 21036 87050 21038
rect 87106 21036 87130 21038
rect 86968 20984 86970 21036
rect 87032 20984 87044 21036
rect 87106 20984 87108 21036
rect 86946 20982 86970 20984
rect 87026 20982 87050 20984
rect 87106 20982 87130 20984
rect 86890 20962 87186 20982
rect 86890 19950 87186 19970
rect 86946 19948 86970 19950
rect 87026 19948 87050 19950
rect 87106 19948 87130 19950
rect 86968 19896 86970 19948
rect 87032 19896 87044 19948
rect 87106 19896 87108 19948
rect 86946 19894 86970 19896
rect 87026 19894 87050 19896
rect 87106 19894 87130 19896
rect 86890 19874 87186 19894
rect 86890 18862 87186 18882
rect 86946 18860 86970 18862
rect 87026 18860 87050 18862
rect 87106 18860 87130 18862
rect 86968 18808 86970 18860
rect 87032 18808 87044 18860
rect 87106 18808 87108 18860
rect 86946 18806 86970 18808
rect 87026 18806 87050 18808
rect 87106 18806 87130 18808
rect 86890 18786 87186 18806
rect 86890 17774 87186 17794
rect 86946 17772 86970 17774
rect 87026 17772 87050 17774
rect 87106 17772 87130 17774
rect 86968 17720 86970 17772
rect 87032 17720 87044 17772
rect 87106 17720 87108 17772
rect 86946 17718 86970 17720
rect 87026 17718 87050 17720
rect 87106 17718 87130 17720
rect 86890 17698 87186 17718
rect 86890 16686 87186 16706
rect 86946 16684 86970 16686
rect 87026 16684 87050 16686
rect 87106 16684 87130 16686
rect 86968 16632 86970 16684
rect 87032 16632 87044 16684
rect 87106 16632 87108 16684
rect 86946 16630 86970 16632
rect 87026 16630 87050 16632
rect 87106 16630 87130 16632
rect 86890 16610 87186 16630
rect 86890 15598 87186 15618
rect 86946 15596 86970 15598
rect 87026 15596 87050 15598
rect 87106 15596 87130 15598
rect 86968 15544 86970 15596
rect 87032 15544 87044 15596
rect 87106 15544 87108 15596
rect 86946 15542 86970 15544
rect 87026 15542 87050 15544
rect 87106 15542 87130 15544
rect 86890 15522 87186 15542
rect 86890 14510 87186 14530
rect 86946 14508 86970 14510
rect 87026 14508 87050 14510
rect 87106 14508 87130 14510
rect 86968 14456 86970 14508
rect 87032 14456 87044 14508
rect 87106 14456 87108 14508
rect 86946 14454 86970 14456
rect 87026 14454 87050 14456
rect 87106 14454 87130 14456
rect 86890 14434 87186 14454
rect 86890 13422 87186 13442
rect 86946 13420 86970 13422
rect 87026 13420 87050 13422
rect 87106 13420 87130 13422
rect 86968 13368 86970 13420
rect 87032 13368 87044 13420
rect 87106 13368 87108 13420
rect 86946 13366 86970 13368
rect 87026 13366 87050 13368
rect 87106 13366 87130 13368
rect 86890 13346 87186 13366
rect 86890 12334 87186 12354
rect 86946 12332 86970 12334
rect 87026 12332 87050 12334
rect 87106 12332 87130 12334
rect 86968 12280 86970 12332
rect 87032 12280 87044 12332
rect 87106 12280 87108 12332
rect 86946 12278 86970 12280
rect 87026 12278 87050 12280
rect 87106 12278 87130 12280
rect 86890 12258 87186 12278
rect 86890 11246 87186 11266
rect 86946 11244 86970 11246
rect 87026 11244 87050 11246
rect 87106 11244 87130 11246
rect 86968 11192 86970 11244
rect 87032 11192 87044 11244
rect 87106 11192 87108 11244
rect 86946 11190 86970 11192
rect 87026 11190 87050 11192
rect 87106 11190 87130 11192
rect 86890 11170 87186 11190
rect 86890 10158 87186 10178
rect 86946 10156 86970 10158
rect 87026 10156 87050 10158
rect 87106 10156 87130 10158
rect 86968 10104 86970 10156
rect 87032 10104 87044 10156
rect 87106 10104 87108 10156
rect 86946 10102 86970 10104
rect 87026 10102 87050 10104
rect 87106 10102 87130 10104
rect 86890 10082 87186 10102
rect 86890 9070 87186 9090
rect 86946 9068 86970 9070
rect 87026 9068 87050 9070
rect 87106 9068 87130 9070
rect 86968 9016 86970 9068
rect 87032 9016 87044 9068
rect 87106 9016 87108 9068
rect 86946 9014 86970 9016
rect 87026 9014 87050 9016
rect 87106 9014 87130 9016
rect 86890 8994 87186 9014
rect 86890 7982 87186 8002
rect 86946 7980 86970 7982
rect 87026 7980 87050 7982
rect 87106 7980 87130 7982
rect 86968 7928 86970 7980
rect 87032 7928 87044 7980
rect 87106 7928 87108 7980
rect 86946 7926 86970 7928
rect 87026 7926 87050 7928
rect 87106 7926 87130 7928
rect 86890 7906 87186 7926
rect 86890 6894 87186 6914
rect 86946 6892 86970 6894
rect 87026 6892 87050 6894
rect 87106 6892 87130 6894
rect 86968 6840 86970 6892
rect 87032 6840 87044 6892
rect 87106 6840 87108 6892
rect 86946 6838 86970 6840
rect 87026 6838 87050 6840
rect 87106 6838 87130 6840
rect 86890 6818 87186 6838
rect 86890 5806 87186 5826
rect 86946 5804 86970 5806
rect 87026 5804 87050 5806
rect 87106 5804 87130 5806
rect 86968 5752 86970 5804
rect 87032 5752 87044 5804
rect 87106 5752 87108 5804
rect 86946 5750 86970 5752
rect 87026 5750 87050 5752
rect 87106 5750 87130 5752
rect 86890 5730 87186 5750
rect 86890 4718 87186 4738
rect 86946 4716 86970 4718
rect 87026 4716 87050 4718
rect 87106 4716 87130 4718
rect 86968 4664 86970 4716
rect 87032 4664 87044 4716
rect 87106 4664 87108 4716
rect 86946 4662 86970 4664
rect 87026 4662 87050 4664
rect 87106 4662 87130 4664
rect 86890 4642 87186 4662
rect 86890 3630 87186 3650
rect 86946 3628 86970 3630
rect 87026 3628 87050 3630
rect 87106 3628 87130 3630
rect 86968 3576 86970 3628
rect 87032 3576 87044 3628
rect 87106 3576 87108 3628
rect 86946 3574 86970 3576
rect 87026 3574 87050 3576
rect 87106 3574 87130 3576
rect 86890 3554 87186 3574
rect 86630 2914 86682 2920
rect 86630 2856 86682 2862
rect 86538 2778 86590 2784
rect 86538 2720 86590 2726
rect 86890 2542 87186 2562
rect 86946 2540 86970 2542
rect 87026 2540 87050 2542
rect 87106 2540 87130 2542
rect 86968 2488 86970 2540
rect 87032 2488 87044 2540
rect 87106 2488 87108 2540
rect 86946 2486 86970 2488
rect 87026 2486 87050 2488
rect 87106 2486 87130 2488
rect 86890 2466 87186 2486
rect 8706 58 8758 64
rect 8706 0 8758 6
rect 85526 58 85578 64
rect 85526 0 85578 6
<< via2 >>
rect 84328 189146 84384 189202
rect 1252 187242 1308 187298
rect 890 186956 946 186958
rect 970 186956 1026 186958
rect 1050 186956 1106 186958
rect 1130 186956 1186 186958
rect 890 186904 916 186956
rect 916 186904 946 186956
rect 970 186904 980 186956
rect 980 186904 1026 186956
rect 1050 186904 1096 186956
rect 1096 186904 1106 186956
rect 1130 186904 1160 186956
rect 1160 186904 1186 186956
rect 890 186902 946 186904
rect 970 186902 1026 186904
rect 1050 186902 1106 186904
rect 1130 186902 1186 186904
rect 890 185868 946 185870
rect 970 185868 1026 185870
rect 1050 185868 1106 185870
rect 1130 185868 1186 185870
rect 890 185816 916 185868
rect 916 185816 946 185868
rect 970 185816 980 185868
rect 980 185816 1026 185868
rect 1050 185816 1096 185868
rect 1096 185816 1106 185868
rect 1130 185816 1160 185868
rect 1160 185816 1186 185868
rect 890 185814 946 185816
rect 970 185814 1026 185816
rect 1050 185814 1106 185816
rect 1130 185814 1186 185816
rect 890 184780 946 184782
rect 970 184780 1026 184782
rect 1050 184780 1106 184782
rect 1130 184780 1186 184782
rect 890 184728 916 184780
rect 916 184728 946 184780
rect 970 184728 980 184780
rect 980 184728 1026 184780
rect 1050 184728 1096 184780
rect 1096 184728 1106 184780
rect 1130 184728 1160 184780
rect 1160 184728 1186 184780
rect 890 184726 946 184728
rect 970 184726 1026 184728
rect 1050 184726 1106 184728
rect 1130 184726 1186 184728
rect 890 183692 946 183694
rect 970 183692 1026 183694
rect 1050 183692 1106 183694
rect 1130 183692 1186 183694
rect 890 183640 916 183692
rect 916 183640 946 183692
rect 970 183640 980 183692
rect 980 183640 1026 183692
rect 1050 183640 1096 183692
rect 1096 183640 1106 183692
rect 1130 183640 1160 183692
rect 1160 183640 1186 183692
rect 890 183638 946 183640
rect 970 183638 1026 183640
rect 1050 183638 1106 183640
rect 1130 183638 1186 183640
rect 890 182604 946 182606
rect 970 182604 1026 182606
rect 1050 182604 1106 182606
rect 1130 182604 1186 182606
rect 890 182552 916 182604
rect 916 182552 946 182604
rect 970 182552 980 182604
rect 980 182552 1026 182604
rect 1050 182552 1096 182604
rect 1096 182552 1106 182604
rect 1130 182552 1160 182604
rect 1160 182552 1186 182604
rect 890 182550 946 182552
rect 970 182550 1026 182552
rect 1050 182550 1106 182552
rect 1130 182550 1186 182552
rect 890 181516 946 181518
rect 970 181516 1026 181518
rect 1050 181516 1106 181518
rect 1130 181516 1186 181518
rect 890 181464 916 181516
rect 916 181464 946 181516
rect 970 181464 980 181516
rect 980 181464 1026 181516
rect 1050 181464 1096 181516
rect 1096 181464 1106 181516
rect 1130 181464 1160 181516
rect 1160 181464 1186 181516
rect 890 181462 946 181464
rect 970 181462 1026 181464
rect 1050 181462 1106 181464
rect 1130 181462 1186 181464
rect 890 180428 946 180430
rect 970 180428 1026 180430
rect 1050 180428 1106 180430
rect 1130 180428 1186 180430
rect 890 180376 916 180428
rect 916 180376 946 180428
rect 970 180376 980 180428
rect 980 180376 1026 180428
rect 1050 180376 1096 180428
rect 1096 180376 1106 180428
rect 1130 180376 1160 180428
rect 1160 180376 1186 180428
rect 890 180374 946 180376
rect 970 180374 1026 180376
rect 1050 180374 1106 180376
rect 1130 180374 1186 180376
rect 890 179340 946 179342
rect 970 179340 1026 179342
rect 1050 179340 1106 179342
rect 1130 179340 1186 179342
rect 890 179288 916 179340
rect 916 179288 946 179340
rect 970 179288 980 179340
rect 980 179288 1026 179340
rect 1050 179288 1096 179340
rect 1096 179288 1106 179340
rect 1130 179288 1160 179340
rect 1160 179288 1186 179340
rect 890 179286 946 179288
rect 970 179286 1026 179288
rect 1050 179286 1106 179288
rect 1130 179286 1186 179288
rect 890 178252 946 178254
rect 970 178252 1026 178254
rect 1050 178252 1106 178254
rect 1130 178252 1186 178254
rect 890 178200 916 178252
rect 916 178200 946 178252
rect 970 178200 980 178252
rect 980 178200 1026 178252
rect 1050 178200 1096 178252
rect 1096 178200 1106 178252
rect 1130 178200 1160 178252
rect 1160 178200 1186 178252
rect 890 178198 946 178200
rect 970 178198 1026 178200
rect 1050 178198 1106 178200
rect 1130 178198 1186 178200
rect 890 177164 946 177166
rect 970 177164 1026 177166
rect 1050 177164 1106 177166
rect 1130 177164 1186 177166
rect 890 177112 916 177164
rect 916 177112 946 177164
rect 970 177112 980 177164
rect 980 177112 1026 177164
rect 1050 177112 1096 177164
rect 1096 177112 1106 177164
rect 1130 177112 1160 177164
rect 1160 177112 1186 177164
rect 890 177110 946 177112
rect 970 177110 1026 177112
rect 1050 177110 1106 177112
rect 1130 177110 1186 177112
rect 890 176076 946 176078
rect 970 176076 1026 176078
rect 1050 176076 1106 176078
rect 1130 176076 1186 176078
rect 890 176024 916 176076
rect 916 176024 946 176076
rect 970 176024 980 176076
rect 980 176024 1026 176076
rect 1050 176024 1096 176076
rect 1096 176024 1106 176076
rect 1130 176024 1160 176076
rect 1160 176024 1186 176076
rect 890 176022 946 176024
rect 970 176022 1026 176024
rect 1050 176022 1106 176024
rect 1130 176022 1186 176024
rect 890 174988 946 174990
rect 970 174988 1026 174990
rect 1050 174988 1106 174990
rect 1130 174988 1186 174990
rect 890 174936 916 174988
rect 916 174936 946 174988
rect 970 174936 980 174988
rect 980 174936 1026 174988
rect 1050 174936 1096 174988
rect 1096 174936 1106 174988
rect 1130 174936 1160 174988
rect 1160 174936 1186 174988
rect 890 174934 946 174936
rect 970 174934 1026 174936
rect 1050 174934 1106 174936
rect 1130 174934 1186 174936
rect 890 173900 946 173902
rect 970 173900 1026 173902
rect 1050 173900 1106 173902
rect 1130 173900 1186 173902
rect 890 173848 916 173900
rect 916 173848 946 173900
rect 970 173848 980 173900
rect 980 173848 1026 173900
rect 1050 173848 1096 173900
rect 1096 173848 1106 173900
rect 1130 173848 1160 173900
rect 1160 173848 1186 173900
rect 890 173846 946 173848
rect 970 173846 1026 173848
rect 1050 173846 1106 173848
rect 1130 173846 1186 173848
rect 890 172812 946 172814
rect 970 172812 1026 172814
rect 1050 172812 1106 172814
rect 1130 172812 1186 172814
rect 890 172760 916 172812
rect 916 172760 946 172812
rect 970 172760 980 172812
rect 980 172760 1026 172812
rect 1050 172760 1096 172812
rect 1096 172760 1106 172812
rect 1130 172760 1160 172812
rect 1160 172760 1186 172812
rect 890 172758 946 172760
rect 970 172758 1026 172760
rect 1050 172758 1106 172760
rect 1130 172758 1186 172760
rect 890 171724 946 171726
rect 970 171724 1026 171726
rect 1050 171724 1106 171726
rect 1130 171724 1186 171726
rect 890 171672 916 171724
rect 916 171672 946 171724
rect 970 171672 980 171724
rect 980 171672 1026 171724
rect 1050 171672 1096 171724
rect 1096 171672 1106 171724
rect 1130 171672 1160 171724
rect 1160 171672 1186 171724
rect 890 171670 946 171672
rect 970 171670 1026 171672
rect 1050 171670 1106 171672
rect 1130 171670 1186 171672
rect 890 170636 946 170638
rect 970 170636 1026 170638
rect 1050 170636 1106 170638
rect 1130 170636 1186 170638
rect 890 170584 916 170636
rect 916 170584 946 170636
rect 970 170584 980 170636
rect 980 170584 1026 170636
rect 1050 170584 1096 170636
rect 1096 170584 1106 170636
rect 1130 170584 1160 170636
rect 1160 170584 1186 170636
rect 890 170582 946 170584
rect 970 170582 1026 170584
rect 1050 170582 1106 170584
rect 1130 170582 1186 170584
rect 890 169548 946 169550
rect 970 169548 1026 169550
rect 1050 169548 1106 169550
rect 1130 169548 1186 169550
rect 890 169496 916 169548
rect 916 169496 946 169548
rect 970 169496 980 169548
rect 980 169496 1026 169548
rect 1050 169496 1096 169548
rect 1096 169496 1106 169548
rect 1130 169496 1160 169548
rect 1160 169496 1186 169548
rect 890 169494 946 169496
rect 970 169494 1026 169496
rect 1050 169494 1106 169496
rect 1130 169494 1186 169496
rect 890 168460 946 168462
rect 970 168460 1026 168462
rect 1050 168460 1106 168462
rect 1130 168460 1186 168462
rect 890 168408 916 168460
rect 916 168408 946 168460
rect 970 168408 980 168460
rect 980 168408 1026 168460
rect 1050 168408 1096 168460
rect 1096 168408 1106 168460
rect 1130 168408 1160 168460
rect 1160 168408 1186 168460
rect 890 168406 946 168408
rect 970 168406 1026 168408
rect 1050 168406 1106 168408
rect 1130 168406 1186 168408
rect 890 167372 946 167374
rect 970 167372 1026 167374
rect 1050 167372 1106 167374
rect 1130 167372 1186 167374
rect 890 167320 916 167372
rect 916 167320 946 167372
rect 970 167320 980 167372
rect 980 167320 1026 167372
rect 1050 167320 1096 167372
rect 1096 167320 1106 167372
rect 1130 167320 1160 167372
rect 1160 167320 1186 167372
rect 890 167318 946 167320
rect 970 167318 1026 167320
rect 1050 167318 1106 167320
rect 1130 167318 1186 167320
rect 890 166284 946 166286
rect 970 166284 1026 166286
rect 1050 166284 1106 166286
rect 1130 166284 1186 166286
rect 890 166232 916 166284
rect 916 166232 946 166284
rect 970 166232 980 166284
rect 980 166232 1026 166284
rect 1050 166232 1096 166284
rect 1096 166232 1106 166284
rect 1130 166232 1160 166284
rect 1160 166232 1186 166284
rect 890 166230 946 166232
rect 970 166230 1026 166232
rect 1050 166230 1106 166232
rect 1130 166230 1186 166232
rect 890 165196 946 165198
rect 970 165196 1026 165198
rect 1050 165196 1106 165198
rect 1130 165196 1186 165198
rect 890 165144 916 165196
rect 916 165144 946 165196
rect 970 165144 980 165196
rect 980 165144 1026 165196
rect 1050 165144 1096 165196
rect 1096 165144 1106 165196
rect 1130 165144 1160 165196
rect 1160 165144 1186 165196
rect 890 165142 946 165144
rect 970 165142 1026 165144
rect 1050 165142 1106 165144
rect 1130 165142 1186 165144
rect 890 164108 946 164110
rect 970 164108 1026 164110
rect 1050 164108 1106 164110
rect 1130 164108 1186 164110
rect 890 164056 916 164108
rect 916 164056 946 164108
rect 970 164056 980 164108
rect 980 164056 1026 164108
rect 1050 164056 1096 164108
rect 1096 164056 1106 164108
rect 1130 164056 1160 164108
rect 1160 164056 1186 164108
rect 890 164054 946 164056
rect 970 164054 1026 164056
rect 1050 164054 1106 164056
rect 1130 164054 1186 164056
rect 890 163020 946 163022
rect 970 163020 1026 163022
rect 1050 163020 1106 163022
rect 1130 163020 1186 163022
rect 890 162968 916 163020
rect 916 162968 946 163020
rect 970 162968 980 163020
rect 980 162968 1026 163020
rect 1050 162968 1096 163020
rect 1096 162968 1106 163020
rect 1130 162968 1160 163020
rect 1160 162968 1186 163020
rect 890 162966 946 162968
rect 970 162966 1026 162968
rect 1050 162966 1106 162968
rect 1130 162966 1186 162968
rect 890 161932 946 161934
rect 970 161932 1026 161934
rect 1050 161932 1106 161934
rect 1130 161932 1186 161934
rect 890 161880 916 161932
rect 916 161880 946 161932
rect 970 161880 980 161932
rect 980 161880 1026 161932
rect 1050 161880 1096 161932
rect 1096 161880 1106 161932
rect 1130 161880 1160 161932
rect 1160 161880 1186 161932
rect 890 161878 946 161880
rect 970 161878 1026 161880
rect 1050 161878 1106 161880
rect 1130 161878 1186 161880
rect 890 160844 946 160846
rect 970 160844 1026 160846
rect 1050 160844 1106 160846
rect 1130 160844 1186 160846
rect 890 160792 916 160844
rect 916 160792 946 160844
rect 970 160792 980 160844
rect 980 160792 1026 160844
rect 1050 160792 1096 160844
rect 1096 160792 1106 160844
rect 1130 160792 1160 160844
rect 1160 160792 1186 160844
rect 890 160790 946 160792
rect 970 160790 1026 160792
rect 1050 160790 1106 160792
rect 1130 160790 1186 160792
rect 890 159756 946 159758
rect 970 159756 1026 159758
rect 1050 159756 1106 159758
rect 1130 159756 1186 159758
rect 890 159704 916 159756
rect 916 159704 946 159756
rect 970 159704 980 159756
rect 980 159704 1026 159756
rect 1050 159704 1096 159756
rect 1096 159704 1106 159756
rect 1130 159704 1160 159756
rect 1160 159704 1186 159756
rect 890 159702 946 159704
rect 970 159702 1026 159704
rect 1050 159702 1106 159704
rect 1130 159702 1186 159704
rect 890 158668 946 158670
rect 970 158668 1026 158670
rect 1050 158668 1106 158670
rect 1130 158668 1186 158670
rect 890 158616 916 158668
rect 916 158616 946 158668
rect 970 158616 980 158668
rect 980 158616 1026 158668
rect 1050 158616 1096 158668
rect 1096 158616 1106 158668
rect 1130 158616 1160 158668
rect 1160 158616 1186 158668
rect 890 158614 946 158616
rect 970 158614 1026 158616
rect 1050 158614 1106 158616
rect 1130 158614 1186 158616
rect 890 157580 946 157582
rect 970 157580 1026 157582
rect 1050 157580 1106 157582
rect 1130 157580 1186 157582
rect 890 157528 916 157580
rect 916 157528 946 157580
rect 970 157528 980 157580
rect 980 157528 1026 157580
rect 1050 157528 1096 157580
rect 1096 157528 1106 157580
rect 1130 157528 1160 157580
rect 1160 157528 1186 157580
rect 890 157526 946 157528
rect 970 157526 1026 157528
rect 1050 157526 1106 157528
rect 1130 157526 1186 157528
rect 890 156492 946 156494
rect 970 156492 1026 156494
rect 1050 156492 1106 156494
rect 1130 156492 1186 156494
rect 890 156440 916 156492
rect 916 156440 946 156492
rect 970 156440 980 156492
rect 980 156440 1026 156492
rect 1050 156440 1096 156492
rect 1096 156440 1106 156492
rect 1130 156440 1160 156492
rect 1160 156440 1186 156492
rect 890 156438 946 156440
rect 970 156438 1026 156440
rect 1050 156438 1106 156440
rect 1130 156438 1186 156440
rect 890 155404 946 155406
rect 970 155404 1026 155406
rect 1050 155404 1106 155406
rect 1130 155404 1186 155406
rect 890 155352 916 155404
rect 916 155352 946 155404
rect 970 155352 980 155404
rect 980 155352 1026 155404
rect 1050 155352 1096 155404
rect 1096 155352 1106 155404
rect 1130 155352 1160 155404
rect 1160 155352 1186 155404
rect 890 155350 946 155352
rect 970 155350 1026 155352
rect 1050 155350 1106 155352
rect 1130 155350 1186 155352
rect 890 154316 946 154318
rect 970 154316 1026 154318
rect 1050 154316 1106 154318
rect 1130 154316 1186 154318
rect 890 154264 916 154316
rect 916 154264 946 154316
rect 970 154264 980 154316
rect 980 154264 1026 154316
rect 1050 154264 1096 154316
rect 1096 154264 1106 154316
rect 1130 154264 1160 154316
rect 1160 154264 1186 154316
rect 890 154262 946 154264
rect 970 154262 1026 154264
rect 1050 154262 1106 154264
rect 1130 154262 1186 154264
rect 890 153228 946 153230
rect 970 153228 1026 153230
rect 1050 153228 1106 153230
rect 1130 153228 1186 153230
rect 890 153176 916 153228
rect 916 153176 946 153228
rect 970 153176 980 153228
rect 980 153176 1026 153228
rect 1050 153176 1096 153228
rect 1096 153176 1106 153228
rect 1130 153176 1160 153228
rect 1160 153176 1186 153228
rect 890 153174 946 153176
rect 970 153174 1026 153176
rect 1050 153174 1106 153176
rect 1130 153174 1186 153176
rect 890 152140 946 152142
rect 970 152140 1026 152142
rect 1050 152140 1106 152142
rect 1130 152140 1186 152142
rect 890 152088 916 152140
rect 916 152088 946 152140
rect 970 152088 980 152140
rect 980 152088 1026 152140
rect 1050 152088 1096 152140
rect 1096 152088 1106 152140
rect 1130 152088 1160 152140
rect 1160 152088 1186 152140
rect 890 152086 946 152088
rect 970 152086 1026 152088
rect 1050 152086 1106 152088
rect 1130 152086 1186 152088
rect 890 151052 946 151054
rect 970 151052 1026 151054
rect 1050 151052 1106 151054
rect 1130 151052 1186 151054
rect 890 151000 916 151052
rect 916 151000 946 151052
rect 970 151000 980 151052
rect 980 151000 1026 151052
rect 1050 151000 1096 151052
rect 1096 151000 1106 151052
rect 1130 151000 1160 151052
rect 1160 151000 1186 151052
rect 890 150998 946 151000
rect 970 150998 1026 151000
rect 1050 150998 1106 151000
rect 1130 150998 1186 151000
rect 890 149964 946 149966
rect 970 149964 1026 149966
rect 1050 149964 1106 149966
rect 1130 149964 1186 149966
rect 890 149912 916 149964
rect 916 149912 946 149964
rect 970 149912 980 149964
rect 980 149912 1026 149964
rect 1050 149912 1096 149964
rect 1096 149912 1106 149964
rect 1130 149912 1160 149964
rect 1160 149912 1186 149964
rect 890 149910 946 149912
rect 970 149910 1026 149912
rect 1050 149910 1106 149912
rect 1130 149910 1186 149912
rect 890 148876 946 148878
rect 970 148876 1026 148878
rect 1050 148876 1106 148878
rect 1130 148876 1186 148878
rect 890 148824 916 148876
rect 916 148824 946 148876
rect 970 148824 980 148876
rect 980 148824 1026 148876
rect 1050 148824 1096 148876
rect 1096 148824 1106 148876
rect 1130 148824 1160 148876
rect 1160 148824 1186 148876
rect 890 148822 946 148824
rect 970 148822 1026 148824
rect 1050 148822 1106 148824
rect 1130 148822 1186 148824
rect 890 147788 946 147790
rect 970 147788 1026 147790
rect 1050 147788 1106 147790
rect 1130 147788 1186 147790
rect 890 147736 916 147788
rect 916 147736 946 147788
rect 970 147736 980 147788
rect 980 147736 1026 147788
rect 1050 147736 1096 147788
rect 1096 147736 1106 147788
rect 1130 147736 1160 147788
rect 1160 147736 1186 147788
rect 890 147734 946 147736
rect 970 147734 1026 147736
rect 1050 147734 1106 147736
rect 1130 147734 1186 147736
rect 890 146700 946 146702
rect 970 146700 1026 146702
rect 1050 146700 1106 146702
rect 1130 146700 1186 146702
rect 890 146648 916 146700
rect 916 146648 946 146700
rect 970 146648 980 146700
rect 980 146648 1026 146700
rect 1050 146648 1096 146700
rect 1096 146648 1106 146700
rect 1130 146648 1160 146700
rect 1160 146648 1186 146700
rect 890 146646 946 146648
rect 970 146646 1026 146648
rect 1050 146646 1106 146648
rect 1130 146646 1186 146648
rect 890 145612 946 145614
rect 970 145612 1026 145614
rect 1050 145612 1106 145614
rect 1130 145612 1186 145614
rect 890 145560 916 145612
rect 916 145560 946 145612
rect 970 145560 980 145612
rect 980 145560 1026 145612
rect 1050 145560 1096 145612
rect 1096 145560 1106 145612
rect 1130 145560 1160 145612
rect 1160 145560 1186 145612
rect 890 145558 946 145560
rect 970 145558 1026 145560
rect 1050 145558 1106 145560
rect 1130 145558 1186 145560
rect 890 144524 946 144526
rect 970 144524 1026 144526
rect 1050 144524 1106 144526
rect 1130 144524 1186 144526
rect 890 144472 916 144524
rect 916 144472 946 144524
rect 970 144472 980 144524
rect 980 144472 1026 144524
rect 1050 144472 1096 144524
rect 1096 144472 1106 144524
rect 1130 144472 1160 144524
rect 1160 144472 1186 144524
rect 890 144470 946 144472
rect 970 144470 1026 144472
rect 1050 144470 1106 144472
rect 1130 144470 1186 144472
rect 890 143436 946 143438
rect 970 143436 1026 143438
rect 1050 143436 1106 143438
rect 1130 143436 1186 143438
rect 890 143384 916 143436
rect 916 143384 946 143436
rect 970 143384 980 143436
rect 980 143384 1026 143436
rect 1050 143384 1096 143436
rect 1096 143384 1106 143436
rect 1130 143384 1160 143436
rect 1160 143384 1186 143436
rect 890 143382 946 143384
rect 970 143382 1026 143384
rect 1050 143382 1106 143384
rect 1130 143382 1186 143384
rect 890 142348 946 142350
rect 970 142348 1026 142350
rect 1050 142348 1106 142350
rect 1130 142348 1186 142350
rect 890 142296 916 142348
rect 916 142296 946 142348
rect 970 142296 980 142348
rect 980 142296 1026 142348
rect 1050 142296 1096 142348
rect 1096 142296 1106 142348
rect 1130 142296 1160 142348
rect 1160 142296 1186 142348
rect 890 142294 946 142296
rect 970 142294 1026 142296
rect 1050 142294 1106 142296
rect 1130 142294 1186 142296
rect 890 141260 946 141262
rect 970 141260 1026 141262
rect 1050 141260 1106 141262
rect 1130 141260 1186 141262
rect 890 141208 916 141260
rect 916 141208 946 141260
rect 970 141208 980 141260
rect 980 141208 1026 141260
rect 1050 141208 1096 141260
rect 1096 141208 1106 141260
rect 1130 141208 1160 141260
rect 1160 141208 1186 141260
rect 890 141206 946 141208
rect 970 141206 1026 141208
rect 1050 141206 1106 141208
rect 1130 141206 1186 141208
rect 890 140172 946 140174
rect 970 140172 1026 140174
rect 1050 140172 1106 140174
rect 1130 140172 1186 140174
rect 890 140120 916 140172
rect 916 140120 946 140172
rect 970 140120 980 140172
rect 980 140120 1026 140172
rect 1050 140120 1096 140172
rect 1096 140120 1106 140172
rect 1130 140120 1160 140172
rect 1160 140120 1186 140172
rect 890 140118 946 140120
rect 970 140118 1026 140120
rect 1050 140118 1106 140120
rect 1130 140118 1186 140120
rect 890 139084 946 139086
rect 970 139084 1026 139086
rect 1050 139084 1106 139086
rect 1130 139084 1186 139086
rect 890 139032 916 139084
rect 916 139032 946 139084
rect 970 139032 980 139084
rect 980 139032 1026 139084
rect 1050 139032 1096 139084
rect 1096 139032 1106 139084
rect 1130 139032 1160 139084
rect 1160 139032 1186 139084
rect 890 139030 946 139032
rect 970 139030 1026 139032
rect 1050 139030 1106 139032
rect 1130 139030 1186 139032
rect 890 137996 946 137998
rect 970 137996 1026 137998
rect 1050 137996 1106 137998
rect 1130 137996 1186 137998
rect 890 137944 916 137996
rect 916 137944 946 137996
rect 970 137944 980 137996
rect 980 137944 1026 137996
rect 1050 137944 1096 137996
rect 1096 137944 1106 137996
rect 1130 137944 1160 137996
rect 1160 137944 1186 137996
rect 890 137942 946 137944
rect 970 137942 1026 137944
rect 1050 137942 1106 137944
rect 1130 137942 1186 137944
rect 890 136908 946 136910
rect 970 136908 1026 136910
rect 1050 136908 1106 136910
rect 1130 136908 1186 136910
rect 890 136856 916 136908
rect 916 136856 946 136908
rect 970 136856 980 136908
rect 980 136856 1026 136908
rect 1050 136856 1096 136908
rect 1096 136856 1106 136908
rect 1130 136856 1160 136908
rect 1160 136856 1186 136908
rect 890 136854 946 136856
rect 970 136854 1026 136856
rect 1050 136854 1106 136856
rect 1130 136854 1186 136856
rect 890 135820 946 135822
rect 970 135820 1026 135822
rect 1050 135820 1106 135822
rect 1130 135820 1186 135822
rect 890 135768 916 135820
rect 916 135768 946 135820
rect 970 135768 980 135820
rect 980 135768 1026 135820
rect 1050 135768 1096 135820
rect 1096 135768 1106 135820
rect 1130 135768 1160 135820
rect 1160 135768 1186 135820
rect 890 135766 946 135768
rect 970 135766 1026 135768
rect 1050 135766 1106 135768
rect 1130 135766 1186 135768
rect 890 134732 946 134734
rect 970 134732 1026 134734
rect 1050 134732 1106 134734
rect 1130 134732 1186 134734
rect 890 134680 916 134732
rect 916 134680 946 134732
rect 970 134680 980 134732
rect 980 134680 1026 134732
rect 1050 134680 1096 134732
rect 1096 134680 1106 134732
rect 1130 134680 1160 134732
rect 1160 134680 1186 134732
rect 890 134678 946 134680
rect 970 134678 1026 134680
rect 1050 134678 1106 134680
rect 1130 134678 1186 134680
rect 890 133644 946 133646
rect 970 133644 1026 133646
rect 1050 133644 1106 133646
rect 1130 133644 1186 133646
rect 890 133592 916 133644
rect 916 133592 946 133644
rect 970 133592 980 133644
rect 980 133592 1026 133644
rect 1050 133592 1096 133644
rect 1096 133592 1106 133644
rect 1130 133592 1160 133644
rect 1160 133592 1186 133644
rect 890 133590 946 133592
rect 970 133590 1026 133592
rect 1050 133590 1106 133592
rect 1130 133590 1186 133592
rect 890 132556 946 132558
rect 970 132556 1026 132558
rect 1050 132556 1106 132558
rect 1130 132556 1186 132558
rect 890 132504 916 132556
rect 916 132504 946 132556
rect 970 132504 980 132556
rect 980 132504 1026 132556
rect 1050 132504 1096 132556
rect 1096 132504 1106 132556
rect 1130 132504 1160 132556
rect 1160 132504 1186 132556
rect 890 132502 946 132504
rect 970 132502 1026 132504
rect 1050 132502 1106 132504
rect 1130 132502 1186 132504
rect 890 131468 946 131470
rect 970 131468 1026 131470
rect 1050 131468 1106 131470
rect 1130 131468 1186 131470
rect 890 131416 916 131468
rect 916 131416 946 131468
rect 970 131416 980 131468
rect 980 131416 1026 131468
rect 1050 131416 1096 131468
rect 1096 131416 1106 131468
rect 1130 131416 1160 131468
rect 1160 131416 1186 131468
rect 890 131414 946 131416
rect 970 131414 1026 131416
rect 1050 131414 1106 131416
rect 1130 131414 1186 131416
rect 890 130380 946 130382
rect 970 130380 1026 130382
rect 1050 130380 1106 130382
rect 1130 130380 1186 130382
rect 890 130328 916 130380
rect 916 130328 946 130380
rect 970 130328 980 130380
rect 980 130328 1026 130380
rect 1050 130328 1096 130380
rect 1096 130328 1106 130380
rect 1130 130328 1160 130380
rect 1160 130328 1186 130380
rect 890 130326 946 130328
rect 970 130326 1026 130328
rect 1050 130326 1106 130328
rect 1130 130326 1186 130328
rect 890 129292 946 129294
rect 970 129292 1026 129294
rect 1050 129292 1106 129294
rect 1130 129292 1186 129294
rect 890 129240 916 129292
rect 916 129240 946 129292
rect 970 129240 980 129292
rect 980 129240 1026 129292
rect 1050 129240 1096 129292
rect 1096 129240 1106 129292
rect 1130 129240 1160 129292
rect 1160 129240 1186 129292
rect 890 129238 946 129240
rect 970 129238 1026 129240
rect 1050 129238 1106 129240
rect 1130 129238 1186 129240
rect 890 128204 946 128206
rect 970 128204 1026 128206
rect 1050 128204 1106 128206
rect 1130 128204 1186 128206
rect 890 128152 916 128204
rect 916 128152 946 128204
rect 970 128152 980 128204
rect 980 128152 1026 128204
rect 1050 128152 1096 128204
rect 1096 128152 1106 128204
rect 1130 128152 1160 128204
rect 1160 128152 1186 128204
rect 890 128150 946 128152
rect 970 128150 1026 128152
rect 1050 128150 1106 128152
rect 1130 128150 1186 128152
rect 890 127116 946 127118
rect 970 127116 1026 127118
rect 1050 127116 1106 127118
rect 1130 127116 1186 127118
rect 890 127064 916 127116
rect 916 127064 946 127116
rect 970 127064 980 127116
rect 980 127064 1026 127116
rect 1050 127064 1096 127116
rect 1096 127064 1106 127116
rect 1130 127064 1160 127116
rect 1160 127064 1186 127116
rect 890 127062 946 127064
rect 970 127062 1026 127064
rect 1050 127062 1106 127064
rect 1130 127062 1186 127064
rect 890 126028 946 126030
rect 970 126028 1026 126030
rect 1050 126028 1106 126030
rect 1130 126028 1186 126030
rect 890 125976 916 126028
rect 916 125976 946 126028
rect 970 125976 980 126028
rect 980 125976 1026 126028
rect 1050 125976 1096 126028
rect 1096 125976 1106 126028
rect 1130 125976 1160 126028
rect 1160 125976 1186 126028
rect 890 125974 946 125976
rect 970 125974 1026 125976
rect 1050 125974 1106 125976
rect 1130 125974 1186 125976
rect 890 124940 946 124942
rect 970 124940 1026 124942
rect 1050 124940 1106 124942
rect 1130 124940 1186 124942
rect 890 124888 916 124940
rect 916 124888 946 124940
rect 970 124888 980 124940
rect 980 124888 1026 124940
rect 1050 124888 1096 124940
rect 1096 124888 1106 124940
rect 1130 124888 1160 124940
rect 1160 124888 1186 124940
rect 890 124886 946 124888
rect 970 124886 1026 124888
rect 1050 124886 1106 124888
rect 1130 124886 1186 124888
rect 890 123852 946 123854
rect 970 123852 1026 123854
rect 1050 123852 1106 123854
rect 1130 123852 1186 123854
rect 890 123800 916 123852
rect 916 123800 946 123852
rect 970 123800 980 123852
rect 980 123800 1026 123852
rect 1050 123800 1096 123852
rect 1096 123800 1106 123852
rect 1130 123800 1160 123852
rect 1160 123800 1186 123852
rect 890 123798 946 123800
rect 970 123798 1026 123800
rect 1050 123798 1106 123800
rect 1130 123798 1186 123800
rect 890 122764 946 122766
rect 970 122764 1026 122766
rect 1050 122764 1106 122766
rect 1130 122764 1186 122766
rect 890 122712 916 122764
rect 916 122712 946 122764
rect 970 122712 980 122764
rect 980 122712 1026 122764
rect 1050 122712 1096 122764
rect 1096 122712 1106 122764
rect 1130 122712 1160 122764
rect 1160 122712 1186 122764
rect 890 122710 946 122712
rect 970 122710 1026 122712
rect 1050 122710 1106 122712
rect 1130 122710 1186 122712
rect 890 121676 946 121678
rect 970 121676 1026 121678
rect 1050 121676 1106 121678
rect 1130 121676 1186 121678
rect 890 121624 916 121676
rect 916 121624 946 121676
rect 970 121624 980 121676
rect 980 121624 1026 121676
rect 1050 121624 1096 121676
rect 1096 121624 1106 121676
rect 1130 121624 1160 121676
rect 1160 121624 1186 121676
rect 890 121622 946 121624
rect 970 121622 1026 121624
rect 1050 121622 1106 121624
rect 1130 121622 1186 121624
rect 890 120588 946 120590
rect 970 120588 1026 120590
rect 1050 120588 1106 120590
rect 1130 120588 1186 120590
rect 890 120536 916 120588
rect 916 120536 946 120588
rect 970 120536 980 120588
rect 980 120536 1026 120588
rect 1050 120536 1096 120588
rect 1096 120536 1106 120588
rect 1130 120536 1160 120588
rect 1160 120536 1186 120588
rect 890 120534 946 120536
rect 970 120534 1026 120536
rect 1050 120534 1106 120536
rect 1130 120534 1186 120536
rect 890 119500 946 119502
rect 970 119500 1026 119502
rect 1050 119500 1106 119502
rect 1130 119500 1186 119502
rect 890 119448 916 119500
rect 916 119448 946 119500
rect 970 119448 980 119500
rect 980 119448 1026 119500
rect 1050 119448 1096 119500
rect 1096 119448 1106 119500
rect 1130 119448 1160 119500
rect 1160 119448 1186 119500
rect 890 119446 946 119448
rect 970 119446 1026 119448
rect 1050 119446 1106 119448
rect 1130 119446 1186 119448
rect 890 118412 946 118414
rect 970 118412 1026 118414
rect 1050 118412 1106 118414
rect 1130 118412 1186 118414
rect 890 118360 916 118412
rect 916 118360 946 118412
rect 970 118360 980 118412
rect 980 118360 1026 118412
rect 1050 118360 1096 118412
rect 1096 118360 1106 118412
rect 1130 118360 1160 118412
rect 1160 118360 1186 118412
rect 890 118358 946 118360
rect 970 118358 1026 118360
rect 1050 118358 1106 118360
rect 1130 118358 1186 118360
rect 890 117324 946 117326
rect 970 117324 1026 117326
rect 1050 117324 1106 117326
rect 1130 117324 1186 117326
rect 890 117272 916 117324
rect 916 117272 946 117324
rect 970 117272 980 117324
rect 980 117272 1026 117324
rect 1050 117272 1096 117324
rect 1096 117272 1106 117324
rect 1130 117272 1160 117324
rect 1160 117272 1186 117324
rect 890 117270 946 117272
rect 970 117270 1026 117272
rect 1050 117270 1106 117272
rect 1130 117270 1186 117272
rect 890 116236 946 116238
rect 970 116236 1026 116238
rect 1050 116236 1106 116238
rect 1130 116236 1186 116238
rect 890 116184 916 116236
rect 916 116184 946 116236
rect 970 116184 980 116236
rect 980 116184 1026 116236
rect 1050 116184 1096 116236
rect 1096 116184 1106 116236
rect 1130 116184 1160 116236
rect 1160 116184 1186 116236
rect 890 116182 946 116184
rect 970 116182 1026 116184
rect 1050 116182 1106 116184
rect 1130 116182 1186 116184
rect 890 115148 946 115150
rect 970 115148 1026 115150
rect 1050 115148 1106 115150
rect 1130 115148 1186 115150
rect 890 115096 916 115148
rect 916 115096 946 115148
rect 970 115096 980 115148
rect 980 115096 1026 115148
rect 1050 115096 1096 115148
rect 1096 115096 1106 115148
rect 1130 115096 1160 115148
rect 1160 115096 1186 115148
rect 890 115094 946 115096
rect 970 115094 1026 115096
rect 1050 115094 1106 115096
rect 1130 115094 1186 115096
rect 890 114060 946 114062
rect 970 114060 1026 114062
rect 1050 114060 1106 114062
rect 1130 114060 1186 114062
rect 890 114008 916 114060
rect 916 114008 946 114060
rect 970 114008 980 114060
rect 980 114008 1026 114060
rect 1050 114008 1096 114060
rect 1096 114008 1106 114060
rect 1130 114008 1160 114060
rect 1160 114008 1186 114060
rect 890 114006 946 114008
rect 970 114006 1026 114008
rect 1050 114006 1106 114008
rect 1130 114006 1186 114008
rect 890 112972 946 112974
rect 970 112972 1026 112974
rect 1050 112972 1106 112974
rect 1130 112972 1186 112974
rect 890 112920 916 112972
rect 916 112920 946 112972
rect 970 112920 980 112972
rect 980 112920 1026 112972
rect 1050 112920 1096 112972
rect 1096 112920 1106 112972
rect 1130 112920 1160 112972
rect 1160 112920 1186 112972
rect 890 112918 946 112920
rect 970 112918 1026 112920
rect 1050 112918 1106 112920
rect 1130 112918 1186 112920
rect 890 111884 946 111886
rect 970 111884 1026 111886
rect 1050 111884 1106 111886
rect 1130 111884 1186 111886
rect 890 111832 916 111884
rect 916 111832 946 111884
rect 970 111832 980 111884
rect 980 111832 1026 111884
rect 1050 111832 1096 111884
rect 1096 111832 1106 111884
rect 1130 111832 1160 111884
rect 1160 111832 1186 111884
rect 890 111830 946 111832
rect 970 111830 1026 111832
rect 1050 111830 1106 111832
rect 1130 111830 1186 111832
rect 890 110796 946 110798
rect 970 110796 1026 110798
rect 1050 110796 1106 110798
rect 1130 110796 1186 110798
rect 890 110744 916 110796
rect 916 110744 946 110796
rect 970 110744 980 110796
rect 980 110744 1026 110796
rect 1050 110744 1096 110796
rect 1096 110744 1106 110796
rect 1130 110744 1160 110796
rect 1160 110744 1186 110796
rect 890 110742 946 110744
rect 970 110742 1026 110744
rect 1050 110742 1106 110744
rect 1130 110742 1186 110744
rect 890 109708 946 109710
rect 970 109708 1026 109710
rect 1050 109708 1106 109710
rect 1130 109708 1186 109710
rect 890 109656 916 109708
rect 916 109656 946 109708
rect 970 109656 980 109708
rect 980 109656 1026 109708
rect 1050 109656 1096 109708
rect 1096 109656 1106 109708
rect 1130 109656 1160 109708
rect 1160 109656 1186 109708
rect 890 109654 946 109656
rect 970 109654 1026 109656
rect 1050 109654 1106 109656
rect 1130 109654 1186 109656
rect 890 108620 946 108622
rect 970 108620 1026 108622
rect 1050 108620 1106 108622
rect 1130 108620 1186 108622
rect 890 108568 916 108620
rect 916 108568 946 108620
rect 970 108568 980 108620
rect 980 108568 1026 108620
rect 1050 108568 1096 108620
rect 1096 108568 1106 108620
rect 1130 108568 1160 108620
rect 1160 108568 1186 108620
rect 890 108566 946 108568
rect 970 108566 1026 108568
rect 1050 108566 1106 108568
rect 1130 108566 1186 108568
rect 890 107532 946 107534
rect 970 107532 1026 107534
rect 1050 107532 1106 107534
rect 1130 107532 1186 107534
rect 890 107480 916 107532
rect 916 107480 946 107532
rect 970 107480 980 107532
rect 980 107480 1026 107532
rect 1050 107480 1096 107532
rect 1096 107480 1106 107532
rect 1130 107480 1160 107532
rect 1160 107480 1186 107532
rect 890 107478 946 107480
rect 970 107478 1026 107480
rect 1050 107478 1106 107480
rect 1130 107478 1186 107480
rect 890 106444 946 106446
rect 970 106444 1026 106446
rect 1050 106444 1106 106446
rect 1130 106444 1186 106446
rect 890 106392 916 106444
rect 916 106392 946 106444
rect 970 106392 980 106444
rect 980 106392 1026 106444
rect 1050 106392 1096 106444
rect 1096 106392 1106 106444
rect 1130 106392 1160 106444
rect 1160 106392 1186 106444
rect 890 106390 946 106392
rect 970 106390 1026 106392
rect 1050 106390 1106 106392
rect 1130 106390 1186 106392
rect 890 105356 946 105358
rect 970 105356 1026 105358
rect 1050 105356 1106 105358
rect 1130 105356 1186 105358
rect 890 105304 916 105356
rect 916 105304 946 105356
rect 970 105304 980 105356
rect 980 105304 1026 105356
rect 1050 105304 1096 105356
rect 1096 105304 1106 105356
rect 1130 105304 1160 105356
rect 1160 105304 1186 105356
rect 890 105302 946 105304
rect 970 105302 1026 105304
rect 1050 105302 1106 105304
rect 1130 105302 1186 105304
rect 890 104268 946 104270
rect 970 104268 1026 104270
rect 1050 104268 1106 104270
rect 1130 104268 1186 104270
rect 890 104216 916 104268
rect 916 104216 946 104268
rect 970 104216 980 104268
rect 980 104216 1026 104268
rect 1050 104216 1096 104268
rect 1096 104216 1106 104268
rect 1130 104216 1160 104268
rect 1160 104216 1186 104268
rect 890 104214 946 104216
rect 970 104214 1026 104216
rect 1050 104214 1106 104216
rect 1130 104214 1186 104216
rect 890 103180 946 103182
rect 970 103180 1026 103182
rect 1050 103180 1106 103182
rect 1130 103180 1186 103182
rect 890 103128 916 103180
rect 916 103128 946 103180
rect 970 103128 980 103180
rect 980 103128 1026 103180
rect 1050 103128 1096 103180
rect 1096 103128 1106 103180
rect 1130 103128 1160 103180
rect 1160 103128 1186 103180
rect 890 103126 946 103128
rect 970 103126 1026 103128
rect 1050 103126 1106 103128
rect 1130 103126 1186 103128
rect 890 102092 946 102094
rect 970 102092 1026 102094
rect 1050 102092 1106 102094
rect 1130 102092 1186 102094
rect 890 102040 916 102092
rect 916 102040 946 102092
rect 970 102040 980 102092
rect 980 102040 1026 102092
rect 1050 102040 1096 102092
rect 1096 102040 1106 102092
rect 1130 102040 1160 102092
rect 1160 102040 1186 102092
rect 890 102038 946 102040
rect 970 102038 1026 102040
rect 1050 102038 1106 102040
rect 1130 102038 1186 102040
rect 890 101004 946 101006
rect 970 101004 1026 101006
rect 1050 101004 1106 101006
rect 1130 101004 1186 101006
rect 890 100952 916 101004
rect 916 100952 946 101004
rect 970 100952 980 101004
rect 980 100952 1026 101004
rect 1050 100952 1096 101004
rect 1096 100952 1106 101004
rect 1130 100952 1160 101004
rect 1160 100952 1186 101004
rect 890 100950 946 100952
rect 970 100950 1026 100952
rect 1050 100950 1106 100952
rect 1130 100950 1186 100952
rect 890 99916 946 99918
rect 970 99916 1026 99918
rect 1050 99916 1106 99918
rect 1130 99916 1186 99918
rect 890 99864 916 99916
rect 916 99864 946 99916
rect 970 99864 980 99916
rect 980 99864 1026 99916
rect 1050 99864 1096 99916
rect 1096 99864 1106 99916
rect 1130 99864 1160 99916
rect 1160 99864 1186 99916
rect 890 99862 946 99864
rect 970 99862 1026 99864
rect 1050 99862 1106 99864
rect 1130 99862 1186 99864
rect 890 98828 946 98830
rect 970 98828 1026 98830
rect 1050 98828 1106 98830
rect 1130 98828 1186 98830
rect 890 98776 916 98828
rect 916 98776 946 98828
rect 970 98776 980 98828
rect 980 98776 1026 98828
rect 1050 98776 1096 98828
rect 1096 98776 1106 98828
rect 1130 98776 1160 98828
rect 1160 98776 1186 98828
rect 890 98774 946 98776
rect 970 98774 1026 98776
rect 1050 98774 1106 98776
rect 1130 98774 1186 98776
rect 890 97740 946 97742
rect 970 97740 1026 97742
rect 1050 97740 1106 97742
rect 1130 97740 1186 97742
rect 890 97688 916 97740
rect 916 97688 946 97740
rect 970 97688 980 97740
rect 980 97688 1026 97740
rect 1050 97688 1096 97740
rect 1096 97688 1106 97740
rect 1130 97688 1160 97740
rect 1160 97688 1186 97740
rect 890 97686 946 97688
rect 970 97686 1026 97688
rect 1050 97686 1106 97688
rect 1130 97686 1186 97688
rect 890 96652 946 96654
rect 970 96652 1026 96654
rect 1050 96652 1106 96654
rect 1130 96652 1186 96654
rect 890 96600 916 96652
rect 916 96600 946 96652
rect 970 96600 980 96652
rect 980 96600 1026 96652
rect 1050 96600 1096 96652
rect 1096 96600 1106 96652
rect 1130 96600 1160 96652
rect 1160 96600 1186 96652
rect 890 96598 946 96600
rect 970 96598 1026 96600
rect 1050 96598 1106 96600
rect 1130 96598 1186 96600
rect 890 95564 946 95566
rect 970 95564 1026 95566
rect 1050 95564 1106 95566
rect 1130 95564 1186 95566
rect 890 95512 916 95564
rect 916 95512 946 95564
rect 970 95512 980 95564
rect 980 95512 1026 95564
rect 1050 95512 1096 95564
rect 1096 95512 1106 95564
rect 1130 95512 1160 95564
rect 1160 95512 1186 95564
rect 890 95510 946 95512
rect 970 95510 1026 95512
rect 1050 95510 1106 95512
rect 1130 95510 1186 95512
rect 890 94476 946 94478
rect 970 94476 1026 94478
rect 1050 94476 1106 94478
rect 1130 94476 1186 94478
rect 890 94424 916 94476
rect 916 94424 946 94476
rect 970 94424 980 94476
rect 980 94424 1026 94476
rect 1050 94424 1096 94476
rect 1096 94424 1106 94476
rect 1130 94424 1160 94476
rect 1160 94424 1186 94476
rect 890 94422 946 94424
rect 970 94422 1026 94424
rect 1050 94422 1106 94424
rect 1130 94422 1186 94424
rect 890 93388 946 93390
rect 970 93388 1026 93390
rect 1050 93388 1106 93390
rect 1130 93388 1186 93390
rect 890 93336 916 93388
rect 916 93336 946 93388
rect 970 93336 980 93388
rect 980 93336 1026 93388
rect 1050 93336 1096 93388
rect 1096 93336 1106 93388
rect 1130 93336 1160 93388
rect 1160 93336 1186 93388
rect 890 93334 946 93336
rect 970 93334 1026 93336
rect 1050 93334 1106 93336
rect 1130 93334 1186 93336
rect 890 92300 946 92302
rect 970 92300 1026 92302
rect 1050 92300 1106 92302
rect 1130 92300 1186 92302
rect 890 92248 916 92300
rect 916 92248 946 92300
rect 970 92248 980 92300
rect 980 92248 1026 92300
rect 1050 92248 1096 92300
rect 1096 92248 1106 92300
rect 1130 92248 1160 92300
rect 1160 92248 1186 92300
rect 890 92246 946 92248
rect 970 92246 1026 92248
rect 1050 92246 1106 92248
rect 1130 92246 1186 92248
rect 890 91212 946 91214
rect 970 91212 1026 91214
rect 1050 91212 1106 91214
rect 1130 91212 1186 91214
rect 890 91160 916 91212
rect 916 91160 946 91212
rect 970 91160 980 91212
rect 980 91160 1026 91212
rect 1050 91160 1096 91212
rect 1096 91160 1106 91212
rect 1130 91160 1160 91212
rect 1160 91160 1186 91212
rect 890 91158 946 91160
rect 970 91158 1026 91160
rect 1050 91158 1106 91160
rect 1130 91158 1186 91160
rect 890 90124 946 90126
rect 970 90124 1026 90126
rect 1050 90124 1106 90126
rect 1130 90124 1186 90126
rect 890 90072 916 90124
rect 916 90072 946 90124
rect 970 90072 980 90124
rect 980 90072 1026 90124
rect 1050 90072 1096 90124
rect 1096 90072 1106 90124
rect 1130 90072 1160 90124
rect 1160 90072 1186 90124
rect 890 90070 946 90072
rect 970 90070 1026 90072
rect 1050 90070 1106 90072
rect 1130 90070 1186 90072
rect 890 89036 946 89038
rect 970 89036 1026 89038
rect 1050 89036 1106 89038
rect 1130 89036 1186 89038
rect 890 88984 916 89036
rect 916 88984 946 89036
rect 970 88984 980 89036
rect 980 88984 1026 89036
rect 1050 88984 1096 89036
rect 1096 88984 1106 89036
rect 1130 88984 1160 89036
rect 1160 88984 1186 89036
rect 890 88982 946 88984
rect 970 88982 1026 88984
rect 1050 88982 1106 88984
rect 1130 88982 1186 88984
rect 890 87948 946 87950
rect 970 87948 1026 87950
rect 1050 87948 1106 87950
rect 1130 87948 1186 87950
rect 890 87896 916 87948
rect 916 87896 946 87948
rect 970 87896 980 87948
rect 980 87896 1026 87948
rect 1050 87896 1096 87948
rect 1096 87896 1106 87948
rect 1130 87896 1160 87948
rect 1160 87896 1186 87948
rect 890 87894 946 87896
rect 970 87894 1026 87896
rect 1050 87894 1106 87896
rect 1130 87894 1186 87896
rect 890 86860 946 86862
rect 970 86860 1026 86862
rect 1050 86860 1106 86862
rect 1130 86860 1186 86862
rect 890 86808 916 86860
rect 916 86808 946 86860
rect 970 86808 980 86860
rect 980 86808 1026 86860
rect 1050 86808 1096 86860
rect 1096 86808 1106 86860
rect 1130 86808 1160 86860
rect 1160 86808 1186 86860
rect 890 86806 946 86808
rect 970 86806 1026 86808
rect 1050 86806 1106 86808
rect 1130 86806 1186 86808
rect 890 85772 946 85774
rect 970 85772 1026 85774
rect 1050 85772 1106 85774
rect 1130 85772 1186 85774
rect 890 85720 916 85772
rect 916 85720 946 85772
rect 970 85720 980 85772
rect 980 85720 1026 85772
rect 1050 85720 1096 85772
rect 1096 85720 1106 85772
rect 1130 85720 1160 85772
rect 1160 85720 1186 85772
rect 890 85718 946 85720
rect 970 85718 1026 85720
rect 1050 85718 1106 85720
rect 1130 85718 1186 85720
rect 890 84684 946 84686
rect 970 84684 1026 84686
rect 1050 84684 1106 84686
rect 1130 84684 1186 84686
rect 890 84632 916 84684
rect 916 84632 946 84684
rect 970 84632 980 84684
rect 980 84632 1026 84684
rect 1050 84632 1096 84684
rect 1096 84632 1106 84684
rect 1130 84632 1160 84684
rect 1160 84632 1186 84684
rect 890 84630 946 84632
rect 970 84630 1026 84632
rect 1050 84630 1106 84632
rect 1130 84630 1186 84632
rect 890 83596 946 83598
rect 970 83596 1026 83598
rect 1050 83596 1106 83598
rect 1130 83596 1186 83598
rect 890 83544 916 83596
rect 916 83544 946 83596
rect 970 83544 980 83596
rect 980 83544 1026 83596
rect 1050 83544 1096 83596
rect 1096 83544 1106 83596
rect 1130 83544 1160 83596
rect 1160 83544 1186 83596
rect 890 83542 946 83544
rect 970 83542 1026 83544
rect 1050 83542 1106 83544
rect 1130 83542 1186 83544
rect 890 82508 946 82510
rect 970 82508 1026 82510
rect 1050 82508 1106 82510
rect 1130 82508 1186 82510
rect 890 82456 916 82508
rect 916 82456 946 82508
rect 970 82456 980 82508
rect 980 82456 1026 82508
rect 1050 82456 1096 82508
rect 1096 82456 1106 82508
rect 1130 82456 1160 82508
rect 1160 82456 1186 82508
rect 890 82454 946 82456
rect 970 82454 1026 82456
rect 1050 82454 1106 82456
rect 1130 82454 1186 82456
rect 890 81420 946 81422
rect 970 81420 1026 81422
rect 1050 81420 1106 81422
rect 1130 81420 1186 81422
rect 890 81368 916 81420
rect 916 81368 946 81420
rect 970 81368 980 81420
rect 980 81368 1026 81420
rect 1050 81368 1096 81420
rect 1096 81368 1106 81420
rect 1130 81368 1160 81420
rect 1160 81368 1186 81420
rect 890 81366 946 81368
rect 970 81366 1026 81368
rect 1050 81366 1106 81368
rect 1130 81366 1186 81368
rect 890 80332 946 80334
rect 970 80332 1026 80334
rect 1050 80332 1106 80334
rect 1130 80332 1186 80334
rect 890 80280 916 80332
rect 916 80280 946 80332
rect 970 80280 980 80332
rect 980 80280 1026 80332
rect 1050 80280 1096 80332
rect 1096 80280 1106 80332
rect 1130 80280 1160 80332
rect 1160 80280 1186 80332
rect 890 80278 946 80280
rect 970 80278 1026 80280
rect 1050 80278 1106 80280
rect 1130 80278 1186 80280
rect 890 79244 946 79246
rect 970 79244 1026 79246
rect 1050 79244 1106 79246
rect 1130 79244 1186 79246
rect 890 79192 916 79244
rect 916 79192 946 79244
rect 970 79192 980 79244
rect 980 79192 1026 79244
rect 1050 79192 1096 79244
rect 1096 79192 1106 79244
rect 1130 79192 1160 79244
rect 1160 79192 1186 79244
rect 890 79190 946 79192
rect 970 79190 1026 79192
rect 1050 79190 1106 79192
rect 1130 79190 1186 79192
rect 890 78156 946 78158
rect 970 78156 1026 78158
rect 1050 78156 1106 78158
rect 1130 78156 1186 78158
rect 890 78104 916 78156
rect 916 78104 946 78156
rect 970 78104 980 78156
rect 980 78104 1026 78156
rect 1050 78104 1096 78156
rect 1096 78104 1106 78156
rect 1130 78104 1160 78156
rect 1160 78104 1186 78156
rect 890 78102 946 78104
rect 970 78102 1026 78104
rect 1050 78102 1106 78104
rect 1130 78102 1186 78104
rect 890 77068 946 77070
rect 970 77068 1026 77070
rect 1050 77068 1106 77070
rect 1130 77068 1186 77070
rect 890 77016 916 77068
rect 916 77016 946 77068
rect 970 77016 980 77068
rect 980 77016 1026 77068
rect 1050 77016 1096 77068
rect 1096 77016 1106 77068
rect 1130 77016 1160 77068
rect 1160 77016 1186 77068
rect 890 77014 946 77016
rect 970 77014 1026 77016
rect 1050 77014 1106 77016
rect 1130 77014 1186 77016
rect 890 75980 946 75982
rect 970 75980 1026 75982
rect 1050 75980 1106 75982
rect 1130 75980 1186 75982
rect 890 75928 916 75980
rect 916 75928 946 75980
rect 970 75928 980 75980
rect 980 75928 1026 75980
rect 1050 75928 1096 75980
rect 1096 75928 1106 75980
rect 1130 75928 1160 75980
rect 1160 75928 1186 75980
rect 890 75926 946 75928
rect 970 75926 1026 75928
rect 1050 75926 1106 75928
rect 1130 75926 1186 75928
rect 890 74892 946 74894
rect 970 74892 1026 74894
rect 1050 74892 1106 74894
rect 1130 74892 1186 74894
rect 890 74840 916 74892
rect 916 74840 946 74892
rect 970 74840 980 74892
rect 980 74840 1026 74892
rect 1050 74840 1096 74892
rect 1096 74840 1106 74892
rect 1130 74840 1160 74892
rect 1160 74840 1186 74892
rect 890 74838 946 74840
rect 970 74838 1026 74840
rect 1050 74838 1106 74840
rect 1130 74838 1186 74840
rect 890 73804 946 73806
rect 970 73804 1026 73806
rect 1050 73804 1106 73806
rect 1130 73804 1186 73806
rect 890 73752 916 73804
rect 916 73752 946 73804
rect 970 73752 980 73804
rect 980 73752 1026 73804
rect 1050 73752 1096 73804
rect 1096 73752 1106 73804
rect 1130 73752 1160 73804
rect 1160 73752 1186 73804
rect 890 73750 946 73752
rect 970 73750 1026 73752
rect 1050 73750 1106 73752
rect 1130 73750 1186 73752
rect 890 72716 946 72718
rect 970 72716 1026 72718
rect 1050 72716 1106 72718
rect 1130 72716 1186 72718
rect 890 72664 916 72716
rect 916 72664 946 72716
rect 970 72664 980 72716
rect 980 72664 1026 72716
rect 1050 72664 1096 72716
rect 1096 72664 1106 72716
rect 1130 72664 1160 72716
rect 1160 72664 1186 72716
rect 890 72662 946 72664
rect 970 72662 1026 72664
rect 1050 72662 1106 72664
rect 1130 72662 1186 72664
rect 890 71628 946 71630
rect 970 71628 1026 71630
rect 1050 71628 1106 71630
rect 1130 71628 1186 71630
rect 890 71576 916 71628
rect 916 71576 946 71628
rect 970 71576 980 71628
rect 980 71576 1026 71628
rect 1050 71576 1096 71628
rect 1096 71576 1106 71628
rect 1130 71576 1160 71628
rect 1160 71576 1186 71628
rect 890 71574 946 71576
rect 970 71574 1026 71576
rect 1050 71574 1106 71576
rect 1130 71574 1186 71576
rect 890 70540 946 70542
rect 970 70540 1026 70542
rect 1050 70540 1106 70542
rect 1130 70540 1186 70542
rect 890 70488 916 70540
rect 916 70488 946 70540
rect 970 70488 980 70540
rect 980 70488 1026 70540
rect 1050 70488 1096 70540
rect 1096 70488 1106 70540
rect 1130 70488 1160 70540
rect 1160 70488 1186 70540
rect 890 70486 946 70488
rect 970 70486 1026 70488
rect 1050 70486 1106 70488
rect 1130 70486 1186 70488
rect 890 69452 946 69454
rect 970 69452 1026 69454
rect 1050 69452 1106 69454
rect 1130 69452 1186 69454
rect 890 69400 916 69452
rect 916 69400 946 69452
rect 970 69400 980 69452
rect 980 69400 1026 69452
rect 1050 69400 1096 69452
rect 1096 69400 1106 69452
rect 1130 69400 1160 69452
rect 1160 69400 1186 69452
rect 890 69398 946 69400
rect 970 69398 1026 69400
rect 1050 69398 1106 69400
rect 1130 69398 1186 69400
rect 890 68364 946 68366
rect 970 68364 1026 68366
rect 1050 68364 1106 68366
rect 1130 68364 1186 68366
rect 890 68312 916 68364
rect 916 68312 946 68364
rect 970 68312 980 68364
rect 980 68312 1026 68364
rect 1050 68312 1096 68364
rect 1096 68312 1106 68364
rect 1130 68312 1160 68364
rect 1160 68312 1186 68364
rect 890 68310 946 68312
rect 970 68310 1026 68312
rect 1050 68310 1106 68312
rect 1130 68310 1186 68312
rect 890 67276 946 67278
rect 970 67276 1026 67278
rect 1050 67276 1106 67278
rect 1130 67276 1186 67278
rect 890 67224 916 67276
rect 916 67224 946 67276
rect 970 67224 980 67276
rect 980 67224 1026 67276
rect 1050 67224 1096 67276
rect 1096 67224 1106 67276
rect 1130 67224 1160 67276
rect 1160 67224 1186 67276
rect 890 67222 946 67224
rect 970 67222 1026 67224
rect 1050 67222 1106 67224
rect 1130 67222 1186 67224
rect 890 66188 946 66190
rect 970 66188 1026 66190
rect 1050 66188 1106 66190
rect 1130 66188 1186 66190
rect 890 66136 916 66188
rect 916 66136 946 66188
rect 970 66136 980 66188
rect 980 66136 1026 66188
rect 1050 66136 1096 66188
rect 1096 66136 1106 66188
rect 1130 66136 1160 66188
rect 1160 66136 1186 66188
rect 890 66134 946 66136
rect 970 66134 1026 66136
rect 1050 66134 1106 66136
rect 1130 66134 1186 66136
rect 890 65100 946 65102
rect 970 65100 1026 65102
rect 1050 65100 1106 65102
rect 1130 65100 1186 65102
rect 890 65048 916 65100
rect 916 65048 946 65100
rect 970 65048 980 65100
rect 980 65048 1026 65100
rect 1050 65048 1096 65100
rect 1096 65048 1106 65100
rect 1130 65048 1160 65100
rect 1160 65048 1186 65100
rect 890 65046 946 65048
rect 970 65046 1026 65048
rect 1050 65046 1106 65048
rect 1130 65046 1186 65048
rect 890 64012 946 64014
rect 970 64012 1026 64014
rect 1050 64012 1106 64014
rect 1130 64012 1186 64014
rect 890 63960 916 64012
rect 916 63960 946 64012
rect 970 63960 980 64012
rect 980 63960 1026 64012
rect 1050 63960 1096 64012
rect 1096 63960 1106 64012
rect 1130 63960 1160 64012
rect 1160 63960 1186 64012
rect 890 63958 946 63960
rect 970 63958 1026 63960
rect 1050 63958 1106 63960
rect 1130 63958 1186 63960
rect 890 62924 946 62926
rect 970 62924 1026 62926
rect 1050 62924 1106 62926
rect 1130 62924 1186 62926
rect 890 62872 916 62924
rect 916 62872 946 62924
rect 970 62872 980 62924
rect 980 62872 1026 62924
rect 1050 62872 1096 62924
rect 1096 62872 1106 62924
rect 1130 62872 1160 62924
rect 1160 62872 1186 62924
rect 890 62870 946 62872
rect 970 62870 1026 62872
rect 1050 62870 1106 62872
rect 1130 62870 1186 62872
rect 890 61836 946 61838
rect 970 61836 1026 61838
rect 1050 61836 1106 61838
rect 1130 61836 1186 61838
rect 890 61784 916 61836
rect 916 61784 946 61836
rect 970 61784 980 61836
rect 980 61784 1026 61836
rect 1050 61784 1096 61836
rect 1096 61784 1106 61836
rect 1130 61784 1160 61836
rect 1160 61784 1186 61836
rect 890 61782 946 61784
rect 970 61782 1026 61784
rect 1050 61782 1106 61784
rect 1130 61782 1186 61784
rect 890 60748 946 60750
rect 970 60748 1026 60750
rect 1050 60748 1106 60750
rect 1130 60748 1186 60750
rect 890 60696 916 60748
rect 916 60696 946 60748
rect 970 60696 980 60748
rect 980 60696 1026 60748
rect 1050 60696 1096 60748
rect 1096 60696 1106 60748
rect 1130 60696 1160 60748
rect 1160 60696 1186 60748
rect 890 60694 946 60696
rect 970 60694 1026 60696
rect 1050 60694 1106 60696
rect 1130 60694 1186 60696
rect 890 59660 946 59662
rect 970 59660 1026 59662
rect 1050 59660 1106 59662
rect 1130 59660 1186 59662
rect 890 59608 916 59660
rect 916 59608 946 59660
rect 970 59608 980 59660
rect 980 59608 1026 59660
rect 1050 59608 1096 59660
rect 1096 59608 1106 59660
rect 1130 59608 1160 59660
rect 1160 59608 1186 59660
rect 890 59606 946 59608
rect 970 59606 1026 59608
rect 1050 59606 1106 59608
rect 1130 59606 1186 59608
rect 890 58572 946 58574
rect 970 58572 1026 58574
rect 1050 58572 1106 58574
rect 1130 58572 1186 58574
rect 890 58520 916 58572
rect 916 58520 946 58572
rect 970 58520 980 58572
rect 980 58520 1026 58572
rect 1050 58520 1096 58572
rect 1096 58520 1106 58572
rect 1130 58520 1160 58572
rect 1160 58520 1186 58572
rect 890 58518 946 58520
rect 970 58518 1026 58520
rect 1050 58518 1106 58520
rect 1130 58518 1186 58520
rect 890 57484 946 57486
rect 970 57484 1026 57486
rect 1050 57484 1106 57486
rect 1130 57484 1186 57486
rect 890 57432 916 57484
rect 916 57432 946 57484
rect 970 57432 980 57484
rect 980 57432 1026 57484
rect 1050 57432 1096 57484
rect 1096 57432 1106 57484
rect 1130 57432 1160 57484
rect 1160 57432 1186 57484
rect 890 57430 946 57432
rect 970 57430 1026 57432
rect 1050 57430 1106 57432
rect 1130 57430 1186 57432
rect 890 56396 946 56398
rect 970 56396 1026 56398
rect 1050 56396 1106 56398
rect 1130 56396 1186 56398
rect 890 56344 916 56396
rect 916 56344 946 56396
rect 970 56344 980 56396
rect 980 56344 1026 56396
rect 1050 56344 1096 56396
rect 1096 56344 1106 56396
rect 1130 56344 1160 56396
rect 1160 56344 1186 56396
rect 890 56342 946 56344
rect 970 56342 1026 56344
rect 1050 56342 1106 56344
rect 1130 56342 1186 56344
rect 890 55308 946 55310
rect 970 55308 1026 55310
rect 1050 55308 1106 55310
rect 1130 55308 1186 55310
rect 890 55256 916 55308
rect 916 55256 946 55308
rect 970 55256 980 55308
rect 980 55256 1026 55308
rect 1050 55256 1096 55308
rect 1096 55256 1106 55308
rect 1130 55256 1160 55308
rect 1160 55256 1186 55308
rect 890 55254 946 55256
rect 970 55254 1026 55256
rect 1050 55254 1106 55256
rect 1130 55254 1186 55256
rect 890 54220 946 54222
rect 970 54220 1026 54222
rect 1050 54220 1106 54222
rect 1130 54220 1186 54222
rect 890 54168 916 54220
rect 916 54168 946 54220
rect 970 54168 980 54220
rect 980 54168 1026 54220
rect 1050 54168 1096 54220
rect 1096 54168 1106 54220
rect 1130 54168 1160 54220
rect 1160 54168 1186 54220
rect 890 54166 946 54168
rect 970 54166 1026 54168
rect 1050 54166 1106 54168
rect 1130 54166 1186 54168
rect 890 53132 946 53134
rect 970 53132 1026 53134
rect 1050 53132 1106 53134
rect 1130 53132 1186 53134
rect 890 53080 916 53132
rect 916 53080 946 53132
rect 970 53080 980 53132
rect 980 53080 1026 53132
rect 1050 53080 1096 53132
rect 1096 53080 1106 53132
rect 1130 53080 1160 53132
rect 1160 53080 1186 53132
rect 890 53078 946 53080
rect 970 53078 1026 53080
rect 1050 53078 1106 53080
rect 1130 53078 1186 53080
rect 890 52044 946 52046
rect 970 52044 1026 52046
rect 1050 52044 1106 52046
rect 1130 52044 1186 52046
rect 890 51992 916 52044
rect 916 51992 946 52044
rect 970 51992 980 52044
rect 980 51992 1026 52044
rect 1050 51992 1096 52044
rect 1096 51992 1106 52044
rect 1130 51992 1160 52044
rect 1160 51992 1186 52044
rect 890 51990 946 51992
rect 970 51990 1026 51992
rect 1050 51990 1106 51992
rect 1130 51990 1186 51992
rect 890 50956 946 50958
rect 970 50956 1026 50958
rect 1050 50956 1106 50958
rect 1130 50956 1186 50958
rect 890 50904 916 50956
rect 916 50904 946 50956
rect 970 50904 980 50956
rect 980 50904 1026 50956
rect 1050 50904 1096 50956
rect 1096 50904 1106 50956
rect 1130 50904 1160 50956
rect 1160 50904 1186 50956
rect 890 50902 946 50904
rect 970 50902 1026 50904
rect 1050 50902 1106 50904
rect 1130 50902 1186 50904
rect 890 49868 946 49870
rect 970 49868 1026 49870
rect 1050 49868 1106 49870
rect 1130 49868 1186 49870
rect 890 49816 916 49868
rect 916 49816 946 49868
rect 970 49816 980 49868
rect 980 49816 1026 49868
rect 1050 49816 1096 49868
rect 1096 49816 1106 49868
rect 1130 49816 1160 49868
rect 1160 49816 1186 49868
rect 890 49814 946 49816
rect 970 49814 1026 49816
rect 1050 49814 1106 49816
rect 1130 49814 1186 49816
rect 890 48780 946 48782
rect 970 48780 1026 48782
rect 1050 48780 1106 48782
rect 1130 48780 1186 48782
rect 890 48728 916 48780
rect 916 48728 946 48780
rect 970 48728 980 48780
rect 980 48728 1026 48780
rect 1050 48728 1096 48780
rect 1096 48728 1106 48780
rect 1130 48728 1160 48780
rect 1160 48728 1186 48780
rect 890 48726 946 48728
rect 970 48726 1026 48728
rect 1050 48726 1106 48728
rect 1130 48726 1186 48728
rect 890 47692 946 47694
rect 970 47692 1026 47694
rect 1050 47692 1106 47694
rect 1130 47692 1186 47694
rect 890 47640 916 47692
rect 916 47640 946 47692
rect 970 47640 980 47692
rect 980 47640 1026 47692
rect 1050 47640 1096 47692
rect 1096 47640 1106 47692
rect 1130 47640 1160 47692
rect 1160 47640 1186 47692
rect 890 47638 946 47640
rect 970 47638 1026 47640
rect 1050 47638 1106 47640
rect 1130 47638 1186 47640
rect 890 46604 946 46606
rect 970 46604 1026 46606
rect 1050 46604 1106 46606
rect 1130 46604 1186 46606
rect 890 46552 916 46604
rect 916 46552 946 46604
rect 970 46552 980 46604
rect 980 46552 1026 46604
rect 1050 46552 1096 46604
rect 1096 46552 1106 46604
rect 1130 46552 1160 46604
rect 1160 46552 1186 46604
rect 890 46550 946 46552
rect 970 46550 1026 46552
rect 1050 46550 1106 46552
rect 1130 46550 1186 46552
rect 890 45516 946 45518
rect 970 45516 1026 45518
rect 1050 45516 1106 45518
rect 1130 45516 1186 45518
rect 890 45464 916 45516
rect 916 45464 946 45516
rect 970 45464 980 45516
rect 980 45464 1026 45516
rect 1050 45464 1096 45516
rect 1096 45464 1106 45516
rect 1130 45464 1160 45516
rect 1160 45464 1186 45516
rect 890 45462 946 45464
rect 970 45462 1026 45464
rect 1050 45462 1106 45464
rect 1130 45462 1186 45464
rect 890 44428 946 44430
rect 970 44428 1026 44430
rect 1050 44428 1106 44430
rect 1130 44428 1186 44430
rect 890 44376 916 44428
rect 916 44376 946 44428
rect 970 44376 980 44428
rect 980 44376 1026 44428
rect 1050 44376 1096 44428
rect 1096 44376 1106 44428
rect 1130 44376 1160 44428
rect 1160 44376 1186 44428
rect 890 44374 946 44376
rect 970 44374 1026 44376
rect 1050 44374 1106 44376
rect 1130 44374 1186 44376
rect 890 43340 946 43342
rect 970 43340 1026 43342
rect 1050 43340 1106 43342
rect 1130 43340 1186 43342
rect 890 43288 916 43340
rect 916 43288 946 43340
rect 970 43288 980 43340
rect 980 43288 1026 43340
rect 1050 43288 1096 43340
rect 1096 43288 1106 43340
rect 1130 43288 1160 43340
rect 1160 43288 1186 43340
rect 890 43286 946 43288
rect 970 43286 1026 43288
rect 1050 43286 1106 43288
rect 1130 43286 1186 43288
rect 890 42252 946 42254
rect 970 42252 1026 42254
rect 1050 42252 1106 42254
rect 1130 42252 1186 42254
rect 890 42200 916 42252
rect 916 42200 946 42252
rect 970 42200 980 42252
rect 980 42200 1026 42252
rect 1050 42200 1096 42252
rect 1096 42200 1106 42252
rect 1130 42200 1160 42252
rect 1160 42200 1186 42252
rect 890 42198 946 42200
rect 970 42198 1026 42200
rect 1050 42198 1106 42200
rect 1130 42198 1186 42200
rect 890 41164 946 41166
rect 970 41164 1026 41166
rect 1050 41164 1106 41166
rect 1130 41164 1186 41166
rect 890 41112 916 41164
rect 916 41112 946 41164
rect 970 41112 980 41164
rect 980 41112 1026 41164
rect 1050 41112 1096 41164
rect 1096 41112 1106 41164
rect 1130 41112 1160 41164
rect 1160 41112 1186 41164
rect 890 41110 946 41112
rect 970 41110 1026 41112
rect 1050 41110 1106 41112
rect 1130 41110 1186 41112
rect 890 40076 946 40078
rect 970 40076 1026 40078
rect 1050 40076 1106 40078
rect 1130 40076 1186 40078
rect 890 40024 916 40076
rect 916 40024 946 40076
rect 970 40024 980 40076
rect 980 40024 1026 40076
rect 1050 40024 1096 40076
rect 1096 40024 1106 40076
rect 1130 40024 1160 40076
rect 1160 40024 1186 40076
rect 890 40022 946 40024
rect 970 40022 1026 40024
rect 1050 40022 1106 40024
rect 1130 40022 1186 40024
rect 890 38988 946 38990
rect 970 38988 1026 38990
rect 1050 38988 1106 38990
rect 1130 38988 1186 38990
rect 890 38936 916 38988
rect 916 38936 946 38988
rect 970 38936 980 38988
rect 980 38936 1026 38988
rect 1050 38936 1096 38988
rect 1096 38936 1106 38988
rect 1130 38936 1160 38988
rect 1160 38936 1186 38988
rect 890 38934 946 38936
rect 970 38934 1026 38936
rect 1050 38934 1106 38936
rect 1130 38934 1186 38936
rect 890 37900 946 37902
rect 970 37900 1026 37902
rect 1050 37900 1106 37902
rect 1130 37900 1186 37902
rect 890 37848 916 37900
rect 916 37848 946 37900
rect 970 37848 980 37900
rect 980 37848 1026 37900
rect 1050 37848 1096 37900
rect 1096 37848 1106 37900
rect 1130 37848 1160 37900
rect 1160 37848 1186 37900
rect 890 37846 946 37848
rect 970 37846 1026 37848
rect 1050 37846 1106 37848
rect 1130 37846 1186 37848
rect 890 36812 946 36814
rect 970 36812 1026 36814
rect 1050 36812 1106 36814
rect 1130 36812 1186 36814
rect 890 36760 916 36812
rect 916 36760 946 36812
rect 970 36760 980 36812
rect 980 36760 1026 36812
rect 1050 36760 1096 36812
rect 1096 36760 1106 36812
rect 1130 36760 1160 36812
rect 1160 36760 1186 36812
rect 890 36758 946 36760
rect 970 36758 1026 36760
rect 1050 36758 1106 36760
rect 1130 36758 1186 36760
rect 890 35724 946 35726
rect 970 35724 1026 35726
rect 1050 35724 1106 35726
rect 1130 35724 1186 35726
rect 890 35672 916 35724
rect 916 35672 946 35724
rect 970 35672 980 35724
rect 980 35672 1026 35724
rect 1050 35672 1096 35724
rect 1096 35672 1106 35724
rect 1130 35672 1160 35724
rect 1160 35672 1186 35724
rect 890 35670 946 35672
rect 970 35670 1026 35672
rect 1050 35670 1106 35672
rect 1130 35670 1186 35672
rect 890 34636 946 34638
rect 970 34636 1026 34638
rect 1050 34636 1106 34638
rect 1130 34636 1186 34638
rect 890 34584 916 34636
rect 916 34584 946 34636
rect 970 34584 980 34636
rect 980 34584 1026 34636
rect 1050 34584 1096 34636
rect 1096 34584 1106 34636
rect 1130 34584 1160 34636
rect 1160 34584 1186 34636
rect 890 34582 946 34584
rect 970 34582 1026 34584
rect 1050 34582 1106 34584
rect 1130 34582 1186 34584
rect 890 33548 946 33550
rect 970 33548 1026 33550
rect 1050 33548 1106 33550
rect 1130 33548 1186 33550
rect 890 33496 916 33548
rect 916 33496 946 33548
rect 970 33496 980 33548
rect 980 33496 1026 33548
rect 1050 33496 1096 33548
rect 1096 33496 1106 33548
rect 1130 33496 1160 33548
rect 1160 33496 1186 33548
rect 890 33494 946 33496
rect 970 33494 1026 33496
rect 1050 33494 1106 33496
rect 1130 33494 1186 33496
rect 890 32460 946 32462
rect 970 32460 1026 32462
rect 1050 32460 1106 32462
rect 1130 32460 1186 32462
rect 890 32408 916 32460
rect 916 32408 946 32460
rect 970 32408 980 32460
rect 980 32408 1026 32460
rect 1050 32408 1096 32460
rect 1096 32408 1106 32460
rect 1130 32408 1160 32460
rect 1160 32408 1186 32460
rect 890 32406 946 32408
rect 970 32406 1026 32408
rect 1050 32406 1106 32408
rect 1130 32406 1186 32408
rect 890 31372 946 31374
rect 970 31372 1026 31374
rect 1050 31372 1106 31374
rect 1130 31372 1186 31374
rect 890 31320 916 31372
rect 916 31320 946 31372
rect 970 31320 980 31372
rect 980 31320 1026 31372
rect 1050 31320 1096 31372
rect 1096 31320 1106 31372
rect 1130 31320 1160 31372
rect 1160 31320 1186 31372
rect 890 31318 946 31320
rect 970 31318 1026 31320
rect 1050 31318 1106 31320
rect 1130 31318 1186 31320
rect 890 30284 946 30286
rect 970 30284 1026 30286
rect 1050 30284 1106 30286
rect 1130 30284 1186 30286
rect 890 30232 916 30284
rect 916 30232 946 30284
rect 970 30232 980 30284
rect 980 30232 1026 30284
rect 1050 30232 1096 30284
rect 1096 30232 1106 30284
rect 1130 30232 1160 30284
rect 1160 30232 1186 30284
rect 890 30230 946 30232
rect 970 30230 1026 30232
rect 1050 30230 1106 30232
rect 1130 30230 1186 30232
rect 890 29196 946 29198
rect 970 29196 1026 29198
rect 1050 29196 1106 29198
rect 1130 29196 1186 29198
rect 890 29144 916 29196
rect 916 29144 946 29196
rect 970 29144 980 29196
rect 980 29144 1026 29196
rect 1050 29144 1096 29196
rect 1096 29144 1106 29196
rect 1130 29144 1160 29196
rect 1160 29144 1186 29196
rect 890 29142 946 29144
rect 970 29142 1026 29144
rect 1050 29142 1106 29144
rect 1130 29142 1186 29144
rect 890 28108 946 28110
rect 970 28108 1026 28110
rect 1050 28108 1106 28110
rect 1130 28108 1186 28110
rect 890 28056 916 28108
rect 916 28056 946 28108
rect 970 28056 980 28108
rect 980 28056 1026 28108
rect 1050 28056 1096 28108
rect 1096 28056 1106 28108
rect 1130 28056 1160 28108
rect 1160 28056 1186 28108
rect 890 28054 946 28056
rect 970 28054 1026 28056
rect 1050 28054 1106 28056
rect 1130 28054 1186 28056
rect 890 27020 946 27022
rect 970 27020 1026 27022
rect 1050 27020 1106 27022
rect 1130 27020 1186 27022
rect 890 26968 916 27020
rect 916 26968 946 27020
rect 970 26968 980 27020
rect 980 26968 1026 27020
rect 1050 26968 1096 27020
rect 1096 26968 1106 27020
rect 1130 26968 1160 27020
rect 1160 26968 1186 27020
rect 890 26966 946 26968
rect 970 26966 1026 26968
rect 1050 26966 1106 26968
rect 1130 26966 1186 26968
rect 890 25932 946 25934
rect 970 25932 1026 25934
rect 1050 25932 1106 25934
rect 1130 25932 1186 25934
rect 890 25880 916 25932
rect 916 25880 946 25932
rect 970 25880 980 25932
rect 980 25880 1026 25932
rect 1050 25880 1096 25932
rect 1096 25880 1106 25932
rect 1130 25880 1160 25932
rect 1160 25880 1186 25932
rect 890 25878 946 25880
rect 970 25878 1026 25880
rect 1050 25878 1106 25880
rect 1130 25878 1186 25880
rect 890 24844 946 24846
rect 970 24844 1026 24846
rect 1050 24844 1106 24846
rect 1130 24844 1186 24846
rect 890 24792 916 24844
rect 916 24792 946 24844
rect 970 24792 980 24844
rect 980 24792 1026 24844
rect 1050 24792 1096 24844
rect 1096 24792 1106 24844
rect 1130 24792 1160 24844
rect 1160 24792 1186 24844
rect 890 24790 946 24792
rect 970 24790 1026 24792
rect 1050 24790 1106 24792
rect 1130 24790 1186 24792
rect 890 23756 946 23758
rect 970 23756 1026 23758
rect 1050 23756 1106 23758
rect 1130 23756 1186 23758
rect 890 23704 916 23756
rect 916 23704 946 23756
rect 970 23704 980 23756
rect 980 23704 1026 23756
rect 1050 23704 1096 23756
rect 1096 23704 1106 23756
rect 1130 23704 1160 23756
rect 1160 23704 1186 23756
rect 890 23702 946 23704
rect 970 23702 1026 23704
rect 1050 23702 1106 23704
rect 1130 23702 1186 23704
rect 890 22668 946 22670
rect 970 22668 1026 22670
rect 1050 22668 1106 22670
rect 1130 22668 1186 22670
rect 890 22616 916 22668
rect 916 22616 946 22668
rect 970 22616 980 22668
rect 980 22616 1026 22668
rect 1050 22616 1096 22668
rect 1096 22616 1106 22668
rect 1130 22616 1160 22668
rect 1160 22616 1186 22668
rect 890 22614 946 22616
rect 970 22614 1026 22616
rect 1050 22614 1106 22616
rect 1130 22614 1186 22616
rect 890 21580 946 21582
rect 970 21580 1026 21582
rect 1050 21580 1106 21582
rect 1130 21580 1186 21582
rect 890 21528 916 21580
rect 916 21528 946 21580
rect 970 21528 980 21580
rect 980 21528 1026 21580
rect 1050 21528 1096 21580
rect 1096 21528 1106 21580
rect 1130 21528 1160 21580
rect 1160 21528 1186 21580
rect 890 21526 946 21528
rect 970 21526 1026 21528
rect 1050 21526 1106 21528
rect 1130 21526 1186 21528
rect 890 20492 946 20494
rect 970 20492 1026 20494
rect 1050 20492 1106 20494
rect 1130 20492 1186 20494
rect 890 20440 916 20492
rect 916 20440 946 20492
rect 970 20440 980 20492
rect 980 20440 1026 20492
rect 1050 20440 1096 20492
rect 1096 20440 1106 20492
rect 1130 20440 1160 20492
rect 1160 20440 1186 20492
rect 890 20438 946 20440
rect 970 20438 1026 20440
rect 1050 20438 1106 20440
rect 1130 20438 1186 20440
rect 890 19404 946 19406
rect 970 19404 1026 19406
rect 1050 19404 1106 19406
rect 1130 19404 1186 19406
rect 890 19352 916 19404
rect 916 19352 946 19404
rect 970 19352 980 19404
rect 980 19352 1026 19404
rect 1050 19352 1096 19404
rect 1096 19352 1106 19404
rect 1130 19352 1160 19404
rect 1160 19352 1186 19404
rect 890 19350 946 19352
rect 970 19350 1026 19352
rect 1050 19350 1106 19352
rect 1130 19350 1186 19352
rect 890 18316 946 18318
rect 970 18316 1026 18318
rect 1050 18316 1106 18318
rect 1130 18316 1186 18318
rect 890 18264 916 18316
rect 916 18264 946 18316
rect 970 18264 980 18316
rect 980 18264 1026 18316
rect 1050 18264 1096 18316
rect 1096 18264 1106 18316
rect 1130 18264 1160 18316
rect 1160 18264 1186 18316
rect 890 18262 946 18264
rect 970 18262 1026 18264
rect 1050 18262 1106 18264
rect 1130 18262 1186 18264
rect 890 17228 946 17230
rect 970 17228 1026 17230
rect 1050 17228 1106 17230
rect 1130 17228 1186 17230
rect 890 17176 916 17228
rect 916 17176 946 17228
rect 970 17176 980 17228
rect 980 17176 1026 17228
rect 1050 17176 1096 17228
rect 1096 17176 1106 17228
rect 1130 17176 1160 17228
rect 1160 17176 1186 17228
rect 890 17174 946 17176
rect 970 17174 1026 17176
rect 1050 17174 1106 17176
rect 1130 17174 1186 17176
rect 890 16140 946 16142
rect 970 16140 1026 16142
rect 1050 16140 1106 16142
rect 1130 16140 1186 16142
rect 890 16088 916 16140
rect 916 16088 946 16140
rect 970 16088 980 16140
rect 980 16088 1026 16140
rect 1050 16088 1096 16140
rect 1096 16088 1106 16140
rect 1130 16088 1160 16140
rect 1160 16088 1186 16140
rect 890 16086 946 16088
rect 970 16086 1026 16088
rect 1050 16086 1106 16088
rect 1130 16086 1186 16088
rect 890 15052 946 15054
rect 970 15052 1026 15054
rect 1050 15052 1106 15054
rect 1130 15052 1186 15054
rect 890 15000 916 15052
rect 916 15000 946 15052
rect 970 15000 980 15052
rect 980 15000 1026 15052
rect 1050 15000 1096 15052
rect 1096 15000 1106 15052
rect 1130 15000 1160 15052
rect 1160 15000 1186 15052
rect 890 14998 946 15000
rect 970 14998 1026 15000
rect 1050 14998 1106 15000
rect 1130 14998 1186 15000
rect 890 13964 946 13966
rect 970 13964 1026 13966
rect 1050 13964 1106 13966
rect 1130 13964 1186 13966
rect 890 13912 916 13964
rect 916 13912 946 13964
rect 970 13912 980 13964
rect 980 13912 1026 13964
rect 1050 13912 1096 13964
rect 1096 13912 1106 13964
rect 1130 13912 1160 13964
rect 1160 13912 1186 13964
rect 890 13910 946 13912
rect 970 13910 1026 13912
rect 1050 13910 1106 13912
rect 1130 13910 1186 13912
rect 890 12876 946 12878
rect 970 12876 1026 12878
rect 1050 12876 1106 12878
rect 1130 12876 1186 12878
rect 890 12824 916 12876
rect 916 12824 946 12876
rect 970 12824 980 12876
rect 980 12824 1026 12876
rect 1050 12824 1096 12876
rect 1096 12824 1106 12876
rect 1130 12824 1160 12876
rect 1160 12824 1186 12876
rect 890 12822 946 12824
rect 970 12822 1026 12824
rect 1050 12822 1106 12824
rect 1130 12822 1186 12824
rect 890 11788 946 11790
rect 970 11788 1026 11790
rect 1050 11788 1106 11790
rect 1130 11788 1186 11790
rect 890 11736 916 11788
rect 916 11736 946 11788
rect 970 11736 980 11788
rect 980 11736 1026 11788
rect 1050 11736 1096 11788
rect 1096 11736 1106 11788
rect 1130 11736 1160 11788
rect 1160 11736 1186 11788
rect 890 11734 946 11736
rect 970 11734 1026 11736
rect 1050 11734 1106 11736
rect 1130 11734 1186 11736
rect 890 10700 946 10702
rect 970 10700 1026 10702
rect 1050 10700 1106 10702
rect 1130 10700 1186 10702
rect 890 10648 916 10700
rect 916 10648 946 10700
rect 970 10648 980 10700
rect 980 10648 1026 10700
rect 1050 10648 1096 10700
rect 1096 10648 1106 10700
rect 1130 10648 1160 10700
rect 1160 10648 1186 10700
rect 890 10646 946 10648
rect 970 10646 1026 10648
rect 1050 10646 1106 10648
rect 1130 10646 1186 10648
rect 890 9612 946 9614
rect 970 9612 1026 9614
rect 1050 9612 1106 9614
rect 1130 9612 1186 9614
rect 890 9560 916 9612
rect 916 9560 946 9612
rect 970 9560 980 9612
rect 980 9560 1026 9612
rect 1050 9560 1096 9612
rect 1096 9560 1106 9612
rect 1130 9560 1160 9612
rect 1160 9560 1186 9612
rect 890 9558 946 9560
rect 970 9558 1026 9560
rect 1050 9558 1106 9560
rect 1130 9558 1186 9560
rect 890 8524 946 8526
rect 970 8524 1026 8526
rect 1050 8524 1106 8526
rect 1130 8524 1186 8526
rect 890 8472 916 8524
rect 916 8472 946 8524
rect 970 8472 980 8524
rect 980 8472 1026 8524
rect 1050 8472 1096 8524
rect 1096 8472 1106 8524
rect 1130 8472 1160 8524
rect 1160 8472 1186 8524
rect 890 8470 946 8472
rect 970 8470 1026 8472
rect 1050 8470 1106 8472
rect 1130 8470 1186 8472
rect 890 7436 946 7438
rect 970 7436 1026 7438
rect 1050 7436 1106 7438
rect 1130 7436 1186 7438
rect 890 7384 916 7436
rect 916 7384 946 7436
rect 970 7384 980 7436
rect 980 7384 1026 7436
rect 1050 7384 1096 7436
rect 1096 7384 1106 7436
rect 1130 7384 1160 7436
rect 1160 7384 1186 7436
rect 890 7382 946 7384
rect 970 7382 1026 7384
rect 1050 7382 1106 7384
rect 1130 7382 1186 7384
rect 890 6348 946 6350
rect 970 6348 1026 6350
rect 1050 6348 1106 6350
rect 1130 6348 1186 6350
rect 890 6296 916 6348
rect 916 6296 946 6348
rect 970 6296 980 6348
rect 980 6296 1026 6348
rect 1050 6296 1096 6348
rect 1096 6296 1106 6348
rect 1130 6296 1160 6348
rect 1160 6296 1186 6348
rect 890 6294 946 6296
rect 970 6294 1026 6296
rect 1050 6294 1106 6296
rect 1130 6294 1186 6296
rect 890 5260 946 5262
rect 970 5260 1026 5262
rect 1050 5260 1106 5262
rect 1130 5260 1186 5262
rect 890 5208 916 5260
rect 916 5208 946 5260
rect 970 5208 980 5260
rect 980 5208 1026 5260
rect 1050 5208 1096 5260
rect 1096 5208 1106 5260
rect 1130 5208 1160 5260
rect 1160 5208 1186 5260
rect 890 5206 946 5208
rect 970 5206 1026 5208
rect 1050 5206 1106 5208
rect 1130 5206 1186 5208
rect 1436 186698 1492 186754
rect 1896 171058 1952 171114
rect 890 4172 946 4174
rect 970 4172 1026 4174
rect 1050 4172 1106 4174
rect 1130 4172 1186 4174
rect 890 4120 916 4172
rect 916 4120 946 4172
rect 970 4120 980 4172
rect 980 4120 1026 4172
rect 1050 4120 1096 4172
rect 1096 4120 1106 4172
rect 1130 4120 1160 4172
rect 1160 4120 1186 4172
rect 890 4118 946 4120
rect 970 4118 1026 4120
rect 1050 4118 1106 4120
rect 1130 4118 1186 4120
rect 890 3084 946 3086
rect 970 3084 1026 3086
rect 1050 3084 1106 3086
rect 1130 3084 1186 3086
rect 890 3032 916 3084
rect 916 3032 946 3084
rect 970 3032 980 3084
rect 980 3032 1026 3084
rect 1050 3032 1096 3084
rect 1096 3032 1106 3084
rect 1130 3032 1160 3084
rect 1160 3032 1186 3084
rect 890 3030 946 3032
rect 970 3030 1026 3032
rect 1050 3030 1106 3032
rect 1130 3030 1186 3032
rect 1344 2826 1400 2882
rect 2264 171058 2320 171114
rect 2172 124718 2174 124738
rect 2174 124718 2226 124738
rect 2226 124718 2228 124738
rect 2172 124682 2228 124718
rect 2172 108090 2228 108146
rect 1804 3234 1860 3290
rect 2540 96938 2596 96994
rect 2890 187500 2946 187502
rect 2970 187500 3026 187502
rect 3050 187500 3106 187502
rect 3130 187500 3186 187502
rect 2890 187448 2916 187500
rect 2916 187448 2946 187500
rect 2970 187448 2980 187500
rect 2980 187448 3026 187500
rect 3050 187448 3096 187500
rect 3096 187448 3106 187500
rect 3130 187448 3160 187500
rect 3160 187448 3186 187500
rect 2890 187446 2946 187448
rect 2970 187446 3026 187448
rect 3050 187446 3106 187448
rect 3130 187446 3186 187448
rect 2890 186412 2946 186414
rect 2970 186412 3026 186414
rect 3050 186412 3106 186414
rect 3130 186412 3186 186414
rect 2890 186360 2916 186412
rect 2916 186360 2946 186412
rect 2970 186360 2980 186412
rect 2980 186360 3026 186412
rect 3050 186360 3096 186412
rect 3096 186360 3106 186412
rect 3130 186360 3160 186412
rect 3160 186360 3186 186412
rect 2890 186358 2946 186360
rect 2970 186358 3026 186360
rect 3050 186358 3106 186360
rect 3130 186358 3186 186360
rect 2890 185324 2946 185326
rect 2970 185324 3026 185326
rect 3050 185324 3106 185326
rect 3130 185324 3186 185326
rect 2890 185272 2916 185324
rect 2916 185272 2946 185324
rect 2970 185272 2980 185324
rect 2980 185272 3026 185324
rect 3050 185272 3096 185324
rect 3096 185272 3106 185324
rect 3130 185272 3160 185324
rect 3160 185272 3186 185324
rect 2890 185270 2946 185272
rect 2970 185270 3026 185272
rect 3050 185270 3106 185272
rect 3130 185270 3186 185272
rect 2890 184236 2946 184238
rect 2970 184236 3026 184238
rect 3050 184236 3106 184238
rect 3130 184236 3186 184238
rect 2890 184184 2916 184236
rect 2916 184184 2946 184236
rect 2970 184184 2980 184236
rect 2980 184184 3026 184236
rect 3050 184184 3096 184236
rect 3096 184184 3106 184236
rect 3130 184184 3160 184236
rect 3160 184184 3186 184236
rect 2890 184182 2946 184184
rect 2970 184182 3026 184184
rect 3050 184182 3106 184184
rect 3130 184182 3186 184184
rect 2890 183148 2946 183150
rect 2970 183148 3026 183150
rect 3050 183148 3106 183150
rect 3130 183148 3186 183150
rect 2890 183096 2916 183148
rect 2916 183096 2946 183148
rect 2970 183096 2980 183148
rect 2980 183096 3026 183148
rect 3050 183096 3096 183148
rect 3096 183096 3106 183148
rect 3130 183096 3160 183148
rect 3160 183096 3186 183148
rect 2890 183094 2946 183096
rect 2970 183094 3026 183096
rect 3050 183094 3106 183096
rect 3130 183094 3186 183096
rect 2890 182060 2946 182062
rect 2970 182060 3026 182062
rect 3050 182060 3106 182062
rect 3130 182060 3186 182062
rect 2890 182008 2916 182060
rect 2916 182008 2946 182060
rect 2970 182008 2980 182060
rect 2980 182008 3026 182060
rect 3050 182008 3096 182060
rect 3096 182008 3106 182060
rect 3130 182008 3160 182060
rect 3160 182008 3186 182060
rect 2890 182006 2946 182008
rect 2970 182006 3026 182008
rect 3050 182006 3106 182008
rect 3130 182006 3186 182008
rect 2890 180972 2946 180974
rect 2970 180972 3026 180974
rect 3050 180972 3106 180974
rect 3130 180972 3186 180974
rect 2890 180920 2916 180972
rect 2916 180920 2946 180972
rect 2970 180920 2980 180972
rect 2980 180920 3026 180972
rect 3050 180920 3096 180972
rect 3096 180920 3106 180972
rect 3130 180920 3160 180972
rect 3160 180920 3186 180972
rect 2890 180918 2946 180920
rect 2970 180918 3026 180920
rect 3050 180918 3106 180920
rect 3130 180918 3186 180920
rect 2890 179884 2946 179886
rect 2970 179884 3026 179886
rect 3050 179884 3106 179886
rect 3130 179884 3186 179886
rect 2890 179832 2916 179884
rect 2916 179832 2946 179884
rect 2970 179832 2980 179884
rect 2980 179832 3026 179884
rect 3050 179832 3096 179884
rect 3096 179832 3106 179884
rect 3130 179832 3160 179884
rect 3160 179832 3186 179884
rect 2890 179830 2946 179832
rect 2970 179830 3026 179832
rect 3050 179830 3106 179832
rect 3130 179830 3186 179832
rect 2890 178796 2946 178798
rect 2970 178796 3026 178798
rect 3050 178796 3106 178798
rect 3130 178796 3186 178798
rect 2890 178744 2916 178796
rect 2916 178744 2946 178796
rect 2970 178744 2980 178796
rect 2980 178744 3026 178796
rect 3050 178744 3096 178796
rect 3096 178744 3106 178796
rect 3130 178744 3160 178796
rect 3160 178744 3186 178796
rect 2890 178742 2946 178744
rect 2970 178742 3026 178744
rect 3050 178742 3106 178744
rect 3130 178742 3186 178744
rect 2890 177708 2946 177710
rect 2970 177708 3026 177710
rect 3050 177708 3106 177710
rect 3130 177708 3186 177710
rect 2890 177656 2916 177708
rect 2916 177656 2946 177708
rect 2970 177656 2980 177708
rect 2980 177656 3026 177708
rect 3050 177656 3096 177708
rect 3096 177656 3106 177708
rect 3130 177656 3160 177708
rect 3160 177656 3186 177708
rect 2890 177654 2946 177656
rect 2970 177654 3026 177656
rect 3050 177654 3106 177656
rect 3130 177654 3186 177656
rect 2890 176620 2946 176622
rect 2970 176620 3026 176622
rect 3050 176620 3106 176622
rect 3130 176620 3186 176622
rect 2890 176568 2916 176620
rect 2916 176568 2946 176620
rect 2970 176568 2980 176620
rect 2980 176568 3026 176620
rect 3050 176568 3096 176620
rect 3096 176568 3106 176620
rect 3130 176568 3160 176620
rect 3160 176568 3186 176620
rect 2890 176566 2946 176568
rect 2970 176566 3026 176568
rect 3050 176566 3106 176568
rect 3130 176566 3186 176568
rect 3276 175682 3332 175738
rect 2890 175532 2946 175534
rect 2970 175532 3026 175534
rect 3050 175532 3106 175534
rect 3130 175532 3186 175534
rect 2890 175480 2916 175532
rect 2916 175480 2946 175532
rect 2970 175480 2980 175532
rect 2980 175480 3026 175532
rect 3050 175480 3096 175532
rect 3096 175480 3106 175532
rect 3130 175480 3160 175532
rect 3160 175480 3186 175532
rect 2890 175478 2946 175480
rect 2970 175478 3026 175480
rect 3050 175478 3106 175480
rect 3130 175478 3186 175480
rect 2890 174444 2946 174446
rect 2970 174444 3026 174446
rect 3050 174444 3106 174446
rect 3130 174444 3186 174446
rect 2890 174392 2916 174444
rect 2916 174392 2946 174444
rect 2970 174392 2980 174444
rect 2980 174392 3026 174444
rect 3050 174392 3096 174444
rect 3096 174392 3106 174444
rect 3130 174392 3160 174444
rect 3160 174392 3186 174444
rect 2890 174390 2946 174392
rect 2970 174390 3026 174392
rect 3050 174390 3106 174392
rect 3130 174390 3186 174392
rect 2890 173356 2946 173358
rect 2970 173356 3026 173358
rect 3050 173356 3106 173358
rect 3130 173356 3186 173358
rect 2890 173304 2916 173356
rect 2916 173304 2946 173356
rect 2970 173304 2980 173356
rect 2980 173304 3026 173356
rect 3050 173304 3096 173356
rect 3096 173304 3106 173356
rect 3130 173304 3160 173356
rect 3160 173304 3186 173356
rect 2890 173302 2946 173304
rect 2970 173302 3026 173304
rect 3050 173302 3106 173304
rect 3130 173302 3186 173304
rect 2890 172268 2946 172270
rect 2970 172268 3026 172270
rect 3050 172268 3106 172270
rect 3130 172268 3186 172270
rect 2890 172216 2916 172268
rect 2916 172216 2946 172268
rect 2970 172216 2980 172268
rect 2980 172216 3026 172268
rect 3050 172216 3096 172268
rect 3096 172216 3106 172268
rect 3130 172216 3160 172268
rect 3160 172216 3186 172268
rect 2890 172214 2946 172216
rect 2970 172214 3026 172216
rect 3050 172214 3106 172216
rect 3130 172214 3186 172216
rect 2890 171180 2946 171182
rect 2970 171180 3026 171182
rect 3050 171180 3106 171182
rect 3130 171180 3186 171182
rect 2890 171128 2916 171180
rect 2916 171128 2946 171180
rect 2970 171128 2980 171180
rect 2980 171128 3026 171180
rect 3050 171128 3096 171180
rect 3096 171128 3106 171180
rect 3130 171128 3160 171180
rect 3160 171128 3186 171180
rect 2890 171126 2946 171128
rect 2970 171126 3026 171128
rect 3050 171126 3106 171128
rect 3130 171126 3186 171128
rect 2890 170092 2946 170094
rect 2970 170092 3026 170094
rect 3050 170092 3106 170094
rect 3130 170092 3186 170094
rect 2890 170040 2916 170092
rect 2916 170040 2946 170092
rect 2970 170040 2980 170092
rect 2980 170040 3026 170092
rect 3050 170040 3096 170092
rect 3096 170040 3106 170092
rect 3130 170040 3160 170092
rect 3160 170040 3186 170092
rect 2890 170038 2946 170040
rect 2970 170038 3026 170040
rect 3050 170038 3106 170040
rect 3130 170038 3186 170040
rect 2890 169004 2946 169006
rect 2970 169004 3026 169006
rect 3050 169004 3106 169006
rect 3130 169004 3186 169006
rect 2890 168952 2916 169004
rect 2916 168952 2946 169004
rect 2970 168952 2980 169004
rect 2980 168952 3026 169004
rect 3050 168952 3096 169004
rect 3096 168952 3106 169004
rect 3130 168952 3160 169004
rect 3160 168952 3186 169004
rect 2890 168950 2946 168952
rect 2970 168950 3026 168952
rect 3050 168950 3106 168952
rect 3130 168950 3186 168952
rect 2890 167916 2946 167918
rect 2970 167916 3026 167918
rect 3050 167916 3106 167918
rect 3130 167916 3186 167918
rect 2890 167864 2916 167916
rect 2916 167864 2946 167916
rect 2970 167864 2980 167916
rect 2980 167864 3026 167916
rect 3050 167864 3096 167916
rect 3096 167864 3106 167916
rect 3130 167864 3160 167916
rect 3160 167864 3186 167916
rect 2890 167862 2946 167864
rect 2970 167862 3026 167864
rect 3050 167862 3106 167864
rect 3130 167862 3186 167864
rect 2890 166828 2946 166830
rect 2970 166828 3026 166830
rect 3050 166828 3106 166830
rect 3130 166828 3186 166830
rect 2890 166776 2916 166828
rect 2916 166776 2946 166828
rect 2970 166776 2980 166828
rect 2980 166776 3026 166828
rect 3050 166776 3096 166828
rect 3096 166776 3106 166828
rect 3130 166776 3160 166828
rect 3160 166776 3186 166828
rect 2890 166774 2946 166776
rect 2970 166774 3026 166776
rect 3050 166774 3106 166776
rect 3130 166774 3186 166776
rect 2890 165740 2946 165742
rect 2970 165740 3026 165742
rect 3050 165740 3106 165742
rect 3130 165740 3186 165742
rect 2890 165688 2916 165740
rect 2916 165688 2946 165740
rect 2970 165688 2980 165740
rect 2980 165688 3026 165740
rect 3050 165688 3096 165740
rect 3096 165688 3106 165740
rect 3130 165688 3160 165740
rect 3160 165688 3186 165740
rect 2890 165686 2946 165688
rect 2970 165686 3026 165688
rect 3050 165686 3106 165688
rect 3130 165686 3186 165688
rect 2890 164652 2946 164654
rect 2970 164652 3026 164654
rect 3050 164652 3106 164654
rect 3130 164652 3186 164654
rect 2890 164600 2916 164652
rect 2916 164600 2946 164652
rect 2970 164600 2980 164652
rect 2980 164600 3026 164652
rect 3050 164600 3096 164652
rect 3096 164600 3106 164652
rect 3130 164600 3160 164652
rect 3160 164600 3186 164652
rect 2890 164598 2946 164600
rect 2970 164598 3026 164600
rect 3050 164598 3106 164600
rect 3130 164598 3186 164600
rect 2890 163564 2946 163566
rect 2970 163564 3026 163566
rect 3050 163564 3106 163566
rect 3130 163564 3186 163566
rect 2890 163512 2916 163564
rect 2916 163512 2946 163564
rect 2970 163512 2980 163564
rect 2980 163512 3026 163564
rect 3050 163512 3096 163564
rect 3096 163512 3106 163564
rect 3130 163512 3160 163564
rect 3160 163512 3186 163564
rect 2890 163510 2946 163512
rect 2970 163510 3026 163512
rect 3050 163510 3106 163512
rect 3130 163510 3186 163512
rect 2890 162476 2946 162478
rect 2970 162476 3026 162478
rect 3050 162476 3106 162478
rect 3130 162476 3186 162478
rect 2890 162424 2916 162476
rect 2916 162424 2946 162476
rect 2970 162424 2980 162476
rect 2980 162424 3026 162476
rect 3050 162424 3096 162476
rect 3096 162424 3106 162476
rect 3130 162424 3160 162476
rect 3160 162424 3186 162476
rect 2890 162422 2946 162424
rect 2970 162422 3026 162424
rect 3050 162422 3106 162424
rect 3130 162422 3186 162424
rect 2890 161388 2946 161390
rect 2970 161388 3026 161390
rect 3050 161388 3106 161390
rect 3130 161388 3186 161390
rect 2890 161336 2916 161388
rect 2916 161336 2946 161388
rect 2970 161336 2980 161388
rect 2980 161336 3026 161388
rect 3050 161336 3096 161388
rect 3096 161336 3106 161388
rect 3130 161336 3160 161388
rect 3160 161336 3186 161388
rect 2890 161334 2946 161336
rect 2970 161334 3026 161336
rect 3050 161334 3106 161336
rect 3130 161334 3186 161336
rect 2890 160300 2946 160302
rect 2970 160300 3026 160302
rect 3050 160300 3106 160302
rect 3130 160300 3186 160302
rect 2890 160248 2916 160300
rect 2916 160248 2946 160300
rect 2970 160248 2980 160300
rect 2980 160248 3026 160300
rect 3050 160248 3096 160300
rect 3096 160248 3106 160300
rect 3130 160248 3160 160300
rect 3160 160248 3186 160300
rect 2890 160246 2946 160248
rect 2970 160246 3026 160248
rect 3050 160246 3106 160248
rect 3130 160246 3186 160248
rect 2890 159212 2946 159214
rect 2970 159212 3026 159214
rect 3050 159212 3106 159214
rect 3130 159212 3186 159214
rect 2890 159160 2916 159212
rect 2916 159160 2946 159212
rect 2970 159160 2980 159212
rect 2980 159160 3026 159212
rect 3050 159160 3096 159212
rect 3096 159160 3106 159212
rect 3130 159160 3160 159212
rect 3160 159160 3186 159212
rect 2890 159158 2946 159160
rect 2970 159158 3026 159160
rect 3050 159158 3106 159160
rect 3130 159158 3186 159160
rect 2890 158124 2946 158126
rect 2970 158124 3026 158126
rect 3050 158124 3106 158126
rect 3130 158124 3186 158126
rect 2890 158072 2916 158124
rect 2916 158072 2946 158124
rect 2970 158072 2980 158124
rect 2980 158072 3026 158124
rect 3050 158072 3096 158124
rect 3096 158072 3106 158124
rect 3130 158072 3160 158124
rect 3160 158072 3186 158124
rect 2890 158070 2946 158072
rect 2970 158070 3026 158072
rect 3050 158070 3106 158072
rect 3130 158070 3186 158072
rect 2890 157036 2946 157038
rect 2970 157036 3026 157038
rect 3050 157036 3106 157038
rect 3130 157036 3186 157038
rect 2890 156984 2916 157036
rect 2916 156984 2946 157036
rect 2970 156984 2980 157036
rect 2980 156984 3026 157036
rect 3050 156984 3096 157036
rect 3096 156984 3106 157036
rect 3130 156984 3160 157036
rect 3160 156984 3186 157036
rect 2890 156982 2946 156984
rect 2970 156982 3026 156984
rect 3050 156982 3106 156984
rect 3130 156982 3186 156984
rect 2890 155948 2946 155950
rect 2970 155948 3026 155950
rect 3050 155948 3106 155950
rect 3130 155948 3186 155950
rect 2890 155896 2916 155948
rect 2916 155896 2946 155948
rect 2970 155896 2980 155948
rect 2980 155896 3026 155948
rect 3050 155896 3096 155948
rect 3096 155896 3106 155948
rect 3130 155896 3160 155948
rect 3160 155896 3186 155948
rect 2890 155894 2946 155896
rect 2970 155894 3026 155896
rect 3050 155894 3106 155896
rect 3130 155894 3186 155896
rect 2890 154860 2946 154862
rect 2970 154860 3026 154862
rect 3050 154860 3106 154862
rect 3130 154860 3186 154862
rect 2890 154808 2916 154860
rect 2916 154808 2946 154860
rect 2970 154808 2980 154860
rect 2980 154808 3026 154860
rect 3050 154808 3096 154860
rect 3096 154808 3106 154860
rect 3130 154808 3160 154860
rect 3160 154808 3186 154860
rect 2890 154806 2946 154808
rect 2970 154806 3026 154808
rect 3050 154806 3106 154808
rect 3130 154806 3186 154808
rect 2890 153772 2946 153774
rect 2970 153772 3026 153774
rect 3050 153772 3106 153774
rect 3130 153772 3186 153774
rect 2890 153720 2916 153772
rect 2916 153720 2946 153772
rect 2970 153720 2980 153772
rect 2980 153720 3026 153772
rect 3050 153720 3096 153772
rect 3096 153720 3106 153772
rect 3130 153720 3160 153772
rect 3160 153720 3186 153772
rect 2890 153718 2946 153720
rect 2970 153718 3026 153720
rect 3050 153718 3106 153720
rect 3130 153718 3186 153720
rect 2890 152684 2946 152686
rect 2970 152684 3026 152686
rect 3050 152684 3106 152686
rect 3130 152684 3186 152686
rect 2890 152632 2916 152684
rect 2916 152632 2946 152684
rect 2970 152632 2980 152684
rect 2980 152632 3026 152684
rect 3050 152632 3096 152684
rect 3096 152632 3106 152684
rect 3130 152632 3160 152684
rect 3160 152632 3186 152684
rect 2890 152630 2946 152632
rect 2970 152630 3026 152632
rect 3050 152630 3106 152632
rect 3130 152630 3186 152632
rect 2890 151596 2946 151598
rect 2970 151596 3026 151598
rect 3050 151596 3106 151598
rect 3130 151596 3186 151598
rect 2890 151544 2916 151596
rect 2916 151544 2946 151596
rect 2970 151544 2980 151596
rect 2980 151544 3026 151596
rect 3050 151544 3096 151596
rect 3096 151544 3106 151596
rect 3130 151544 3160 151596
rect 3160 151544 3186 151596
rect 2890 151542 2946 151544
rect 2970 151542 3026 151544
rect 3050 151542 3106 151544
rect 3130 151542 3186 151544
rect 2890 150508 2946 150510
rect 2970 150508 3026 150510
rect 3050 150508 3106 150510
rect 3130 150508 3186 150510
rect 2890 150456 2916 150508
rect 2916 150456 2946 150508
rect 2970 150456 2980 150508
rect 2980 150456 3026 150508
rect 3050 150456 3096 150508
rect 3096 150456 3106 150508
rect 3130 150456 3160 150508
rect 3160 150456 3186 150508
rect 2890 150454 2946 150456
rect 2970 150454 3026 150456
rect 3050 150454 3106 150456
rect 3130 150454 3186 150456
rect 2890 149420 2946 149422
rect 2970 149420 3026 149422
rect 3050 149420 3106 149422
rect 3130 149420 3186 149422
rect 2890 149368 2916 149420
rect 2916 149368 2946 149420
rect 2970 149368 2980 149420
rect 2980 149368 3026 149420
rect 3050 149368 3096 149420
rect 3096 149368 3106 149420
rect 3130 149368 3160 149420
rect 3160 149368 3186 149420
rect 2890 149366 2946 149368
rect 2970 149366 3026 149368
rect 3050 149366 3106 149368
rect 3130 149366 3186 149368
rect 2890 148332 2946 148334
rect 2970 148332 3026 148334
rect 3050 148332 3106 148334
rect 3130 148332 3186 148334
rect 2890 148280 2916 148332
rect 2916 148280 2946 148332
rect 2970 148280 2980 148332
rect 2980 148280 3026 148332
rect 3050 148280 3096 148332
rect 3096 148280 3106 148332
rect 3130 148280 3160 148332
rect 3160 148280 3186 148332
rect 2890 148278 2946 148280
rect 2970 148278 3026 148280
rect 3050 148278 3106 148280
rect 3130 148278 3186 148280
rect 2890 147244 2946 147246
rect 2970 147244 3026 147246
rect 3050 147244 3106 147246
rect 3130 147244 3186 147246
rect 2890 147192 2916 147244
rect 2916 147192 2946 147244
rect 2970 147192 2980 147244
rect 2980 147192 3026 147244
rect 3050 147192 3096 147244
rect 3096 147192 3106 147244
rect 3130 147192 3160 147244
rect 3160 147192 3186 147244
rect 2890 147190 2946 147192
rect 2970 147190 3026 147192
rect 3050 147190 3106 147192
rect 3130 147190 3186 147192
rect 2890 146156 2946 146158
rect 2970 146156 3026 146158
rect 3050 146156 3106 146158
rect 3130 146156 3186 146158
rect 2890 146104 2916 146156
rect 2916 146104 2946 146156
rect 2970 146104 2980 146156
rect 2980 146104 3026 146156
rect 3050 146104 3096 146156
rect 3096 146104 3106 146156
rect 3130 146104 3160 146156
rect 3160 146104 3186 146156
rect 2890 146102 2946 146104
rect 2970 146102 3026 146104
rect 3050 146102 3106 146104
rect 3130 146102 3186 146104
rect 2890 145068 2946 145070
rect 2970 145068 3026 145070
rect 3050 145068 3106 145070
rect 3130 145068 3186 145070
rect 2890 145016 2916 145068
rect 2916 145016 2946 145068
rect 2970 145016 2980 145068
rect 2980 145016 3026 145068
rect 3050 145016 3096 145068
rect 3096 145016 3106 145068
rect 3130 145016 3160 145068
rect 3160 145016 3186 145068
rect 2890 145014 2946 145016
rect 2970 145014 3026 145016
rect 3050 145014 3106 145016
rect 3130 145014 3186 145016
rect 2890 143980 2946 143982
rect 2970 143980 3026 143982
rect 3050 143980 3106 143982
rect 3130 143980 3186 143982
rect 2890 143928 2916 143980
rect 2916 143928 2946 143980
rect 2970 143928 2980 143980
rect 2980 143928 3026 143980
rect 3050 143928 3096 143980
rect 3096 143928 3106 143980
rect 3130 143928 3160 143980
rect 3160 143928 3186 143980
rect 2890 143926 2946 143928
rect 2970 143926 3026 143928
rect 3050 143926 3106 143928
rect 3130 143926 3186 143928
rect 2890 142892 2946 142894
rect 2970 142892 3026 142894
rect 3050 142892 3106 142894
rect 3130 142892 3186 142894
rect 2890 142840 2916 142892
rect 2916 142840 2946 142892
rect 2970 142840 2980 142892
rect 2980 142840 3026 142892
rect 3050 142840 3096 142892
rect 3096 142840 3106 142892
rect 3130 142840 3160 142892
rect 3160 142840 3186 142892
rect 2890 142838 2946 142840
rect 2970 142838 3026 142840
rect 3050 142838 3106 142840
rect 3130 142838 3186 142840
rect 2890 141804 2946 141806
rect 2970 141804 3026 141806
rect 3050 141804 3106 141806
rect 3130 141804 3186 141806
rect 2890 141752 2916 141804
rect 2916 141752 2946 141804
rect 2970 141752 2980 141804
rect 2980 141752 3026 141804
rect 3050 141752 3096 141804
rect 3096 141752 3106 141804
rect 3130 141752 3160 141804
rect 3160 141752 3186 141804
rect 2890 141750 2946 141752
rect 2970 141750 3026 141752
rect 3050 141750 3106 141752
rect 3130 141750 3186 141752
rect 2890 140716 2946 140718
rect 2970 140716 3026 140718
rect 3050 140716 3106 140718
rect 3130 140716 3186 140718
rect 2890 140664 2916 140716
rect 2916 140664 2946 140716
rect 2970 140664 2980 140716
rect 2980 140664 3026 140716
rect 3050 140664 3096 140716
rect 3096 140664 3106 140716
rect 3130 140664 3160 140716
rect 3160 140664 3186 140716
rect 2890 140662 2946 140664
rect 2970 140662 3026 140664
rect 3050 140662 3106 140664
rect 3130 140662 3186 140664
rect 2890 139628 2946 139630
rect 2970 139628 3026 139630
rect 3050 139628 3106 139630
rect 3130 139628 3186 139630
rect 2890 139576 2916 139628
rect 2916 139576 2946 139628
rect 2970 139576 2980 139628
rect 2980 139576 3026 139628
rect 3050 139576 3096 139628
rect 3096 139576 3106 139628
rect 3130 139576 3160 139628
rect 3160 139576 3186 139628
rect 2890 139574 2946 139576
rect 2970 139574 3026 139576
rect 3050 139574 3106 139576
rect 3130 139574 3186 139576
rect 2890 138540 2946 138542
rect 2970 138540 3026 138542
rect 3050 138540 3106 138542
rect 3130 138540 3186 138542
rect 2890 138488 2916 138540
rect 2916 138488 2946 138540
rect 2970 138488 2980 138540
rect 2980 138488 3026 138540
rect 3050 138488 3096 138540
rect 3096 138488 3106 138540
rect 3130 138488 3160 138540
rect 3160 138488 3186 138540
rect 2890 138486 2946 138488
rect 2970 138486 3026 138488
rect 3050 138486 3106 138488
rect 3130 138486 3186 138488
rect 2890 137452 2946 137454
rect 2970 137452 3026 137454
rect 3050 137452 3106 137454
rect 3130 137452 3186 137454
rect 2890 137400 2916 137452
rect 2916 137400 2946 137452
rect 2970 137400 2980 137452
rect 2980 137400 3026 137452
rect 3050 137400 3096 137452
rect 3096 137400 3106 137452
rect 3130 137400 3160 137452
rect 3160 137400 3186 137452
rect 2890 137398 2946 137400
rect 2970 137398 3026 137400
rect 3050 137398 3106 137400
rect 3130 137398 3186 137400
rect 2890 136364 2946 136366
rect 2970 136364 3026 136366
rect 3050 136364 3106 136366
rect 3130 136364 3186 136366
rect 2890 136312 2916 136364
rect 2916 136312 2946 136364
rect 2970 136312 2980 136364
rect 2980 136312 3026 136364
rect 3050 136312 3096 136364
rect 3096 136312 3106 136364
rect 3130 136312 3160 136364
rect 3160 136312 3186 136364
rect 2890 136310 2946 136312
rect 2970 136310 3026 136312
rect 3050 136310 3106 136312
rect 3130 136310 3186 136312
rect 2890 135276 2946 135278
rect 2970 135276 3026 135278
rect 3050 135276 3106 135278
rect 3130 135276 3186 135278
rect 2890 135224 2916 135276
rect 2916 135224 2946 135276
rect 2970 135224 2980 135276
rect 2980 135224 3026 135276
rect 3050 135224 3096 135276
rect 3096 135224 3106 135276
rect 3130 135224 3160 135276
rect 3160 135224 3186 135276
rect 2890 135222 2946 135224
rect 2970 135222 3026 135224
rect 3050 135222 3106 135224
rect 3130 135222 3186 135224
rect 2890 134188 2946 134190
rect 2970 134188 3026 134190
rect 3050 134188 3106 134190
rect 3130 134188 3186 134190
rect 2890 134136 2916 134188
rect 2916 134136 2946 134188
rect 2970 134136 2980 134188
rect 2980 134136 3026 134188
rect 3050 134136 3096 134188
rect 3096 134136 3106 134188
rect 3130 134136 3160 134188
rect 3160 134136 3186 134188
rect 2890 134134 2946 134136
rect 2970 134134 3026 134136
rect 3050 134134 3106 134136
rect 3130 134134 3186 134136
rect 2890 133100 2946 133102
rect 2970 133100 3026 133102
rect 3050 133100 3106 133102
rect 3130 133100 3186 133102
rect 2890 133048 2916 133100
rect 2916 133048 2946 133100
rect 2970 133048 2980 133100
rect 2980 133048 3026 133100
rect 3050 133048 3096 133100
rect 3096 133048 3106 133100
rect 3130 133048 3160 133100
rect 3160 133048 3186 133100
rect 2890 133046 2946 133048
rect 2970 133046 3026 133048
rect 3050 133046 3106 133048
rect 3130 133046 3186 133048
rect 2890 132012 2946 132014
rect 2970 132012 3026 132014
rect 3050 132012 3106 132014
rect 3130 132012 3186 132014
rect 2890 131960 2916 132012
rect 2916 131960 2946 132012
rect 2970 131960 2980 132012
rect 2980 131960 3026 132012
rect 3050 131960 3096 132012
rect 3096 131960 3106 132012
rect 3130 131960 3160 132012
rect 3160 131960 3186 132012
rect 2890 131958 2946 131960
rect 2970 131958 3026 131960
rect 3050 131958 3106 131960
rect 3130 131958 3186 131960
rect 2890 130924 2946 130926
rect 2970 130924 3026 130926
rect 3050 130924 3106 130926
rect 3130 130924 3186 130926
rect 2890 130872 2916 130924
rect 2916 130872 2946 130924
rect 2970 130872 2980 130924
rect 2980 130872 3026 130924
rect 3050 130872 3096 130924
rect 3096 130872 3106 130924
rect 3130 130872 3160 130924
rect 3160 130872 3186 130924
rect 2890 130870 2946 130872
rect 2970 130870 3026 130872
rect 3050 130870 3106 130872
rect 3130 130870 3186 130872
rect 2890 129836 2946 129838
rect 2970 129836 3026 129838
rect 3050 129836 3106 129838
rect 3130 129836 3186 129838
rect 2890 129784 2916 129836
rect 2916 129784 2946 129836
rect 2970 129784 2980 129836
rect 2980 129784 3026 129836
rect 3050 129784 3096 129836
rect 3096 129784 3106 129836
rect 3130 129784 3160 129836
rect 3160 129784 3186 129836
rect 2890 129782 2946 129784
rect 2970 129782 3026 129784
rect 3050 129782 3106 129784
rect 3130 129782 3186 129784
rect 2890 128748 2946 128750
rect 2970 128748 3026 128750
rect 3050 128748 3106 128750
rect 3130 128748 3186 128750
rect 2890 128696 2916 128748
rect 2916 128696 2946 128748
rect 2970 128696 2980 128748
rect 2980 128696 3026 128748
rect 3050 128696 3096 128748
rect 3096 128696 3106 128748
rect 3130 128696 3160 128748
rect 3160 128696 3186 128748
rect 2890 128694 2946 128696
rect 2970 128694 3026 128696
rect 3050 128694 3106 128696
rect 3130 128694 3186 128696
rect 2890 127660 2946 127662
rect 2970 127660 3026 127662
rect 3050 127660 3106 127662
rect 3130 127660 3186 127662
rect 2890 127608 2916 127660
rect 2916 127608 2946 127660
rect 2970 127608 2980 127660
rect 2980 127608 3026 127660
rect 3050 127608 3096 127660
rect 3096 127608 3106 127660
rect 3130 127608 3160 127660
rect 3160 127608 3186 127660
rect 2890 127606 2946 127608
rect 2970 127606 3026 127608
rect 3050 127606 3106 127608
rect 3130 127606 3186 127608
rect 2890 126572 2946 126574
rect 2970 126572 3026 126574
rect 3050 126572 3106 126574
rect 3130 126572 3186 126574
rect 2890 126520 2916 126572
rect 2916 126520 2946 126572
rect 2970 126520 2980 126572
rect 2980 126520 3026 126572
rect 3050 126520 3096 126572
rect 3096 126520 3106 126572
rect 3130 126520 3160 126572
rect 3160 126520 3186 126572
rect 2890 126518 2946 126520
rect 2970 126518 3026 126520
rect 3050 126518 3106 126520
rect 3130 126518 3186 126520
rect 2890 125484 2946 125486
rect 2970 125484 3026 125486
rect 3050 125484 3106 125486
rect 3130 125484 3186 125486
rect 2890 125432 2916 125484
rect 2916 125432 2946 125484
rect 2970 125432 2980 125484
rect 2980 125432 3026 125484
rect 3050 125432 3096 125484
rect 3096 125432 3106 125484
rect 3130 125432 3160 125484
rect 3160 125432 3186 125484
rect 2890 125430 2946 125432
rect 2970 125430 3026 125432
rect 3050 125430 3106 125432
rect 3130 125430 3186 125432
rect 2890 124396 2946 124398
rect 2970 124396 3026 124398
rect 3050 124396 3106 124398
rect 3130 124396 3186 124398
rect 2890 124344 2916 124396
rect 2916 124344 2946 124396
rect 2970 124344 2980 124396
rect 2980 124344 3026 124396
rect 3050 124344 3096 124396
rect 3096 124344 3106 124396
rect 3130 124344 3160 124396
rect 3160 124344 3186 124396
rect 2890 124342 2946 124344
rect 2970 124342 3026 124344
rect 3050 124342 3106 124344
rect 3130 124342 3186 124344
rect 2890 123308 2946 123310
rect 2970 123308 3026 123310
rect 3050 123308 3106 123310
rect 3130 123308 3186 123310
rect 2890 123256 2916 123308
rect 2916 123256 2946 123308
rect 2970 123256 2980 123308
rect 2980 123256 3026 123308
rect 3050 123256 3096 123308
rect 3096 123256 3106 123308
rect 3130 123256 3160 123308
rect 3160 123256 3186 123308
rect 2890 123254 2946 123256
rect 2970 123254 3026 123256
rect 3050 123254 3106 123256
rect 3130 123254 3186 123256
rect 2890 122220 2946 122222
rect 2970 122220 3026 122222
rect 3050 122220 3106 122222
rect 3130 122220 3186 122222
rect 2890 122168 2916 122220
rect 2916 122168 2946 122220
rect 2970 122168 2980 122220
rect 2980 122168 3026 122220
rect 3050 122168 3096 122220
rect 3096 122168 3106 122220
rect 3130 122168 3160 122220
rect 3160 122168 3186 122220
rect 2890 122166 2946 122168
rect 2970 122166 3026 122168
rect 3050 122166 3106 122168
rect 3130 122166 3186 122168
rect 2890 121132 2946 121134
rect 2970 121132 3026 121134
rect 3050 121132 3106 121134
rect 3130 121132 3186 121134
rect 2890 121080 2916 121132
rect 2916 121080 2946 121132
rect 2970 121080 2980 121132
rect 2980 121080 3026 121132
rect 3050 121080 3096 121132
rect 3096 121080 3106 121132
rect 3130 121080 3160 121132
rect 3160 121080 3186 121132
rect 2890 121078 2946 121080
rect 2970 121078 3026 121080
rect 3050 121078 3106 121080
rect 3130 121078 3186 121080
rect 2890 120044 2946 120046
rect 2970 120044 3026 120046
rect 3050 120044 3106 120046
rect 3130 120044 3186 120046
rect 2890 119992 2916 120044
rect 2916 119992 2946 120044
rect 2970 119992 2980 120044
rect 2980 119992 3026 120044
rect 3050 119992 3096 120044
rect 3096 119992 3106 120044
rect 3130 119992 3160 120044
rect 3160 119992 3186 120044
rect 2890 119990 2946 119992
rect 2970 119990 3026 119992
rect 3050 119990 3106 119992
rect 3130 119990 3186 119992
rect 2890 118956 2946 118958
rect 2970 118956 3026 118958
rect 3050 118956 3106 118958
rect 3130 118956 3186 118958
rect 2890 118904 2916 118956
rect 2916 118904 2946 118956
rect 2970 118904 2980 118956
rect 2980 118904 3026 118956
rect 3050 118904 3096 118956
rect 3096 118904 3106 118956
rect 3130 118904 3160 118956
rect 3160 118904 3186 118956
rect 2890 118902 2946 118904
rect 2970 118902 3026 118904
rect 3050 118902 3106 118904
rect 3130 118902 3186 118904
rect 2890 117868 2946 117870
rect 2970 117868 3026 117870
rect 3050 117868 3106 117870
rect 3130 117868 3186 117870
rect 2890 117816 2916 117868
rect 2916 117816 2946 117868
rect 2970 117816 2980 117868
rect 2980 117816 3026 117868
rect 3050 117816 3096 117868
rect 3096 117816 3106 117868
rect 3130 117816 3160 117868
rect 3160 117816 3186 117868
rect 2890 117814 2946 117816
rect 2970 117814 3026 117816
rect 3050 117814 3106 117816
rect 3130 117814 3186 117816
rect 2890 116780 2946 116782
rect 2970 116780 3026 116782
rect 3050 116780 3106 116782
rect 3130 116780 3186 116782
rect 2890 116728 2916 116780
rect 2916 116728 2946 116780
rect 2970 116728 2980 116780
rect 2980 116728 3026 116780
rect 3050 116728 3096 116780
rect 3096 116728 3106 116780
rect 3130 116728 3160 116780
rect 3160 116728 3186 116780
rect 2890 116726 2946 116728
rect 2970 116726 3026 116728
rect 3050 116726 3106 116728
rect 3130 116726 3186 116728
rect 2890 115692 2946 115694
rect 2970 115692 3026 115694
rect 3050 115692 3106 115694
rect 3130 115692 3186 115694
rect 2890 115640 2916 115692
rect 2916 115640 2946 115692
rect 2970 115640 2980 115692
rect 2980 115640 3026 115692
rect 3050 115640 3096 115692
rect 3096 115640 3106 115692
rect 3130 115640 3160 115692
rect 3160 115640 3186 115692
rect 2890 115638 2946 115640
rect 2970 115638 3026 115640
rect 3050 115638 3106 115640
rect 3130 115638 3186 115640
rect 2890 114604 2946 114606
rect 2970 114604 3026 114606
rect 3050 114604 3106 114606
rect 3130 114604 3186 114606
rect 2890 114552 2916 114604
rect 2916 114552 2946 114604
rect 2970 114552 2980 114604
rect 2980 114552 3026 114604
rect 3050 114552 3096 114604
rect 3096 114552 3106 114604
rect 3130 114552 3160 114604
rect 3160 114552 3186 114604
rect 2890 114550 2946 114552
rect 2970 114550 3026 114552
rect 3050 114550 3106 114552
rect 3130 114550 3186 114552
rect 2890 113516 2946 113518
rect 2970 113516 3026 113518
rect 3050 113516 3106 113518
rect 3130 113516 3186 113518
rect 2890 113464 2916 113516
rect 2916 113464 2946 113516
rect 2970 113464 2980 113516
rect 2980 113464 3026 113516
rect 3050 113464 3096 113516
rect 3096 113464 3106 113516
rect 3130 113464 3160 113516
rect 3160 113464 3186 113516
rect 2890 113462 2946 113464
rect 2970 113462 3026 113464
rect 3050 113462 3106 113464
rect 3130 113462 3186 113464
rect 2890 112428 2946 112430
rect 2970 112428 3026 112430
rect 3050 112428 3106 112430
rect 3130 112428 3186 112430
rect 2890 112376 2916 112428
rect 2916 112376 2946 112428
rect 2970 112376 2980 112428
rect 2980 112376 3026 112428
rect 3050 112376 3096 112428
rect 3096 112376 3106 112428
rect 3130 112376 3160 112428
rect 3160 112376 3186 112428
rect 2890 112374 2946 112376
rect 2970 112374 3026 112376
rect 3050 112374 3106 112376
rect 3130 112374 3186 112376
rect 2890 111340 2946 111342
rect 2970 111340 3026 111342
rect 3050 111340 3106 111342
rect 3130 111340 3186 111342
rect 2890 111288 2916 111340
rect 2916 111288 2946 111340
rect 2970 111288 2980 111340
rect 2980 111288 3026 111340
rect 3050 111288 3096 111340
rect 3096 111288 3106 111340
rect 3130 111288 3160 111340
rect 3160 111288 3186 111340
rect 2890 111286 2946 111288
rect 2970 111286 3026 111288
rect 3050 111286 3106 111288
rect 3130 111286 3186 111288
rect 2890 110252 2946 110254
rect 2970 110252 3026 110254
rect 3050 110252 3106 110254
rect 3130 110252 3186 110254
rect 2890 110200 2916 110252
rect 2916 110200 2946 110252
rect 2970 110200 2980 110252
rect 2980 110200 3026 110252
rect 3050 110200 3096 110252
rect 3096 110200 3106 110252
rect 3130 110200 3160 110252
rect 3160 110200 3186 110252
rect 2890 110198 2946 110200
rect 2970 110198 3026 110200
rect 3050 110198 3106 110200
rect 3130 110198 3186 110200
rect 2890 109164 2946 109166
rect 2970 109164 3026 109166
rect 3050 109164 3106 109166
rect 3130 109164 3186 109166
rect 2890 109112 2916 109164
rect 2916 109112 2946 109164
rect 2970 109112 2980 109164
rect 2980 109112 3026 109164
rect 3050 109112 3096 109164
rect 3096 109112 3106 109164
rect 3130 109112 3160 109164
rect 3160 109112 3186 109164
rect 2890 109110 2946 109112
rect 2970 109110 3026 109112
rect 3050 109110 3106 109112
rect 3130 109110 3186 109112
rect 2890 108076 2946 108078
rect 2970 108076 3026 108078
rect 3050 108076 3106 108078
rect 3130 108076 3186 108078
rect 2890 108024 2916 108076
rect 2916 108024 2946 108076
rect 2970 108024 2980 108076
rect 2980 108024 3026 108076
rect 3050 108024 3096 108076
rect 3096 108024 3106 108076
rect 3130 108024 3160 108076
rect 3160 108024 3186 108076
rect 2890 108022 2946 108024
rect 2970 108022 3026 108024
rect 3050 108022 3106 108024
rect 3130 108022 3186 108024
rect 2890 106988 2946 106990
rect 2970 106988 3026 106990
rect 3050 106988 3106 106990
rect 3130 106988 3186 106990
rect 2890 106936 2916 106988
rect 2916 106936 2946 106988
rect 2970 106936 2980 106988
rect 2980 106936 3026 106988
rect 3050 106936 3096 106988
rect 3096 106936 3106 106988
rect 3130 106936 3160 106988
rect 3160 106936 3186 106988
rect 2890 106934 2946 106936
rect 2970 106934 3026 106936
rect 3050 106934 3106 106936
rect 3130 106934 3186 106936
rect 2890 105900 2946 105902
rect 2970 105900 3026 105902
rect 3050 105900 3106 105902
rect 3130 105900 3186 105902
rect 2890 105848 2916 105900
rect 2916 105848 2946 105900
rect 2970 105848 2980 105900
rect 2980 105848 3026 105900
rect 3050 105848 3096 105900
rect 3096 105848 3106 105900
rect 3130 105848 3160 105900
rect 3160 105848 3186 105900
rect 2890 105846 2946 105848
rect 2970 105846 3026 105848
rect 3050 105846 3106 105848
rect 3130 105846 3186 105848
rect 2890 104812 2946 104814
rect 2970 104812 3026 104814
rect 3050 104812 3106 104814
rect 3130 104812 3186 104814
rect 2890 104760 2916 104812
rect 2916 104760 2946 104812
rect 2970 104760 2980 104812
rect 2980 104760 3026 104812
rect 3050 104760 3096 104812
rect 3096 104760 3106 104812
rect 3130 104760 3160 104812
rect 3160 104760 3186 104812
rect 2890 104758 2946 104760
rect 2970 104758 3026 104760
rect 3050 104758 3106 104760
rect 3130 104758 3186 104760
rect 2890 103724 2946 103726
rect 2970 103724 3026 103726
rect 3050 103724 3106 103726
rect 3130 103724 3186 103726
rect 2890 103672 2916 103724
rect 2916 103672 2946 103724
rect 2970 103672 2980 103724
rect 2980 103672 3026 103724
rect 3050 103672 3096 103724
rect 3096 103672 3106 103724
rect 3130 103672 3160 103724
rect 3160 103672 3186 103724
rect 2890 103670 2946 103672
rect 2970 103670 3026 103672
rect 3050 103670 3106 103672
rect 3130 103670 3186 103672
rect 2890 102636 2946 102638
rect 2970 102636 3026 102638
rect 3050 102636 3106 102638
rect 3130 102636 3186 102638
rect 2890 102584 2916 102636
rect 2916 102584 2946 102636
rect 2970 102584 2980 102636
rect 2980 102584 3026 102636
rect 3050 102584 3096 102636
rect 3096 102584 3106 102636
rect 3130 102584 3160 102636
rect 3160 102584 3186 102636
rect 2890 102582 2946 102584
rect 2970 102582 3026 102584
rect 3050 102582 3106 102584
rect 3130 102582 3186 102584
rect 2890 101548 2946 101550
rect 2970 101548 3026 101550
rect 3050 101548 3106 101550
rect 3130 101548 3186 101550
rect 2890 101496 2916 101548
rect 2916 101496 2946 101548
rect 2970 101496 2980 101548
rect 2980 101496 3026 101548
rect 3050 101496 3096 101548
rect 3096 101496 3106 101548
rect 3130 101496 3160 101548
rect 3160 101496 3186 101548
rect 2890 101494 2946 101496
rect 2970 101494 3026 101496
rect 3050 101494 3106 101496
rect 3130 101494 3186 101496
rect 2890 100460 2946 100462
rect 2970 100460 3026 100462
rect 3050 100460 3106 100462
rect 3130 100460 3186 100462
rect 2890 100408 2916 100460
rect 2916 100408 2946 100460
rect 2970 100408 2980 100460
rect 2980 100408 3026 100460
rect 3050 100408 3096 100460
rect 3096 100408 3106 100460
rect 3130 100408 3160 100460
rect 3160 100408 3186 100460
rect 2890 100406 2946 100408
rect 2970 100406 3026 100408
rect 3050 100406 3106 100408
rect 3130 100406 3186 100408
rect 2890 99372 2946 99374
rect 2970 99372 3026 99374
rect 3050 99372 3106 99374
rect 3130 99372 3186 99374
rect 2890 99320 2916 99372
rect 2916 99320 2946 99372
rect 2970 99320 2980 99372
rect 2980 99320 3026 99372
rect 3050 99320 3096 99372
rect 3096 99320 3106 99372
rect 3130 99320 3160 99372
rect 3160 99320 3186 99372
rect 2890 99318 2946 99320
rect 2970 99318 3026 99320
rect 3050 99318 3106 99320
rect 3130 99318 3186 99320
rect 2890 98284 2946 98286
rect 2970 98284 3026 98286
rect 3050 98284 3106 98286
rect 3130 98284 3186 98286
rect 2890 98232 2916 98284
rect 2916 98232 2946 98284
rect 2970 98232 2980 98284
rect 2980 98232 3026 98284
rect 3050 98232 3096 98284
rect 3096 98232 3106 98284
rect 3130 98232 3160 98284
rect 3160 98232 3186 98284
rect 2890 98230 2946 98232
rect 2970 98230 3026 98232
rect 3050 98230 3106 98232
rect 3130 98230 3186 98232
rect 890 1996 946 1998
rect 970 1996 1026 1998
rect 1050 1996 1106 1998
rect 1130 1996 1186 1998
rect 890 1944 916 1996
rect 916 1944 946 1996
rect 970 1944 980 1996
rect 980 1944 1026 1996
rect 1050 1944 1096 1996
rect 1096 1944 1106 1996
rect 1130 1944 1160 1996
rect 1160 1944 1186 1996
rect 890 1942 946 1944
rect 970 1942 1026 1944
rect 1050 1942 1106 1944
rect 1130 1942 1186 1944
rect 2890 97196 2946 97198
rect 2970 97196 3026 97198
rect 3050 97196 3106 97198
rect 3130 97196 3186 97198
rect 2890 97144 2916 97196
rect 2916 97144 2946 97196
rect 2970 97144 2980 97196
rect 2980 97144 3026 97196
rect 3050 97144 3096 97196
rect 3096 97144 3106 97196
rect 3130 97144 3160 97196
rect 3160 97144 3186 97196
rect 2890 97142 2946 97144
rect 2970 97142 3026 97144
rect 3050 97142 3106 97144
rect 3130 97142 3186 97144
rect 3000 96702 3002 96722
rect 3002 96702 3054 96722
rect 3054 96702 3056 96722
rect 3000 96666 3056 96702
rect 3184 96294 3186 96314
rect 3186 96294 3238 96314
rect 3238 96294 3240 96314
rect 3184 96258 3240 96294
rect 2890 96108 2946 96110
rect 2970 96108 3026 96110
rect 3050 96108 3106 96110
rect 3130 96108 3186 96110
rect 2890 96056 2916 96108
rect 2916 96056 2946 96108
rect 2970 96056 2980 96108
rect 2980 96056 3026 96108
rect 3050 96056 3096 96108
rect 3096 96056 3106 96108
rect 3130 96056 3160 96108
rect 3160 96056 3186 96108
rect 2890 96054 2946 96056
rect 2970 96054 3026 96056
rect 3050 96054 3106 96056
rect 3130 96054 3186 96056
rect 2890 95020 2946 95022
rect 2970 95020 3026 95022
rect 3050 95020 3106 95022
rect 3130 95020 3186 95022
rect 2890 94968 2916 95020
rect 2916 94968 2946 95020
rect 2970 94968 2980 95020
rect 2980 94968 3026 95020
rect 3050 94968 3096 95020
rect 3096 94968 3106 95020
rect 3130 94968 3160 95020
rect 3160 94968 3186 95020
rect 2890 94966 2946 94968
rect 2970 94966 3026 94968
rect 3050 94966 3106 94968
rect 3130 94966 3186 94968
rect 2890 93932 2946 93934
rect 2970 93932 3026 93934
rect 3050 93932 3106 93934
rect 3130 93932 3186 93934
rect 2890 93880 2916 93932
rect 2916 93880 2946 93932
rect 2970 93880 2980 93932
rect 2980 93880 3026 93932
rect 3050 93880 3096 93932
rect 3096 93880 3106 93932
rect 3130 93880 3160 93932
rect 3160 93880 3186 93932
rect 2890 93878 2946 93880
rect 2970 93878 3026 93880
rect 3050 93878 3106 93880
rect 3130 93878 3186 93880
rect 2890 92844 2946 92846
rect 2970 92844 3026 92846
rect 3050 92844 3106 92846
rect 3130 92844 3186 92846
rect 2890 92792 2916 92844
rect 2916 92792 2946 92844
rect 2970 92792 2980 92844
rect 2980 92792 3026 92844
rect 3050 92792 3096 92844
rect 3096 92792 3106 92844
rect 3130 92792 3160 92844
rect 3160 92792 3186 92844
rect 2890 92790 2946 92792
rect 2970 92790 3026 92792
rect 3050 92790 3106 92792
rect 3130 92790 3186 92792
rect 2890 91756 2946 91758
rect 2970 91756 3026 91758
rect 3050 91756 3106 91758
rect 3130 91756 3186 91758
rect 2890 91704 2916 91756
rect 2916 91704 2946 91756
rect 2970 91704 2980 91756
rect 2980 91704 3026 91756
rect 3050 91704 3096 91756
rect 3096 91704 3106 91756
rect 3130 91704 3160 91756
rect 3160 91704 3186 91756
rect 2890 91702 2946 91704
rect 2970 91702 3026 91704
rect 3050 91702 3106 91704
rect 3130 91702 3186 91704
rect 2890 90668 2946 90670
rect 2970 90668 3026 90670
rect 3050 90668 3106 90670
rect 3130 90668 3186 90670
rect 2890 90616 2916 90668
rect 2916 90616 2946 90668
rect 2970 90616 2980 90668
rect 2980 90616 3026 90668
rect 3050 90616 3096 90668
rect 3096 90616 3106 90668
rect 3130 90616 3160 90668
rect 3160 90616 3186 90668
rect 2890 90614 2946 90616
rect 2970 90614 3026 90616
rect 3050 90614 3106 90616
rect 3130 90614 3186 90616
rect 2890 89580 2946 89582
rect 2970 89580 3026 89582
rect 3050 89580 3106 89582
rect 3130 89580 3186 89582
rect 2890 89528 2916 89580
rect 2916 89528 2946 89580
rect 2970 89528 2980 89580
rect 2980 89528 3026 89580
rect 3050 89528 3096 89580
rect 3096 89528 3106 89580
rect 3130 89528 3160 89580
rect 3160 89528 3186 89580
rect 2890 89526 2946 89528
rect 2970 89526 3026 89528
rect 3050 89526 3106 89528
rect 3130 89526 3186 89528
rect 2448 2962 2504 3018
rect 2890 88492 2946 88494
rect 2970 88492 3026 88494
rect 3050 88492 3106 88494
rect 3130 88492 3186 88494
rect 2890 88440 2916 88492
rect 2916 88440 2946 88492
rect 2970 88440 2980 88492
rect 2980 88440 3026 88492
rect 3050 88440 3096 88492
rect 3096 88440 3106 88492
rect 3130 88440 3160 88492
rect 3160 88440 3186 88492
rect 2890 88438 2946 88440
rect 2970 88438 3026 88440
rect 3050 88438 3106 88440
rect 3130 88438 3186 88440
rect 2890 87404 2946 87406
rect 2970 87404 3026 87406
rect 3050 87404 3106 87406
rect 3130 87404 3186 87406
rect 2890 87352 2916 87404
rect 2916 87352 2946 87404
rect 2970 87352 2980 87404
rect 2980 87352 3026 87404
rect 3050 87352 3096 87404
rect 3096 87352 3106 87404
rect 3130 87352 3160 87404
rect 3160 87352 3186 87404
rect 2890 87350 2946 87352
rect 2970 87350 3026 87352
rect 3050 87350 3106 87352
rect 3130 87350 3186 87352
rect 2890 86316 2946 86318
rect 2970 86316 3026 86318
rect 3050 86316 3106 86318
rect 3130 86316 3186 86318
rect 2890 86264 2916 86316
rect 2916 86264 2946 86316
rect 2970 86264 2980 86316
rect 2980 86264 3026 86316
rect 3050 86264 3096 86316
rect 3096 86264 3106 86316
rect 3130 86264 3160 86316
rect 3160 86264 3186 86316
rect 2890 86262 2946 86264
rect 2970 86262 3026 86264
rect 3050 86262 3106 86264
rect 3130 86262 3186 86264
rect 2890 85228 2946 85230
rect 2970 85228 3026 85230
rect 3050 85228 3106 85230
rect 3130 85228 3186 85230
rect 2890 85176 2916 85228
rect 2916 85176 2946 85228
rect 2970 85176 2980 85228
rect 2980 85176 3026 85228
rect 3050 85176 3096 85228
rect 3096 85176 3106 85228
rect 3130 85176 3160 85228
rect 3160 85176 3186 85228
rect 2890 85174 2946 85176
rect 2970 85174 3026 85176
rect 3050 85174 3106 85176
rect 3130 85174 3186 85176
rect 2890 84140 2946 84142
rect 2970 84140 3026 84142
rect 3050 84140 3106 84142
rect 3130 84140 3186 84142
rect 2890 84088 2916 84140
rect 2916 84088 2946 84140
rect 2970 84088 2980 84140
rect 2980 84088 3026 84140
rect 3050 84088 3096 84140
rect 3096 84088 3106 84140
rect 3130 84088 3160 84140
rect 3160 84088 3186 84140
rect 2890 84086 2946 84088
rect 2970 84086 3026 84088
rect 3050 84086 3106 84088
rect 3130 84086 3186 84088
rect 2890 83052 2946 83054
rect 2970 83052 3026 83054
rect 3050 83052 3106 83054
rect 3130 83052 3186 83054
rect 2890 83000 2916 83052
rect 2916 83000 2946 83052
rect 2970 83000 2980 83052
rect 2980 83000 3026 83052
rect 3050 83000 3096 83052
rect 3096 83000 3106 83052
rect 3130 83000 3160 83052
rect 3160 83000 3186 83052
rect 2890 82998 2946 83000
rect 2970 82998 3026 83000
rect 3050 82998 3106 83000
rect 3130 82998 3186 83000
rect 3920 182774 3976 182810
rect 3920 182754 3922 182774
rect 3922 182754 3974 182774
rect 3974 182754 3976 182774
rect 3552 181686 3608 181722
rect 3552 181666 3554 181686
rect 3554 181666 3606 181686
rect 3606 181666 3608 181686
rect 3552 179898 3608 179954
rect 3644 176770 3700 176826
rect 3644 174050 3700 174106
rect 3460 114774 3516 114810
rect 3460 114754 3462 114774
rect 3462 114754 3514 114774
rect 3514 114754 3516 114774
rect 3276 81978 3332 82034
rect 2890 81964 2946 81966
rect 2970 81964 3026 81966
rect 3050 81964 3106 81966
rect 3130 81964 3186 81966
rect 2890 81912 2916 81964
rect 2916 81912 2946 81964
rect 2970 81912 2980 81964
rect 2980 81912 3026 81964
rect 3050 81912 3096 81964
rect 3096 81912 3106 81964
rect 3130 81912 3160 81964
rect 3160 81912 3186 81964
rect 2890 81910 2946 81912
rect 2970 81910 3026 81912
rect 3050 81910 3106 81912
rect 3130 81910 3186 81912
rect 2890 80876 2946 80878
rect 2970 80876 3026 80878
rect 3050 80876 3106 80878
rect 3130 80876 3186 80878
rect 2890 80824 2916 80876
rect 2916 80824 2946 80876
rect 2970 80824 2980 80876
rect 2980 80824 3026 80876
rect 3050 80824 3096 80876
rect 3096 80824 3106 80876
rect 3130 80824 3160 80876
rect 3160 80824 3186 80876
rect 2890 80822 2946 80824
rect 2970 80822 3026 80824
rect 3050 80822 3106 80824
rect 3130 80822 3186 80824
rect 2890 79788 2946 79790
rect 2970 79788 3026 79790
rect 3050 79788 3106 79790
rect 3130 79788 3186 79790
rect 2890 79736 2916 79788
rect 2916 79736 2946 79788
rect 2970 79736 2980 79788
rect 2980 79736 3026 79788
rect 3050 79736 3096 79788
rect 3096 79736 3106 79788
rect 3130 79736 3160 79788
rect 3160 79736 3186 79788
rect 2890 79734 2946 79736
rect 2970 79734 3026 79736
rect 3050 79734 3106 79736
rect 3130 79734 3186 79736
rect 2890 78700 2946 78702
rect 2970 78700 3026 78702
rect 3050 78700 3106 78702
rect 3130 78700 3186 78702
rect 2890 78648 2916 78700
rect 2916 78648 2946 78700
rect 2970 78648 2980 78700
rect 2980 78648 3026 78700
rect 3050 78648 3096 78700
rect 3096 78648 3106 78700
rect 3130 78648 3160 78700
rect 3160 78648 3186 78700
rect 2890 78646 2946 78648
rect 2970 78646 3026 78648
rect 3050 78646 3106 78648
rect 3130 78646 3186 78648
rect 2890 77612 2946 77614
rect 2970 77612 3026 77614
rect 3050 77612 3106 77614
rect 3130 77612 3186 77614
rect 2890 77560 2916 77612
rect 2916 77560 2946 77612
rect 2970 77560 2980 77612
rect 2980 77560 3026 77612
rect 3050 77560 3096 77612
rect 3096 77560 3106 77612
rect 3130 77560 3160 77612
rect 3160 77560 3186 77612
rect 2890 77558 2946 77560
rect 2970 77558 3026 77560
rect 3050 77558 3106 77560
rect 3130 77558 3186 77560
rect 2890 76524 2946 76526
rect 2970 76524 3026 76526
rect 3050 76524 3106 76526
rect 3130 76524 3186 76526
rect 2890 76472 2916 76524
rect 2916 76472 2946 76524
rect 2970 76472 2980 76524
rect 2980 76472 3026 76524
rect 3050 76472 3096 76524
rect 3096 76472 3106 76524
rect 3130 76472 3160 76524
rect 3160 76472 3186 76524
rect 2890 76470 2946 76472
rect 2970 76470 3026 76472
rect 3050 76470 3106 76472
rect 3130 76470 3186 76472
rect 2890 75436 2946 75438
rect 2970 75436 3026 75438
rect 3050 75436 3106 75438
rect 3130 75436 3186 75438
rect 2890 75384 2916 75436
rect 2916 75384 2946 75436
rect 2970 75384 2980 75436
rect 2980 75384 3026 75436
rect 3050 75384 3096 75436
rect 3096 75384 3106 75436
rect 3130 75384 3160 75436
rect 3160 75384 3186 75436
rect 2890 75382 2946 75384
rect 2970 75382 3026 75384
rect 3050 75382 3106 75384
rect 3130 75382 3186 75384
rect 2890 74348 2946 74350
rect 2970 74348 3026 74350
rect 3050 74348 3106 74350
rect 3130 74348 3186 74350
rect 2890 74296 2916 74348
rect 2916 74296 2946 74348
rect 2970 74296 2980 74348
rect 2980 74296 3026 74348
rect 3050 74296 3096 74348
rect 3096 74296 3106 74348
rect 3130 74296 3160 74348
rect 3160 74296 3186 74348
rect 2890 74294 2946 74296
rect 2970 74294 3026 74296
rect 3050 74294 3106 74296
rect 3130 74294 3186 74296
rect 2890 73260 2946 73262
rect 2970 73260 3026 73262
rect 3050 73260 3106 73262
rect 3130 73260 3186 73262
rect 2890 73208 2916 73260
rect 2916 73208 2946 73260
rect 2970 73208 2980 73260
rect 2980 73208 3026 73260
rect 3050 73208 3096 73260
rect 3096 73208 3106 73260
rect 3130 73208 3160 73260
rect 3160 73208 3186 73260
rect 2890 73206 2946 73208
rect 2970 73206 3026 73208
rect 3050 73206 3106 73208
rect 3130 73206 3186 73208
rect 2890 72172 2946 72174
rect 2970 72172 3026 72174
rect 3050 72172 3106 72174
rect 3130 72172 3186 72174
rect 2890 72120 2916 72172
rect 2916 72120 2946 72172
rect 2970 72120 2980 72172
rect 2980 72120 3026 72172
rect 3050 72120 3096 72172
rect 3096 72120 3106 72172
rect 3130 72120 3160 72172
rect 3160 72120 3186 72172
rect 2890 72118 2946 72120
rect 2970 72118 3026 72120
rect 3050 72118 3106 72120
rect 3130 72118 3186 72120
rect 2890 71084 2946 71086
rect 2970 71084 3026 71086
rect 3050 71084 3106 71086
rect 3130 71084 3186 71086
rect 2890 71032 2916 71084
rect 2916 71032 2946 71084
rect 2970 71032 2980 71084
rect 2980 71032 3026 71084
rect 3050 71032 3096 71084
rect 3096 71032 3106 71084
rect 3130 71032 3160 71084
rect 3160 71032 3186 71084
rect 2890 71030 2946 71032
rect 2970 71030 3026 71032
rect 3050 71030 3106 71032
rect 3130 71030 3186 71032
rect 2890 69996 2946 69998
rect 2970 69996 3026 69998
rect 3050 69996 3106 69998
rect 3130 69996 3186 69998
rect 2890 69944 2916 69996
rect 2916 69944 2946 69996
rect 2970 69944 2980 69996
rect 2980 69944 3026 69996
rect 3050 69944 3096 69996
rect 3096 69944 3106 69996
rect 3130 69944 3160 69996
rect 3160 69944 3186 69996
rect 2890 69942 2946 69944
rect 2970 69942 3026 69944
rect 3050 69942 3106 69944
rect 3130 69942 3186 69944
rect 2890 68908 2946 68910
rect 2970 68908 3026 68910
rect 3050 68908 3106 68910
rect 3130 68908 3186 68910
rect 2890 68856 2916 68908
rect 2916 68856 2946 68908
rect 2970 68856 2980 68908
rect 2980 68856 3026 68908
rect 3050 68856 3096 68908
rect 3096 68856 3106 68908
rect 3130 68856 3160 68908
rect 3160 68856 3186 68908
rect 2890 68854 2946 68856
rect 2970 68854 3026 68856
rect 3050 68854 3106 68856
rect 3130 68854 3186 68856
rect 2890 67820 2946 67822
rect 2970 67820 3026 67822
rect 3050 67820 3106 67822
rect 3130 67820 3186 67822
rect 2890 67768 2916 67820
rect 2916 67768 2946 67820
rect 2970 67768 2980 67820
rect 2980 67768 3026 67820
rect 3050 67768 3096 67820
rect 3096 67768 3106 67820
rect 3130 67768 3160 67820
rect 3160 67768 3186 67820
rect 2890 67766 2946 67768
rect 2970 67766 3026 67768
rect 3050 67766 3106 67768
rect 3130 67766 3186 67768
rect 2890 66732 2946 66734
rect 2970 66732 3026 66734
rect 3050 66732 3106 66734
rect 3130 66732 3186 66734
rect 2890 66680 2916 66732
rect 2916 66680 2946 66732
rect 2970 66680 2980 66732
rect 2980 66680 3026 66732
rect 3050 66680 3096 66732
rect 3096 66680 3106 66732
rect 3130 66680 3160 66732
rect 3160 66680 3186 66732
rect 2890 66678 2946 66680
rect 2970 66678 3026 66680
rect 3050 66678 3106 66680
rect 3130 66678 3186 66680
rect 2890 65644 2946 65646
rect 2970 65644 3026 65646
rect 3050 65644 3106 65646
rect 3130 65644 3186 65646
rect 2890 65592 2916 65644
rect 2916 65592 2946 65644
rect 2970 65592 2980 65644
rect 2980 65592 3026 65644
rect 3050 65592 3096 65644
rect 3096 65592 3106 65644
rect 3130 65592 3160 65644
rect 3160 65592 3186 65644
rect 2890 65590 2946 65592
rect 2970 65590 3026 65592
rect 3050 65590 3106 65592
rect 3130 65590 3186 65592
rect 2890 64556 2946 64558
rect 2970 64556 3026 64558
rect 3050 64556 3106 64558
rect 3130 64556 3186 64558
rect 2890 64504 2916 64556
rect 2916 64504 2946 64556
rect 2970 64504 2980 64556
rect 2980 64504 3026 64556
rect 3050 64504 3096 64556
rect 3096 64504 3106 64556
rect 3130 64504 3160 64556
rect 3160 64504 3186 64556
rect 2890 64502 2946 64504
rect 2970 64502 3026 64504
rect 3050 64502 3106 64504
rect 3130 64502 3186 64504
rect 2890 63468 2946 63470
rect 2970 63468 3026 63470
rect 3050 63468 3106 63470
rect 3130 63468 3186 63470
rect 2890 63416 2916 63468
rect 2916 63416 2946 63468
rect 2970 63416 2980 63468
rect 2980 63416 3026 63468
rect 3050 63416 3096 63468
rect 3096 63416 3106 63468
rect 3130 63416 3160 63468
rect 3160 63416 3186 63468
rect 2890 63414 2946 63416
rect 2970 63414 3026 63416
rect 3050 63414 3106 63416
rect 3130 63414 3186 63416
rect 2890 62380 2946 62382
rect 2970 62380 3026 62382
rect 3050 62380 3106 62382
rect 3130 62380 3186 62382
rect 2890 62328 2916 62380
rect 2916 62328 2946 62380
rect 2970 62328 2980 62380
rect 2980 62328 3026 62380
rect 3050 62328 3096 62380
rect 3096 62328 3106 62380
rect 3130 62328 3160 62380
rect 3160 62328 3186 62380
rect 2890 62326 2946 62328
rect 2970 62326 3026 62328
rect 3050 62326 3106 62328
rect 3130 62326 3186 62328
rect 2890 61292 2946 61294
rect 2970 61292 3026 61294
rect 3050 61292 3106 61294
rect 3130 61292 3186 61294
rect 2890 61240 2916 61292
rect 2916 61240 2946 61292
rect 2970 61240 2980 61292
rect 2980 61240 3026 61292
rect 3050 61240 3096 61292
rect 3096 61240 3106 61292
rect 3130 61240 3160 61292
rect 3160 61240 3186 61292
rect 2890 61238 2946 61240
rect 2970 61238 3026 61240
rect 3050 61238 3106 61240
rect 3130 61238 3186 61240
rect 2890 60204 2946 60206
rect 2970 60204 3026 60206
rect 3050 60204 3106 60206
rect 3130 60204 3186 60206
rect 2890 60152 2916 60204
rect 2916 60152 2946 60204
rect 2970 60152 2980 60204
rect 2980 60152 3026 60204
rect 3050 60152 3096 60204
rect 3096 60152 3106 60204
rect 3130 60152 3160 60204
rect 3160 60152 3186 60204
rect 2890 60150 2946 60152
rect 2970 60150 3026 60152
rect 3050 60150 3106 60152
rect 3130 60150 3186 60152
rect 2890 59116 2946 59118
rect 2970 59116 3026 59118
rect 3050 59116 3106 59118
rect 3130 59116 3186 59118
rect 2890 59064 2916 59116
rect 2916 59064 2946 59116
rect 2970 59064 2980 59116
rect 2980 59064 3026 59116
rect 3050 59064 3096 59116
rect 3096 59064 3106 59116
rect 3130 59064 3160 59116
rect 3160 59064 3186 59116
rect 2890 59062 2946 59064
rect 2970 59062 3026 59064
rect 3050 59062 3106 59064
rect 3130 59062 3186 59064
rect 2890 58028 2946 58030
rect 2970 58028 3026 58030
rect 3050 58028 3106 58030
rect 3130 58028 3186 58030
rect 2890 57976 2916 58028
rect 2916 57976 2946 58028
rect 2970 57976 2980 58028
rect 2980 57976 3026 58028
rect 3050 57976 3096 58028
rect 3096 57976 3106 58028
rect 3130 57976 3160 58028
rect 3160 57976 3186 58028
rect 2890 57974 2946 57976
rect 2970 57974 3026 57976
rect 3050 57974 3106 57976
rect 3130 57974 3186 57976
rect 2890 56940 2946 56942
rect 2970 56940 3026 56942
rect 3050 56940 3106 56942
rect 3130 56940 3186 56942
rect 2890 56888 2916 56940
rect 2916 56888 2946 56940
rect 2970 56888 2980 56940
rect 2980 56888 3026 56940
rect 3050 56888 3096 56940
rect 3096 56888 3106 56940
rect 3130 56888 3160 56940
rect 3160 56888 3186 56940
rect 2890 56886 2946 56888
rect 2970 56886 3026 56888
rect 3050 56886 3106 56888
rect 3130 56886 3186 56888
rect 2890 55852 2946 55854
rect 2970 55852 3026 55854
rect 3050 55852 3106 55854
rect 3130 55852 3186 55854
rect 2890 55800 2916 55852
rect 2916 55800 2946 55852
rect 2970 55800 2980 55852
rect 2980 55800 3026 55852
rect 3050 55800 3096 55852
rect 3096 55800 3106 55852
rect 3130 55800 3160 55852
rect 3160 55800 3186 55852
rect 2890 55798 2946 55800
rect 2970 55798 3026 55800
rect 3050 55798 3106 55800
rect 3130 55798 3186 55800
rect 2890 54764 2946 54766
rect 2970 54764 3026 54766
rect 3050 54764 3106 54766
rect 3130 54764 3186 54766
rect 2890 54712 2916 54764
rect 2916 54712 2946 54764
rect 2970 54712 2980 54764
rect 2980 54712 3026 54764
rect 3050 54712 3096 54764
rect 3096 54712 3106 54764
rect 3130 54712 3160 54764
rect 3160 54712 3186 54764
rect 2890 54710 2946 54712
rect 2970 54710 3026 54712
rect 3050 54710 3106 54712
rect 3130 54710 3186 54712
rect 2890 53676 2946 53678
rect 2970 53676 3026 53678
rect 3050 53676 3106 53678
rect 3130 53676 3186 53678
rect 2890 53624 2916 53676
rect 2916 53624 2946 53676
rect 2970 53624 2980 53676
rect 2980 53624 3026 53676
rect 3050 53624 3096 53676
rect 3096 53624 3106 53676
rect 3130 53624 3160 53676
rect 3160 53624 3186 53676
rect 2890 53622 2946 53624
rect 2970 53622 3026 53624
rect 3050 53622 3106 53624
rect 3130 53622 3186 53624
rect 2890 52588 2946 52590
rect 2970 52588 3026 52590
rect 3050 52588 3106 52590
rect 3130 52588 3186 52590
rect 2890 52536 2916 52588
rect 2916 52536 2946 52588
rect 2970 52536 2980 52588
rect 2980 52536 3026 52588
rect 3050 52536 3096 52588
rect 3096 52536 3106 52588
rect 3130 52536 3160 52588
rect 3160 52536 3186 52588
rect 2890 52534 2946 52536
rect 2970 52534 3026 52536
rect 3050 52534 3106 52536
rect 3130 52534 3186 52536
rect 2890 51500 2946 51502
rect 2970 51500 3026 51502
rect 3050 51500 3106 51502
rect 3130 51500 3186 51502
rect 2890 51448 2916 51500
rect 2916 51448 2946 51500
rect 2970 51448 2980 51500
rect 2980 51448 3026 51500
rect 3050 51448 3096 51500
rect 3096 51448 3106 51500
rect 3130 51448 3160 51500
rect 3160 51448 3186 51500
rect 2890 51446 2946 51448
rect 2970 51446 3026 51448
rect 3050 51446 3106 51448
rect 3130 51446 3186 51448
rect 2890 50412 2946 50414
rect 2970 50412 3026 50414
rect 3050 50412 3106 50414
rect 3130 50412 3186 50414
rect 2890 50360 2916 50412
rect 2916 50360 2946 50412
rect 2970 50360 2980 50412
rect 2980 50360 3026 50412
rect 3050 50360 3096 50412
rect 3096 50360 3106 50412
rect 3130 50360 3160 50412
rect 3160 50360 3186 50412
rect 2890 50358 2946 50360
rect 2970 50358 3026 50360
rect 3050 50358 3106 50360
rect 3130 50358 3186 50360
rect 2890 49324 2946 49326
rect 2970 49324 3026 49326
rect 3050 49324 3106 49326
rect 3130 49324 3186 49326
rect 2890 49272 2916 49324
rect 2916 49272 2946 49324
rect 2970 49272 2980 49324
rect 2980 49272 3026 49324
rect 3050 49272 3096 49324
rect 3096 49272 3106 49324
rect 3130 49272 3160 49324
rect 3160 49272 3186 49324
rect 2890 49270 2946 49272
rect 2970 49270 3026 49272
rect 3050 49270 3106 49272
rect 3130 49270 3186 49272
rect 2890 48236 2946 48238
rect 2970 48236 3026 48238
rect 3050 48236 3106 48238
rect 3130 48236 3186 48238
rect 2890 48184 2916 48236
rect 2916 48184 2946 48236
rect 2970 48184 2980 48236
rect 2980 48184 3026 48236
rect 3050 48184 3096 48236
rect 3096 48184 3106 48236
rect 3130 48184 3160 48236
rect 3160 48184 3186 48236
rect 2890 48182 2946 48184
rect 2970 48182 3026 48184
rect 3050 48182 3106 48184
rect 3130 48182 3186 48184
rect 2890 47148 2946 47150
rect 2970 47148 3026 47150
rect 3050 47148 3106 47150
rect 3130 47148 3186 47150
rect 2890 47096 2916 47148
rect 2916 47096 2946 47148
rect 2970 47096 2980 47148
rect 2980 47096 3026 47148
rect 3050 47096 3096 47148
rect 3096 47096 3106 47148
rect 3130 47096 3160 47148
rect 3160 47096 3186 47148
rect 2890 47094 2946 47096
rect 2970 47094 3026 47096
rect 3050 47094 3106 47096
rect 3130 47094 3186 47096
rect 2890 46060 2946 46062
rect 2970 46060 3026 46062
rect 3050 46060 3106 46062
rect 3130 46060 3186 46062
rect 2890 46008 2916 46060
rect 2916 46008 2946 46060
rect 2970 46008 2980 46060
rect 2980 46008 3026 46060
rect 3050 46008 3096 46060
rect 3096 46008 3106 46060
rect 3130 46008 3160 46060
rect 3160 46008 3186 46060
rect 2890 46006 2946 46008
rect 2970 46006 3026 46008
rect 3050 46006 3106 46008
rect 3130 46006 3186 46008
rect 2890 44972 2946 44974
rect 2970 44972 3026 44974
rect 3050 44972 3106 44974
rect 3130 44972 3186 44974
rect 2890 44920 2916 44972
rect 2916 44920 2946 44972
rect 2970 44920 2980 44972
rect 2980 44920 3026 44972
rect 3050 44920 3096 44972
rect 3096 44920 3106 44972
rect 3130 44920 3160 44972
rect 3160 44920 3186 44972
rect 2890 44918 2946 44920
rect 2970 44918 3026 44920
rect 3050 44918 3106 44920
rect 3130 44918 3186 44920
rect 2890 43884 2946 43886
rect 2970 43884 3026 43886
rect 3050 43884 3106 43886
rect 3130 43884 3186 43886
rect 2890 43832 2916 43884
rect 2916 43832 2946 43884
rect 2970 43832 2980 43884
rect 2980 43832 3026 43884
rect 3050 43832 3096 43884
rect 3096 43832 3106 43884
rect 3130 43832 3160 43884
rect 3160 43832 3186 43884
rect 2890 43830 2946 43832
rect 2970 43830 3026 43832
rect 3050 43830 3106 43832
rect 3130 43830 3186 43832
rect 2890 42796 2946 42798
rect 2970 42796 3026 42798
rect 3050 42796 3106 42798
rect 3130 42796 3186 42798
rect 2890 42744 2916 42796
rect 2916 42744 2946 42796
rect 2970 42744 2980 42796
rect 2980 42744 3026 42796
rect 3050 42744 3096 42796
rect 3096 42744 3106 42796
rect 3130 42744 3160 42796
rect 3160 42744 3186 42796
rect 2890 42742 2946 42744
rect 2970 42742 3026 42744
rect 3050 42742 3106 42744
rect 3130 42742 3186 42744
rect 2890 41708 2946 41710
rect 2970 41708 3026 41710
rect 3050 41708 3106 41710
rect 3130 41708 3186 41710
rect 2890 41656 2916 41708
rect 2916 41656 2946 41708
rect 2970 41656 2980 41708
rect 2980 41656 3026 41708
rect 3050 41656 3096 41708
rect 3096 41656 3106 41708
rect 3130 41656 3160 41708
rect 3160 41656 3186 41708
rect 2890 41654 2946 41656
rect 2970 41654 3026 41656
rect 3050 41654 3106 41656
rect 3130 41654 3186 41656
rect 2890 40620 2946 40622
rect 2970 40620 3026 40622
rect 3050 40620 3106 40622
rect 3130 40620 3186 40622
rect 2890 40568 2916 40620
rect 2916 40568 2946 40620
rect 2970 40568 2980 40620
rect 2980 40568 3026 40620
rect 3050 40568 3096 40620
rect 3096 40568 3106 40620
rect 3130 40568 3160 40620
rect 3160 40568 3186 40620
rect 2890 40566 2946 40568
rect 2970 40566 3026 40568
rect 3050 40566 3106 40568
rect 3130 40566 3186 40568
rect 2890 39532 2946 39534
rect 2970 39532 3026 39534
rect 3050 39532 3106 39534
rect 3130 39532 3186 39534
rect 2890 39480 2916 39532
rect 2916 39480 2946 39532
rect 2970 39480 2980 39532
rect 2980 39480 3026 39532
rect 3050 39480 3096 39532
rect 3096 39480 3106 39532
rect 3130 39480 3160 39532
rect 3160 39480 3186 39532
rect 2890 39478 2946 39480
rect 2970 39478 3026 39480
rect 3050 39478 3106 39480
rect 3130 39478 3186 39480
rect 2890 38444 2946 38446
rect 2970 38444 3026 38446
rect 3050 38444 3106 38446
rect 3130 38444 3186 38446
rect 2890 38392 2916 38444
rect 2916 38392 2946 38444
rect 2970 38392 2980 38444
rect 2980 38392 3026 38444
rect 3050 38392 3096 38444
rect 3096 38392 3106 38444
rect 3130 38392 3160 38444
rect 3160 38392 3186 38444
rect 2890 38390 2946 38392
rect 2970 38390 3026 38392
rect 3050 38390 3106 38392
rect 3130 38390 3186 38392
rect 2890 37356 2946 37358
rect 2970 37356 3026 37358
rect 3050 37356 3106 37358
rect 3130 37356 3186 37358
rect 2890 37304 2916 37356
rect 2916 37304 2946 37356
rect 2970 37304 2980 37356
rect 2980 37304 3026 37356
rect 3050 37304 3096 37356
rect 3096 37304 3106 37356
rect 3130 37304 3160 37356
rect 3160 37304 3186 37356
rect 2890 37302 2946 37304
rect 2970 37302 3026 37304
rect 3050 37302 3106 37304
rect 3130 37302 3186 37304
rect 2890 36268 2946 36270
rect 2970 36268 3026 36270
rect 3050 36268 3106 36270
rect 3130 36268 3186 36270
rect 2890 36216 2916 36268
rect 2916 36216 2946 36268
rect 2970 36216 2980 36268
rect 2980 36216 3026 36268
rect 3050 36216 3096 36268
rect 3096 36216 3106 36268
rect 3130 36216 3160 36268
rect 3160 36216 3186 36268
rect 2890 36214 2946 36216
rect 2970 36214 3026 36216
rect 3050 36214 3106 36216
rect 3130 36214 3186 36216
rect 2890 35180 2946 35182
rect 2970 35180 3026 35182
rect 3050 35180 3106 35182
rect 3130 35180 3186 35182
rect 2890 35128 2916 35180
rect 2916 35128 2946 35180
rect 2970 35128 2980 35180
rect 2980 35128 3026 35180
rect 3050 35128 3096 35180
rect 3096 35128 3106 35180
rect 3130 35128 3160 35180
rect 3160 35128 3186 35180
rect 2890 35126 2946 35128
rect 2970 35126 3026 35128
rect 3050 35126 3106 35128
rect 3130 35126 3186 35128
rect 3276 34514 3332 34570
rect 2890 34092 2946 34094
rect 2970 34092 3026 34094
rect 3050 34092 3106 34094
rect 3130 34092 3186 34094
rect 2890 34040 2916 34092
rect 2916 34040 2946 34092
rect 2970 34040 2980 34092
rect 2980 34040 3026 34092
rect 3050 34040 3096 34092
rect 3096 34040 3106 34092
rect 3130 34040 3160 34092
rect 3160 34040 3186 34092
rect 2890 34038 2946 34040
rect 2970 34038 3026 34040
rect 3050 34038 3106 34040
rect 3130 34038 3186 34040
rect 2890 33004 2946 33006
rect 2970 33004 3026 33006
rect 3050 33004 3106 33006
rect 3130 33004 3186 33006
rect 2890 32952 2916 33004
rect 2916 32952 2946 33004
rect 2970 32952 2980 33004
rect 2980 32952 3026 33004
rect 3050 32952 3096 33004
rect 3096 32952 3106 33004
rect 3130 32952 3160 33004
rect 3160 32952 3186 33004
rect 2890 32950 2946 32952
rect 2970 32950 3026 32952
rect 3050 32950 3106 32952
rect 3130 32950 3186 32952
rect 2890 31916 2946 31918
rect 2970 31916 3026 31918
rect 3050 31916 3106 31918
rect 3130 31916 3186 31918
rect 2890 31864 2916 31916
rect 2916 31864 2946 31916
rect 2970 31864 2980 31916
rect 2980 31864 3026 31916
rect 3050 31864 3096 31916
rect 3096 31864 3106 31916
rect 3130 31864 3160 31916
rect 3160 31864 3186 31916
rect 2890 31862 2946 31864
rect 2970 31862 3026 31864
rect 3050 31862 3106 31864
rect 3130 31862 3186 31864
rect 2890 30828 2946 30830
rect 2970 30828 3026 30830
rect 3050 30828 3106 30830
rect 3130 30828 3186 30830
rect 2890 30776 2916 30828
rect 2916 30776 2946 30828
rect 2970 30776 2980 30828
rect 2980 30776 3026 30828
rect 3050 30776 3096 30828
rect 3096 30776 3106 30828
rect 3130 30776 3160 30828
rect 3160 30776 3186 30828
rect 2890 30774 2946 30776
rect 2970 30774 3026 30776
rect 3050 30774 3106 30776
rect 3130 30774 3186 30776
rect 2890 29740 2946 29742
rect 2970 29740 3026 29742
rect 3050 29740 3106 29742
rect 3130 29740 3186 29742
rect 2890 29688 2916 29740
rect 2916 29688 2946 29740
rect 2970 29688 2980 29740
rect 2980 29688 3026 29740
rect 3050 29688 3096 29740
rect 3096 29688 3106 29740
rect 3130 29688 3160 29740
rect 3160 29688 3186 29740
rect 2890 29686 2946 29688
rect 2970 29686 3026 29688
rect 3050 29686 3106 29688
rect 3130 29686 3186 29688
rect 2890 28652 2946 28654
rect 2970 28652 3026 28654
rect 3050 28652 3106 28654
rect 3130 28652 3186 28654
rect 2890 28600 2916 28652
rect 2916 28600 2946 28652
rect 2970 28600 2980 28652
rect 2980 28600 3026 28652
rect 3050 28600 3096 28652
rect 3096 28600 3106 28652
rect 3130 28600 3160 28652
rect 3160 28600 3186 28652
rect 2890 28598 2946 28600
rect 2970 28598 3026 28600
rect 3050 28598 3106 28600
rect 3130 28598 3186 28600
rect 2890 27564 2946 27566
rect 2970 27564 3026 27566
rect 3050 27564 3106 27566
rect 3130 27564 3186 27566
rect 2890 27512 2916 27564
rect 2916 27512 2946 27564
rect 2970 27512 2980 27564
rect 2980 27512 3026 27564
rect 3050 27512 3096 27564
rect 3096 27512 3106 27564
rect 3130 27512 3160 27564
rect 3160 27512 3186 27564
rect 2890 27510 2946 27512
rect 2970 27510 3026 27512
rect 3050 27510 3106 27512
rect 3130 27510 3186 27512
rect 2890 26476 2946 26478
rect 2970 26476 3026 26478
rect 3050 26476 3106 26478
rect 3130 26476 3186 26478
rect 2890 26424 2916 26476
rect 2916 26424 2946 26476
rect 2970 26424 2980 26476
rect 2980 26424 3026 26476
rect 3050 26424 3096 26476
rect 3096 26424 3106 26476
rect 3130 26424 3160 26476
rect 3160 26424 3186 26476
rect 2890 26422 2946 26424
rect 2970 26422 3026 26424
rect 3050 26422 3106 26424
rect 3130 26422 3186 26424
rect 3368 25558 3424 25594
rect 3368 25538 3370 25558
rect 3370 25538 3422 25558
rect 3422 25538 3424 25558
rect 2890 25388 2946 25390
rect 2970 25388 3026 25390
rect 3050 25388 3106 25390
rect 3130 25388 3186 25390
rect 2890 25336 2916 25388
rect 2916 25336 2946 25388
rect 2970 25336 2980 25388
rect 2980 25336 3026 25388
rect 3050 25336 3096 25388
rect 3096 25336 3106 25388
rect 3130 25336 3160 25388
rect 3160 25336 3186 25388
rect 2890 25334 2946 25336
rect 2970 25334 3026 25336
rect 3050 25334 3106 25336
rect 3130 25334 3186 25336
rect 2890 24300 2946 24302
rect 2970 24300 3026 24302
rect 3050 24300 3106 24302
rect 3130 24300 3186 24302
rect 2890 24248 2916 24300
rect 2916 24248 2946 24300
rect 2970 24248 2980 24300
rect 2980 24248 3026 24300
rect 3050 24248 3096 24300
rect 3096 24248 3106 24300
rect 3130 24248 3160 24300
rect 3160 24248 3186 24300
rect 2890 24246 2946 24248
rect 2970 24246 3026 24248
rect 3050 24246 3106 24248
rect 3130 24246 3186 24248
rect 2890 23212 2946 23214
rect 2970 23212 3026 23214
rect 3050 23212 3106 23214
rect 3130 23212 3186 23214
rect 2890 23160 2916 23212
rect 2916 23160 2946 23212
rect 2970 23160 2980 23212
rect 2980 23160 3026 23212
rect 3050 23160 3096 23212
rect 3096 23160 3106 23212
rect 3130 23160 3160 23212
rect 3160 23160 3186 23212
rect 2890 23158 2946 23160
rect 2970 23158 3026 23160
rect 3050 23158 3106 23160
rect 3130 23158 3186 23160
rect 2890 22124 2946 22126
rect 2970 22124 3026 22126
rect 3050 22124 3106 22126
rect 3130 22124 3186 22126
rect 2890 22072 2916 22124
rect 2916 22072 2946 22124
rect 2970 22072 2980 22124
rect 2980 22072 3026 22124
rect 3050 22072 3096 22124
rect 3096 22072 3106 22124
rect 3130 22072 3160 22124
rect 3160 22072 3186 22124
rect 2890 22070 2946 22072
rect 2970 22070 3026 22072
rect 3050 22070 3106 22072
rect 3130 22070 3186 22072
rect 2890 21036 2946 21038
rect 2970 21036 3026 21038
rect 3050 21036 3106 21038
rect 3130 21036 3186 21038
rect 2890 20984 2916 21036
rect 2916 20984 2946 21036
rect 2970 20984 2980 21036
rect 2980 20984 3026 21036
rect 3050 20984 3096 21036
rect 3096 20984 3106 21036
rect 3130 20984 3160 21036
rect 3160 20984 3186 21036
rect 2890 20982 2946 20984
rect 2970 20982 3026 20984
rect 3050 20982 3106 20984
rect 3130 20982 3186 20984
rect 2890 19948 2946 19950
rect 2970 19948 3026 19950
rect 3050 19948 3106 19950
rect 3130 19948 3186 19950
rect 2890 19896 2916 19948
rect 2916 19896 2946 19948
rect 2970 19896 2980 19948
rect 2980 19896 3026 19948
rect 3050 19896 3096 19948
rect 3096 19896 3106 19948
rect 3130 19896 3160 19948
rect 3160 19896 3186 19948
rect 2890 19894 2946 19896
rect 2970 19894 3026 19896
rect 3050 19894 3106 19896
rect 3130 19894 3186 19896
rect 2890 18860 2946 18862
rect 2970 18860 3026 18862
rect 3050 18860 3106 18862
rect 3130 18860 3186 18862
rect 2890 18808 2916 18860
rect 2916 18808 2946 18860
rect 2970 18808 2980 18860
rect 2980 18808 3026 18860
rect 3050 18808 3096 18860
rect 3096 18808 3106 18860
rect 3130 18808 3160 18860
rect 3160 18808 3186 18860
rect 2890 18806 2946 18808
rect 2970 18806 3026 18808
rect 3050 18806 3106 18808
rect 3130 18806 3186 18808
rect 2890 17772 2946 17774
rect 2970 17772 3026 17774
rect 3050 17772 3106 17774
rect 3130 17772 3186 17774
rect 2890 17720 2916 17772
rect 2916 17720 2946 17772
rect 2970 17720 2980 17772
rect 2980 17720 3026 17772
rect 3050 17720 3096 17772
rect 3096 17720 3106 17772
rect 3130 17720 3160 17772
rect 3160 17720 3186 17772
rect 2890 17718 2946 17720
rect 2970 17718 3026 17720
rect 3050 17718 3106 17720
rect 3130 17718 3186 17720
rect 3552 83102 3554 83122
rect 3554 83102 3606 83122
rect 3606 83102 3608 83122
rect 3552 83066 3608 83102
rect 3460 16970 3516 17026
rect 2890 16684 2946 16686
rect 2970 16684 3026 16686
rect 3050 16684 3106 16686
rect 3130 16684 3186 16686
rect 2890 16632 2916 16684
rect 2916 16632 2946 16684
rect 2970 16632 2980 16684
rect 2980 16632 3026 16684
rect 3050 16632 3096 16684
rect 3096 16632 3106 16684
rect 3130 16632 3160 16684
rect 3160 16632 3186 16684
rect 2890 16630 2946 16632
rect 2970 16630 3026 16632
rect 3050 16630 3106 16632
rect 3130 16630 3186 16632
rect 3460 16562 3516 16618
rect 2890 15596 2946 15598
rect 2970 15596 3026 15598
rect 3050 15596 3106 15598
rect 3130 15596 3186 15598
rect 2890 15544 2916 15596
rect 2916 15544 2946 15596
rect 2970 15544 2980 15596
rect 2980 15544 3026 15596
rect 3050 15544 3096 15596
rect 3096 15544 3106 15596
rect 3130 15544 3160 15596
rect 3160 15544 3186 15596
rect 2890 15542 2946 15544
rect 2970 15542 3026 15544
rect 3050 15542 3106 15544
rect 3130 15542 3186 15544
rect 2890 14508 2946 14510
rect 2970 14508 3026 14510
rect 3050 14508 3106 14510
rect 3130 14508 3186 14510
rect 2890 14456 2916 14508
rect 2916 14456 2946 14508
rect 2970 14456 2980 14508
rect 2980 14456 3026 14508
rect 3050 14456 3096 14508
rect 3096 14456 3106 14508
rect 3130 14456 3160 14508
rect 3160 14456 3186 14508
rect 2890 14454 2946 14456
rect 2970 14454 3026 14456
rect 3050 14454 3106 14456
rect 3130 14454 3186 14456
rect 2890 13420 2946 13422
rect 2970 13420 3026 13422
rect 3050 13420 3106 13422
rect 3130 13420 3186 13422
rect 2890 13368 2916 13420
rect 2916 13368 2946 13420
rect 2970 13368 2980 13420
rect 2980 13368 3026 13420
rect 3050 13368 3096 13420
rect 3096 13368 3106 13420
rect 3130 13368 3160 13420
rect 3160 13368 3186 13420
rect 2890 13366 2946 13368
rect 2970 13366 3026 13368
rect 3050 13366 3106 13368
rect 3130 13366 3186 13368
rect 2890 12332 2946 12334
rect 2970 12332 3026 12334
rect 3050 12332 3106 12334
rect 3130 12332 3186 12334
rect 2890 12280 2916 12332
rect 2916 12280 2946 12332
rect 2970 12280 2980 12332
rect 2980 12280 3026 12332
rect 3050 12280 3096 12332
rect 3096 12280 3106 12332
rect 3130 12280 3160 12332
rect 3160 12280 3186 12332
rect 2890 12278 2946 12280
rect 2970 12278 3026 12280
rect 3050 12278 3106 12280
rect 3130 12278 3186 12280
rect 2890 11244 2946 11246
rect 2970 11244 3026 11246
rect 3050 11244 3106 11246
rect 3130 11244 3186 11246
rect 2890 11192 2916 11244
rect 2916 11192 2946 11244
rect 2970 11192 2980 11244
rect 2980 11192 3026 11244
rect 3050 11192 3096 11244
rect 3096 11192 3106 11244
rect 3130 11192 3160 11244
rect 3160 11192 3186 11244
rect 2890 11190 2946 11192
rect 2970 11190 3026 11192
rect 3050 11190 3106 11192
rect 3130 11190 3186 11192
rect 2890 10156 2946 10158
rect 2970 10156 3026 10158
rect 3050 10156 3106 10158
rect 3130 10156 3186 10158
rect 2890 10104 2916 10156
rect 2916 10104 2946 10156
rect 2970 10104 2980 10156
rect 2980 10104 3026 10156
rect 3050 10104 3096 10156
rect 3096 10104 3106 10156
rect 3130 10104 3160 10156
rect 3160 10104 3186 10156
rect 2890 10102 2946 10104
rect 2970 10102 3026 10104
rect 3050 10102 3106 10104
rect 3130 10102 3186 10104
rect 2890 9068 2946 9070
rect 2970 9068 3026 9070
rect 3050 9068 3106 9070
rect 3130 9068 3186 9070
rect 2890 9016 2916 9068
rect 2916 9016 2946 9068
rect 2970 9016 2980 9068
rect 2980 9016 3026 9068
rect 3050 9016 3096 9068
rect 3096 9016 3106 9068
rect 3130 9016 3160 9068
rect 3160 9016 3186 9068
rect 2890 9014 2946 9016
rect 2970 9014 3026 9016
rect 3050 9014 3106 9016
rect 3130 9014 3186 9016
rect 2890 7980 2946 7982
rect 2970 7980 3026 7982
rect 3050 7980 3106 7982
rect 3130 7980 3186 7982
rect 2890 7928 2916 7980
rect 2916 7928 2946 7980
rect 2970 7928 2980 7980
rect 2980 7928 3026 7980
rect 3050 7928 3096 7980
rect 3096 7928 3106 7980
rect 3130 7928 3160 7980
rect 3160 7928 3186 7980
rect 2890 7926 2946 7928
rect 2970 7926 3026 7928
rect 3050 7926 3106 7928
rect 3130 7926 3186 7928
rect 2890 6892 2946 6894
rect 2970 6892 3026 6894
rect 3050 6892 3106 6894
rect 3130 6892 3186 6894
rect 2890 6840 2916 6892
rect 2916 6840 2946 6892
rect 2970 6840 2980 6892
rect 2980 6840 3026 6892
rect 3050 6840 3096 6892
rect 3096 6840 3106 6892
rect 3130 6840 3160 6892
rect 3160 6840 3186 6892
rect 2890 6838 2946 6840
rect 2970 6838 3026 6840
rect 3050 6838 3106 6840
rect 3130 6838 3186 6840
rect 2890 5804 2946 5806
rect 2970 5804 3026 5806
rect 3050 5804 3106 5806
rect 3130 5804 3186 5806
rect 2890 5752 2916 5804
rect 2916 5752 2946 5804
rect 2970 5752 2980 5804
rect 2980 5752 3026 5804
rect 3050 5752 3096 5804
rect 3096 5752 3106 5804
rect 3130 5752 3160 5804
rect 3160 5752 3186 5804
rect 2890 5750 2946 5752
rect 2970 5750 3026 5752
rect 3050 5750 3106 5752
rect 3130 5750 3186 5752
rect 2890 4716 2946 4718
rect 2970 4716 3026 4718
rect 3050 4716 3106 4718
rect 3130 4716 3186 4718
rect 2890 4664 2916 4716
rect 2916 4664 2946 4716
rect 2970 4664 2980 4716
rect 2980 4664 3026 4716
rect 3050 4664 3096 4716
rect 3096 4664 3106 4716
rect 3130 4664 3160 4716
rect 3160 4664 3186 4716
rect 2890 4662 2946 4664
rect 2970 4662 3026 4664
rect 3050 4662 3106 4664
rect 3130 4662 3186 4664
rect 2908 4222 2910 4242
rect 2910 4222 2962 4242
rect 2962 4222 2964 4242
rect 2908 4186 2964 4222
rect 2890 3628 2946 3630
rect 2970 3628 3026 3630
rect 3050 3628 3106 3630
rect 3130 3628 3186 3630
rect 2890 3576 2916 3628
rect 2916 3576 2946 3628
rect 2970 3576 2980 3628
rect 2980 3576 3026 3628
rect 3050 3576 3096 3628
rect 3096 3576 3106 3628
rect 3130 3576 3160 3628
rect 3160 3576 3186 3628
rect 2890 3574 2946 3576
rect 2970 3574 3026 3576
rect 3050 3574 3106 3576
rect 3130 3574 3186 3576
rect 3276 3526 3332 3562
rect 3276 3506 3278 3526
rect 3278 3506 3330 3526
rect 3330 3506 3332 3526
rect 3000 3098 3056 3154
rect 2724 2710 2780 2746
rect 2724 2690 2726 2710
rect 2726 2690 2778 2710
rect 2778 2690 2780 2710
rect 2890 2540 2946 2542
rect 2970 2540 3026 2542
rect 3050 2540 3106 2542
rect 3130 2540 3186 2542
rect 2890 2488 2916 2540
rect 2916 2488 2946 2540
rect 2970 2488 2980 2540
rect 2980 2488 3026 2540
rect 3050 2488 3096 2540
rect 3096 2488 3106 2540
rect 3130 2488 3160 2540
rect 3160 2488 3186 2540
rect 2890 2486 2946 2488
rect 2970 2486 3026 2488
rect 3050 2486 3106 2488
rect 3130 2486 3186 2488
rect 3828 179898 3884 179954
rect 3736 146714 3792 146770
rect 3736 88778 3792 88834
rect 3736 87554 3792 87610
rect 3644 79938 3700 79994
rect 4012 178846 4014 178866
rect 4014 178846 4066 178866
rect 4066 178846 4068 178866
rect 4012 178810 4068 178846
rect 4012 146714 4068 146770
rect 3920 88506 3976 88562
rect 3828 63074 3884 63130
rect 4104 98334 4106 98354
rect 4106 98334 4158 98354
rect 4158 98334 4160 98354
rect 4104 98298 4160 98334
rect 4104 98182 4160 98218
rect 4104 98162 4106 98182
rect 4106 98162 4158 98182
rect 4158 98162 4160 98182
rect 4104 96394 4160 96450
rect 4288 116422 4290 116442
rect 4290 116422 4342 116442
rect 4342 116422 4344 116442
rect 4288 116386 4344 116422
rect 4472 98298 4528 98354
rect 4196 96258 4252 96314
rect 4288 95034 4344 95090
rect 4104 88542 4106 88562
rect 4106 88542 4158 88562
rect 4158 88542 4160 88562
rect 4104 88506 4160 88542
rect 4012 84698 4068 84754
rect 3736 62938 3792 62994
rect 3644 5158 3700 5194
rect 3644 5138 3646 5158
rect 3646 5138 3698 5158
rect 3698 5138 3700 5158
rect 3460 1466 3516 1522
rect 3920 34514 3976 34570
rect 3920 25538 3976 25594
rect 3828 22818 3884 22874
rect 3736 1738 3792 1794
rect 4196 85922 4252 85978
rect 4012 2010 4068 2066
rect 4288 20542 4290 20562
rect 4290 20542 4342 20562
rect 4342 20542 4344 20562
rect 4288 20506 4344 20542
rect 4196 1874 4252 1930
rect 4380 4614 4436 4650
rect 4380 4594 4382 4614
rect 4382 4594 4434 4614
rect 4434 4594 4436 4614
rect 4380 3234 4436 3290
rect 4380 2690 4436 2746
rect 4748 2554 4804 2610
rect 5576 151782 5578 151802
rect 5578 151782 5630 151802
rect 5630 151782 5632 151802
rect 5576 151746 5632 151782
rect 5208 96666 5264 96722
rect 81752 187922 81808 187978
rect 85156 187922 85212 187978
rect 82488 151746 82544 151802
rect 14592 96802 14648 96858
rect 28484 96802 28540 96858
rect 22136 96666 22192 96722
rect 25264 96666 25320 96722
rect 28944 96686 29000 96722
rect 28944 96666 28946 96686
rect 28946 96666 28998 96686
rect 28998 96666 29000 96686
rect 29956 96666 30012 96722
rect 35016 96666 35072 96722
rect 36856 96666 36912 96722
rect 37040 96686 37096 96722
rect 37040 96666 37042 96686
rect 37042 96666 37094 96686
rect 37094 96666 37096 96686
rect 15696 96530 15752 96586
rect 24712 96530 24768 96586
rect 24988 96278 25044 96314
rect 33636 96394 33692 96450
rect 24988 96258 24990 96278
rect 24990 96258 25042 96278
rect 25042 96258 25044 96278
rect 18364 96006 18420 96042
rect 18364 95986 18366 96006
rect 18366 95986 18418 96006
rect 18418 95986 18420 96006
rect 23424 95986 23480 96042
rect 14040 95850 14096 95906
rect 16984 95850 17040 95906
rect 23976 95870 24032 95906
rect 23976 95850 23978 95870
rect 23978 95850 24030 95870
rect 24030 95850 24032 95870
rect 19836 95714 19892 95770
rect 16984 95442 17040 95498
rect 20756 95342 20758 95362
rect 20758 95342 20810 95362
rect 20810 95342 20812 95362
rect 20756 95306 20812 95342
rect 27196 95578 27252 95634
rect 24436 95190 24492 95226
rect 24436 95170 24438 95190
rect 24438 95170 24490 95190
rect 24490 95170 24492 95190
rect 25724 95170 25780 95226
rect 26644 95170 26700 95226
rect 8152 95070 8154 95090
rect 8154 95070 8206 95090
rect 8206 95070 8208 95090
rect 8152 95034 8208 95070
rect 11832 95034 11888 95090
rect 11096 94898 11152 94954
rect 23332 94898 23388 94954
rect 25908 94918 25964 94954
rect 25908 94898 25910 94918
rect 25910 94898 25962 94918
rect 25962 94898 25964 94918
rect 18180 94762 18236 94818
rect 19836 94762 19892 94818
rect 20848 94762 20904 94818
rect 5300 27986 5356 28042
rect 18272 94354 18328 94410
rect 26000 94782 26056 94818
rect 26000 94762 26002 94782
rect 26002 94762 26054 94782
rect 26054 94762 26056 94782
rect 24620 94082 24676 94138
rect 27288 94646 27344 94682
rect 27288 94626 27290 94646
rect 27290 94626 27342 94646
rect 27342 94626 27344 94646
rect 28392 94102 28448 94138
rect 28392 94082 28394 94102
rect 28394 94082 28446 94102
rect 28446 94082 28448 94102
rect 38144 96122 38200 96178
rect 34464 95170 34520 95226
rect 31152 95034 31208 95090
rect 35660 95170 35716 95226
rect 36212 95170 36268 95226
rect 48724 96938 48780 96994
rect 55532 96938 55588 96994
rect 46608 96802 46664 96858
rect 51024 96802 51080 96858
rect 48724 96666 48780 96722
rect 48908 96686 48964 96722
rect 48908 96666 48910 96686
rect 48910 96666 48962 96686
rect 48962 96666 48964 96686
rect 50196 96666 50252 96722
rect 46608 96530 46664 96586
rect 37500 95170 37556 95226
rect 38604 95170 38660 95226
rect 41824 95170 41880 95226
rect 43756 95170 43812 95226
rect 44492 95170 44548 95226
rect 36304 95034 36360 95090
rect 37316 95054 37372 95090
rect 37316 95034 37318 95054
rect 37318 95034 37370 95054
rect 37370 95034 37372 95054
rect 38788 95034 38844 95090
rect 43940 95034 43996 95090
rect 35016 94898 35072 94954
rect 29772 94374 29828 94410
rect 29772 94354 29774 94374
rect 29774 94354 29826 94374
rect 29826 94354 29828 94374
rect 32440 94626 32496 94682
rect 31060 93946 31116 94002
rect 30692 93810 30748 93866
rect 29680 93402 29736 93458
rect 27196 93266 27252 93322
rect 32348 93810 32404 93866
rect 33636 93810 33692 93866
rect 34924 93810 34980 93866
rect 36212 93810 36268 93866
rect 36304 93674 36360 93730
rect 38052 93538 38108 93594
rect 38236 93538 38292 93594
rect 40076 94490 40132 94546
rect 38880 93810 38936 93866
rect 41456 94510 41512 94546
rect 41456 94490 41458 94510
rect 41458 94490 41510 94510
rect 41510 94490 41512 94510
rect 42652 94510 42708 94546
rect 42652 94490 42654 94510
rect 42654 94490 42706 94510
rect 42706 94490 42708 94510
rect 41272 94354 41328 94410
rect 41732 94354 41788 94410
rect 43940 94354 43996 94410
rect 45228 94354 45284 94410
rect 42652 94082 42708 94138
rect 42744 93810 42800 93866
rect 47620 96122 47676 96178
rect 46516 95170 46572 95226
rect 47804 95170 47860 95226
rect 48724 95190 48780 95226
rect 48724 95170 48726 95190
rect 48726 95170 48778 95190
rect 48778 95170 48780 95190
rect 50196 95170 50252 95226
rect 49092 95070 49094 95090
rect 49094 95070 49146 95090
rect 49146 95070 49148 95090
rect 49092 95034 49148 95070
rect 50380 95034 50436 95090
rect 51484 95578 51540 95634
rect 51576 95170 51632 95226
rect 55532 96394 55588 96450
rect 50288 94782 50344 94818
rect 50288 94762 50290 94782
rect 50290 94762 50342 94782
rect 50342 94762 50344 94782
rect 49092 94626 49148 94682
rect 51668 94374 51724 94410
rect 51668 94354 51670 94374
rect 51670 94354 51722 94374
rect 51722 94354 51724 94374
rect 46148 93946 46204 94002
rect 48816 92994 48872 93050
rect 52956 94646 53012 94682
rect 52956 94626 52958 94646
rect 52958 94626 53010 94646
rect 53010 94626 53012 94646
rect 56636 95170 56692 95226
rect 54244 95034 54300 95090
rect 54152 94762 54208 94818
rect 57924 95170 57980 95226
rect 59396 95206 59398 95226
rect 59398 95206 59450 95226
rect 59450 95206 59452 95226
rect 59396 95170 59452 95206
rect 58108 95034 58164 95090
rect 56360 94354 56416 94410
rect 54152 93946 54208 94002
rect 53692 93810 53748 93866
rect 56912 94218 56968 94274
rect 56912 92722 56968 92778
rect 77980 96938 78036 96994
rect 64548 96666 64604 96722
rect 66572 96666 66628 96722
rect 73472 96666 73528 96722
rect 64916 96530 64972 96586
rect 62064 96430 62066 96450
rect 62066 96430 62118 96450
rect 62118 96430 62120 96450
rect 62064 96394 62120 96430
rect 61788 95170 61844 95226
rect 62432 96122 62488 96178
rect 61972 94218 62028 94274
rect 77980 96530 78036 96586
rect 73564 96394 73620 96450
rect 62800 95170 62856 95226
rect 66480 95070 66482 95090
rect 66482 95070 66534 95090
rect 66534 95070 66536 95090
rect 66480 95034 66536 95070
rect 68504 94490 68560 94546
rect 66480 94390 66482 94410
rect 66482 94390 66534 94410
rect 66534 94390 66536 94410
rect 66480 94354 66536 94390
rect 55348 92606 55404 92642
rect 55348 92586 55350 92606
rect 55350 92586 55402 92606
rect 55402 92586 55404 92606
rect 60500 92586 60556 92642
rect 70988 94490 71044 94546
rect 70988 94390 70990 94410
rect 70990 94390 71042 94410
rect 71042 94390 71044 94410
rect 70988 94354 71044 94390
rect 80096 95714 80152 95770
rect 81476 96666 81532 96722
rect 81660 95850 81716 95906
rect 80096 94898 80152 94954
rect 81844 95986 81900 96042
rect 86890 187500 86946 187502
rect 86970 187500 87026 187502
rect 87050 187500 87106 187502
rect 87130 187500 87186 187502
rect 86890 187448 86916 187500
rect 86916 187448 86946 187500
rect 86970 187448 86980 187500
rect 86980 187448 87026 187500
rect 87050 187448 87096 187500
rect 87096 187448 87106 187500
rect 87130 187448 87160 187500
rect 87160 187448 87186 187500
rect 86890 187446 86946 187448
rect 86970 187446 87026 187448
rect 87050 187446 87106 187448
rect 87130 187446 87186 187448
rect 84236 187378 84292 187434
rect 83960 180714 84016 180770
rect 83776 176770 83832 176826
rect 83316 165346 83372 165402
rect 83224 150658 83280 150714
rect 83316 136106 83372 136162
rect 82488 96122 82544 96178
rect 83224 95306 83280 95362
rect 83592 130122 83648 130178
rect 82672 94626 82728 94682
rect 78440 93810 78496 93866
rect 80096 92722 80152 92778
rect 73748 92586 73804 92642
rect 81752 94354 81808 94410
rect 81844 93674 81900 93730
rect 81660 93538 81716 93594
rect 81384 93130 81440 93186
rect 82488 93402 82544 93458
rect 82120 93266 82176 93322
rect 82304 92994 82360 93050
rect 5760 29482 5816 29538
rect 81476 3234 81532 3290
rect 7876 2454 7878 2474
rect 7878 2454 7930 2474
rect 7930 2454 7932 2474
rect 7876 2418 7932 2454
rect 19744 2826 19800 2882
rect 22136 2826 22192 2882
rect 23976 2862 23978 2882
rect 23978 2862 24030 2882
rect 24030 2862 24032 2882
rect 23976 2826 24032 2862
rect 25080 2826 25136 2882
rect 27472 2846 27528 2882
rect 27472 2826 27474 2846
rect 27474 2826 27526 2846
rect 27526 2826 27528 2846
rect 19468 2590 19470 2610
rect 19470 2590 19522 2610
rect 19522 2590 19524 2610
rect 19468 2554 19524 2590
rect 24620 2590 24622 2610
rect 24622 2590 24674 2610
rect 24674 2590 24676 2610
rect 24620 2554 24676 2590
rect 31060 2826 31116 2882
rect 33728 2826 33784 2882
rect 26000 2454 26002 2474
rect 26002 2454 26054 2474
rect 26054 2454 26056 2474
rect 26000 2418 26056 2454
rect 18272 2282 18328 2338
rect 28392 2282 28448 2338
rect 19376 2146 19432 2202
rect 19560 2146 19616 2202
rect 26368 2146 26424 2202
rect 8704 1602 8760 1658
rect 22412 1602 22468 1658
rect 24712 1602 24768 1658
rect 29220 1602 29276 1658
rect 33084 1330 33140 1386
rect 11648 922 11704 978
rect 11832 922 11888 978
rect 14408 958 14410 978
rect 14410 958 14462 978
rect 14462 958 14464 978
rect 14408 922 14464 958
rect 16984 922 17040 978
rect 18088 922 18144 978
rect 18916 922 18972 978
rect 20848 922 20904 978
rect 21308 942 21364 978
rect 21308 922 21310 942
rect 21310 922 21362 942
rect 21362 922 21364 942
rect 23424 922 23480 978
rect 24252 922 24308 978
rect 28300 922 28356 978
rect 29404 958 29406 978
rect 29406 958 29458 978
rect 29458 958 29460 978
rect 29404 922 29460 958
rect 31060 922 31116 978
rect 31888 922 31944 978
rect 32900 922 32956 978
rect 34740 922 34796 978
rect 20756 650 20812 706
rect 29864 670 29920 706
rect 29864 650 29866 670
rect 29866 650 29918 670
rect 29918 650 29920 670
rect 32440 534 32496 570
rect 36948 2826 37004 2882
rect 38788 2846 38844 2882
rect 38788 2826 38790 2846
rect 38790 2826 38842 2846
rect 38842 2826 38844 2846
rect 41364 2826 41420 2882
rect 35016 2166 35072 2202
rect 35016 2146 35018 2166
rect 35018 2146 35070 2166
rect 35070 2146 35072 2166
rect 36304 1602 36360 1658
rect 36488 1602 36544 1658
rect 36488 1330 36544 1386
rect 81384 3098 81440 3154
rect 50196 2554 50252 2610
rect 53692 2554 53748 2610
rect 78072 2690 78128 2746
rect 41824 2146 41880 2202
rect 35292 922 35348 978
rect 38328 922 38384 978
rect 32440 514 32442 534
rect 32442 514 32494 534
rect 32494 514 32496 534
rect 38052 378 38108 434
rect 45228 2146 45284 2202
rect 46700 2146 46756 2202
rect 47896 2146 47952 2202
rect 49828 2146 49884 2202
rect 50012 2146 50068 2202
rect 42284 1350 42340 1386
rect 42284 1330 42286 1350
rect 42286 1330 42338 1350
rect 42338 1330 42340 1350
rect 42468 1330 42524 1386
rect 50012 1330 50068 1386
rect 78072 2418 78128 2474
rect 54244 2282 54300 2338
rect 80740 1602 80796 1658
rect 51484 1330 51540 1386
rect 80740 1330 80796 1386
rect 40076 922 40132 978
rect 43940 922 43996 978
rect 46148 922 46204 978
rect 50472 922 50528 978
rect 81292 2690 81348 2746
rect 81292 242 81348 298
rect 81752 786 81808 842
rect 83868 175818 83924 175874
rect 84236 182346 84292 182402
rect 84604 186970 84660 187026
rect 84144 179490 84200 179546
rect 84144 174730 84200 174786
rect 84052 173506 84108 173562
rect 83960 157866 84016 157922
rect 83960 149570 84016 149626
rect 83960 148482 84016 148538
rect 83960 146986 84016 147042
rect 83960 145762 84016 145818
rect 83960 144674 84016 144730
rect 83960 121826 84016 121882
rect 83960 115842 84016 115898
rect 83960 109334 84016 109370
rect 83960 109314 83962 109334
rect 83962 109314 84014 109334
rect 84014 109314 84016 109334
rect 83960 108226 84016 108282
rect 83960 107274 84016 107330
rect 83776 97618 83832 97674
rect 83500 96802 83556 96858
rect 83224 94490 83280 94546
rect 83316 76130 83372 76186
rect 83132 63074 83188 63130
rect 83132 62938 83188 62994
rect 83316 61578 83372 61634
rect 82856 43626 82912 43682
rect 83040 43626 83096 43682
rect 83132 38730 83188 38786
rect 83040 37642 83096 37698
rect 82672 28122 82728 28178
rect 82672 24314 82728 24370
rect 82672 24178 82728 24234
rect 82488 17786 82544 17842
rect 82764 17786 82820 17842
rect 82672 15338 82728 15394
rect 82580 8830 82636 8866
rect 82580 8810 82582 8830
rect 82582 8810 82634 8830
rect 82634 8810 82636 8830
rect 82764 8810 82820 8866
rect 82488 8538 82544 8594
rect 82672 6090 82728 6146
rect 82764 3778 82820 3834
rect 82672 2982 82728 3018
rect 82672 2962 82674 2982
rect 82674 2962 82726 2982
rect 82726 2962 82728 2982
rect 82580 1738 82636 1794
rect 83224 27850 83280 27906
rect 83408 53282 83464 53338
rect 82764 514 82820 570
rect 83592 96258 83648 96314
rect 83592 51786 83648 51842
rect 83500 28122 83556 28178
rect 83500 25674 83556 25730
rect 83500 17786 83556 17842
rect 83500 8810 83556 8866
rect 83776 97074 83832 97130
rect 83776 96838 83778 96858
rect 83778 96838 83830 96858
rect 83830 96838 83832 96858
rect 83776 96802 83832 96838
rect 84420 164938 84476 164994
rect 84236 164394 84292 164450
rect 84420 164258 84476 164314
rect 84328 162626 84384 162682
rect 84604 181938 84660 181994
rect 84604 178538 84660 178594
rect 84890 186956 84946 186958
rect 84970 186956 85026 186958
rect 85050 186956 85106 186958
rect 85130 186956 85186 186958
rect 84890 186904 84916 186956
rect 84916 186904 84946 186956
rect 84970 186904 84980 186956
rect 84980 186904 85026 186956
rect 85050 186904 85096 186956
rect 85096 186904 85106 186956
rect 85130 186904 85160 186956
rect 85160 186904 85186 186956
rect 84890 186902 84946 186904
rect 84970 186902 85026 186904
rect 85050 186902 85106 186904
rect 85130 186902 85186 186904
rect 85156 186718 85212 186754
rect 85156 186698 85158 186718
rect 85158 186698 85210 186718
rect 85210 186698 85212 186718
rect 86890 186412 86946 186414
rect 86970 186412 87026 186414
rect 87050 186412 87106 186414
rect 87130 186412 87186 186414
rect 86890 186360 86916 186412
rect 86916 186360 86946 186412
rect 86970 186360 86980 186412
rect 86980 186360 87026 186412
rect 87050 186360 87096 186412
rect 87096 186360 87106 186412
rect 87130 186360 87160 186412
rect 87160 186360 87186 186412
rect 86890 186358 86946 186360
rect 86970 186358 87026 186360
rect 87050 186358 87106 186360
rect 87130 186358 87186 186360
rect 84890 185868 84946 185870
rect 84970 185868 85026 185870
rect 85050 185868 85106 185870
rect 85130 185868 85186 185870
rect 84890 185816 84916 185868
rect 84916 185816 84946 185868
rect 84970 185816 84980 185868
rect 84980 185816 85026 185868
rect 85050 185816 85096 185868
rect 85096 185816 85106 185868
rect 85130 185816 85160 185868
rect 85160 185816 85186 185868
rect 84890 185814 84946 185816
rect 84970 185814 85026 185816
rect 85050 185814 85106 185816
rect 85130 185814 85186 185816
rect 84788 185474 84844 185530
rect 84604 164802 84660 164858
rect 84604 160450 84660 160506
rect 84328 159362 84384 159418
rect 84420 155554 84476 155610
rect 84512 152970 84568 153026
rect 86890 185324 86946 185326
rect 86970 185324 87026 185326
rect 87050 185324 87106 185326
rect 87130 185324 87186 185326
rect 86890 185272 86916 185324
rect 86916 185272 86946 185324
rect 86970 185272 86980 185324
rect 86980 185272 87026 185324
rect 87050 185272 87096 185324
rect 87096 185272 87106 185324
rect 87130 185272 87160 185324
rect 87160 185272 87186 185324
rect 86890 185270 86946 185272
rect 86970 185270 87026 185272
rect 87050 185270 87106 185272
rect 87130 185270 87186 185272
rect 84890 184780 84946 184782
rect 84970 184780 85026 184782
rect 85050 184780 85106 184782
rect 85130 184780 85186 184782
rect 84890 184728 84916 184780
rect 84916 184728 84946 184780
rect 84970 184728 84980 184780
rect 84980 184728 85026 184780
rect 85050 184728 85096 184780
rect 85096 184728 85106 184780
rect 85130 184728 85160 184780
rect 85160 184728 85186 184780
rect 84890 184726 84946 184728
rect 84970 184726 85026 184728
rect 85050 184726 85106 184728
rect 85130 184726 85186 184728
rect 86890 184236 86946 184238
rect 86970 184236 87026 184238
rect 87050 184236 87106 184238
rect 87130 184236 87186 184238
rect 86890 184184 86916 184236
rect 86916 184184 86946 184236
rect 86970 184184 86980 184236
rect 86980 184184 87026 184236
rect 87050 184184 87096 184236
rect 87096 184184 87106 184236
rect 87130 184184 87160 184236
rect 87160 184184 87186 184236
rect 86890 184182 86946 184184
rect 86970 184182 87026 184184
rect 87050 184182 87106 184184
rect 87130 184182 87186 184184
rect 84890 183692 84946 183694
rect 84970 183692 85026 183694
rect 85050 183692 85106 183694
rect 85130 183692 85186 183694
rect 84890 183640 84916 183692
rect 84916 183640 84946 183692
rect 84970 183640 84980 183692
rect 84980 183640 85026 183692
rect 85050 183640 85096 183692
rect 85096 183640 85106 183692
rect 85130 183640 85160 183692
rect 85160 183640 85186 183692
rect 84890 183638 84946 183640
rect 84970 183638 85026 183640
rect 85050 183638 85106 183640
rect 85130 183638 85186 183640
rect 86890 183148 86946 183150
rect 86970 183148 87026 183150
rect 87050 183148 87106 183150
rect 87130 183148 87186 183150
rect 86890 183096 86916 183148
rect 86916 183096 86946 183148
rect 86970 183096 86980 183148
rect 86980 183096 87026 183148
rect 87050 183096 87096 183148
rect 87096 183096 87106 183148
rect 87130 183096 87160 183148
rect 87160 183096 87186 183148
rect 86890 183094 86946 183096
rect 86970 183094 87026 183096
rect 87050 183094 87106 183096
rect 87130 183094 87186 183096
rect 84890 182604 84946 182606
rect 84970 182604 85026 182606
rect 85050 182604 85106 182606
rect 85130 182604 85186 182606
rect 84890 182552 84916 182604
rect 84916 182552 84946 182604
rect 84970 182552 84980 182604
rect 84980 182552 85026 182604
rect 85050 182552 85096 182604
rect 85096 182552 85106 182604
rect 85130 182552 85160 182604
rect 85160 182552 85186 182604
rect 84890 182550 84946 182552
rect 84970 182550 85026 182552
rect 85050 182550 85106 182552
rect 85130 182550 85186 182552
rect 86890 182060 86946 182062
rect 86970 182060 87026 182062
rect 87050 182060 87106 182062
rect 87130 182060 87186 182062
rect 86890 182008 86916 182060
rect 86916 182008 86946 182060
rect 86970 182008 86980 182060
rect 86980 182008 87026 182060
rect 87050 182008 87096 182060
rect 87096 182008 87106 182060
rect 87130 182008 87160 182060
rect 87160 182008 87186 182060
rect 86890 182006 86946 182008
rect 86970 182006 87026 182008
rect 87050 182006 87106 182008
rect 87130 182006 87186 182008
rect 84890 181516 84946 181518
rect 84970 181516 85026 181518
rect 85050 181516 85106 181518
rect 85130 181516 85186 181518
rect 84890 181464 84916 181516
rect 84916 181464 84946 181516
rect 84970 181464 84980 181516
rect 84980 181464 85026 181516
rect 85050 181464 85096 181516
rect 85096 181464 85106 181516
rect 85130 181464 85160 181516
rect 85160 181464 85186 181516
rect 84890 181462 84946 181464
rect 84970 181462 85026 181464
rect 85050 181462 85106 181464
rect 85130 181462 85186 181464
rect 86890 180972 86946 180974
rect 86970 180972 87026 180974
rect 87050 180972 87106 180974
rect 87130 180972 87186 180974
rect 86890 180920 86916 180972
rect 86916 180920 86946 180972
rect 86970 180920 86980 180972
rect 86980 180920 87026 180972
rect 87050 180920 87096 180972
rect 87096 180920 87106 180972
rect 87130 180920 87160 180972
rect 87160 180920 87186 180972
rect 86890 180918 86946 180920
rect 86970 180918 87026 180920
rect 87050 180918 87106 180920
rect 87130 180918 87186 180920
rect 84890 180428 84946 180430
rect 84970 180428 85026 180430
rect 85050 180428 85106 180430
rect 85130 180428 85186 180430
rect 84890 180376 84916 180428
rect 84916 180376 84946 180428
rect 84970 180376 84980 180428
rect 84980 180376 85026 180428
rect 85050 180376 85096 180428
rect 85096 180376 85106 180428
rect 85130 180376 85160 180428
rect 85160 180376 85186 180428
rect 84890 180374 84946 180376
rect 84970 180374 85026 180376
rect 85050 180374 85106 180376
rect 85130 180374 85186 180376
rect 86890 179884 86946 179886
rect 86970 179884 87026 179886
rect 87050 179884 87106 179886
rect 87130 179884 87186 179886
rect 86890 179832 86916 179884
rect 86916 179832 86946 179884
rect 86970 179832 86980 179884
rect 86980 179832 87026 179884
rect 87050 179832 87096 179884
rect 87096 179832 87106 179884
rect 87130 179832 87160 179884
rect 87160 179832 87186 179884
rect 86890 179830 86946 179832
rect 86970 179830 87026 179832
rect 87050 179830 87106 179832
rect 87130 179830 87186 179832
rect 84890 179340 84946 179342
rect 84970 179340 85026 179342
rect 85050 179340 85106 179342
rect 85130 179340 85186 179342
rect 84890 179288 84916 179340
rect 84916 179288 84946 179340
rect 84970 179288 84980 179340
rect 84980 179288 85026 179340
rect 85050 179288 85096 179340
rect 85096 179288 85106 179340
rect 85130 179288 85160 179340
rect 85160 179288 85186 179340
rect 84890 179286 84946 179288
rect 84970 179286 85026 179288
rect 85050 179286 85106 179288
rect 85130 179286 85186 179288
rect 86890 178796 86946 178798
rect 86970 178796 87026 178798
rect 87050 178796 87106 178798
rect 87130 178796 87186 178798
rect 86890 178744 86916 178796
rect 86916 178744 86946 178796
rect 86970 178744 86980 178796
rect 86980 178744 87026 178796
rect 87050 178744 87096 178796
rect 87096 178744 87106 178796
rect 87130 178744 87160 178796
rect 87160 178744 87186 178796
rect 86890 178742 86946 178744
rect 86970 178742 87026 178744
rect 87050 178742 87106 178744
rect 87130 178742 87186 178744
rect 84890 178252 84946 178254
rect 84970 178252 85026 178254
rect 85050 178252 85106 178254
rect 85130 178252 85186 178254
rect 84890 178200 84916 178252
rect 84916 178200 84946 178252
rect 84970 178200 84980 178252
rect 84980 178200 85026 178252
rect 85050 178200 85096 178252
rect 85096 178200 85106 178252
rect 85130 178200 85160 178252
rect 85160 178200 85186 178252
rect 84890 178198 84946 178200
rect 84970 178198 85026 178200
rect 85050 178198 85106 178200
rect 85130 178198 85186 178200
rect 86890 177708 86946 177710
rect 86970 177708 87026 177710
rect 87050 177708 87106 177710
rect 87130 177708 87186 177710
rect 86890 177656 86916 177708
rect 86916 177656 86946 177708
rect 86970 177656 86980 177708
rect 86980 177656 87026 177708
rect 87050 177656 87096 177708
rect 87096 177656 87106 177708
rect 87130 177656 87160 177708
rect 87160 177656 87186 177708
rect 86890 177654 86946 177656
rect 86970 177654 87026 177656
rect 87050 177654 87106 177656
rect 87130 177654 87186 177656
rect 84890 177164 84946 177166
rect 84970 177164 85026 177166
rect 85050 177164 85106 177166
rect 85130 177164 85186 177166
rect 84890 177112 84916 177164
rect 84916 177112 84946 177164
rect 84970 177112 84980 177164
rect 84980 177112 85026 177164
rect 85050 177112 85096 177164
rect 85096 177112 85106 177164
rect 85130 177112 85160 177164
rect 85160 177112 85186 177164
rect 84890 177110 84946 177112
rect 84970 177110 85026 177112
rect 85050 177110 85106 177112
rect 85130 177110 85186 177112
rect 86890 176620 86946 176622
rect 86970 176620 87026 176622
rect 87050 176620 87106 176622
rect 87130 176620 87186 176622
rect 86890 176568 86916 176620
rect 86916 176568 86946 176620
rect 86970 176568 86980 176620
rect 86980 176568 87026 176620
rect 87050 176568 87096 176620
rect 87096 176568 87106 176620
rect 87130 176568 87160 176620
rect 87160 176568 87186 176620
rect 86890 176566 86946 176568
rect 86970 176566 87026 176568
rect 87050 176566 87106 176568
rect 87130 176566 87186 176568
rect 84890 176076 84946 176078
rect 84970 176076 85026 176078
rect 85050 176076 85106 176078
rect 85130 176076 85186 176078
rect 84890 176024 84916 176076
rect 84916 176024 84946 176076
rect 84970 176024 84980 176076
rect 84980 176024 85026 176076
rect 85050 176024 85096 176076
rect 85096 176024 85106 176076
rect 85130 176024 85160 176076
rect 85160 176024 85186 176076
rect 84890 176022 84946 176024
rect 84970 176022 85026 176024
rect 85050 176022 85106 176024
rect 85130 176022 85186 176024
rect 86890 175532 86946 175534
rect 86970 175532 87026 175534
rect 87050 175532 87106 175534
rect 87130 175532 87186 175534
rect 86890 175480 86916 175532
rect 86916 175480 86946 175532
rect 86970 175480 86980 175532
rect 86980 175480 87026 175532
rect 87050 175480 87096 175532
rect 87096 175480 87106 175532
rect 87130 175480 87160 175532
rect 87160 175480 87186 175532
rect 86890 175478 86946 175480
rect 86970 175478 87026 175480
rect 87050 175478 87106 175480
rect 87130 175478 87186 175480
rect 84890 174988 84946 174990
rect 84970 174988 85026 174990
rect 85050 174988 85106 174990
rect 85130 174988 85186 174990
rect 84890 174936 84916 174988
rect 84916 174936 84946 174988
rect 84970 174936 84980 174988
rect 84980 174936 85026 174988
rect 85050 174936 85096 174988
rect 85096 174936 85106 174988
rect 85130 174936 85160 174988
rect 85160 174936 85186 174988
rect 84890 174934 84946 174936
rect 84970 174934 85026 174936
rect 85050 174934 85106 174936
rect 85130 174934 85186 174936
rect 86890 174444 86946 174446
rect 86970 174444 87026 174446
rect 87050 174444 87106 174446
rect 87130 174444 87186 174446
rect 86890 174392 86916 174444
rect 86916 174392 86946 174444
rect 86970 174392 86980 174444
rect 86980 174392 87026 174444
rect 87050 174392 87096 174444
rect 87096 174392 87106 174444
rect 87130 174392 87160 174444
rect 87160 174392 87186 174444
rect 86890 174390 86946 174392
rect 86970 174390 87026 174392
rect 87050 174390 87106 174392
rect 87130 174390 87186 174392
rect 84890 173900 84946 173902
rect 84970 173900 85026 173902
rect 85050 173900 85106 173902
rect 85130 173900 85186 173902
rect 84890 173848 84916 173900
rect 84916 173848 84946 173900
rect 84970 173848 84980 173900
rect 84980 173848 85026 173900
rect 85050 173848 85096 173900
rect 85096 173848 85106 173900
rect 85130 173848 85160 173900
rect 85160 173848 85186 173900
rect 84890 173846 84946 173848
rect 84970 173846 85026 173848
rect 85050 173846 85106 173848
rect 85130 173846 85186 173848
rect 86890 173356 86946 173358
rect 86970 173356 87026 173358
rect 87050 173356 87106 173358
rect 87130 173356 87186 173358
rect 86890 173304 86916 173356
rect 86916 173304 86946 173356
rect 86970 173304 86980 173356
rect 86980 173304 87026 173356
rect 87050 173304 87096 173356
rect 87096 173304 87106 173356
rect 87130 173304 87160 173356
rect 87160 173304 87186 173356
rect 86890 173302 86946 173304
rect 86970 173302 87026 173304
rect 87050 173302 87106 173304
rect 87130 173302 87186 173304
rect 84890 172812 84946 172814
rect 84970 172812 85026 172814
rect 85050 172812 85106 172814
rect 85130 172812 85186 172814
rect 84890 172760 84916 172812
rect 84916 172760 84946 172812
rect 84970 172760 84980 172812
rect 84980 172760 85026 172812
rect 85050 172760 85096 172812
rect 85096 172760 85106 172812
rect 85130 172760 85160 172812
rect 85160 172760 85186 172812
rect 84890 172758 84946 172760
rect 84970 172758 85026 172760
rect 85050 172758 85106 172760
rect 85130 172758 85186 172760
rect 86890 172268 86946 172270
rect 86970 172268 87026 172270
rect 87050 172268 87106 172270
rect 87130 172268 87186 172270
rect 86890 172216 86916 172268
rect 86916 172216 86946 172268
rect 86970 172216 86980 172268
rect 86980 172216 87026 172268
rect 87050 172216 87096 172268
rect 87096 172216 87106 172268
rect 87130 172216 87160 172268
rect 87160 172216 87186 172268
rect 86890 172214 86946 172216
rect 86970 172214 87026 172216
rect 87050 172214 87106 172216
rect 87130 172214 87186 172216
rect 84890 171724 84946 171726
rect 84970 171724 85026 171726
rect 85050 171724 85106 171726
rect 85130 171724 85186 171726
rect 84890 171672 84916 171724
rect 84916 171672 84946 171724
rect 84970 171672 84980 171724
rect 84980 171672 85026 171724
rect 85050 171672 85096 171724
rect 85096 171672 85106 171724
rect 85130 171672 85160 171724
rect 85160 171672 85186 171724
rect 84890 171670 84946 171672
rect 84970 171670 85026 171672
rect 85050 171670 85106 171672
rect 85130 171670 85186 171672
rect 86890 171180 86946 171182
rect 86970 171180 87026 171182
rect 87050 171180 87106 171182
rect 87130 171180 87186 171182
rect 86890 171128 86916 171180
rect 86916 171128 86946 171180
rect 86970 171128 86980 171180
rect 86980 171128 87026 171180
rect 87050 171128 87096 171180
rect 87096 171128 87106 171180
rect 87130 171128 87160 171180
rect 87160 171128 87186 171180
rect 86890 171126 86946 171128
rect 86970 171126 87026 171128
rect 87050 171126 87106 171128
rect 87130 171126 87186 171128
rect 84788 170922 84844 170978
rect 84696 151882 84752 151938
rect 84236 143722 84292 143778
rect 84512 142090 84568 142146
rect 84236 138282 84292 138338
rect 84420 133794 84476 133850
rect 84328 132842 84384 132898
rect 84236 131754 84292 131810
rect 84236 125226 84292 125282
rect 84604 139778 84660 139834
rect 84512 127810 84568 127866
rect 84420 124138 84476 124194
rect 84420 122914 84476 122970
rect 84236 120194 84292 120250
rect 84328 118154 84384 118210
rect 84236 116930 84292 116986
rect 84328 114754 84384 114810
rect 84328 113258 84384 113314
rect 84236 106186 84292 106242
rect 84144 102378 84200 102434
rect 83776 96294 83778 96314
rect 83778 96294 83830 96314
rect 83830 96294 83832 96314
rect 83776 96258 83832 96294
rect 84144 97094 84200 97130
rect 84144 97074 84146 97094
rect 84146 97074 84198 97094
rect 84198 97074 84200 97094
rect 84328 97890 84384 97946
rect 84144 96666 84200 96722
rect 84144 94490 84200 94546
rect 84696 135018 84752 135074
rect 84890 170636 84946 170638
rect 84970 170636 85026 170638
rect 85050 170636 85106 170638
rect 85130 170636 85186 170638
rect 84890 170584 84916 170636
rect 84916 170584 84946 170636
rect 84970 170584 84980 170636
rect 84980 170584 85026 170636
rect 85050 170584 85096 170636
rect 85096 170584 85106 170636
rect 85130 170584 85160 170636
rect 85160 170584 85186 170636
rect 84890 170582 84946 170584
rect 84970 170582 85026 170584
rect 85050 170582 85106 170584
rect 85130 170582 85186 170584
rect 86890 170092 86946 170094
rect 86970 170092 87026 170094
rect 87050 170092 87106 170094
rect 87130 170092 87186 170094
rect 86890 170040 86916 170092
rect 86916 170040 86946 170092
rect 86970 170040 86980 170092
rect 86980 170040 87026 170092
rect 87050 170040 87096 170092
rect 87096 170040 87106 170092
rect 87130 170040 87160 170092
rect 87160 170040 87186 170092
rect 86890 170038 86946 170040
rect 86970 170038 87026 170040
rect 87050 170038 87106 170040
rect 87130 170038 87186 170040
rect 84890 169548 84946 169550
rect 84970 169548 85026 169550
rect 85050 169548 85106 169550
rect 85130 169548 85186 169550
rect 84890 169496 84916 169548
rect 84916 169496 84946 169548
rect 84970 169496 84980 169548
rect 84980 169496 85026 169548
rect 85050 169496 85096 169548
rect 85096 169496 85106 169548
rect 85130 169496 85160 169548
rect 85160 169496 85186 169548
rect 84890 169494 84946 169496
rect 84970 169494 85026 169496
rect 85050 169494 85106 169496
rect 85130 169494 85186 169496
rect 86890 169004 86946 169006
rect 86970 169004 87026 169006
rect 87050 169004 87106 169006
rect 87130 169004 87186 169006
rect 86890 168952 86916 169004
rect 86916 168952 86946 169004
rect 86970 168952 86980 169004
rect 86980 168952 87026 169004
rect 87050 168952 87096 169004
rect 87096 168952 87106 169004
rect 87130 168952 87160 169004
rect 87160 168952 87186 169004
rect 86890 168950 86946 168952
rect 86970 168950 87026 168952
rect 87050 168950 87106 168952
rect 87130 168950 87186 168952
rect 84890 168460 84946 168462
rect 84970 168460 85026 168462
rect 85050 168460 85106 168462
rect 85130 168460 85186 168462
rect 84890 168408 84916 168460
rect 84916 168408 84946 168460
rect 84970 168408 84980 168460
rect 84980 168408 85026 168460
rect 85050 168408 85096 168460
rect 85096 168408 85106 168460
rect 85130 168408 85160 168460
rect 85160 168408 85186 168460
rect 84890 168406 84946 168408
rect 84970 168406 85026 168408
rect 85050 168406 85106 168408
rect 85130 168406 85186 168408
rect 86890 167916 86946 167918
rect 86970 167916 87026 167918
rect 87050 167916 87106 167918
rect 87130 167916 87186 167918
rect 86890 167864 86916 167916
rect 86916 167864 86946 167916
rect 86970 167864 86980 167916
rect 86980 167864 87026 167916
rect 87050 167864 87096 167916
rect 87096 167864 87106 167916
rect 87130 167864 87160 167916
rect 87160 167864 87186 167916
rect 86890 167862 86946 167864
rect 86970 167862 87026 167864
rect 87050 167862 87106 167864
rect 87130 167862 87186 167864
rect 84890 167372 84946 167374
rect 84970 167372 85026 167374
rect 85050 167372 85106 167374
rect 85130 167372 85186 167374
rect 84890 167320 84916 167372
rect 84916 167320 84946 167372
rect 84970 167320 84980 167372
rect 84980 167320 85026 167372
rect 85050 167320 85096 167372
rect 85096 167320 85106 167372
rect 85130 167320 85160 167372
rect 85160 167320 85186 167372
rect 84890 167318 84946 167320
rect 84970 167318 85026 167320
rect 85050 167318 85106 167320
rect 85130 167318 85186 167320
rect 86890 166828 86946 166830
rect 86970 166828 87026 166830
rect 87050 166828 87106 166830
rect 87130 166828 87186 166830
rect 86890 166776 86916 166828
rect 86916 166776 86946 166828
rect 86970 166776 86980 166828
rect 86980 166776 87026 166828
rect 87050 166776 87096 166828
rect 87096 166776 87106 166828
rect 87130 166776 87160 166828
rect 87160 166776 87186 166828
rect 86890 166774 86946 166776
rect 86970 166774 87026 166776
rect 87050 166774 87106 166776
rect 87130 166774 87186 166776
rect 84890 166284 84946 166286
rect 84970 166284 85026 166286
rect 85050 166284 85106 166286
rect 85130 166284 85186 166286
rect 84890 166232 84916 166284
rect 84916 166232 84946 166284
rect 84970 166232 84980 166284
rect 84980 166232 85026 166284
rect 85050 166232 85096 166284
rect 85096 166232 85106 166284
rect 85130 166232 85160 166284
rect 85160 166232 85186 166284
rect 84890 166230 84946 166232
rect 84970 166230 85026 166232
rect 85050 166230 85106 166232
rect 85130 166230 85186 166232
rect 86890 165740 86946 165742
rect 86970 165740 87026 165742
rect 87050 165740 87106 165742
rect 87130 165740 87186 165742
rect 86890 165688 86916 165740
rect 86916 165688 86946 165740
rect 86970 165688 86980 165740
rect 86980 165688 87026 165740
rect 87050 165688 87096 165740
rect 87096 165688 87106 165740
rect 87130 165688 87160 165740
rect 87160 165688 87186 165740
rect 86890 165686 86946 165688
rect 86970 165686 87026 165688
rect 87050 165686 87106 165688
rect 87130 165686 87186 165688
rect 84890 165196 84946 165198
rect 84970 165196 85026 165198
rect 85050 165196 85106 165198
rect 85130 165196 85186 165198
rect 84890 165144 84916 165196
rect 84916 165144 84946 165196
rect 84970 165144 84980 165196
rect 84980 165144 85026 165196
rect 85050 165144 85096 165196
rect 85096 165144 85106 165196
rect 85130 165144 85160 165196
rect 85160 165144 85186 165196
rect 84890 165142 84946 165144
rect 84970 165142 85026 165144
rect 85050 165142 85106 165144
rect 85130 165142 85186 165144
rect 86890 164652 86946 164654
rect 86970 164652 87026 164654
rect 87050 164652 87106 164654
rect 87130 164652 87186 164654
rect 86890 164600 86916 164652
rect 86916 164600 86946 164652
rect 86970 164600 86980 164652
rect 86980 164600 87026 164652
rect 87050 164600 87096 164652
rect 87096 164600 87106 164652
rect 87130 164600 87160 164652
rect 87160 164600 87186 164652
rect 86890 164598 86946 164600
rect 86970 164598 87026 164600
rect 87050 164598 87106 164600
rect 87130 164598 87186 164600
rect 84890 164108 84946 164110
rect 84970 164108 85026 164110
rect 85050 164108 85106 164110
rect 85130 164108 85186 164110
rect 84890 164056 84916 164108
rect 84916 164056 84946 164108
rect 84970 164056 84980 164108
rect 84980 164056 85026 164108
rect 85050 164056 85096 164108
rect 85096 164056 85106 164108
rect 85130 164056 85160 164108
rect 85160 164056 85186 164108
rect 84890 164054 84946 164056
rect 84970 164054 85026 164056
rect 85050 164054 85106 164056
rect 85130 164054 85186 164056
rect 85156 163886 85158 163906
rect 85158 163886 85210 163906
rect 85210 163886 85212 163906
rect 85156 163850 85212 163886
rect 84890 163020 84946 163022
rect 84970 163020 85026 163022
rect 85050 163020 85106 163022
rect 85130 163020 85186 163022
rect 84890 162968 84916 163020
rect 84916 162968 84946 163020
rect 84970 162968 84980 163020
rect 84980 162968 85026 163020
rect 85050 162968 85096 163020
rect 85096 162968 85106 163020
rect 85130 162968 85160 163020
rect 85160 162968 85186 163020
rect 84890 162966 84946 162968
rect 84970 162966 85026 162968
rect 85050 162966 85106 162968
rect 85130 162966 85186 162968
rect 86890 163564 86946 163566
rect 86970 163564 87026 163566
rect 87050 163564 87106 163566
rect 87130 163564 87186 163566
rect 86890 163512 86916 163564
rect 86916 163512 86946 163564
rect 86970 163512 86980 163564
rect 86980 163512 87026 163564
rect 87050 163512 87096 163564
rect 87096 163512 87106 163564
rect 87130 163512 87160 163564
rect 87160 163512 87186 163564
rect 86890 163510 86946 163512
rect 86970 163510 87026 163512
rect 87050 163510 87106 163512
rect 87130 163510 87186 163512
rect 86890 162476 86946 162478
rect 86970 162476 87026 162478
rect 87050 162476 87106 162478
rect 87130 162476 87186 162478
rect 86890 162424 86916 162476
rect 86916 162424 86946 162476
rect 86970 162424 86980 162476
rect 86980 162424 87026 162476
rect 87050 162424 87096 162476
rect 87096 162424 87106 162476
rect 87130 162424 87160 162476
rect 87160 162424 87186 162476
rect 86890 162422 86946 162424
rect 86970 162422 87026 162424
rect 87050 162422 87106 162424
rect 87130 162422 87186 162424
rect 84890 161932 84946 161934
rect 84970 161932 85026 161934
rect 85050 161932 85106 161934
rect 85130 161932 85186 161934
rect 84890 161880 84916 161932
rect 84916 161880 84946 161932
rect 84970 161880 84980 161932
rect 84980 161880 85026 161932
rect 85050 161880 85096 161932
rect 85096 161880 85106 161932
rect 85130 161880 85160 161932
rect 85160 161880 85186 161932
rect 84890 161878 84946 161880
rect 84970 161878 85026 161880
rect 85050 161878 85106 161880
rect 85130 161878 85186 161880
rect 85156 161538 85212 161594
rect 86890 161388 86946 161390
rect 86970 161388 87026 161390
rect 87050 161388 87106 161390
rect 87130 161388 87186 161390
rect 86890 161336 86916 161388
rect 86916 161336 86946 161388
rect 86970 161336 86980 161388
rect 86980 161336 87026 161388
rect 87050 161336 87096 161388
rect 87096 161336 87106 161388
rect 87130 161336 87160 161388
rect 87160 161336 87186 161388
rect 86890 161334 86946 161336
rect 86970 161334 87026 161336
rect 87050 161334 87106 161336
rect 87130 161334 87186 161336
rect 84890 160844 84946 160846
rect 84970 160844 85026 160846
rect 85050 160844 85106 160846
rect 85130 160844 85186 160846
rect 84890 160792 84916 160844
rect 84916 160792 84946 160844
rect 84970 160792 84980 160844
rect 84980 160792 85026 160844
rect 85050 160792 85096 160844
rect 85096 160792 85106 160844
rect 85130 160792 85160 160844
rect 85160 160792 85186 160844
rect 84890 160790 84946 160792
rect 84970 160790 85026 160792
rect 85050 160790 85106 160792
rect 85130 160790 85186 160792
rect 84890 159756 84946 159758
rect 84970 159756 85026 159758
rect 85050 159756 85106 159758
rect 85130 159756 85186 159758
rect 84890 159704 84916 159756
rect 84916 159704 84946 159756
rect 84970 159704 84980 159756
rect 84980 159704 85026 159756
rect 85050 159704 85096 159756
rect 85096 159704 85106 159756
rect 85130 159704 85160 159756
rect 85160 159704 85186 159756
rect 84890 159702 84946 159704
rect 84970 159702 85026 159704
rect 85050 159702 85106 159704
rect 85130 159702 85186 159704
rect 84890 158668 84946 158670
rect 84970 158668 85026 158670
rect 85050 158668 85106 158670
rect 85130 158668 85186 158670
rect 84890 158616 84916 158668
rect 84916 158616 84946 158668
rect 84970 158616 84980 158668
rect 84980 158616 85026 158668
rect 85050 158616 85096 158668
rect 85096 158616 85106 158668
rect 85130 158616 85160 158668
rect 85160 158616 85186 158668
rect 84890 158614 84946 158616
rect 84970 158614 85026 158616
rect 85050 158614 85106 158616
rect 85130 158614 85186 158616
rect 84890 157580 84946 157582
rect 84970 157580 85026 157582
rect 85050 157580 85106 157582
rect 85130 157580 85186 157582
rect 84890 157528 84916 157580
rect 84916 157528 84946 157580
rect 84970 157528 84980 157580
rect 84980 157528 85026 157580
rect 85050 157528 85096 157580
rect 85096 157528 85106 157580
rect 85130 157528 85160 157580
rect 85160 157528 85186 157580
rect 84890 157526 84946 157528
rect 84970 157526 85026 157528
rect 85050 157526 85106 157528
rect 85130 157526 85186 157528
rect 85064 156642 85120 156698
rect 84890 156492 84946 156494
rect 84970 156492 85026 156494
rect 85050 156492 85106 156494
rect 85130 156492 85186 156494
rect 84890 156440 84916 156492
rect 84916 156440 84946 156492
rect 84970 156440 84980 156492
rect 84980 156440 85026 156492
rect 85050 156440 85096 156492
rect 85096 156440 85106 156492
rect 85130 156440 85160 156492
rect 85160 156440 85186 156492
rect 84890 156438 84946 156440
rect 84970 156438 85026 156440
rect 85050 156438 85106 156440
rect 85130 156438 85186 156440
rect 84890 155404 84946 155406
rect 84970 155404 85026 155406
rect 85050 155404 85106 155406
rect 85130 155404 85186 155406
rect 84890 155352 84916 155404
rect 84916 155352 84946 155404
rect 84970 155352 84980 155404
rect 84980 155352 85026 155404
rect 85050 155352 85096 155404
rect 85096 155352 85106 155404
rect 85130 155352 85160 155404
rect 85160 155352 85186 155404
rect 84890 155350 84946 155352
rect 84970 155350 85026 155352
rect 85050 155350 85106 155352
rect 85130 155350 85186 155352
rect 84890 154316 84946 154318
rect 84970 154316 85026 154318
rect 85050 154316 85106 154318
rect 85130 154316 85186 154318
rect 84890 154264 84916 154316
rect 84916 154264 84946 154316
rect 84970 154264 84980 154316
rect 84980 154264 85026 154316
rect 85050 154264 85096 154316
rect 85096 154264 85106 154316
rect 85130 154264 85160 154316
rect 85160 154264 85186 154316
rect 84890 154262 84946 154264
rect 84970 154262 85026 154264
rect 85050 154262 85106 154264
rect 85130 154262 85186 154264
rect 86890 160300 86946 160302
rect 86970 160300 87026 160302
rect 87050 160300 87106 160302
rect 87130 160300 87186 160302
rect 86890 160248 86916 160300
rect 86916 160248 86946 160300
rect 86970 160248 86980 160300
rect 86980 160248 87026 160300
rect 87050 160248 87096 160300
rect 87096 160248 87106 160300
rect 87130 160248 87160 160300
rect 87160 160248 87186 160300
rect 86890 160246 86946 160248
rect 86970 160246 87026 160248
rect 87050 160246 87106 160248
rect 87130 160246 87186 160248
rect 86890 159212 86946 159214
rect 86970 159212 87026 159214
rect 87050 159212 87106 159214
rect 87130 159212 87186 159214
rect 86890 159160 86916 159212
rect 86916 159160 86946 159212
rect 86970 159160 86980 159212
rect 86980 159160 87026 159212
rect 87050 159160 87096 159212
rect 87096 159160 87106 159212
rect 87130 159160 87160 159212
rect 87160 159160 87186 159212
rect 86890 159158 86946 159160
rect 86970 159158 87026 159160
rect 87050 159158 87106 159160
rect 87130 159158 87186 159160
rect 86890 158124 86946 158126
rect 86970 158124 87026 158126
rect 87050 158124 87106 158126
rect 87130 158124 87186 158126
rect 86890 158072 86916 158124
rect 86916 158072 86946 158124
rect 86970 158072 86980 158124
rect 86980 158072 87026 158124
rect 87050 158072 87096 158124
rect 87096 158072 87106 158124
rect 87130 158072 87160 158124
rect 87160 158072 87186 158124
rect 86890 158070 86946 158072
rect 86970 158070 87026 158072
rect 87050 158070 87106 158072
rect 87130 158070 87186 158072
rect 86890 157036 86946 157038
rect 86970 157036 87026 157038
rect 87050 157036 87106 157038
rect 87130 157036 87186 157038
rect 86890 156984 86916 157036
rect 86916 156984 86946 157036
rect 86970 156984 86980 157036
rect 86980 156984 87026 157036
rect 87050 156984 87096 157036
rect 87096 156984 87106 157036
rect 87130 156984 87160 157036
rect 87160 156984 87186 157036
rect 86890 156982 86946 156984
rect 86970 156982 87026 156984
rect 87050 156982 87106 156984
rect 87130 156982 87186 156984
rect 86890 155948 86946 155950
rect 86970 155948 87026 155950
rect 87050 155948 87106 155950
rect 87130 155948 87186 155950
rect 86890 155896 86916 155948
rect 86916 155896 86946 155948
rect 86970 155896 86980 155948
rect 86980 155896 87026 155948
rect 87050 155896 87096 155948
rect 87096 155896 87106 155948
rect 87130 155896 87160 155948
rect 87160 155896 87186 155948
rect 86890 155894 86946 155896
rect 86970 155894 87026 155896
rect 87050 155894 87106 155896
rect 87130 155894 87186 155896
rect 86890 154860 86946 154862
rect 86970 154860 87026 154862
rect 87050 154860 87106 154862
rect 87130 154860 87186 154862
rect 86890 154808 86916 154860
rect 86916 154808 86946 154860
rect 86970 154808 86980 154860
rect 86980 154808 87026 154860
rect 87050 154808 87096 154860
rect 87096 154808 87106 154860
rect 87130 154808 87160 154860
rect 87160 154808 87186 154860
rect 86890 154806 86946 154808
rect 86970 154806 87026 154808
rect 87050 154806 87106 154808
rect 87130 154806 87186 154808
rect 85340 154194 85396 154250
rect 86890 153772 86946 153774
rect 86970 153772 87026 153774
rect 87050 153772 87106 153774
rect 87130 153772 87186 153774
rect 86890 153720 86916 153772
rect 86916 153720 86946 153772
rect 86970 153720 86980 153772
rect 86980 153720 87026 153772
rect 87050 153720 87096 153772
rect 87096 153720 87106 153772
rect 87130 153720 87160 153772
rect 87160 153720 87186 153772
rect 86890 153718 86946 153720
rect 86970 153718 87026 153720
rect 87050 153718 87106 153720
rect 87130 153718 87186 153720
rect 84890 153228 84946 153230
rect 84970 153228 85026 153230
rect 85050 153228 85106 153230
rect 85130 153228 85186 153230
rect 84890 153176 84916 153228
rect 84916 153176 84946 153228
rect 84970 153176 84980 153228
rect 84980 153176 85026 153228
rect 85050 153176 85096 153228
rect 85096 153176 85106 153228
rect 85130 153176 85160 153228
rect 85160 153176 85186 153228
rect 84890 153174 84946 153176
rect 84970 153174 85026 153176
rect 85050 153174 85106 153176
rect 85130 153174 85186 153176
rect 86890 152684 86946 152686
rect 86970 152684 87026 152686
rect 87050 152684 87106 152686
rect 87130 152684 87186 152686
rect 86890 152632 86916 152684
rect 86916 152632 86946 152684
rect 86970 152632 86980 152684
rect 86980 152632 87026 152684
rect 87050 152632 87096 152684
rect 87096 152632 87106 152684
rect 87130 152632 87160 152684
rect 87160 152632 87186 152684
rect 86890 152630 86946 152632
rect 86970 152630 87026 152632
rect 87050 152630 87106 152632
rect 87130 152630 87186 152632
rect 84890 152140 84946 152142
rect 84970 152140 85026 152142
rect 85050 152140 85106 152142
rect 85130 152140 85186 152142
rect 84890 152088 84916 152140
rect 84916 152088 84946 152140
rect 84970 152088 84980 152140
rect 84980 152088 85026 152140
rect 85050 152088 85096 152140
rect 85096 152088 85106 152140
rect 85130 152088 85160 152140
rect 85160 152088 85186 152140
rect 84890 152086 84946 152088
rect 84970 152086 85026 152088
rect 85050 152086 85106 152088
rect 85130 152086 85186 152088
rect 86890 151596 86946 151598
rect 86970 151596 87026 151598
rect 87050 151596 87106 151598
rect 87130 151596 87186 151598
rect 86890 151544 86916 151596
rect 86916 151544 86946 151596
rect 86970 151544 86980 151596
rect 86980 151544 87026 151596
rect 87050 151544 87096 151596
rect 87096 151544 87106 151596
rect 87130 151544 87160 151596
rect 87160 151544 87186 151596
rect 86890 151542 86946 151544
rect 86970 151542 87026 151544
rect 87050 151542 87106 151544
rect 87130 151542 87186 151544
rect 84890 151052 84946 151054
rect 84970 151052 85026 151054
rect 85050 151052 85106 151054
rect 85130 151052 85186 151054
rect 84890 151000 84916 151052
rect 84916 151000 84946 151052
rect 84970 151000 84980 151052
rect 84980 151000 85026 151052
rect 85050 151000 85096 151052
rect 85096 151000 85106 151052
rect 85130 151000 85160 151052
rect 85160 151000 85186 151052
rect 84890 150998 84946 151000
rect 84970 150998 85026 151000
rect 85050 150998 85106 151000
rect 85130 150998 85186 151000
rect 86890 150508 86946 150510
rect 86970 150508 87026 150510
rect 87050 150508 87106 150510
rect 87130 150508 87186 150510
rect 86890 150456 86916 150508
rect 86916 150456 86946 150508
rect 86970 150456 86980 150508
rect 86980 150456 87026 150508
rect 87050 150456 87096 150508
rect 87096 150456 87106 150508
rect 87130 150456 87160 150508
rect 87160 150456 87186 150508
rect 86890 150454 86946 150456
rect 86970 150454 87026 150456
rect 87050 150454 87106 150456
rect 87130 150454 87186 150456
rect 84890 149964 84946 149966
rect 84970 149964 85026 149966
rect 85050 149964 85106 149966
rect 85130 149964 85186 149966
rect 84890 149912 84916 149964
rect 84916 149912 84946 149964
rect 84970 149912 84980 149964
rect 84980 149912 85026 149964
rect 85050 149912 85096 149964
rect 85096 149912 85106 149964
rect 85130 149912 85160 149964
rect 85160 149912 85186 149964
rect 84890 149910 84946 149912
rect 84970 149910 85026 149912
rect 85050 149910 85106 149912
rect 85130 149910 85186 149912
rect 86890 149420 86946 149422
rect 86970 149420 87026 149422
rect 87050 149420 87106 149422
rect 87130 149420 87186 149422
rect 86890 149368 86916 149420
rect 86916 149368 86946 149420
rect 86970 149368 86980 149420
rect 86980 149368 87026 149420
rect 87050 149368 87096 149420
rect 87096 149368 87106 149420
rect 87130 149368 87160 149420
rect 87160 149368 87186 149420
rect 86890 149366 86946 149368
rect 86970 149366 87026 149368
rect 87050 149366 87106 149368
rect 87130 149366 87186 149368
rect 84890 148876 84946 148878
rect 84970 148876 85026 148878
rect 85050 148876 85106 148878
rect 85130 148876 85186 148878
rect 84890 148824 84916 148876
rect 84916 148824 84946 148876
rect 84970 148824 84980 148876
rect 84980 148824 85026 148876
rect 85050 148824 85096 148876
rect 85096 148824 85106 148876
rect 85130 148824 85160 148876
rect 85160 148824 85186 148876
rect 84890 148822 84946 148824
rect 84970 148822 85026 148824
rect 85050 148822 85106 148824
rect 85130 148822 85186 148824
rect 86890 148332 86946 148334
rect 86970 148332 87026 148334
rect 87050 148332 87106 148334
rect 87130 148332 87186 148334
rect 86890 148280 86916 148332
rect 86916 148280 86946 148332
rect 86970 148280 86980 148332
rect 86980 148280 87026 148332
rect 87050 148280 87096 148332
rect 87096 148280 87106 148332
rect 87130 148280 87160 148332
rect 87160 148280 87186 148332
rect 86890 148278 86946 148280
rect 86970 148278 87026 148280
rect 87050 148278 87106 148280
rect 87130 148278 87186 148280
rect 84890 147788 84946 147790
rect 84970 147788 85026 147790
rect 85050 147788 85106 147790
rect 85130 147788 85186 147790
rect 84890 147736 84916 147788
rect 84916 147736 84946 147788
rect 84970 147736 84980 147788
rect 84980 147736 85026 147788
rect 85050 147736 85096 147788
rect 85096 147736 85106 147788
rect 85130 147736 85160 147788
rect 85160 147736 85186 147788
rect 84890 147734 84946 147736
rect 84970 147734 85026 147736
rect 85050 147734 85106 147736
rect 85130 147734 85186 147736
rect 86890 147244 86946 147246
rect 86970 147244 87026 147246
rect 87050 147244 87106 147246
rect 87130 147244 87186 147246
rect 86890 147192 86916 147244
rect 86916 147192 86946 147244
rect 86970 147192 86980 147244
rect 86980 147192 87026 147244
rect 87050 147192 87096 147244
rect 87096 147192 87106 147244
rect 87130 147192 87160 147244
rect 87160 147192 87186 147244
rect 86890 147190 86946 147192
rect 86970 147190 87026 147192
rect 87050 147190 87106 147192
rect 87130 147190 87186 147192
rect 84890 146700 84946 146702
rect 84970 146700 85026 146702
rect 85050 146700 85106 146702
rect 85130 146700 85186 146702
rect 84890 146648 84916 146700
rect 84916 146648 84946 146700
rect 84970 146648 84980 146700
rect 84980 146648 85026 146700
rect 85050 146648 85096 146700
rect 85096 146648 85106 146700
rect 85130 146648 85160 146700
rect 85160 146648 85186 146700
rect 84890 146646 84946 146648
rect 84970 146646 85026 146648
rect 85050 146646 85106 146648
rect 85130 146646 85186 146648
rect 86890 146156 86946 146158
rect 86970 146156 87026 146158
rect 87050 146156 87106 146158
rect 87130 146156 87186 146158
rect 86890 146104 86916 146156
rect 86916 146104 86946 146156
rect 86970 146104 86980 146156
rect 86980 146104 87026 146156
rect 87050 146104 87096 146156
rect 87096 146104 87106 146156
rect 87130 146104 87160 146156
rect 87160 146104 87186 146156
rect 86890 146102 86946 146104
rect 86970 146102 87026 146104
rect 87050 146102 87106 146104
rect 87130 146102 87186 146104
rect 84890 145612 84946 145614
rect 84970 145612 85026 145614
rect 85050 145612 85106 145614
rect 85130 145612 85186 145614
rect 84890 145560 84916 145612
rect 84916 145560 84946 145612
rect 84970 145560 84980 145612
rect 84980 145560 85026 145612
rect 85050 145560 85096 145612
rect 85096 145560 85106 145612
rect 85130 145560 85160 145612
rect 85160 145560 85186 145612
rect 84890 145558 84946 145560
rect 84970 145558 85026 145560
rect 85050 145558 85106 145560
rect 85130 145558 85186 145560
rect 86890 145068 86946 145070
rect 86970 145068 87026 145070
rect 87050 145068 87106 145070
rect 87130 145068 87186 145070
rect 86890 145016 86916 145068
rect 86916 145016 86946 145068
rect 86970 145016 86980 145068
rect 86980 145016 87026 145068
rect 87050 145016 87096 145068
rect 87096 145016 87106 145068
rect 87130 145016 87160 145068
rect 87160 145016 87186 145068
rect 86890 145014 86946 145016
rect 86970 145014 87026 145016
rect 87050 145014 87106 145016
rect 87130 145014 87186 145016
rect 84890 144524 84946 144526
rect 84970 144524 85026 144526
rect 85050 144524 85106 144526
rect 85130 144524 85186 144526
rect 84890 144472 84916 144524
rect 84916 144472 84946 144524
rect 84970 144472 84980 144524
rect 84980 144472 85026 144524
rect 85050 144472 85096 144524
rect 85096 144472 85106 144524
rect 85130 144472 85160 144524
rect 85160 144472 85186 144524
rect 84890 144470 84946 144472
rect 84970 144470 85026 144472
rect 85050 144470 85106 144472
rect 85130 144470 85186 144472
rect 86890 143980 86946 143982
rect 86970 143980 87026 143982
rect 87050 143980 87106 143982
rect 87130 143980 87186 143982
rect 86890 143928 86916 143980
rect 86916 143928 86946 143980
rect 86970 143928 86980 143980
rect 86980 143928 87026 143980
rect 87050 143928 87096 143980
rect 87096 143928 87106 143980
rect 87130 143928 87160 143980
rect 87160 143928 87186 143980
rect 86890 143926 86946 143928
rect 86970 143926 87026 143928
rect 87050 143926 87106 143928
rect 87130 143926 87186 143928
rect 84890 143436 84946 143438
rect 84970 143436 85026 143438
rect 85050 143436 85106 143438
rect 85130 143436 85186 143438
rect 84890 143384 84916 143436
rect 84916 143384 84946 143436
rect 84970 143384 84980 143436
rect 84980 143384 85026 143436
rect 85050 143384 85096 143436
rect 85096 143384 85106 143436
rect 85130 143384 85160 143436
rect 85160 143384 85186 143436
rect 84890 143382 84946 143384
rect 84970 143382 85026 143384
rect 85050 143382 85106 143384
rect 85130 143382 85186 143384
rect 86890 142892 86946 142894
rect 86970 142892 87026 142894
rect 87050 142892 87106 142894
rect 87130 142892 87186 142894
rect 86890 142840 86916 142892
rect 86916 142840 86946 142892
rect 86970 142840 86980 142892
rect 86980 142840 87026 142892
rect 87050 142840 87096 142892
rect 87096 142840 87106 142892
rect 87130 142840 87160 142892
rect 87160 142840 87186 142892
rect 86890 142838 86946 142840
rect 86970 142838 87026 142840
rect 87050 142838 87106 142840
rect 87130 142838 87186 142840
rect 84890 142348 84946 142350
rect 84970 142348 85026 142350
rect 85050 142348 85106 142350
rect 85130 142348 85186 142350
rect 84890 142296 84916 142348
rect 84916 142296 84946 142348
rect 84970 142296 84980 142348
rect 84980 142296 85026 142348
rect 85050 142296 85096 142348
rect 85096 142296 85106 142348
rect 85130 142296 85160 142348
rect 85160 142296 85186 142348
rect 84890 142294 84946 142296
rect 84970 142294 85026 142296
rect 85050 142294 85106 142296
rect 85130 142294 85186 142296
rect 86890 141804 86946 141806
rect 86970 141804 87026 141806
rect 87050 141804 87106 141806
rect 87130 141804 87186 141806
rect 86890 141752 86916 141804
rect 86916 141752 86946 141804
rect 86970 141752 86980 141804
rect 86980 141752 87026 141804
rect 87050 141752 87096 141804
rect 87096 141752 87106 141804
rect 87130 141752 87160 141804
rect 87160 141752 87186 141804
rect 86890 141750 86946 141752
rect 86970 141750 87026 141752
rect 87050 141750 87106 141752
rect 87130 141750 87186 141752
rect 84890 141260 84946 141262
rect 84970 141260 85026 141262
rect 85050 141260 85106 141262
rect 85130 141260 85186 141262
rect 84890 141208 84916 141260
rect 84916 141208 84946 141260
rect 84970 141208 84980 141260
rect 84980 141208 85026 141260
rect 85050 141208 85096 141260
rect 85096 141208 85106 141260
rect 85130 141208 85160 141260
rect 85160 141208 85186 141260
rect 84890 141206 84946 141208
rect 84970 141206 85026 141208
rect 85050 141206 85106 141208
rect 85130 141206 85186 141208
rect 86890 140716 86946 140718
rect 86970 140716 87026 140718
rect 87050 140716 87106 140718
rect 87130 140716 87186 140718
rect 86890 140664 86916 140716
rect 86916 140664 86946 140716
rect 86970 140664 86980 140716
rect 86980 140664 87026 140716
rect 87050 140664 87096 140716
rect 87096 140664 87106 140716
rect 87130 140664 87160 140716
rect 87160 140664 87186 140716
rect 86890 140662 86946 140664
rect 86970 140662 87026 140664
rect 87050 140662 87106 140664
rect 87130 140662 87186 140664
rect 84890 140172 84946 140174
rect 84970 140172 85026 140174
rect 85050 140172 85106 140174
rect 85130 140172 85186 140174
rect 84890 140120 84916 140172
rect 84916 140120 84946 140172
rect 84970 140120 84980 140172
rect 84980 140120 85026 140172
rect 85050 140120 85096 140172
rect 85096 140120 85106 140172
rect 85130 140120 85160 140172
rect 85160 140120 85186 140172
rect 84890 140118 84946 140120
rect 84970 140118 85026 140120
rect 85050 140118 85106 140120
rect 85130 140118 85186 140120
rect 86890 139628 86946 139630
rect 86970 139628 87026 139630
rect 87050 139628 87106 139630
rect 87130 139628 87186 139630
rect 86890 139576 86916 139628
rect 86916 139576 86946 139628
rect 86970 139576 86980 139628
rect 86980 139576 87026 139628
rect 87050 139576 87096 139628
rect 87096 139576 87106 139628
rect 87130 139576 87160 139628
rect 87160 139576 87186 139628
rect 86890 139574 86946 139576
rect 86970 139574 87026 139576
rect 87050 139574 87106 139576
rect 87130 139574 87186 139576
rect 84890 139084 84946 139086
rect 84970 139084 85026 139086
rect 85050 139084 85106 139086
rect 85130 139084 85186 139086
rect 84890 139032 84916 139084
rect 84916 139032 84946 139084
rect 84970 139032 84980 139084
rect 84980 139032 85026 139084
rect 85050 139032 85096 139084
rect 85096 139032 85106 139084
rect 85130 139032 85160 139084
rect 85160 139032 85186 139084
rect 84890 139030 84946 139032
rect 84970 139030 85026 139032
rect 85050 139030 85106 139032
rect 85130 139030 85186 139032
rect 86890 138540 86946 138542
rect 86970 138540 87026 138542
rect 87050 138540 87106 138542
rect 87130 138540 87186 138542
rect 86890 138488 86916 138540
rect 86916 138488 86946 138540
rect 86970 138488 86980 138540
rect 86980 138488 87026 138540
rect 87050 138488 87096 138540
rect 87096 138488 87106 138540
rect 87130 138488 87160 138540
rect 87160 138488 87186 138540
rect 86890 138486 86946 138488
rect 86970 138486 87026 138488
rect 87050 138486 87106 138488
rect 87130 138486 87186 138488
rect 84890 137996 84946 137998
rect 84970 137996 85026 137998
rect 85050 137996 85106 137998
rect 85130 137996 85186 137998
rect 84890 137944 84916 137996
rect 84916 137944 84946 137996
rect 84970 137944 84980 137996
rect 84980 137944 85026 137996
rect 85050 137944 85096 137996
rect 85096 137944 85106 137996
rect 85130 137944 85160 137996
rect 85160 137944 85186 137996
rect 84890 137942 84946 137944
rect 84970 137942 85026 137944
rect 85050 137942 85106 137944
rect 85130 137942 85186 137944
rect 86890 137452 86946 137454
rect 86970 137452 87026 137454
rect 87050 137452 87106 137454
rect 87130 137452 87186 137454
rect 86890 137400 86916 137452
rect 86916 137400 86946 137452
rect 86970 137400 86980 137452
rect 86980 137400 87026 137452
rect 87050 137400 87096 137452
rect 87096 137400 87106 137452
rect 87130 137400 87160 137452
rect 87160 137400 87186 137452
rect 86890 137398 86946 137400
rect 86970 137398 87026 137400
rect 87050 137398 87106 137400
rect 87130 137398 87186 137400
rect 85800 137194 85856 137250
rect 84890 136908 84946 136910
rect 84970 136908 85026 136910
rect 85050 136908 85106 136910
rect 85130 136908 85186 136910
rect 84890 136856 84916 136908
rect 84916 136856 84946 136908
rect 84970 136856 84980 136908
rect 84980 136856 85026 136908
rect 85050 136856 85096 136908
rect 85096 136856 85106 136908
rect 85130 136856 85160 136908
rect 85160 136856 85186 136908
rect 84890 136854 84946 136856
rect 84970 136854 85026 136856
rect 85050 136854 85106 136856
rect 85130 136854 85186 136856
rect 84890 135820 84946 135822
rect 84970 135820 85026 135822
rect 85050 135820 85106 135822
rect 85130 135820 85186 135822
rect 84890 135768 84916 135820
rect 84916 135768 84946 135820
rect 84970 135768 84980 135820
rect 84980 135768 85026 135820
rect 85050 135768 85096 135820
rect 85096 135768 85106 135820
rect 85130 135768 85160 135820
rect 85160 135768 85186 135820
rect 84890 135766 84946 135768
rect 84970 135766 85026 135768
rect 85050 135766 85106 135768
rect 85130 135766 85186 135768
rect 84890 134732 84946 134734
rect 84970 134732 85026 134734
rect 85050 134732 85106 134734
rect 85130 134732 85186 134734
rect 84890 134680 84916 134732
rect 84916 134680 84946 134732
rect 84970 134680 84980 134732
rect 84980 134680 85026 134732
rect 85050 134680 85096 134732
rect 85096 134680 85106 134732
rect 85130 134680 85160 134732
rect 85160 134680 85186 134732
rect 84890 134678 84946 134680
rect 84970 134678 85026 134680
rect 85050 134678 85106 134680
rect 85130 134678 85186 134680
rect 84890 133644 84946 133646
rect 84970 133644 85026 133646
rect 85050 133644 85106 133646
rect 85130 133644 85186 133646
rect 84890 133592 84916 133644
rect 84916 133592 84946 133644
rect 84970 133592 84980 133644
rect 84980 133592 85026 133644
rect 85050 133592 85096 133644
rect 85096 133592 85106 133644
rect 85130 133592 85160 133644
rect 85160 133592 85186 133644
rect 84890 133590 84946 133592
rect 84970 133590 85026 133592
rect 85050 133590 85106 133592
rect 85130 133590 85186 133592
rect 84890 132556 84946 132558
rect 84970 132556 85026 132558
rect 85050 132556 85106 132558
rect 85130 132556 85186 132558
rect 84890 132504 84916 132556
rect 84916 132504 84946 132556
rect 84970 132504 84980 132556
rect 84980 132504 85026 132556
rect 85050 132504 85096 132556
rect 85096 132504 85106 132556
rect 85130 132504 85160 132556
rect 85160 132504 85186 132556
rect 84890 132502 84946 132504
rect 84970 132502 85026 132504
rect 85050 132502 85106 132504
rect 85130 132502 85186 132504
rect 84890 131468 84946 131470
rect 84970 131468 85026 131470
rect 85050 131468 85106 131470
rect 85130 131468 85186 131470
rect 84890 131416 84916 131468
rect 84916 131416 84946 131468
rect 84970 131416 84980 131468
rect 84980 131416 85026 131468
rect 85050 131416 85096 131468
rect 85096 131416 85106 131468
rect 85130 131416 85160 131468
rect 85160 131416 85186 131468
rect 84890 131414 84946 131416
rect 84970 131414 85026 131416
rect 85050 131414 85106 131416
rect 85130 131414 85186 131416
rect 84890 130380 84946 130382
rect 84970 130380 85026 130382
rect 85050 130380 85106 130382
rect 85130 130380 85186 130382
rect 84890 130328 84916 130380
rect 84916 130328 84946 130380
rect 84970 130328 84980 130380
rect 84980 130328 85026 130380
rect 85050 130328 85096 130380
rect 85096 130328 85106 130380
rect 85130 130328 85160 130380
rect 85160 130328 85186 130380
rect 84890 130326 84946 130328
rect 84970 130326 85026 130328
rect 85050 130326 85106 130328
rect 85130 130326 85186 130328
rect 84890 129292 84946 129294
rect 84970 129292 85026 129294
rect 85050 129292 85106 129294
rect 85130 129292 85186 129294
rect 84890 129240 84916 129292
rect 84916 129240 84946 129292
rect 84970 129240 84980 129292
rect 84980 129240 85026 129292
rect 85050 129240 85096 129292
rect 85096 129240 85106 129292
rect 85130 129240 85160 129292
rect 85160 129240 85186 129292
rect 84890 129238 84946 129240
rect 84970 129238 85026 129240
rect 85050 129238 85106 129240
rect 85130 129238 85186 129240
rect 84890 128204 84946 128206
rect 84970 128204 85026 128206
rect 85050 128204 85106 128206
rect 85130 128204 85186 128206
rect 84890 128152 84916 128204
rect 84916 128152 84946 128204
rect 84970 128152 84980 128204
rect 84980 128152 85026 128204
rect 85050 128152 85096 128204
rect 85096 128152 85106 128204
rect 85130 128152 85160 128204
rect 85160 128152 85186 128204
rect 84890 128150 84946 128152
rect 84970 128150 85026 128152
rect 85050 128150 85106 128152
rect 85130 128150 85186 128152
rect 84890 127116 84946 127118
rect 84970 127116 85026 127118
rect 85050 127116 85106 127118
rect 85130 127116 85186 127118
rect 84890 127064 84916 127116
rect 84916 127064 84946 127116
rect 84970 127064 84980 127116
rect 84980 127064 85026 127116
rect 85050 127064 85096 127116
rect 85096 127064 85106 127116
rect 85130 127064 85160 127116
rect 85160 127064 85186 127116
rect 84890 127062 84946 127064
rect 84970 127062 85026 127064
rect 85050 127062 85106 127064
rect 85130 127062 85186 127064
rect 84890 126028 84946 126030
rect 84970 126028 85026 126030
rect 85050 126028 85106 126030
rect 85130 126028 85186 126030
rect 84890 125976 84916 126028
rect 84916 125976 84946 126028
rect 84970 125976 84980 126028
rect 84980 125976 85026 126028
rect 85050 125976 85096 126028
rect 85096 125976 85106 126028
rect 85130 125976 85160 126028
rect 85160 125976 85186 126028
rect 84890 125974 84946 125976
rect 84970 125974 85026 125976
rect 85050 125974 85106 125976
rect 85130 125974 85186 125976
rect 84890 124940 84946 124942
rect 84970 124940 85026 124942
rect 85050 124940 85106 124942
rect 85130 124940 85186 124942
rect 84890 124888 84916 124940
rect 84916 124888 84946 124940
rect 84970 124888 84980 124940
rect 84980 124888 85026 124940
rect 85050 124888 85096 124940
rect 85096 124888 85106 124940
rect 85130 124888 85160 124940
rect 85160 124888 85186 124940
rect 84890 124886 84946 124888
rect 84970 124886 85026 124888
rect 85050 124886 85106 124888
rect 85130 124886 85186 124888
rect 84890 123852 84946 123854
rect 84970 123852 85026 123854
rect 85050 123852 85106 123854
rect 85130 123852 85186 123854
rect 84890 123800 84916 123852
rect 84916 123800 84946 123852
rect 84970 123800 84980 123852
rect 84980 123800 85026 123852
rect 85050 123800 85096 123852
rect 85096 123800 85106 123852
rect 85130 123800 85160 123852
rect 85160 123800 85186 123852
rect 84890 123798 84946 123800
rect 84970 123798 85026 123800
rect 85050 123798 85106 123800
rect 85130 123798 85186 123800
rect 84890 122764 84946 122766
rect 84970 122764 85026 122766
rect 85050 122764 85106 122766
rect 85130 122764 85186 122766
rect 84890 122712 84916 122764
rect 84916 122712 84946 122764
rect 84970 122712 84980 122764
rect 84980 122712 85026 122764
rect 85050 122712 85096 122764
rect 85096 122712 85106 122764
rect 85130 122712 85160 122764
rect 85160 122712 85186 122764
rect 84890 122710 84946 122712
rect 84970 122710 85026 122712
rect 85050 122710 85106 122712
rect 85130 122710 85186 122712
rect 84890 121676 84946 121678
rect 84970 121676 85026 121678
rect 85050 121676 85106 121678
rect 85130 121676 85186 121678
rect 84890 121624 84916 121676
rect 84916 121624 84946 121676
rect 84970 121624 84980 121676
rect 84980 121624 85026 121676
rect 85050 121624 85096 121676
rect 85096 121624 85106 121676
rect 85130 121624 85160 121676
rect 85160 121624 85186 121676
rect 84890 121622 84946 121624
rect 84970 121622 85026 121624
rect 85050 121622 85106 121624
rect 85130 121622 85186 121624
rect 84890 120588 84946 120590
rect 84970 120588 85026 120590
rect 85050 120588 85106 120590
rect 85130 120588 85186 120590
rect 84890 120536 84916 120588
rect 84916 120536 84946 120588
rect 84970 120536 84980 120588
rect 84980 120536 85026 120588
rect 85050 120536 85096 120588
rect 85096 120536 85106 120588
rect 85130 120536 85160 120588
rect 85160 120536 85186 120588
rect 84890 120534 84946 120536
rect 84970 120534 85026 120536
rect 85050 120534 85106 120536
rect 85130 120534 85186 120536
rect 84890 119500 84946 119502
rect 84970 119500 85026 119502
rect 85050 119500 85106 119502
rect 85130 119500 85186 119502
rect 84890 119448 84916 119500
rect 84916 119448 84946 119500
rect 84970 119448 84980 119500
rect 84980 119448 85026 119500
rect 85050 119448 85096 119500
rect 85096 119448 85106 119500
rect 85130 119448 85160 119500
rect 85160 119448 85186 119500
rect 84890 119446 84946 119448
rect 84970 119446 85026 119448
rect 85050 119446 85106 119448
rect 85130 119446 85186 119448
rect 85340 119398 85396 119434
rect 85340 119378 85342 119398
rect 85342 119378 85394 119398
rect 85394 119378 85396 119398
rect 84890 118412 84946 118414
rect 84970 118412 85026 118414
rect 85050 118412 85106 118414
rect 85130 118412 85186 118414
rect 84890 118360 84916 118412
rect 84916 118360 84946 118412
rect 84970 118360 84980 118412
rect 84980 118360 85026 118412
rect 85050 118360 85096 118412
rect 85096 118360 85106 118412
rect 85130 118360 85160 118412
rect 85160 118360 85186 118412
rect 84890 118358 84946 118360
rect 84970 118358 85026 118360
rect 85050 118358 85106 118360
rect 85130 118358 85186 118360
rect 84890 117324 84946 117326
rect 84970 117324 85026 117326
rect 85050 117324 85106 117326
rect 85130 117324 85186 117326
rect 84890 117272 84916 117324
rect 84916 117272 84946 117324
rect 84970 117272 84980 117324
rect 84980 117272 85026 117324
rect 85050 117272 85096 117324
rect 85096 117272 85106 117324
rect 85130 117272 85160 117324
rect 85160 117272 85186 117324
rect 84890 117270 84946 117272
rect 84970 117270 85026 117272
rect 85050 117270 85106 117272
rect 85130 117270 85186 117272
rect 84890 116236 84946 116238
rect 84970 116236 85026 116238
rect 85050 116236 85106 116238
rect 85130 116236 85186 116238
rect 84890 116184 84916 116236
rect 84916 116184 84946 116236
rect 84970 116184 84980 116236
rect 84980 116184 85026 116236
rect 85050 116184 85096 116236
rect 85096 116184 85106 116236
rect 85130 116184 85160 116236
rect 85160 116184 85186 116236
rect 84890 116182 84946 116184
rect 84970 116182 85026 116184
rect 85050 116182 85106 116184
rect 85130 116182 85186 116184
rect 84890 115148 84946 115150
rect 84970 115148 85026 115150
rect 85050 115148 85106 115150
rect 85130 115148 85186 115150
rect 84890 115096 84916 115148
rect 84916 115096 84946 115148
rect 84970 115096 84980 115148
rect 84980 115096 85026 115148
rect 85050 115096 85096 115148
rect 85096 115096 85106 115148
rect 85130 115096 85160 115148
rect 85160 115096 85186 115148
rect 84890 115094 84946 115096
rect 84970 115094 85026 115096
rect 85050 115094 85106 115096
rect 85130 115094 85186 115096
rect 84890 114060 84946 114062
rect 84970 114060 85026 114062
rect 85050 114060 85106 114062
rect 85130 114060 85186 114062
rect 84890 114008 84916 114060
rect 84916 114008 84946 114060
rect 84970 114008 84980 114060
rect 84980 114008 85026 114060
rect 85050 114008 85096 114060
rect 85096 114008 85106 114060
rect 85130 114008 85160 114060
rect 85160 114008 85186 114060
rect 84890 114006 84946 114008
rect 84970 114006 85026 114008
rect 85050 114006 85106 114008
rect 85130 114006 85186 114008
rect 84890 112972 84946 112974
rect 84970 112972 85026 112974
rect 85050 112972 85106 112974
rect 85130 112972 85186 112974
rect 84890 112920 84916 112972
rect 84916 112920 84946 112972
rect 84970 112920 84980 112972
rect 84980 112920 85026 112972
rect 85050 112920 85096 112972
rect 85096 112920 85106 112972
rect 85130 112920 85160 112972
rect 85160 112920 85186 112972
rect 84890 112918 84946 112920
rect 84970 112918 85026 112920
rect 85050 112918 85106 112920
rect 85130 112918 85186 112920
rect 84880 112170 84936 112226
rect 84890 111884 84946 111886
rect 84970 111884 85026 111886
rect 85050 111884 85106 111886
rect 85130 111884 85186 111886
rect 84890 111832 84916 111884
rect 84916 111832 84946 111884
rect 84970 111832 84980 111884
rect 84980 111832 85026 111884
rect 85050 111832 85096 111884
rect 85096 111832 85106 111884
rect 85130 111832 85160 111884
rect 85160 111832 85186 111884
rect 84890 111830 84946 111832
rect 84970 111830 85026 111832
rect 85050 111830 85106 111832
rect 85130 111830 85186 111832
rect 84890 110796 84946 110798
rect 84970 110796 85026 110798
rect 85050 110796 85106 110798
rect 85130 110796 85186 110798
rect 84890 110744 84916 110796
rect 84916 110744 84946 110796
rect 84970 110744 84980 110796
rect 84980 110744 85026 110796
rect 85050 110744 85096 110796
rect 85096 110744 85106 110796
rect 85130 110744 85160 110796
rect 85160 110744 85186 110796
rect 84890 110742 84946 110744
rect 84970 110742 85026 110744
rect 85050 110742 85106 110744
rect 85130 110742 85186 110744
rect 84890 109708 84946 109710
rect 84970 109708 85026 109710
rect 85050 109708 85106 109710
rect 85130 109708 85186 109710
rect 84890 109656 84916 109708
rect 84916 109656 84946 109708
rect 84970 109656 84980 109708
rect 84980 109656 85026 109708
rect 85050 109656 85096 109708
rect 85096 109656 85106 109708
rect 85130 109656 85160 109708
rect 85160 109656 85186 109708
rect 84890 109654 84946 109656
rect 84970 109654 85026 109656
rect 85050 109654 85106 109656
rect 85130 109654 85186 109656
rect 84890 108620 84946 108622
rect 84970 108620 85026 108622
rect 85050 108620 85106 108622
rect 85130 108620 85186 108622
rect 84890 108568 84916 108620
rect 84916 108568 84946 108620
rect 84970 108568 84980 108620
rect 84980 108568 85026 108620
rect 85050 108568 85096 108620
rect 85096 108568 85106 108620
rect 85130 108568 85160 108620
rect 85160 108568 85186 108620
rect 84890 108566 84946 108568
rect 84970 108566 85026 108568
rect 85050 108566 85106 108568
rect 85130 108566 85186 108568
rect 84890 107532 84946 107534
rect 84970 107532 85026 107534
rect 85050 107532 85106 107534
rect 85130 107532 85186 107534
rect 84890 107480 84916 107532
rect 84916 107480 84946 107532
rect 84970 107480 84980 107532
rect 84980 107480 85026 107532
rect 85050 107480 85096 107532
rect 85096 107480 85106 107532
rect 85130 107480 85160 107532
rect 85160 107480 85186 107532
rect 84890 107478 84946 107480
rect 84970 107478 85026 107480
rect 85050 107478 85106 107480
rect 85130 107478 85186 107480
rect 84890 106444 84946 106446
rect 84970 106444 85026 106446
rect 85050 106444 85106 106446
rect 85130 106444 85186 106446
rect 84890 106392 84916 106444
rect 84916 106392 84946 106444
rect 84970 106392 84980 106444
rect 84980 106392 85026 106444
rect 85050 106392 85096 106444
rect 85096 106392 85106 106444
rect 85130 106392 85160 106444
rect 85160 106392 85186 106444
rect 84890 106390 84946 106392
rect 84970 106390 85026 106392
rect 85050 106390 85106 106392
rect 85130 106390 85186 106392
rect 84890 105356 84946 105358
rect 84970 105356 85026 105358
rect 85050 105356 85106 105358
rect 85130 105356 85186 105358
rect 84890 105304 84916 105356
rect 84916 105304 84946 105356
rect 84970 105304 84980 105356
rect 84980 105304 85026 105356
rect 85050 105304 85096 105356
rect 85096 105304 85106 105356
rect 85130 105304 85160 105356
rect 85160 105304 85186 105356
rect 84890 105302 84946 105304
rect 84970 105302 85026 105304
rect 85050 105302 85106 105304
rect 85130 105302 85186 105304
rect 84890 104268 84946 104270
rect 84970 104268 85026 104270
rect 85050 104268 85106 104270
rect 85130 104268 85186 104270
rect 84890 104216 84916 104268
rect 84916 104216 84946 104268
rect 84970 104216 84980 104268
rect 84980 104216 85026 104268
rect 85050 104216 85096 104268
rect 85096 104216 85106 104268
rect 85130 104216 85160 104268
rect 85160 104216 85186 104268
rect 84890 104214 84946 104216
rect 84970 104214 85026 104216
rect 85050 104214 85106 104216
rect 85130 104214 85186 104216
rect 84890 103180 84946 103182
rect 84970 103180 85026 103182
rect 85050 103180 85106 103182
rect 85130 103180 85186 103182
rect 84890 103128 84916 103180
rect 84916 103128 84946 103180
rect 84970 103128 84980 103180
rect 84980 103128 85026 103180
rect 85050 103128 85096 103180
rect 85096 103128 85106 103180
rect 85130 103128 85160 103180
rect 85160 103128 85186 103180
rect 84890 103126 84946 103128
rect 84970 103126 85026 103128
rect 85050 103126 85106 103128
rect 85130 103126 85186 103128
rect 84890 102092 84946 102094
rect 84970 102092 85026 102094
rect 85050 102092 85106 102094
rect 85130 102092 85186 102094
rect 84890 102040 84916 102092
rect 84916 102040 84946 102092
rect 84970 102040 84980 102092
rect 84980 102040 85026 102092
rect 85050 102040 85096 102092
rect 85096 102040 85106 102092
rect 85130 102040 85160 102092
rect 85160 102040 85186 102092
rect 84890 102038 84946 102040
rect 84970 102038 85026 102040
rect 85050 102038 85106 102040
rect 85130 102038 85186 102040
rect 84890 101004 84946 101006
rect 84970 101004 85026 101006
rect 85050 101004 85106 101006
rect 85130 101004 85186 101006
rect 84890 100952 84916 101004
rect 84916 100952 84946 101004
rect 84970 100952 84980 101004
rect 84980 100952 85026 101004
rect 85050 100952 85096 101004
rect 85096 100952 85106 101004
rect 85130 100952 85160 101004
rect 85160 100952 85186 101004
rect 84890 100950 84946 100952
rect 84970 100950 85026 100952
rect 85050 100950 85106 100952
rect 85130 100950 85186 100952
rect 84696 100066 84752 100122
rect 84604 98978 84660 99034
rect 84512 95442 84568 95498
rect 84890 99916 84946 99918
rect 84970 99916 85026 99918
rect 85050 99916 85106 99918
rect 85130 99916 85186 99918
rect 84890 99864 84916 99916
rect 84916 99864 84946 99916
rect 84970 99864 84980 99916
rect 84980 99864 85026 99916
rect 85050 99864 85096 99916
rect 85096 99864 85106 99916
rect 85130 99864 85160 99916
rect 85160 99864 85186 99916
rect 84890 99862 84946 99864
rect 84970 99862 85026 99864
rect 85050 99862 85106 99864
rect 85130 99862 85186 99864
rect 85708 101290 85764 101346
rect 84890 98828 84946 98830
rect 84970 98828 85026 98830
rect 85050 98828 85106 98830
rect 85130 98828 85186 98830
rect 84890 98776 84916 98828
rect 84916 98776 84946 98828
rect 84970 98776 84980 98828
rect 84980 98776 85026 98828
rect 85050 98776 85096 98828
rect 85096 98776 85106 98828
rect 85130 98776 85160 98828
rect 85160 98776 85186 98828
rect 84890 98774 84946 98776
rect 84970 98774 85026 98776
rect 85050 98774 85106 98776
rect 85130 98774 85186 98776
rect 84890 97740 84946 97742
rect 84970 97740 85026 97742
rect 85050 97740 85106 97742
rect 85130 97740 85186 97742
rect 84890 97688 84916 97740
rect 84916 97688 84946 97740
rect 84970 97688 84980 97740
rect 84980 97688 85026 97740
rect 85050 97688 85096 97740
rect 85096 97688 85106 97740
rect 85130 97688 85160 97740
rect 85160 97688 85186 97740
rect 84890 97686 84946 97688
rect 84970 97686 85026 97688
rect 85050 97686 85106 97688
rect 85130 97686 85186 97688
rect 84890 96652 84946 96654
rect 84970 96652 85026 96654
rect 85050 96652 85106 96654
rect 85130 96652 85186 96654
rect 84890 96600 84916 96652
rect 84916 96600 84946 96652
rect 84970 96600 84980 96652
rect 84980 96600 85026 96652
rect 85050 96600 85096 96652
rect 85096 96600 85106 96652
rect 85130 96600 85160 96652
rect 85160 96600 85186 96652
rect 84890 96598 84946 96600
rect 84970 96598 85026 96600
rect 85050 96598 85106 96600
rect 85130 96598 85186 96600
rect 85340 96802 85396 96858
rect 85432 96530 85488 96586
rect 84890 95564 84946 95566
rect 84970 95564 85026 95566
rect 85050 95564 85106 95566
rect 85130 95564 85186 95566
rect 84890 95512 84916 95564
rect 84916 95512 84946 95564
rect 84970 95512 84980 95564
rect 84980 95512 85026 95564
rect 85050 95512 85096 95564
rect 85096 95512 85106 95564
rect 85130 95512 85160 95564
rect 85160 95512 85186 95564
rect 84890 95510 84946 95512
rect 84970 95510 85026 95512
rect 85050 95510 85106 95512
rect 85130 95510 85186 95512
rect 85156 95306 85212 95362
rect 86890 136364 86946 136366
rect 86970 136364 87026 136366
rect 87050 136364 87106 136366
rect 87130 136364 87186 136366
rect 86890 136312 86916 136364
rect 86916 136312 86946 136364
rect 86970 136312 86980 136364
rect 86980 136312 87026 136364
rect 87050 136312 87096 136364
rect 87096 136312 87106 136364
rect 87130 136312 87160 136364
rect 87160 136312 87186 136364
rect 86890 136310 86946 136312
rect 86970 136310 87026 136312
rect 87050 136310 87106 136312
rect 87130 136310 87186 136312
rect 86890 135276 86946 135278
rect 86970 135276 87026 135278
rect 87050 135276 87106 135278
rect 87130 135276 87186 135278
rect 86890 135224 86916 135276
rect 86916 135224 86946 135276
rect 86970 135224 86980 135276
rect 86980 135224 87026 135276
rect 87050 135224 87096 135276
rect 87096 135224 87106 135276
rect 87130 135224 87160 135276
rect 87160 135224 87186 135276
rect 86890 135222 86946 135224
rect 86970 135222 87026 135224
rect 87050 135222 87106 135224
rect 87130 135222 87186 135224
rect 86890 134188 86946 134190
rect 86970 134188 87026 134190
rect 87050 134188 87106 134190
rect 87130 134188 87186 134190
rect 86890 134136 86916 134188
rect 86916 134136 86946 134188
rect 86970 134136 86980 134188
rect 86980 134136 87026 134188
rect 87050 134136 87096 134188
rect 87096 134136 87106 134188
rect 87130 134136 87160 134188
rect 87160 134136 87186 134188
rect 86890 134134 86946 134136
rect 86970 134134 87026 134136
rect 87050 134134 87106 134136
rect 87130 134134 87186 134136
rect 86890 133100 86946 133102
rect 86970 133100 87026 133102
rect 87050 133100 87106 133102
rect 87130 133100 87186 133102
rect 86890 133048 86916 133100
rect 86916 133048 86946 133100
rect 86970 133048 86980 133100
rect 86980 133048 87026 133100
rect 87050 133048 87096 133100
rect 87096 133048 87106 133100
rect 87130 133048 87160 133100
rect 87160 133048 87186 133100
rect 86890 133046 86946 133048
rect 86970 133046 87026 133048
rect 87050 133046 87106 133048
rect 87130 133046 87186 133048
rect 86890 132012 86946 132014
rect 86970 132012 87026 132014
rect 87050 132012 87106 132014
rect 87130 132012 87186 132014
rect 86890 131960 86916 132012
rect 86916 131960 86946 132012
rect 86970 131960 86980 132012
rect 86980 131960 87026 132012
rect 87050 131960 87096 132012
rect 87096 131960 87106 132012
rect 87130 131960 87160 132012
rect 87160 131960 87186 132012
rect 86890 131958 86946 131960
rect 86970 131958 87026 131960
rect 87050 131958 87106 131960
rect 87130 131958 87186 131960
rect 86890 130924 86946 130926
rect 86970 130924 87026 130926
rect 87050 130924 87106 130926
rect 87130 130924 87186 130926
rect 86890 130872 86916 130924
rect 86916 130872 86946 130924
rect 86970 130872 86980 130924
rect 86980 130872 87026 130924
rect 87050 130872 87096 130924
rect 87096 130872 87106 130924
rect 87130 130872 87160 130924
rect 87160 130872 87186 130924
rect 86890 130870 86946 130872
rect 86970 130870 87026 130872
rect 87050 130870 87106 130872
rect 87130 130870 87186 130872
rect 86890 129836 86946 129838
rect 86970 129836 87026 129838
rect 87050 129836 87106 129838
rect 87130 129836 87186 129838
rect 86890 129784 86916 129836
rect 86916 129784 86946 129836
rect 86970 129784 86980 129836
rect 86980 129784 87026 129836
rect 87050 129784 87096 129836
rect 87096 129784 87106 129836
rect 87130 129784 87160 129836
rect 87160 129784 87186 129836
rect 86890 129782 86946 129784
rect 86970 129782 87026 129784
rect 87050 129782 87106 129784
rect 87130 129782 87186 129784
rect 85892 129034 85948 129090
rect 86890 128748 86946 128750
rect 86970 128748 87026 128750
rect 87050 128748 87106 128750
rect 87130 128748 87186 128750
rect 86890 128696 86916 128748
rect 86916 128696 86946 128748
rect 86970 128696 86980 128748
rect 86980 128696 87026 128748
rect 87050 128696 87096 128748
rect 87096 128696 87106 128748
rect 87130 128696 87160 128748
rect 87160 128696 87186 128748
rect 86890 128694 86946 128696
rect 86970 128694 87026 128696
rect 87050 128694 87106 128696
rect 87130 128694 87186 128696
rect 86890 127660 86946 127662
rect 86970 127660 87026 127662
rect 87050 127660 87106 127662
rect 87130 127660 87186 127662
rect 86890 127608 86916 127660
rect 86916 127608 86946 127660
rect 86970 127608 86980 127660
rect 86980 127608 87026 127660
rect 87050 127608 87096 127660
rect 87096 127608 87106 127660
rect 87130 127608 87160 127660
rect 87160 127608 87186 127660
rect 86890 127606 86946 127608
rect 86970 127606 87026 127608
rect 87050 127606 87106 127608
rect 87130 127606 87186 127608
rect 86890 126572 86946 126574
rect 86970 126572 87026 126574
rect 87050 126572 87106 126574
rect 87130 126572 87186 126574
rect 86890 126520 86916 126572
rect 86916 126520 86946 126572
rect 86970 126520 86980 126572
rect 86980 126520 87026 126572
rect 87050 126520 87096 126572
rect 87096 126520 87106 126572
rect 87130 126520 87160 126572
rect 87160 126520 87186 126572
rect 86890 126518 86946 126520
rect 86970 126518 87026 126520
rect 87050 126518 87106 126520
rect 87130 126518 87186 126520
rect 85984 126314 86040 126370
rect 86890 125484 86946 125486
rect 86970 125484 87026 125486
rect 87050 125484 87106 125486
rect 87130 125484 87186 125486
rect 86890 125432 86916 125484
rect 86916 125432 86946 125484
rect 86970 125432 86980 125484
rect 86980 125432 87026 125484
rect 87050 125432 87096 125484
rect 87096 125432 87106 125484
rect 87130 125432 87160 125484
rect 87160 125432 87186 125484
rect 86890 125430 86946 125432
rect 86970 125430 87026 125432
rect 87050 125430 87106 125432
rect 87130 125430 87186 125432
rect 86890 124396 86946 124398
rect 86970 124396 87026 124398
rect 87050 124396 87106 124398
rect 87130 124396 87186 124398
rect 86890 124344 86916 124396
rect 86916 124344 86946 124396
rect 86970 124344 86980 124396
rect 86980 124344 87026 124396
rect 87050 124344 87096 124396
rect 87096 124344 87106 124396
rect 87130 124344 87160 124396
rect 87160 124344 87186 124396
rect 86890 124342 86946 124344
rect 86970 124342 87026 124344
rect 87050 124342 87106 124344
rect 87130 124342 87186 124344
rect 86890 123308 86946 123310
rect 86970 123308 87026 123310
rect 87050 123308 87106 123310
rect 87130 123308 87186 123310
rect 86890 123256 86916 123308
rect 86916 123256 86946 123308
rect 86970 123256 86980 123308
rect 86980 123256 87026 123308
rect 87050 123256 87096 123308
rect 87096 123256 87106 123308
rect 87130 123256 87160 123308
rect 87160 123256 87186 123308
rect 86890 123254 86946 123256
rect 86970 123254 87026 123256
rect 87050 123254 87106 123256
rect 87130 123254 87186 123256
rect 86890 122220 86946 122222
rect 86970 122220 87026 122222
rect 87050 122220 87106 122222
rect 87130 122220 87186 122222
rect 86890 122168 86916 122220
rect 86916 122168 86946 122220
rect 86970 122168 86980 122220
rect 86980 122168 87026 122220
rect 87050 122168 87096 122220
rect 87096 122168 87106 122220
rect 87130 122168 87160 122220
rect 87160 122168 87186 122220
rect 86890 122166 86946 122168
rect 86970 122166 87026 122168
rect 87050 122166 87106 122168
rect 87130 122166 87186 122168
rect 86890 121132 86946 121134
rect 86970 121132 87026 121134
rect 87050 121132 87106 121134
rect 87130 121132 87186 121134
rect 86890 121080 86916 121132
rect 86916 121080 86946 121132
rect 86970 121080 86980 121132
rect 86980 121080 87026 121132
rect 87050 121080 87096 121132
rect 87096 121080 87106 121132
rect 87130 121080 87160 121132
rect 87160 121080 87186 121132
rect 86890 121078 86946 121080
rect 86970 121078 87026 121080
rect 87050 121078 87106 121080
rect 87130 121078 87186 121080
rect 86890 120044 86946 120046
rect 86970 120044 87026 120046
rect 87050 120044 87106 120046
rect 87130 120044 87186 120046
rect 86890 119992 86916 120044
rect 86916 119992 86946 120044
rect 86970 119992 86980 120044
rect 86980 119992 87026 120044
rect 87050 119992 87096 120044
rect 87096 119992 87106 120044
rect 87130 119992 87160 120044
rect 87160 119992 87186 120044
rect 86890 119990 86946 119992
rect 86970 119990 87026 119992
rect 87050 119990 87106 119992
rect 87130 119990 87186 119992
rect 86890 118956 86946 118958
rect 86970 118956 87026 118958
rect 87050 118956 87106 118958
rect 87130 118956 87186 118958
rect 86890 118904 86916 118956
rect 86916 118904 86946 118956
rect 86970 118904 86980 118956
rect 86980 118904 87026 118956
rect 87050 118904 87096 118956
rect 87096 118904 87106 118956
rect 87130 118904 87160 118956
rect 87160 118904 87186 118956
rect 86890 118902 86946 118904
rect 86970 118902 87026 118904
rect 87050 118902 87106 118904
rect 87130 118902 87186 118904
rect 86890 117868 86946 117870
rect 86970 117868 87026 117870
rect 87050 117868 87106 117870
rect 87130 117868 87186 117870
rect 86890 117816 86916 117868
rect 86916 117816 86946 117868
rect 86970 117816 86980 117868
rect 86980 117816 87026 117868
rect 87050 117816 87096 117868
rect 87096 117816 87106 117868
rect 87130 117816 87160 117868
rect 87160 117816 87186 117868
rect 86890 117814 86946 117816
rect 86970 117814 87026 117816
rect 87050 117814 87106 117816
rect 87130 117814 87186 117816
rect 86890 116780 86946 116782
rect 86970 116780 87026 116782
rect 87050 116780 87106 116782
rect 87130 116780 87186 116782
rect 86890 116728 86916 116780
rect 86916 116728 86946 116780
rect 86970 116728 86980 116780
rect 86980 116728 87026 116780
rect 87050 116728 87096 116780
rect 87096 116728 87106 116780
rect 87130 116728 87160 116780
rect 87160 116728 87186 116780
rect 86890 116726 86946 116728
rect 86970 116726 87026 116728
rect 87050 116726 87106 116728
rect 87130 116726 87186 116728
rect 86890 115692 86946 115694
rect 86970 115692 87026 115694
rect 87050 115692 87106 115694
rect 87130 115692 87186 115694
rect 86890 115640 86916 115692
rect 86916 115640 86946 115692
rect 86970 115640 86980 115692
rect 86980 115640 87026 115692
rect 87050 115640 87096 115692
rect 87096 115640 87106 115692
rect 87130 115640 87160 115692
rect 87160 115640 87186 115692
rect 86890 115638 86946 115640
rect 86970 115638 87026 115640
rect 87050 115638 87106 115640
rect 87130 115638 87186 115640
rect 86890 114604 86946 114606
rect 86970 114604 87026 114606
rect 87050 114604 87106 114606
rect 87130 114604 87186 114606
rect 86890 114552 86916 114604
rect 86916 114552 86946 114604
rect 86970 114552 86980 114604
rect 86980 114552 87026 114604
rect 87050 114552 87096 114604
rect 87096 114552 87106 114604
rect 87130 114552 87160 114604
rect 87160 114552 87186 114604
rect 86890 114550 86946 114552
rect 86970 114550 87026 114552
rect 87050 114550 87106 114552
rect 87130 114550 87186 114552
rect 86890 113516 86946 113518
rect 86970 113516 87026 113518
rect 87050 113516 87106 113518
rect 87130 113516 87186 113518
rect 86890 113464 86916 113516
rect 86916 113464 86946 113516
rect 86970 113464 86980 113516
rect 86980 113464 87026 113516
rect 87050 113464 87096 113516
rect 87096 113464 87106 113516
rect 87130 113464 87160 113516
rect 87160 113464 87186 113516
rect 86890 113462 86946 113464
rect 86970 113462 87026 113464
rect 87050 113462 87106 113464
rect 87130 113462 87186 113464
rect 86890 112428 86946 112430
rect 86970 112428 87026 112430
rect 87050 112428 87106 112430
rect 87130 112428 87186 112430
rect 86890 112376 86916 112428
rect 86916 112376 86946 112428
rect 86970 112376 86980 112428
rect 86980 112376 87026 112428
rect 87050 112376 87096 112428
rect 87096 112376 87106 112428
rect 87130 112376 87160 112428
rect 87160 112376 87186 112428
rect 86890 112374 86946 112376
rect 86970 112374 87026 112376
rect 87050 112374 87106 112376
rect 87130 112374 87186 112376
rect 86890 111340 86946 111342
rect 86970 111340 87026 111342
rect 87050 111340 87106 111342
rect 87130 111340 87186 111342
rect 86890 111288 86916 111340
rect 86916 111288 86946 111340
rect 86970 111288 86980 111340
rect 86980 111288 87026 111340
rect 87050 111288 87096 111340
rect 87096 111288 87106 111340
rect 87130 111288 87160 111340
rect 87160 111288 87186 111340
rect 86890 111286 86946 111288
rect 86970 111286 87026 111288
rect 87050 111286 87106 111288
rect 87130 111286 87186 111288
rect 86076 110946 86132 111002
rect 86890 110252 86946 110254
rect 86970 110252 87026 110254
rect 87050 110252 87106 110254
rect 87130 110252 87186 110254
rect 86890 110200 86916 110252
rect 86916 110200 86946 110252
rect 86970 110200 86980 110252
rect 86980 110200 87026 110252
rect 87050 110200 87096 110252
rect 87096 110200 87106 110252
rect 87130 110200 87160 110252
rect 87160 110200 87186 110252
rect 86890 110198 86946 110200
rect 86970 110198 87026 110200
rect 87050 110198 87106 110200
rect 87130 110198 87186 110200
rect 86890 109164 86946 109166
rect 86970 109164 87026 109166
rect 87050 109164 87106 109166
rect 87130 109164 87186 109166
rect 86890 109112 86916 109164
rect 86916 109112 86946 109164
rect 86970 109112 86980 109164
rect 86980 109112 87026 109164
rect 87050 109112 87096 109164
rect 87096 109112 87106 109164
rect 87130 109112 87160 109164
rect 87160 109112 87186 109164
rect 86890 109110 86946 109112
rect 86970 109110 87026 109112
rect 87050 109110 87106 109112
rect 87130 109110 87186 109112
rect 86890 108076 86946 108078
rect 86970 108076 87026 108078
rect 87050 108076 87106 108078
rect 87130 108076 87186 108078
rect 86890 108024 86916 108076
rect 86916 108024 86946 108076
rect 86970 108024 86980 108076
rect 86980 108024 87026 108076
rect 87050 108024 87096 108076
rect 87096 108024 87106 108076
rect 87130 108024 87160 108076
rect 87160 108024 87186 108076
rect 86890 108022 86946 108024
rect 86970 108022 87026 108024
rect 87050 108022 87106 108024
rect 87130 108022 87186 108024
rect 86890 106988 86946 106990
rect 86970 106988 87026 106990
rect 87050 106988 87106 106990
rect 87130 106988 87186 106990
rect 86890 106936 86916 106988
rect 86916 106936 86946 106988
rect 86970 106936 86980 106988
rect 86980 106936 87026 106988
rect 87050 106936 87096 106988
rect 87096 106936 87106 106988
rect 87130 106936 87160 106988
rect 87160 106936 87186 106988
rect 86890 106934 86946 106936
rect 86970 106934 87026 106936
rect 87050 106934 87106 106936
rect 87130 106934 87186 106936
rect 86890 105900 86946 105902
rect 86970 105900 87026 105902
rect 87050 105900 87106 105902
rect 87130 105900 87186 105902
rect 86890 105848 86916 105900
rect 86916 105848 86946 105900
rect 86970 105848 86980 105900
rect 86980 105848 87026 105900
rect 87050 105848 87096 105900
rect 87096 105848 87106 105900
rect 87130 105848 87160 105900
rect 87160 105848 87186 105900
rect 86890 105846 86946 105848
rect 86970 105846 87026 105848
rect 87050 105846 87106 105848
rect 87130 105846 87186 105848
rect 86168 104962 86224 105018
rect 85892 94762 85948 94818
rect 84890 94476 84946 94478
rect 84970 94476 85026 94478
rect 85050 94476 85106 94478
rect 85130 94476 85186 94478
rect 84890 94424 84916 94476
rect 84916 94424 84946 94476
rect 84970 94424 84980 94476
rect 84980 94424 85026 94476
rect 85050 94424 85096 94476
rect 85096 94424 85106 94476
rect 85130 94424 85160 94476
rect 85160 94424 85186 94476
rect 84890 94422 84946 94424
rect 84970 94422 85026 94424
rect 85050 94422 85106 94424
rect 85130 94422 85186 94424
rect 83868 93946 83924 94002
rect 83684 30434 83740 30490
rect 83500 2590 83502 2610
rect 83502 2590 83554 2610
rect 83554 2590 83556 2610
rect 83500 2554 83556 2590
rect 83500 2282 83556 2338
rect 83960 91806 83962 91826
rect 83962 91806 84014 91826
rect 84014 91806 84016 91826
rect 83960 91770 84016 91806
rect 83868 46890 83924 46946
rect 84052 90818 84108 90874
rect 84144 89322 84200 89378
rect 84788 94082 84844 94138
rect 86890 104812 86946 104814
rect 86970 104812 87026 104814
rect 87050 104812 87106 104814
rect 87130 104812 87186 104814
rect 86890 104760 86916 104812
rect 86916 104760 86946 104812
rect 86970 104760 86980 104812
rect 86980 104760 87026 104812
rect 87050 104760 87096 104812
rect 87096 104760 87106 104812
rect 87130 104760 87160 104812
rect 87160 104760 87186 104812
rect 86890 104758 86946 104760
rect 86970 104758 87026 104760
rect 87050 104758 87106 104760
rect 87130 104758 87186 104760
rect 86890 103724 86946 103726
rect 86970 103724 87026 103726
rect 87050 103724 87106 103726
rect 87130 103724 87186 103726
rect 86890 103672 86916 103724
rect 86916 103672 86946 103724
rect 86970 103672 86980 103724
rect 86980 103672 87026 103724
rect 87050 103672 87096 103724
rect 87096 103672 87106 103724
rect 87130 103672 87160 103724
rect 87160 103672 87186 103724
rect 86890 103670 86946 103672
rect 86970 103670 87026 103672
rect 87050 103670 87106 103672
rect 87130 103670 87186 103672
rect 86260 103466 86316 103522
rect 86890 102636 86946 102638
rect 86970 102636 87026 102638
rect 87050 102636 87106 102638
rect 87130 102636 87186 102638
rect 86890 102584 86916 102636
rect 86916 102584 86946 102636
rect 86970 102584 86980 102636
rect 86980 102584 87026 102636
rect 87050 102584 87096 102636
rect 87096 102584 87106 102636
rect 87130 102584 87160 102636
rect 87160 102584 87186 102636
rect 86890 102582 86946 102584
rect 86970 102582 87026 102584
rect 87050 102582 87106 102584
rect 87130 102582 87186 102584
rect 86890 101548 86946 101550
rect 86970 101548 87026 101550
rect 87050 101548 87106 101550
rect 87130 101548 87186 101550
rect 86890 101496 86916 101548
rect 86916 101496 86946 101548
rect 86970 101496 86980 101548
rect 86980 101496 87026 101548
rect 87050 101496 87096 101548
rect 87096 101496 87106 101548
rect 87130 101496 87160 101548
rect 87160 101496 87186 101548
rect 86890 101494 86946 101496
rect 86970 101494 87026 101496
rect 87050 101494 87106 101496
rect 87130 101494 87186 101496
rect 86890 100460 86946 100462
rect 86970 100460 87026 100462
rect 87050 100460 87106 100462
rect 87130 100460 87186 100462
rect 86890 100408 86916 100460
rect 86916 100408 86946 100460
rect 86970 100408 86980 100460
rect 86980 100408 87026 100460
rect 87050 100408 87096 100460
rect 87096 100408 87106 100460
rect 87130 100408 87160 100460
rect 87160 100408 87186 100460
rect 86890 100406 86946 100408
rect 86970 100406 87026 100408
rect 87050 100406 87106 100408
rect 87130 100406 87186 100408
rect 86890 99372 86946 99374
rect 86970 99372 87026 99374
rect 87050 99372 87106 99374
rect 87130 99372 87186 99374
rect 86890 99320 86916 99372
rect 86916 99320 86946 99372
rect 86970 99320 86980 99372
rect 86980 99320 87026 99372
rect 87050 99320 87096 99372
rect 87096 99320 87106 99372
rect 87130 99320 87160 99372
rect 87160 99320 87186 99372
rect 86890 99318 86946 99320
rect 86970 99318 87026 99320
rect 87050 99318 87106 99320
rect 87130 99318 87186 99320
rect 86890 98284 86946 98286
rect 86970 98284 87026 98286
rect 87050 98284 87106 98286
rect 87130 98284 87186 98286
rect 86890 98232 86916 98284
rect 86916 98232 86946 98284
rect 86970 98232 86980 98284
rect 86980 98232 87026 98284
rect 87050 98232 87096 98284
rect 87096 98232 87106 98284
rect 87130 98232 87160 98284
rect 87160 98232 87186 98284
rect 86890 98230 86946 98232
rect 86970 98230 87026 98232
rect 87050 98230 87106 98232
rect 87130 98230 87186 98232
rect 86890 97196 86946 97198
rect 86970 97196 87026 97198
rect 87050 97196 87106 97198
rect 87130 97196 87186 97198
rect 86890 97144 86916 97196
rect 86916 97144 86946 97196
rect 86970 97144 86980 97196
rect 86980 97144 87026 97196
rect 87050 97144 87096 97196
rect 87096 97144 87106 97196
rect 87130 97144 87160 97196
rect 87160 97144 87186 97196
rect 86890 97142 86946 97144
rect 86970 97142 87026 97144
rect 87050 97142 87106 97144
rect 87130 97142 87186 97144
rect 86168 93946 86224 94002
rect 84420 88098 84476 88154
rect 84328 85922 84384 85978
rect 84236 84426 84292 84482
rect 84512 83338 84568 83394
rect 84420 82114 84476 82170
rect 84890 93388 84946 93390
rect 84970 93388 85026 93390
rect 85050 93388 85106 93390
rect 85130 93388 85186 93390
rect 84890 93336 84916 93388
rect 84916 93336 84946 93388
rect 84970 93336 84980 93388
rect 84980 93336 85026 93388
rect 85050 93336 85096 93388
rect 85096 93336 85106 93388
rect 85130 93336 85160 93388
rect 85160 93336 85186 93388
rect 84890 93334 84946 93336
rect 84970 93334 85026 93336
rect 85050 93334 85106 93336
rect 85130 93334 85186 93336
rect 85156 92994 85212 93050
rect 84696 87010 84752 87066
rect 84890 92300 84946 92302
rect 84970 92300 85026 92302
rect 85050 92300 85106 92302
rect 85130 92300 85186 92302
rect 84890 92248 84916 92300
rect 84916 92248 84946 92300
rect 84970 92248 84980 92300
rect 84980 92248 85026 92300
rect 85050 92248 85096 92300
rect 85096 92248 85106 92300
rect 85130 92248 85160 92300
rect 85160 92248 85186 92300
rect 84890 92246 84946 92248
rect 84970 92246 85026 92248
rect 85050 92246 85106 92248
rect 85130 92246 85186 92248
rect 85156 91906 85212 91962
rect 84890 91212 84946 91214
rect 84970 91212 85026 91214
rect 85050 91212 85106 91214
rect 85130 91212 85186 91214
rect 84890 91160 84916 91212
rect 84916 91160 84946 91212
rect 84970 91160 84980 91212
rect 84980 91160 85026 91212
rect 85050 91160 85096 91212
rect 85096 91160 85106 91212
rect 85130 91160 85160 91212
rect 85160 91160 85186 91212
rect 84890 91158 84946 91160
rect 84970 91158 85026 91160
rect 85050 91158 85106 91160
rect 85130 91158 85186 91160
rect 84890 90124 84946 90126
rect 84970 90124 85026 90126
rect 85050 90124 85106 90126
rect 85130 90124 85186 90126
rect 84890 90072 84916 90124
rect 84916 90072 84946 90124
rect 84970 90072 84980 90124
rect 84980 90072 85026 90124
rect 85050 90072 85096 90124
rect 85096 90072 85106 90124
rect 85130 90072 85160 90124
rect 85160 90072 85186 90124
rect 84890 90070 84946 90072
rect 84970 90070 85026 90072
rect 85050 90070 85106 90072
rect 85130 90070 85186 90072
rect 84890 89036 84946 89038
rect 84970 89036 85026 89038
rect 85050 89036 85106 89038
rect 85130 89036 85186 89038
rect 84890 88984 84916 89036
rect 84916 88984 84946 89036
rect 84970 88984 84980 89036
rect 84980 88984 85026 89036
rect 85050 88984 85096 89036
rect 85096 88984 85106 89036
rect 85130 88984 85160 89036
rect 85160 88984 85186 89036
rect 84890 88982 84946 88984
rect 84970 88982 85026 88984
rect 85050 88982 85106 88984
rect 85130 88982 85186 88984
rect 84890 87948 84946 87950
rect 84970 87948 85026 87950
rect 85050 87948 85106 87950
rect 85130 87948 85186 87950
rect 84890 87896 84916 87948
rect 84916 87896 84946 87948
rect 84970 87896 84980 87948
rect 84980 87896 85026 87948
rect 85050 87896 85096 87948
rect 85096 87896 85106 87948
rect 85130 87896 85160 87948
rect 85160 87896 85186 87948
rect 84890 87894 84946 87896
rect 84970 87894 85026 87896
rect 85050 87894 85106 87896
rect 85130 87894 85186 87896
rect 84890 86860 84946 86862
rect 84970 86860 85026 86862
rect 85050 86860 85106 86862
rect 85130 86860 85186 86862
rect 84890 86808 84916 86860
rect 84916 86808 84946 86860
rect 84970 86808 84980 86860
rect 84980 86808 85026 86860
rect 85050 86808 85096 86860
rect 85096 86808 85106 86860
rect 85130 86808 85160 86860
rect 85160 86808 85186 86860
rect 84890 86806 84946 86808
rect 84970 86806 85026 86808
rect 85050 86806 85106 86808
rect 85130 86806 85186 86808
rect 84890 85772 84946 85774
rect 84970 85772 85026 85774
rect 85050 85772 85106 85774
rect 85130 85772 85186 85774
rect 84890 85720 84916 85772
rect 84916 85720 84946 85772
rect 84970 85720 84980 85772
rect 84980 85720 85026 85772
rect 85050 85720 85096 85772
rect 85096 85720 85106 85772
rect 85130 85720 85160 85772
rect 85160 85720 85186 85772
rect 84890 85718 84946 85720
rect 84970 85718 85026 85720
rect 85050 85718 85106 85720
rect 85130 85718 85186 85720
rect 84890 84684 84946 84686
rect 84970 84684 85026 84686
rect 85050 84684 85106 84686
rect 85130 84684 85186 84686
rect 84890 84632 84916 84684
rect 84916 84632 84946 84684
rect 84970 84632 84980 84684
rect 84980 84632 85026 84684
rect 85050 84632 85096 84684
rect 85096 84632 85106 84684
rect 85130 84632 85160 84684
rect 85160 84632 85186 84684
rect 84890 84630 84946 84632
rect 84970 84630 85026 84632
rect 85050 84630 85106 84632
rect 85130 84630 85186 84632
rect 84890 83596 84946 83598
rect 84970 83596 85026 83598
rect 85050 83596 85106 83598
rect 85130 83596 85186 83598
rect 84890 83544 84916 83596
rect 84916 83544 84946 83596
rect 84970 83544 84980 83596
rect 84980 83544 85026 83596
rect 85050 83544 85096 83596
rect 85096 83544 85106 83596
rect 85130 83544 85160 83596
rect 85160 83544 85186 83596
rect 84890 83542 84946 83544
rect 84970 83542 85026 83544
rect 85050 83542 85106 83544
rect 85130 83542 85186 83544
rect 84890 82508 84946 82510
rect 84970 82508 85026 82510
rect 85050 82508 85106 82510
rect 85130 82508 85186 82510
rect 84890 82456 84916 82508
rect 84916 82456 84946 82508
rect 84970 82456 84980 82508
rect 84980 82456 85026 82508
rect 85050 82456 85096 82508
rect 85096 82456 85106 82508
rect 85130 82456 85160 82508
rect 85160 82456 85186 82508
rect 84890 82454 84946 82456
rect 84970 82454 85026 82456
rect 85050 82454 85106 82456
rect 85130 82454 85186 82456
rect 84890 81420 84946 81422
rect 84970 81420 85026 81422
rect 85050 81420 85106 81422
rect 85130 81420 85186 81422
rect 84890 81368 84916 81420
rect 84916 81368 84946 81420
rect 84970 81368 84980 81420
rect 84980 81368 85026 81420
rect 85050 81368 85096 81420
rect 85096 81368 85106 81420
rect 85130 81368 85160 81420
rect 85160 81368 85186 81420
rect 84890 81366 84946 81368
rect 84970 81366 85026 81368
rect 85050 81366 85106 81368
rect 85130 81366 85186 81368
rect 84788 80618 84844 80674
rect 84890 80332 84946 80334
rect 84970 80332 85026 80334
rect 85050 80332 85106 80334
rect 85130 80332 85186 80334
rect 84890 80280 84916 80332
rect 84916 80280 84946 80332
rect 84970 80280 84980 80332
rect 84980 80280 85026 80332
rect 85050 80280 85096 80332
rect 85096 80280 85106 80332
rect 85130 80280 85160 80332
rect 85160 80280 85186 80332
rect 84890 80278 84946 80280
rect 84970 80278 85026 80280
rect 85050 80278 85106 80280
rect 85130 80278 85186 80280
rect 84604 79938 84660 79994
rect 84890 79244 84946 79246
rect 84970 79244 85026 79246
rect 85050 79244 85106 79246
rect 85130 79244 85186 79246
rect 84890 79192 84916 79244
rect 84916 79192 84946 79244
rect 84970 79192 84980 79244
rect 84980 79192 85026 79244
rect 85050 79192 85096 79244
rect 85096 79192 85106 79244
rect 85130 79192 85160 79244
rect 85160 79192 85186 79244
rect 84890 79190 84946 79192
rect 84970 79190 85026 79192
rect 85050 79190 85106 79192
rect 85130 79190 85186 79192
rect 84236 78442 84292 78498
rect 84144 77218 84200 77274
rect 84890 78156 84946 78158
rect 84970 78156 85026 78158
rect 85050 78156 85106 78158
rect 85130 78156 85186 78158
rect 84890 78104 84916 78156
rect 84916 78104 84946 78156
rect 84970 78104 84980 78156
rect 84980 78104 85026 78156
rect 85050 78104 85096 78156
rect 85096 78104 85106 78156
rect 85130 78104 85160 78156
rect 85160 78104 85186 78156
rect 84890 78102 84946 78104
rect 84970 78102 85026 78104
rect 85050 78102 85106 78104
rect 85130 78102 85186 78104
rect 84890 77068 84946 77070
rect 84970 77068 85026 77070
rect 85050 77068 85106 77070
rect 85130 77068 85186 77070
rect 84890 77016 84916 77068
rect 84916 77016 84946 77068
rect 84970 77016 84980 77068
rect 84980 77016 85026 77068
rect 85050 77016 85096 77068
rect 85096 77016 85106 77068
rect 85130 77016 85160 77068
rect 85160 77016 85186 77068
rect 84890 77014 84946 77016
rect 84970 77014 85026 77016
rect 85050 77014 85106 77016
rect 85130 77014 85186 77016
rect 84890 75980 84946 75982
rect 84970 75980 85026 75982
rect 85050 75980 85106 75982
rect 85130 75980 85186 75982
rect 84890 75928 84916 75980
rect 84916 75928 84946 75980
rect 84970 75928 84980 75980
rect 84980 75928 85026 75980
rect 85050 75928 85096 75980
rect 85096 75928 85106 75980
rect 85130 75928 85160 75980
rect 85160 75928 85186 75980
rect 84890 75926 84946 75928
rect 84970 75926 85026 75928
rect 85050 75926 85106 75928
rect 85130 75926 85186 75928
rect 84788 75042 84844 75098
rect 84328 70146 84384 70202
rect 84890 74892 84946 74894
rect 84970 74892 85026 74894
rect 85050 74892 85106 74894
rect 85130 74892 85186 74894
rect 84890 74840 84916 74892
rect 84916 74840 84946 74892
rect 84970 74840 84980 74892
rect 84980 74840 85026 74892
rect 85050 74840 85096 74892
rect 85096 74840 85106 74892
rect 85130 74840 85160 74892
rect 85160 74840 85186 74892
rect 84890 74838 84946 74840
rect 84970 74838 85026 74840
rect 85050 74838 85106 74840
rect 85130 74838 85186 74840
rect 84880 73954 84936 74010
rect 84890 73804 84946 73806
rect 84970 73804 85026 73806
rect 85050 73804 85106 73806
rect 85130 73804 85186 73806
rect 84890 73752 84916 73804
rect 84916 73752 84946 73804
rect 84970 73752 84980 73804
rect 84980 73752 85026 73804
rect 85050 73752 85096 73804
rect 85096 73752 85106 73804
rect 85130 73752 85160 73804
rect 85160 73752 85186 73804
rect 84890 73750 84946 73752
rect 84970 73750 85026 73752
rect 85050 73750 85106 73752
rect 85130 73750 85186 73752
rect 84696 72458 84752 72514
rect 84604 71234 84660 71290
rect 84420 69058 84476 69114
rect 84890 72716 84946 72718
rect 84970 72716 85026 72718
rect 85050 72716 85106 72718
rect 85130 72716 85186 72718
rect 84890 72664 84916 72716
rect 84916 72664 84946 72716
rect 84970 72664 84980 72716
rect 84980 72664 85026 72716
rect 85050 72664 85096 72716
rect 85096 72664 85106 72716
rect 85130 72664 85160 72716
rect 85160 72664 85186 72716
rect 84890 72662 84946 72664
rect 84970 72662 85026 72664
rect 85050 72662 85106 72664
rect 85130 72662 85186 72664
rect 84890 71628 84946 71630
rect 84970 71628 85026 71630
rect 85050 71628 85106 71630
rect 85130 71628 85186 71630
rect 84890 71576 84916 71628
rect 84916 71576 84946 71628
rect 84970 71576 84980 71628
rect 84980 71576 85026 71628
rect 85050 71576 85096 71628
rect 85096 71576 85106 71628
rect 85130 71576 85160 71628
rect 85160 71576 85186 71628
rect 84890 71574 84946 71576
rect 84970 71574 85026 71576
rect 85050 71574 85106 71576
rect 85130 71574 85186 71576
rect 84890 70540 84946 70542
rect 84970 70540 85026 70542
rect 85050 70540 85106 70542
rect 85130 70540 85186 70542
rect 84890 70488 84916 70540
rect 84916 70488 84946 70540
rect 84970 70488 84980 70540
rect 84980 70488 85026 70540
rect 85050 70488 85096 70540
rect 85096 70488 85106 70540
rect 85130 70488 85160 70540
rect 85160 70488 85186 70540
rect 84890 70486 84946 70488
rect 84970 70486 85026 70488
rect 85050 70486 85106 70488
rect 85130 70486 85186 70488
rect 84890 69452 84946 69454
rect 84970 69452 85026 69454
rect 85050 69452 85106 69454
rect 85130 69452 85186 69454
rect 84890 69400 84916 69452
rect 84916 69400 84946 69452
rect 84970 69400 84980 69452
rect 84980 69400 85026 69452
rect 85050 69400 85096 69452
rect 85096 69400 85106 69452
rect 85130 69400 85160 69452
rect 85160 69400 85186 69452
rect 84890 69398 84946 69400
rect 84970 69398 85026 69400
rect 85050 69398 85106 69400
rect 85130 69398 85186 69400
rect 84890 68364 84946 68366
rect 84970 68364 85026 68366
rect 85050 68364 85106 68366
rect 85130 68364 85186 68366
rect 84890 68312 84916 68364
rect 84916 68312 84946 68364
rect 84970 68312 84980 68364
rect 84980 68312 85026 68364
rect 85050 68312 85096 68364
rect 85096 68312 85106 68364
rect 85130 68312 85160 68364
rect 85160 68312 85186 68364
rect 84890 68310 84946 68312
rect 84970 68310 85026 68312
rect 85050 68310 85106 68312
rect 85130 68310 85186 68312
rect 84788 67970 84844 68026
rect 84890 67276 84946 67278
rect 84970 67276 85026 67278
rect 85050 67276 85106 67278
rect 85130 67276 85186 67278
rect 84890 67224 84916 67276
rect 84916 67224 84946 67276
rect 84970 67224 84980 67276
rect 84980 67224 85026 67276
rect 85050 67224 85096 67276
rect 85096 67224 85106 67276
rect 85130 67224 85160 67276
rect 85160 67224 85186 67276
rect 84890 67222 84946 67224
rect 84970 67222 85026 67224
rect 85050 67222 85106 67224
rect 85130 67222 85186 67224
rect 85156 66474 85212 66530
rect 84890 66188 84946 66190
rect 84970 66188 85026 66190
rect 85050 66188 85106 66190
rect 85130 66188 85186 66190
rect 84890 66136 84916 66188
rect 84916 66136 84946 66188
rect 84970 66136 84980 66188
rect 84980 66136 85026 66188
rect 85050 66136 85096 66188
rect 85096 66136 85106 66188
rect 85130 66136 85160 66188
rect 85160 66136 85186 66188
rect 84890 66134 84946 66136
rect 84970 66134 85026 66136
rect 85050 66134 85106 66136
rect 85130 66134 85186 66136
rect 84604 65250 84660 65306
rect 84052 60490 84108 60546
rect 84420 55594 84476 55650
rect 84052 55186 84108 55242
rect 84328 45122 84384 45178
rect 84144 42402 84200 42458
rect 84236 41314 84292 41370
rect 84144 31522 84200 31578
rect 84052 31422 84054 31442
rect 84054 31422 84106 31442
rect 84106 31422 84108 31442
rect 84052 31386 84108 31422
rect 84052 29910 84108 29946
rect 84052 29890 84054 29910
rect 84054 29890 84106 29910
rect 84106 29890 84108 29910
rect 83960 23362 84016 23418
rect 83960 23090 84016 23146
rect 84144 28702 84146 28722
rect 84146 28702 84198 28722
rect 84198 28702 84200 28722
rect 84144 28666 84200 28702
rect 84236 27070 84238 27090
rect 84238 27070 84290 27090
rect 84290 27070 84292 27090
rect 84236 27034 84292 27070
rect 84512 54370 84568 54426
rect 84328 26762 84384 26818
rect 84236 23906 84292 23962
rect 83960 18466 84016 18522
rect 83868 17786 83924 17842
rect 84236 19554 84292 19610
rect 84144 17378 84200 17434
rect 84420 20778 84476 20834
rect 84236 14794 84292 14850
rect 84052 13570 84108 13626
rect 83960 12482 84016 12538
rect 84144 9898 84200 9954
rect 83960 8674 84016 8730
rect 83776 4070 83832 4106
rect 83776 4050 83778 4070
rect 83778 4050 83830 4070
rect 83830 4050 83832 4070
rect 83776 2826 83832 2882
rect 84144 5002 84200 5058
rect 84052 3914 84108 3970
rect 83960 2418 84016 2474
rect 84236 2554 84292 2610
rect 84144 2010 84200 2066
rect 83960 1466 84016 1522
rect 83960 414 83962 434
rect 83962 414 84014 434
rect 84014 414 84016 434
rect 83960 378 84016 414
rect 81200 106 81256 162
rect 84890 65100 84946 65102
rect 84970 65100 85026 65102
rect 85050 65100 85106 65102
rect 85130 65100 85186 65102
rect 84890 65048 84916 65100
rect 84916 65048 84946 65100
rect 84970 65048 84980 65100
rect 84980 65048 85026 65100
rect 85050 65048 85096 65100
rect 85096 65048 85106 65100
rect 85130 65048 85160 65100
rect 85160 65048 85186 65100
rect 84890 65046 84946 65048
rect 84970 65046 85026 65048
rect 85050 65046 85106 65048
rect 85130 65046 85186 65048
rect 84890 64012 84946 64014
rect 84970 64012 85026 64014
rect 85050 64012 85106 64014
rect 85130 64012 85186 64014
rect 84890 63960 84916 64012
rect 84916 63960 84946 64012
rect 84970 63960 84980 64012
rect 84980 63960 85026 64012
rect 85050 63960 85096 64012
rect 85096 63960 85106 64012
rect 85130 63960 85160 64012
rect 85160 63960 85186 64012
rect 84890 63958 84946 63960
rect 84970 63958 85026 63960
rect 85050 63958 85106 63960
rect 85130 63958 85186 63960
rect 84696 63754 84752 63810
rect 84890 62924 84946 62926
rect 84970 62924 85026 62926
rect 85050 62924 85106 62926
rect 85130 62924 85186 62926
rect 84890 62872 84916 62924
rect 84916 62872 84946 62924
rect 84970 62872 84980 62924
rect 84980 62872 85026 62924
rect 85050 62872 85096 62924
rect 85096 62872 85106 62924
rect 85130 62872 85160 62924
rect 85160 62872 85186 62924
rect 84890 62870 84946 62872
rect 84970 62870 85026 62872
rect 85050 62870 85106 62872
rect 85130 62870 85186 62872
rect 84788 62666 84844 62722
rect 84890 61836 84946 61838
rect 84970 61836 85026 61838
rect 85050 61836 85106 61838
rect 85130 61836 85186 61838
rect 84890 61784 84916 61836
rect 84916 61784 84946 61836
rect 84970 61784 84980 61836
rect 84980 61784 85026 61836
rect 85050 61784 85096 61836
rect 85096 61784 85106 61836
rect 85130 61784 85160 61836
rect 85160 61784 85186 61836
rect 84890 61782 84946 61784
rect 84970 61782 85026 61784
rect 85050 61782 85106 61784
rect 85130 61782 85186 61784
rect 84890 60748 84946 60750
rect 84970 60748 85026 60750
rect 85050 60748 85106 60750
rect 85130 60748 85186 60750
rect 84890 60696 84916 60748
rect 84916 60696 84946 60748
rect 84970 60696 84980 60748
rect 84980 60696 85026 60748
rect 85050 60696 85096 60748
rect 85096 60696 85106 60748
rect 85130 60696 85160 60748
rect 85160 60696 85186 60748
rect 84890 60694 84946 60696
rect 84970 60694 85026 60696
rect 85050 60694 85106 60696
rect 85130 60694 85186 60696
rect 84890 59660 84946 59662
rect 84970 59660 85026 59662
rect 85050 59660 85106 59662
rect 85130 59660 85186 59662
rect 84890 59608 84916 59660
rect 84916 59608 84946 59660
rect 84970 59608 84980 59660
rect 84980 59608 85026 59660
rect 85050 59608 85096 59660
rect 85096 59608 85106 59660
rect 85130 59608 85160 59660
rect 85160 59608 85186 59660
rect 84890 59606 84946 59608
rect 84970 59606 85026 59608
rect 85050 59606 85106 59608
rect 85130 59606 85186 59608
rect 84890 58572 84946 58574
rect 84970 58572 85026 58574
rect 85050 58572 85106 58574
rect 85130 58572 85186 58574
rect 84890 58520 84916 58572
rect 84916 58520 84946 58572
rect 84970 58520 84980 58572
rect 84980 58520 85026 58572
rect 85050 58520 85096 58572
rect 85096 58520 85106 58572
rect 85130 58520 85160 58572
rect 85160 58520 85186 58572
rect 84890 58518 84946 58520
rect 84970 58518 85026 58520
rect 85050 58518 85106 58520
rect 85130 58518 85186 58520
rect 84890 57484 84946 57486
rect 84970 57484 85026 57486
rect 85050 57484 85106 57486
rect 85130 57484 85186 57486
rect 84890 57432 84916 57484
rect 84916 57432 84946 57484
rect 84970 57432 84980 57484
rect 84980 57432 85026 57484
rect 85050 57432 85096 57484
rect 85096 57432 85106 57484
rect 85130 57432 85160 57484
rect 85160 57432 85186 57484
rect 84890 57430 84946 57432
rect 84970 57430 85026 57432
rect 85050 57430 85106 57432
rect 85130 57430 85186 57432
rect 84788 56682 84844 56738
rect 84890 56396 84946 56398
rect 84970 56396 85026 56398
rect 85050 56396 85106 56398
rect 85130 56396 85186 56398
rect 84890 56344 84916 56396
rect 84916 56344 84946 56396
rect 84970 56344 84980 56396
rect 84980 56344 85026 56396
rect 85050 56344 85096 56396
rect 85096 56344 85106 56396
rect 85130 56344 85160 56396
rect 85160 56344 85186 56396
rect 84890 56342 84946 56344
rect 84970 56342 85026 56344
rect 85050 56342 85106 56344
rect 85130 56342 85186 56344
rect 84890 55308 84946 55310
rect 84970 55308 85026 55310
rect 85050 55308 85106 55310
rect 85130 55308 85186 55310
rect 84890 55256 84916 55308
rect 84916 55256 84946 55308
rect 84970 55256 84980 55308
rect 84980 55256 85026 55308
rect 85050 55256 85096 55308
rect 85096 55256 85106 55308
rect 85130 55256 85160 55308
rect 85160 55256 85186 55308
rect 84890 55254 84946 55256
rect 84970 55254 85026 55256
rect 85050 55254 85106 55256
rect 85130 55254 85186 55256
rect 84890 54220 84946 54222
rect 84970 54220 85026 54222
rect 85050 54220 85106 54222
rect 85130 54220 85186 54222
rect 84890 54168 84916 54220
rect 84916 54168 84946 54220
rect 84970 54168 84980 54220
rect 84980 54168 85026 54220
rect 85050 54168 85096 54220
rect 85096 54168 85106 54220
rect 85130 54168 85160 54220
rect 85160 54168 85186 54220
rect 84890 54166 84946 54168
rect 84970 54166 85026 54168
rect 85050 54166 85106 54168
rect 85130 54166 85186 54168
rect 84890 53132 84946 53134
rect 84970 53132 85026 53134
rect 85050 53132 85106 53134
rect 85130 53132 85186 53134
rect 84890 53080 84916 53132
rect 84916 53080 84946 53132
rect 84970 53080 84980 53132
rect 84980 53080 85026 53132
rect 85050 53080 85096 53132
rect 85096 53080 85106 53132
rect 85130 53080 85160 53132
rect 85160 53080 85186 53132
rect 84890 53078 84946 53080
rect 84970 53078 85026 53080
rect 85050 53078 85106 53080
rect 85130 53078 85186 53080
rect 84890 52044 84946 52046
rect 84970 52044 85026 52046
rect 85050 52044 85106 52046
rect 85130 52044 85186 52046
rect 84890 51992 84916 52044
rect 84916 51992 84946 52044
rect 84970 51992 84980 52044
rect 84980 51992 85026 52044
rect 85050 51992 85096 52044
rect 85096 51992 85106 52044
rect 85130 51992 85160 52044
rect 85160 51992 85186 52044
rect 84890 51990 84946 51992
rect 84970 51990 85026 51992
rect 85050 51990 85106 51992
rect 85130 51990 85186 51992
rect 84890 50956 84946 50958
rect 84970 50956 85026 50958
rect 85050 50956 85106 50958
rect 85130 50956 85186 50958
rect 84890 50904 84916 50956
rect 84916 50904 84946 50956
rect 84970 50904 84980 50956
rect 84980 50904 85026 50956
rect 85050 50904 85096 50956
rect 85096 50904 85106 50956
rect 85130 50904 85160 50956
rect 85160 50904 85186 50956
rect 84890 50902 84946 50904
rect 84970 50902 85026 50904
rect 85050 50902 85106 50904
rect 85130 50902 85186 50904
rect 85156 50698 85212 50754
rect 84890 49868 84946 49870
rect 84970 49868 85026 49870
rect 85050 49868 85106 49870
rect 85130 49868 85186 49870
rect 84890 49816 84916 49868
rect 84916 49816 84946 49868
rect 84970 49816 84980 49868
rect 84980 49816 85026 49868
rect 85050 49816 85096 49868
rect 85096 49816 85106 49868
rect 85130 49816 85160 49868
rect 85160 49816 85186 49868
rect 84890 49814 84946 49816
rect 84970 49814 85026 49816
rect 85050 49814 85106 49816
rect 85130 49814 85186 49816
rect 84788 49610 84844 49666
rect 84890 48780 84946 48782
rect 84970 48780 85026 48782
rect 85050 48780 85106 48782
rect 85130 48780 85186 48782
rect 84890 48728 84916 48780
rect 84916 48728 84946 48780
rect 84970 48728 84980 48780
rect 84980 48728 85026 48780
rect 85050 48728 85096 48780
rect 85096 48728 85106 48780
rect 85130 48728 85160 48780
rect 85160 48728 85186 48780
rect 84890 48726 84946 48728
rect 84970 48726 85026 48728
rect 85050 48726 85106 48728
rect 85130 48726 85186 48728
rect 84890 47692 84946 47694
rect 84970 47692 85026 47694
rect 85050 47692 85106 47694
rect 85130 47692 85186 47694
rect 84890 47640 84916 47692
rect 84916 47640 84946 47692
rect 84970 47640 84980 47692
rect 84980 47640 85026 47692
rect 85050 47640 85096 47692
rect 85096 47640 85106 47692
rect 85130 47640 85160 47692
rect 85160 47640 85186 47692
rect 84890 47638 84946 47640
rect 84970 47638 85026 47640
rect 85050 47638 85106 47640
rect 85130 47638 85186 47640
rect 84890 46604 84946 46606
rect 84970 46604 85026 46606
rect 85050 46604 85106 46606
rect 85130 46604 85186 46606
rect 84890 46552 84916 46604
rect 84916 46552 84946 46604
rect 84970 46552 84980 46604
rect 84980 46552 85026 46604
rect 85050 46552 85096 46604
rect 85096 46552 85106 46604
rect 85130 46552 85160 46604
rect 85160 46552 85186 46604
rect 84890 46550 84946 46552
rect 84970 46550 85026 46552
rect 85050 46550 85106 46552
rect 85130 46550 85186 46552
rect 84890 45516 84946 45518
rect 84970 45516 85026 45518
rect 85050 45516 85106 45518
rect 85130 45516 85186 45518
rect 84890 45464 84916 45516
rect 84916 45464 84946 45516
rect 84970 45464 84980 45516
rect 84980 45464 85026 45516
rect 85050 45464 85096 45516
rect 85096 45464 85106 45516
rect 85130 45464 85160 45516
rect 85160 45464 85186 45516
rect 84890 45462 84946 45464
rect 84970 45462 85026 45464
rect 85050 45462 85106 45464
rect 85130 45462 85186 45464
rect 84890 44428 84946 44430
rect 84970 44428 85026 44430
rect 85050 44428 85106 44430
rect 85130 44428 85186 44430
rect 84890 44376 84916 44428
rect 84916 44376 84946 44428
rect 84970 44376 84980 44428
rect 84980 44376 85026 44428
rect 85050 44376 85096 44428
rect 85096 44376 85106 44428
rect 85130 44376 85160 44428
rect 85160 44376 85186 44428
rect 84890 44374 84946 44376
rect 84970 44374 85026 44376
rect 85050 44374 85106 44376
rect 85130 44374 85186 44376
rect 85156 43646 85212 43682
rect 85156 43626 85158 43646
rect 85158 43626 85210 43646
rect 85210 43626 85212 43646
rect 84890 43340 84946 43342
rect 84970 43340 85026 43342
rect 85050 43340 85106 43342
rect 85130 43340 85186 43342
rect 84890 43288 84916 43340
rect 84916 43288 84946 43340
rect 84970 43288 84980 43340
rect 84980 43288 85026 43340
rect 85050 43288 85096 43340
rect 85096 43288 85106 43340
rect 85130 43288 85160 43340
rect 85160 43288 85186 43340
rect 84890 43286 84946 43288
rect 84970 43286 85026 43288
rect 85050 43286 85106 43288
rect 85130 43286 85186 43288
rect 84890 42252 84946 42254
rect 84970 42252 85026 42254
rect 85050 42252 85106 42254
rect 85130 42252 85186 42254
rect 84890 42200 84916 42252
rect 84916 42200 84946 42252
rect 84970 42200 84980 42252
rect 84980 42200 85026 42252
rect 85050 42200 85096 42252
rect 85096 42200 85106 42252
rect 85130 42200 85160 42252
rect 85160 42200 85186 42252
rect 84890 42198 84946 42200
rect 84970 42198 85026 42200
rect 85050 42198 85106 42200
rect 85130 42198 85186 42200
rect 84890 41164 84946 41166
rect 84970 41164 85026 41166
rect 85050 41164 85106 41166
rect 85130 41164 85186 41166
rect 84890 41112 84916 41164
rect 84916 41112 84946 41164
rect 84970 41112 84980 41164
rect 84980 41112 85026 41164
rect 85050 41112 85096 41164
rect 85096 41112 85106 41164
rect 85130 41112 85160 41164
rect 85160 41112 85186 41164
rect 84890 41110 84946 41112
rect 84970 41110 85026 41112
rect 85050 41110 85106 41112
rect 85130 41110 85186 41112
rect 84890 40076 84946 40078
rect 84970 40076 85026 40078
rect 85050 40076 85106 40078
rect 85130 40076 85186 40078
rect 84890 40024 84916 40076
rect 84916 40024 84946 40076
rect 84970 40024 84980 40076
rect 84980 40024 85026 40076
rect 85050 40024 85096 40076
rect 85096 40024 85106 40076
rect 85130 40024 85160 40076
rect 85160 40024 85186 40076
rect 84890 40022 84946 40024
rect 84970 40022 85026 40024
rect 85050 40022 85106 40024
rect 85130 40022 85186 40024
rect 84788 39818 84844 39874
rect 84890 38988 84946 38990
rect 84970 38988 85026 38990
rect 85050 38988 85106 38990
rect 85130 38988 85186 38990
rect 84890 38936 84916 38988
rect 84916 38936 84946 38988
rect 84970 38936 84980 38988
rect 84980 38936 85026 38988
rect 85050 38936 85096 38988
rect 85096 38936 85106 38988
rect 85130 38936 85160 38988
rect 85160 38936 85186 38988
rect 84890 38934 84946 38936
rect 84970 38934 85026 38936
rect 85050 38934 85106 38936
rect 85130 38934 85186 38936
rect 84890 37900 84946 37902
rect 84970 37900 85026 37902
rect 85050 37900 85106 37902
rect 85130 37900 85186 37902
rect 84890 37848 84916 37900
rect 84916 37848 84946 37900
rect 84970 37848 84980 37900
rect 84980 37848 85026 37900
rect 85050 37848 85096 37900
rect 85096 37848 85106 37900
rect 85130 37848 85160 37900
rect 85160 37848 85186 37900
rect 84890 37846 84946 37848
rect 84970 37846 85026 37848
rect 85050 37846 85106 37848
rect 85130 37846 85186 37848
rect 84890 36812 84946 36814
rect 84970 36812 85026 36814
rect 85050 36812 85106 36814
rect 85130 36812 85186 36814
rect 84890 36760 84916 36812
rect 84916 36760 84946 36812
rect 84970 36760 84980 36812
rect 84980 36760 85026 36812
rect 85050 36760 85096 36812
rect 85096 36760 85106 36812
rect 85130 36760 85160 36812
rect 85160 36760 85186 36812
rect 84890 36758 84946 36760
rect 84970 36758 85026 36760
rect 85050 36758 85106 36760
rect 85130 36758 85186 36760
rect 84788 36418 84844 36474
rect 84890 35724 84946 35726
rect 84970 35724 85026 35726
rect 85050 35724 85106 35726
rect 85130 35724 85186 35726
rect 84890 35672 84916 35724
rect 84916 35672 84946 35724
rect 84970 35672 84980 35724
rect 84980 35672 85026 35724
rect 85050 35672 85096 35724
rect 85096 35672 85106 35724
rect 85130 35672 85160 35724
rect 85160 35672 85186 35724
rect 84890 35670 84946 35672
rect 84970 35670 85026 35672
rect 85050 35670 85106 35672
rect 85130 35670 85186 35672
rect 84890 34636 84946 34638
rect 84970 34636 85026 34638
rect 85050 34636 85106 34638
rect 85130 34636 85186 34638
rect 84890 34584 84916 34636
rect 84916 34584 84946 34636
rect 84970 34584 84980 34636
rect 84980 34584 85026 34636
rect 85050 34584 85096 34636
rect 85096 34584 85106 34636
rect 85130 34584 85160 34636
rect 85160 34584 85186 34636
rect 84890 34582 84946 34584
rect 84970 34582 85026 34584
rect 85050 34582 85106 34584
rect 85130 34582 85186 34584
rect 84890 33548 84946 33550
rect 84970 33548 85026 33550
rect 85050 33548 85106 33550
rect 85130 33548 85186 33550
rect 84890 33496 84916 33548
rect 84916 33496 84946 33548
rect 84970 33496 84980 33548
rect 84980 33496 85026 33548
rect 85050 33496 85096 33548
rect 85096 33496 85106 33548
rect 85130 33496 85160 33548
rect 85160 33496 85186 33548
rect 84890 33494 84946 33496
rect 84970 33494 85026 33496
rect 85050 33494 85106 33496
rect 85130 33494 85186 33496
rect 84890 32460 84946 32462
rect 84970 32460 85026 32462
rect 85050 32460 85106 32462
rect 85130 32460 85186 32462
rect 84890 32408 84916 32460
rect 84916 32408 84946 32460
rect 84970 32408 84980 32460
rect 84980 32408 85026 32460
rect 85050 32408 85096 32460
rect 85096 32408 85106 32460
rect 85130 32408 85160 32460
rect 85160 32408 85186 32460
rect 84890 32406 84946 32408
rect 84970 32406 85026 32408
rect 85050 32406 85106 32408
rect 85130 32406 85186 32408
rect 84890 31372 84946 31374
rect 84970 31372 85026 31374
rect 85050 31372 85106 31374
rect 85130 31372 85186 31374
rect 84890 31320 84916 31372
rect 84916 31320 84946 31372
rect 84970 31320 84980 31372
rect 84980 31320 85026 31372
rect 85050 31320 85096 31372
rect 85096 31320 85106 31372
rect 85130 31320 85160 31372
rect 85160 31320 85186 31372
rect 84890 31318 84946 31320
rect 84970 31318 85026 31320
rect 85050 31318 85106 31320
rect 85130 31318 85186 31320
rect 84890 30284 84946 30286
rect 84970 30284 85026 30286
rect 85050 30284 85106 30286
rect 85130 30284 85186 30286
rect 84890 30232 84916 30284
rect 84916 30232 84946 30284
rect 84970 30232 84980 30284
rect 84980 30232 85026 30284
rect 85050 30232 85096 30284
rect 85096 30232 85106 30284
rect 85130 30232 85160 30284
rect 85160 30232 85186 30284
rect 84890 30230 84946 30232
rect 84970 30230 85026 30232
rect 85050 30230 85106 30232
rect 85130 30230 85186 30232
rect 84696 29346 84752 29402
rect 84890 29196 84946 29198
rect 84970 29196 85026 29198
rect 85050 29196 85106 29198
rect 85130 29196 85186 29198
rect 84890 29144 84916 29196
rect 84916 29144 84946 29196
rect 84970 29144 84980 29196
rect 84980 29144 85026 29196
rect 85050 29144 85096 29196
rect 85096 29144 85106 29196
rect 85130 29144 85160 29196
rect 85160 29144 85186 29196
rect 84890 29142 84946 29144
rect 84970 29142 85026 29144
rect 85050 29142 85106 29144
rect 85130 29142 85186 29144
rect 84696 28938 84752 28994
rect 84604 28258 84660 28314
rect 84890 28108 84946 28110
rect 84970 28108 85026 28110
rect 85050 28108 85106 28110
rect 85130 28108 85186 28110
rect 84890 28056 84916 28108
rect 84916 28056 84946 28108
rect 84970 28056 84980 28108
rect 84980 28056 85026 28108
rect 85050 28056 85096 28108
rect 85096 28056 85106 28108
rect 85130 28056 85160 28108
rect 85160 28056 85186 28108
rect 84890 28054 84946 28056
rect 84970 28054 85026 28056
rect 85050 28054 85106 28056
rect 85130 28054 85186 28056
rect 84604 24450 84660 24506
rect 84890 27020 84946 27022
rect 84970 27020 85026 27022
rect 85050 27020 85106 27022
rect 85130 27020 85186 27022
rect 84890 26968 84916 27020
rect 84916 26968 84946 27020
rect 84970 26968 84980 27020
rect 84980 26968 85026 27020
rect 85050 26968 85096 27020
rect 85096 26968 85106 27020
rect 85130 26968 85160 27020
rect 85160 26968 85186 27020
rect 84890 26966 84946 26968
rect 84970 26966 85026 26968
rect 85050 26966 85106 26968
rect 85130 26966 85186 26968
rect 84890 25932 84946 25934
rect 84970 25932 85026 25934
rect 85050 25932 85106 25934
rect 85130 25932 85186 25934
rect 84890 25880 84916 25932
rect 84916 25880 84946 25932
rect 84970 25880 84980 25932
rect 84980 25880 85026 25932
rect 85050 25880 85096 25932
rect 85096 25880 85106 25932
rect 85130 25880 85160 25932
rect 85160 25880 85186 25932
rect 84890 25878 84946 25880
rect 84970 25878 85026 25880
rect 85050 25878 85106 25880
rect 85130 25878 85186 25880
rect 84880 25574 84882 25594
rect 84882 25574 84934 25594
rect 84934 25574 84936 25594
rect 84880 25538 84936 25574
rect 84890 24844 84946 24846
rect 84970 24844 85026 24846
rect 85050 24844 85106 24846
rect 85130 24844 85186 24846
rect 84890 24792 84916 24844
rect 84916 24792 84946 24844
rect 84970 24792 84980 24844
rect 84980 24792 85026 24844
rect 85050 24792 85096 24844
rect 85096 24792 85106 24844
rect 85130 24792 85160 24844
rect 85160 24792 85186 24844
rect 84890 24790 84946 24792
rect 84970 24790 85026 24792
rect 85050 24790 85106 24792
rect 85130 24790 85186 24792
rect 84696 24178 84752 24234
rect 84890 23756 84946 23758
rect 84970 23756 85026 23758
rect 85050 23756 85106 23758
rect 85130 23756 85186 23758
rect 84890 23704 84916 23756
rect 84916 23704 84946 23756
rect 84970 23704 84980 23756
rect 84980 23704 85026 23756
rect 85050 23704 85096 23756
rect 85096 23704 85106 23756
rect 85130 23704 85160 23756
rect 85160 23704 85186 23756
rect 84890 23702 84946 23704
rect 84970 23702 85026 23704
rect 85050 23702 85106 23704
rect 85130 23702 85186 23704
rect 84890 22668 84946 22670
rect 84970 22668 85026 22670
rect 85050 22668 85106 22670
rect 85130 22668 85186 22670
rect 84890 22616 84916 22668
rect 84916 22616 84946 22668
rect 84970 22616 84980 22668
rect 84980 22616 85026 22668
rect 85050 22616 85096 22668
rect 85096 22616 85106 22668
rect 85130 22616 85160 22668
rect 85160 22616 85186 22668
rect 84890 22614 84946 22616
rect 84970 22614 85026 22616
rect 85050 22614 85106 22616
rect 85130 22614 85186 22616
rect 84890 21580 84946 21582
rect 84970 21580 85026 21582
rect 85050 21580 85106 21582
rect 85130 21580 85186 21582
rect 84890 21528 84916 21580
rect 84916 21528 84946 21580
rect 84970 21528 84980 21580
rect 84980 21528 85026 21580
rect 85050 21528 85096 21580
rect 85096 21528 85106 21580
rect 85130 21528 85160 21580
rect 85160 21528 85186 21580
rect 84890 21526 84946 21528
rect 84970 21526 85026 21528
rect 85050 21526 85106 21528
rect 85130 21526 85186 21528
rect 84890 20492 84946 20494
rect 84970 20492 85026 20494
rect 85050 20492 85106 20494
rect 85130 20492 85186 20494
rect 84890 20440 84916 20492
rect 84916 20440 84946 20492
rect 84970 20440 84980 20492
rect 84980 20440 85026 20492
rect 85050 20440 85096 20492
rect 85096 20440 85106 20492
rect 85130 20440 85160 20492
rect 85160 20440 85186 20492
rect 84890 20438 84946 20440
rect 84970 20438 85026 20440
rect 85050 20438 85106 20440
rect 85130 20438 85186 20440
rect 84890 19404 84946 19406
rect 84970 19404 85026 19406
rect 85050 19404 85106 19406
rect 85130 19404 85186 19406
rect 84890 19352 84916 19404
rect 84916 19352 84946 19404
rect 84970 19352 84980 19404
rect 84980 19352 85026 19404
rect 85050 19352 85096 19404
rect 85096 19352 85106 19404
rect 85130 19352 85160 19404
rect 85160 19352 85186 19404
rect 84890 19350 84946 19352
rect 84970 19350 85026 19352
rect 85050 19350 85106 19352
rect 85130 19350 85186 19352
rect 84890 18316 84946 18318
rect 84970 18316 85026 18318
rect 85050 18316 85106 18318
rect 85130 18316 85186 18318
rect 84890 18264 84916 18316
rect 84916 18264 84946 18316
rect 84970 18264 84980 18316
rect 84980 18264 85026 18316
rect 85050 18264 85096 18316
rect 85096 18264 85106 18316
rect 85130 18264 85160 18316
rect 85160 18264 85186 18316
rect 84890 18262 84946 18264
rect 84970 18262 85026 18264
rect 85050 18262 85106 18264
rect 85130 18262 85186 18264
rect 84890 17228 84946 17230
rect 84970 17228 85026 17230
rect 85050 17228 85106 17230
rect 85130 17228 85186 17230
rect 84890 17176 84916 17228
rect 84916 17176 84946 17228
rect 84970 17176 84980 17228
rect 84980 17176 85026 17228
rect 85050 17176 85096 17228
rect 85096 17176 85106 17228
rect 85130 17176 85160 17228
rect 85160 17176 85186 17228
rect 84890 17174 84946 17176
rect 84970 17174 85026 17176
rect 85050 17174 85106 17176
rect 85130 17174 85186 17176
rect 84880 16290 84936 16346
rect 84890 16140 84946 16142
rect 84970 16140 85026 16142
rect 85050 16140 85106 16142
rect 85130 16140 85186 16142
rect 84890 16088 84916 16140
rect 84916 16088 84946 16140
rect 84970 16088 84980 16140
rect 84980 16088 85026 16140
rect 85050 16088 85096 16140
rect 85096 16088 85106 16140
rect 85130 16088 85160 16140
rect 85160 16088 85186 16140
rect 84890 16086 84946 16088
rect 84970 16086 85026 16088
rect 85050 16086 85106 16088
rect 85130 16086 85186 16088
rect 84890 15052 84946 15054
rect 84970 15052 85026 15054
rect 85050 15052 85106 15054
rect 85130 15052 85186 15054
rect 84890 15000 84916 15052
rect 84916 15000 84946 15052
rect 84970 15000 84980 15052
rect 84980 15000 85026 15052
rect 85050 15000 85096 15052
rect 85096 15000 85106 15052
rect 85130 15000 85160 15052
rect 85160 15000 85186 15052
rect 84890 14998 84946 15000
rect 84970 14998 85026 15000
rect 85050 14998 85106 15000
rect 85130 14998 85186 15000
rect 84890 13964 84946 13966
rect 84970 13964 85026 13966
rect 85050 13964 85106 13966
rect 85130 13964 85186 13966
rect 84890 13912 84916 13964
rect 84916 13912 84946 13964
rect 84970 13912 84980 13964
rect 84980 13912 85026 13964
rect 85050 13912 85096 13964
rect 85096 13912 85106 13964
rect 85130 13912 85160 13964
rect 85160 13912 85186 13964
rect 84890 13910 84946 13912
rect 84970 13910 85026 13912
rect 85050 13910 85106 13912
rect 85130 13910 85186 13912
rect 84890 12876 84946 12878
rect 84970 12876 85026 12878
rect 85050 12876 85106 12878
rect 85130 12876 85186 12878
rect 84890 12824 84916 12876
rect 84916 12824 84946 12876
rect 84970 12824 84980 12876
rect 84980 12824 85026 12876
rect 85050 12824 85096 12876
rect 85096 12824 85106 12876
rect 85130 12824 85160 12876
rect 85160 12824 85186 12876
rect 84890 12822 84946 12824
rect 84970 12822 85026 12824
rect 85050 12822 85106 12824
rect 85130 12822 85186 12824
rect 84890 11788 84946 11790
rect 84970 11788 85026 11790
rect 85050 11788 85106 11790
rect 85130 11788 85186 11790
rect 84890 11736 84916 11788
rect 84916 11736 84946 11788
rect 84970 11736 84980 11788
rect 84980 11736 85026 11788
rect 85050 11736 85096 11788
rect 85096 11736 85106 11788
rect 85130 11736 85160 11788
rect 85160 11736 85186 11788
rect 84890 11734 84946 11736
rect 84970 11734 85026 11736
rect 85050 11734 85106 11736
rect 85130 11734 85186 11736
rect 84890 10700 84946 10702
rect 84970 10700 85026 10702
rect 85050 10700 85106 10702
rect 85130 10700 85186 10702
rect 84890 10648 84916 10700
rect 84916 10648 84946 10700
rect 84970 10648 84980 10700
rect 84980 10648 85026 10700
rect 85050 10648 85096 10700
rect 85096 10648 85106 10700
rect 85130 10648 85160 10700
rect 85160 10648 85186 10700
rect 84890 10646 84946 10648
rect 84970 10646 85026 10648
rect 85050 10646 85106 10648
rect 85130 10646 85186 10648
rect 84890 9612 84946 9614
rect 84970 9612 85026 9614
rect 85050 9612 85106 9614
rect 85130 9612 85186 9614
rect 84890 9560 84916 9612
rect 84916 9560 84946 9612
rect 84970 9560 84980 9612
rect 84980 9560 85026 9612
rect 85050 9560 85096 9612
rect 85096 9560 85106 9612
rect 85130 9560 85160 9612
rect 85160 9560 85186 9612
rect 84890 9558 84946 9560
rect 84970 9558 85026 9560
rect 85050 9558 85106 9560
rect 85130 9558 85186 9560
rect 84890 8524 84946 8526
rect 84970 8524 85026 8526
rect 85050 8524 85106 8526
rect 85130 8524 85186 8526
rect 84890 8472 84916 8524
rect 84916 8472 84946 8524
rect 84970 8472 84980 8524
rect 84980 8472 85026 8524
rect 85050 8472 85096 8524
rect 85096 8472 85106 8524
rect 85130 8472 85160 8524
rect 85160 8472 85186 8524
rect 84890 8470 84946 8472
rect 84970 8470 85026 8472
rect 85050 8470 85106 8472
rect 85130 8470 85186 8472
rect 85064 7606 85120 7642
rect 85064 7586 85066 7606
rect 85066 7586 85118 7606
rect 85118 7586 85120 7606
rect 84890 7436 84946 7438
rect 84970 7436 85026 7438
rect 85050 7436 85106 7438
rect 85130 7436 85186 7438
rect 84890 7384 84916 7436
rect 84916 7384 84946 7436
rect 84970 7384 84980 7436
rect 84980 7384 85026 7436
rect 85050 7384 85096 7436
rect 85096 7384 85106 7436
rect 85130 7384 85160 7436
rect 85160 7384 85186 7436
rect 84890 7382 84946 7384
rect 84970 7382 85026 7384
rect 85050 7382 85106 7384
rect 85130 7382 85186 7384
rect 84512 6498 84568 6554
rect 84512 1874 84568 1930
rect 84890 6348 84946 6350
rect 84970 6348 85026 6350
rect 85050 6348 85106 6350
rect 85130 6348 85186 6350
rect 84890 6296 84916 6348
rect 84916 6296 84946 6348
rect 84970 6296 84980 6348
rect 84980 6296 85026 6348
rect 85050 6296 85096 6348
rect 85096 6296 85106 6348
rect 85130 6296 85160 6348
rect 85160 6296 85186 6348
rect 84890 6294 84946 6296
rect 84970 6294 85026 6296
rect 85050 6294 85106 6296
rect 85130 6294 85186 6296
rect 84890 5260 84946 5262
rect 84970 5260 85026 5262
rect 85050 5260 85106 5262
rect 85130 5260 85186 5262
rect 84890 5208 84916 5260
rect 84916 5208 84946 5260
rect 84970 5208 84980 5260
rect 84980 5208 85026 5260
rect 85050 5208 85096 5260
rect 85096 5208 85106 5260
rect 85130 5208 85160 5260
rect 85160 5208 85186 5260
rect 84890 5206 84946 5208
rect 84970 5206 85026 5208
rect 85050 5206 85106 5208
rect 85130 5206 85186 5208
rect 84890 4172 84946 4174
rect 84970 4172 85026 4174
rect 85050 4172 85106 4174
rect 85130 4172 85186 4174
rect 84890 4120 84916 4172
rect 84916 4120 84946 4172
rect 84970 4120 84980 4172
rect 84980 4120 85026 4172
rect 85050 4120 85096 4172
rect 85096 4120 85106 4172
rect 85130 4120 85160 4172
rect 85160 4120 85186 4172
rect 84890 4118 84946 4120
rect 84970 4118 85026 4120
rect 85050 4118 85106 4120
rect 85130 4118 85186 4120
rect 84890 3084 84946 3086
rect 84970 3084 85026 3086
rect 85050 3084 85106 3086
rect 85130 3084 85186 3086
rect 84890 3032 84916 3084
rect 84916 3032 84946 3084
rect 84970 3032 84980 3084
rect 84980 3032 85026 3084
rect 85050 3032 85096 3084
rect 85096 3032 85106 3084
rect 85130 3032 85160 3084
rect 85160 3032 85186 3084
rect 84890 3030 84946 3032
rect 84970 3030 85026 3032
rect 85050 3030 85106 3032
rect 85130 3030 85186 3032
rect 85800 48386 85856 48442
rect 85524 19590 85526 19610
rect 85526 19590 85578 19610
rect 85578 19590 85580 19610
rect 85524 19554 85580 19590
rect 84890 1996 84946 1998
rect 84970 1996 85026 1998
rect 85050 1996 85106 1998
rect 85130 1996 85186 1998
rect 84890 1944 84916 1996
rect 84916 1944 84946 1996
rect 84970 1944 84980 1996
rect 84980 1944 85026 1996
rect 85050 1944 85096 1996
rect 85096 1944 85106 1996
rect 85130 1944 85160 1996
rect 85160 1944 85186 1996
rect 84890 1942 84946 1944
rect 84970 1942 85026 1944
rect 85050 1942 85106 1944
rect 85130 1942 85186 1944
rect 85892 45802 85948 45858
rect 85984 10986 86040 11042
rect 86890 96108 86946 96110
rect 86970 96108 87026 96110
rect 87050 96108 87106 96110
rect 87130 96108 87186 96110
rect 86890 96056 86916 96108
rect 86916 96056 86946 96108
rect 86970 96056 86980 96108
rect 86980 96056 87026 96108
rect 87050 96056 87096 96108
rect 87096 96056 87106 96108
rect 87130 96056 87160 96108
rect 87160 96056 87186 96108
rect 86890 96054 86946 96056
rect 86970 96054 87026 96056
rect 87050 96054 87106 96056
rect 87130 96054 87186 96056
rect 86890 95020 86946 95022
rect 86970 95020 87026 95022
rect 87050 95020 87106 95022
rect 87130 95020 87186 95022
rect 86890 94968 86916 95020
rect 86916 94968 86946 95020
rect 86970 94968 86980 95020
rect 86980 94968 87026 95020
rect 87050 94968 87096 95020
rect 87096 94968 87106 95020
rect 87130 94968 87160 95020
rect 87160 94968 87186 95020
rect 86890 94966 86946 94968
rect 86970 94966 87026 94968
rect 87050 94966 87106 94968
rect 87130 94966 87186 94968
rect 86890 93932 86946 93934
rect 86970 93932 87026 93934
rect 87050 93932 87106 93934
rect 87130 93932 87186 93934
rect 86890 93880 86916 93932
rect 86916 93880 86946 93932
rect 86970 93880 86980 93932
rect 86980 93880 87026 93932
rect 87050 93880 87096 93932
rect 87096 93880 87106 93932
rect 87130 93880 87160 93932
rect 87160 93880 87186 93932
rect 86890 93878 86946 93880
rect 86970 93878 87026 93880
rect 87050 93878 87106 93880
rect 87130 93878 87186 93880
rect 86890 92844 86946 92846
rect 86970 92844 87026 92846
rect 87050 92844 87106 92846
rect 87130 92844 87186 92846
rect 86890 92792 86916 92844
rect 86916 92792 86946 92844
rect 86970 92792 86980 92844
rect 86980 92792 87026 92844
rect 87050 92792 87096 92844
rect 87096 92792 87106 92844
rect 87130 92792 87160 92844
rect 87160 92792 87186 92844
rect 86890 92790 86946 92792
rect 86970 92790 87026 92792
rect 87050 92790 87106 92792
rect 87130 92790 87186 92792
rect 86890 91756 86946 91758
rect 86970 91756 87026 91758
rect 87050 91756 87106 91758
rect 87130 91756 87186 91758
rect 86890 91704 86916 91756
rect 86916 91704 86946 91756
rect 86970 91704 86980 91756
rect 86980 91704 87026 91756
rect 87050 91704 87096 91756
rect 87096 91704 87106 91756
rect 87130 91704 87160 91756
rect 87160 91704 87186 91756
rect 86890 91702 86946 91704
rect 86970 91702 87026 91704
rect 87050 91702 87106 91704
rect 87130 91702 87186 91704
rect 86890 90668 86946 90670
rect 86970 90668 87026 90670
rect 87050 90668 87106 90670
rect 87130 90668 87186 90670
rect 86890 90616 86916 90668
rect 86916 90616 86946 90668
rect 86970 90616 86980 90668
rect 86980 90616 87026 90668
rect 87050 90616 87096 90668
rect 87096 90616 87106 90668
rect 87130 90616 87160 90668
rect 87160 90616 87186 90668
rect 86890 90614 86946 90616
rect 86970 90614 87026 90616
rect 87050 90614 87106 90616
rect 87130 90614 87186 90616
rect 86890 89580 86946 89582
rect 86970 89580 87026 89582
rect 87050 89580 87106 89582
rect 87130 89580 87186 89582
rect 86890 89528 86916 89580
rect 86916 89528 86946 89580
rect 86970 89528 86980 89580
rect 86980 89528 87026 89580
rect 87050 89528 87096 89580
rect 87096 89528 87106 89580
rect 87130 89528 87160 89580
rect 87160 89528 87186 89580
rect 86890 89526 86946 89528
rect 86970 89526 87026 89528
rect 87050 89526 87106 89528
rect 87130 89526 87186 89528
rect 86890 88492 86946 88494
rect 86970 88492 87026 88494
rect 87050 88492 87106 88494
rect 87130 88492 87186 88494
rect 86890 88440 86916 88492
rect 86916 88440 86946 88492
rect 86970 88440 86980 88492
rect 86980 88440 87026 88492
rect 87050 88440 87096 88492
rect 87096 88440 87106 88492
rect 87130 88440 87160 88492
rect 87160 88440 87186 88492
rect 86890 88438 86946 88440
rect 86970 88438 87026 88440
rect 87050 88438 87106 88440
rect 87130 88438 87186 88440
rect 86890 87404 86946 87406
rect 86970 87404 87026 87406
rect 87050 87404 87106 87406
rect 87130 87404 87186 87406
rect 86890 87352 86916 87404
rect 86916 87352 86946 87404
rect 86970 87352 86980 87404
rect 86980 87352 87026 87404
rect 87050 87352 87096 87404
rect 87096 87352 87106 87404
rect 87130 87352 87160 87404
rect 87160 87352 87186 87404
rect 86890 87350 86946 87352
rect 86970 87350 87026 87352
rect 87050 87350 87106 87352
rect 87130 87350 87186 87352
rect 86890 86316 86946 86318
rect 86970 86316 87026 86318
rect 87050 86316 87106 86318
rect 87130 86316 87186 86318
rect 86890 86264 86916 86316
rect 86916 86264 86946 86316
rect 86970 86264 86980 86316
rect 86980 86264 87026 86316
rect 87050 86264 87096 86316
rect 87096 86264 87106 86316
rect 87130 86264 87160 86316
rect 87160 86264 87186 86316
rect 86890 86262 86946 86264
rect 86970 86262 87026 86264
rect 87050 86262 87106 86264
rect 87130 86262 87186 86264
rect 86890 85228 86946 85230
rect 86970 85228 87026 85230
rect 87050 85228 87106 85230
rect 87130 85228 87186 85230
rect 86890 85176 86916 85228
rect 86916 85176 86946 85228
rect 86970 85176 86980 85228
rect 86980 85176 87026 85228
rect 87050 85176 87096 85228
rect 87096 85176 87106 85228
rect 87130 85176 87160 85228
rect 87160 85176 87186 85228
rect 86890 85174 86946 85176
rect 86970 85174 87026 85176
rect 87050 85174 87106 85176
rect 87130 85174 87186 85176
rect 86890 84140 86946 84142
rect 86970 84140 87026 84142
rect 87050 84140 87106 84142
rect 87130 84140 87186 84142
rect 86890 84088 86916 84140
rect 86916 84088 86946 84140
rect 86970 84088 86980 84140
rect 86980 84088 87026 84140
rect 87050 84088 87096 84140
rect 87096 84088 87106 84140
rect 87130 84088 87160 84140
rect 87160 84088 87186 84140
rect 86890 84086 86946 84088
rect 86970 84086 87026 84088
rect 87050 84086 87106 84088
rect 87130 84086 87186 84088
rect 86890 83052 86946 83054
rect 86970 83052 87026 83054
rect 87050 83052 87106 83054
rect 87130 83052 87186 83054
rect 86890 83000 86916 83052
rect 86916 83000 86946 83052
rect 86970 83000 86980 83052
rect 86980 83000 87026 83052
rect 87050 83000 87096 83052
rect 87096 83000 87106 83052
rect 87130 83000 87160 83052
rect 87160 83000 87186 83052
rect 86890 82998 86946 83000
rect 86970 82998 87026 83000
rect 87050 82998 87106 83000
rect 87130 82998 87186 83000
rect 86890 81964 86946 81966
rect 86970 81964 87026 81966
rect 87050 81964 87106 81966
rect 87130 81964 87186 81966
rect 86890 81912 86916 81964
rect 86916 81912 86946 81964
rect 86970 81912 86980 81964
rect 86980 81912 87026 81964
rect 87050 81912 87096 81964
rect 87096 81912 87106 81964
rect 87130 81912 87160 81964
rect 87160 81912 87186 81964
rect 86890 81910 86946 81912
rect 86970 81910 87026 81912
rect 87050 81910 87106 81912
rect 87130 81910 87186 81912
rect 86890 80876 86946 80878
rect 86970 80876 87026 80878
rect 87050 80876 87106 80878
rect 87130 80876 87186 80878
rect 86890 80824 86916 80876
rect 86916 80824 86946 80876
rect 86970 80824 86980 80876
rect 86980 80824 87026 80876
rect 87050 80824 87096 80876
rect 87096 80824 87106 80876
rect 87130 80824 87160 80876
rect 87160 80824 87186 80876
rect 86890 80822 86946 80824
rect 86970 80822 87026 80824
rect 87050 80822 87106 80824
rect 87130 80822 87186 80824
rect 86890 79788 86946 79790
rect 86970 79788 87026 79790
rect 87050 79788 87106 79790
rect 87130 79788 87186 79790
rect 86890 79736 86916 79788
rect 86916 79736 86946 79788
rect 86970 79736 86980 79788
rect 86980 79736 87026 79788
rect 87050 79736 87096 79788
rect 87096 79736 87106 79788
rect 87130 79736 87160 79788
rect 87160 79736 87186 79788
rect 86890 79734 86946 79736
rect 86970 79734 87026 79736
rect 87050 79734 87106 79736
rect 87130 79734 87186 79736
rect 86890 78700 86946 78702
rect 86970 78700 87026 78702
rect 87050 78700 87106 78702
rect 87130 78700 87186 78702
rect 86890 78648 86916 78700
rect 86916 78648 86946 78700
rect 86970 78648 86980 78700
rect 86980 78648 87026 78700
rect 87050 78648 87096 78700
rect 87096 78648 87106 78700
rect 87130 78648 87160 78700
rect 87160 78648 87186 78700
rect 86890 78646 86946 78648
rect 86970 78646 87026 78648
rect 87050 78646 87106 78648
rect 87130 78646 87186 78648
rect 86890 77612 86946 77614
rect 86970 77612 87026 77614
rect 87050 77612 87106 77614
rect 87130 77612 87186 77614
rect 86890 77560 86916 77612
rect 86916 77560 86946 77612
rect 86970 77560 86980 77612
rect 86980 77560 87026 77612
rect 87050 77560 87096 77612
rect 87096 77560 87106 77612
rect 87130 77560 87160 77612
rect 87160 77560 87186 77612
rect 86890 77558 86946 77560
rect 86970 77558 87026 77560
rect 87050 77558 87106 77560
rect 87130 77558 87186 77560
rect 86890 76524 86946 76526
rect 86970 76524 87026 76526
rect 87050 76524 87106 76526
rect 87130 76524 87186 76526
rect 86890 76472 86916 76524
rect 86916 76472 86946 76524
rect 86970 76472 86980 76524
rect 86980 76472 87026 76524
rect 87050 76472 87096 76524
rect 87096 76472 87106 76524
rect 87130 76472 87160 76524
rect 87160 76472 87186 76524
rect 86890 76470 86946 76472
rect 86970 76470 87026 76472
rect 87050 76470 87106 76472
rect 87130 76470 87186 76472
rect 86890 75436 86946 75438
rect 86970 75436 87026 75438
rect 87050 75436 87106 75438
rect 87130 75436 87186 75438
rect 86890 75384 86916 75436
rect 86916 75384 86946 75436
rect 86970 75384 86980 75436
rect 86980 75384 87026 75436
rect 87050 75384 87096 75436
rect 87096 75384 87106 75436
rect 87130 75384 87160 75436
rect 87160 75384 87186 75436
rect 86890 75382 86946 75384
rect 86970 75382 87026 75384
rect 87050 75382 87106 75384
rect 87130 75382 87186 75384
rect 86890 74348 86946 74350
rect 86970 74348 87026 74350
rect 87050 74348 87106 74350
rect 87130 74348 87186 74350
rect 86890 74296 86916 74348
rect 86916 74296 86946 74348
rect 86970 74296 86980 74348
rect 86980 74296 87026 74348
rect 87050 74296 87096 74348
rect 87096 74296 87106 74348
rect 87130 74296 87160 74348
rect 87160 74296 87186 74348
rect 86890 74294 86946 74296
rect 86970 74294 87026 74296
rect 87050 74294 87106 74296
rect 87130 74294 87186 74296
rect 86890 73260 86946 73262
rect 86970 73260 87026 73262
rect 87050 73260 87106 73262
rect 87130 73260 87186 73262
rect 86890 73208 86916 73260
rect 86916 73208 86946 73260
rect 86970 73208 86980 73260
rect 86980 73208 87026 73260
rect 87050 73208 87096 73260
rect 87096 73208 87106 73260
rect 87130 73208 87160 73260
rect 87160 73208 87186 73260
rect 86890 73206 86946 73208
rect 86970 73206 87026 73208
rect 87050 73206 87106 73208
rect 87130 73206 87186 73208
rect 86890 72172 86946 72174
rect 86970 72172 87026 72174
rect 87050 72172 87106 72174
rect 87130 72172 87186 72174
rect 86890 72120 86916 72172
rect 86916 72120 86946 72172
rect 86970 72120 86980 72172
rect 86980 72120 87026 72172
rect 87050 72120 87096 72172
rect 87096 72120 87106 72172
rect 87130 72120 87160 72172
rect 87160 72120 87186 72172
rect 86890 72118 86946 72120
rect 86970 72118 87026 72120
rect 87050 72118 87106 72120
rect 87130 72118 87186 72120
rect 86890 71084 86946 71086
rect 86970 71084 87026 71086
rect 87050 71084 87106 71086
rect 87130 71084 87186 71086
rect 86890 71032 86916 71084
rect 86916 71032 86946 71084
rect 86970 71032 86980 71084
rect 86980 71032 87026 71084
rect 87050 71032 87096 71084
rect 87096 71032 87106 71084
rect 87130 71032 87160 71084
rect 87160 71032 87186 71084
rect 86890 71030 86946 71032
rect 86970 71030 87026 71032
rect 87050 71030 87106 71032
rect 87130 71030 87186 71032
rect 86890 69996 86946 69998
rect 86970 69996 87026 69998
rect 87050 69996 87106 69998
rect 87130 69996 87186 69998
rect 86890 69944 86916 69996
rect 86916 69944 86946 69996
rect 86970 69944 86980 69996
rect 86980 69944 87026 69996
rect 87050 69944 87096 69996
rect 87096 69944 87106 69996
rect 87130 69944 87160 69996
rect 87160 69944 87186 69996
rect 86890 69942 86946 69944
rect 86970 69942 87026 69944
rect 87050 69942 87106 69944
rect 87130 69942 87186 69944
rect 86890 68908 86946 68910
rect 86970 68908 87026 68910
rect 87050 68908 87106 68910
rect 87130 68908 87186 68910
rect 86890 68856 86916 68908
rect 86916 68856 86946 68908
rect 86970 68856 86980 68908
rect 86980 68856 87026 68908
rect 87050 68856 87096 68908
rect 87096 68856 87106 68908
rect 87130 68856 87160 68908
rect 87160 68856 87186 68908
rect 86890 68854 86946 68856
rect 86970 68854 87026 68856
rect 87050 68854 87106 68856
rect 87130 68854 87186 68856
rect 86890 67820 86946 67822
rect 86970 67820 87026 67822
rect 87050 67820 87106 67822
rect 87130 67820 87186 67822
rect 86890 67768 86916 67820
rect 86916 67768 86946 67820
rect 86970 67768 86980 67820
rect 86980 67768 87026 67820
rect 87050 67768 87096 67820
rect 87096 67768 87106 67820
rect 87130 67768 87160 67820
rect 87160 67768 87186 67820
rect 86890 67766 86946 67768
rect 86970 67766 87026 67768
rect 87050 67766 87106 67768
rect 87130 67766 87186 67768
rect 86890 66732 86946 66734
rect 86970 66732 87026 66734
rect 87050 66732 87106 66734
rect 87130 66732 87186 66734
rect 86890 66680 86916 66732
rect 86916 66680 86946 66732
rect 86970 66680 86980 66732
rect 86980 66680 87026 66732
rect 87050 66680 87096 66732
rect 87096 66680 87106 66732
rect 87130 66680 87160 66732
rect 87160 66680 87186 66732
rect 86890 66678 86946 66680
rect 86970 66678 87026 66680
rect 87050 66678 87106 66680
rect 87130 66678 87186 66680
rect 86890 65644 86946 65646
rect 86970 65644 87026 65646
rect 87050 65644 87106 65646
rect 87130 65644 87186 65646
rect 86890 65592 86916 65644
rect 86916 65592 86946 65644
rect 86970 65592 86980 65644
rect 86980 65592 87026 65644
rect 87050 65592 87096 65644
rect 87096 65592 87106 65644
rect 87130 65592 87160 65644
rect 87160 65592 87186 65644
rect 86890 65590 86946 65592
rect 86970 65590 87026 65592
rect 87050 65590 87106 65592
rect 87130 65590 87186 65592
rect 86890 64556 86946 64558
rect 86970 64556 87026 64558
rect 87050 64556 87106 64558
rect 87130 64556 87186 64558
rect 86890 64504 86916 64556
rect 86916 64504 86946 64556
rect 86970 64504 86980 64556
rect 86980 64504 87026 64556
rect 87050 64504 87096 64556
rect 87096 64504 87106 64556
rect 87130 64504 87160 64556
rect 87160 64504 87186 64556
rect 86890 64502 86946 64504
rect 86970 64502 87026 64504
rect 87050 64502 87106 64504
rect 87130 64502 87186 64504
rect 86890 63468 86946 63470
rect 86970 63468 87026 63470
rect 87050 63468 87106 63470
rect 87130 63468 87186 63470
rect 86890 63416 86916 63468
rect 86916 63416 86946 63468
rect 86970 63416 86980 63468
rect 86980 63416 87026 63468
rect 87050 63416 87096 63468
rect 87096 63416 87106 63468
rect 87130 63416 87160 63468
rect 87160 63416 87186 63468
rect 86890 63414 86946 63416
rect 86970 63414 87026 63416
rect 87050 63414 87106 63416
rect 87130 63414 87186 63416
rect 86890 62380 86946 62382
rect 86970 62380 87026 62382
rect 87050 62380 87106 62382
rect 87130 62380 87186 62382
rect 86890 62328 86916 62380
rect 86916 62328 86946 62380
rect 86970 62328 86980 62380
rect 86980 62328 87026 62380
rect 87050 62328 87096 62380
rect 87096 62328 87106 62380
rect 87130 62328 87160 62380
rect 87160 62328 87186 62380
rect 86890 62326 86946 62328
rect 86970 62326 87026 62328
rect 87050 62326 87106 62328
rect 87130 62326 87186 62328
rect 86890 61292 86946 61294
rect 86970 61292 87026 61294
rect 87050 61292 87106 61294
rect 87130 61292 87186 61294
rect 86890 61240 86916 61292
rect 86916 61240 86946 61292
rect 86970 61240 86980 61292
rect 86980 61240 87026 61292
rect 87050 61240 87096 61292
rect 87096 61240 87106 61292
rect 87130 61240 87160 61292
rect 87160 61240 87186 61292
rect 86890 61238 86946 61240
rect 86970 61238 87026 61240
rect 87050 61238 87106 61240
rect 87130 61238 87186 61240
rect 86890 60204 86946 60206
rect 86970 60204 87026 60206
rect 87050 60204 87106 60206
rect 87130 60204 87186 60206
rect 86890 60152 86916 60204
rect 86916 60152 86946 60204
rect 86970 60152 86980 60204
rect 86980 60152 87026 60204
rect 87050 60152 87096 60204
rect 87096 60152 87106 60204
rect 87130 60152 87160 60204
rect 87160 60152 87186 60204
rect 86890 60150 86946 60152
rect 86970 60150 87026 60152
rect 87050 60150 87106 60152
rect 87130 60150 87186 60152
rect 86890 59116 86946 59118
rect 86970 59116 87026 59118
rect 87050 59116 87106 59118
rect 87130 59116 87186 59118
rect 86890 59064 86916 59116
rect 86916 59064 86946 59116
rect 86970 59064 86980 59116
rect 86980 59064 87026 59116
rect 87050 59064 87096 59116
rect 87096 59064 87106 59116
rect 87130 59064 87160 59116
rect 87160 59064 87186 59116
rect 86890 59062 86946 59064
rect 86970 59062 87026 59064
rect 87050 59062 87106 59064
rect 87130 59062 87186 59064
rect 86890 58028 86946 58030
rect 86970 58028 87026 58030
rect 87050 58028 87106 58030
rect 87130 58028 87186 58030
rect 86890 57976 86916 58028
rect 86916 57976 86946 58028
rect 86970 57976 86980 58028
rect 86980 57976 87026 58028
rect 87050 57976 87096 58028
rect 87096 57976 87106 58028
rect 87130 57976 87160 58028
rect 87160 57976 87186 58028
rect 86890 57974 86946 57976
rect 86970 57974 87026 57976
rect 87050 57974 87106 57976
rect 87130 57974 87186 57976
rect 86890 56940 86946 56942
rect 86970 56940 87026 56942
rect 87050 56940 87106 56942
rect 87130 56940 87186 56942
rect 86890 56888 86916 56940
rect 86916 56888 86946 56940
rect 86970 56888 86980 56940
rect 86980 56888 87026 56940
rect 87050 56888 87096 56940
rect 87096 56888 87106 56940
rect 87130 56888 87160 56940
rect 87160 56888 87186 56940
rect 86890 56886 86946 56888
rect 86970 56886 87026 56888
rect 87050 56886 87106 56888
rect 87130 56886 87186 56888
rect 86890 55852 86946 55854
rect 86970 55852 87026 55854
rect 87050 55852 87106 55854
rect 87130 55852 87186 55854
rect 86890 55800 86916 55852
rect 86916 55800 86946 55852
rect 86970 55800 86980 55852
rect 86980 55800 87026 55852
rect 87050 55800 87096 55852
rect 87096 55800 87106 55852
rect 87130 55800 87160 55852
rect 87160 55800 87186 55852
rect 86890 55798 86946 55800
rect 86970 55798 87026 55800
rect 87050 55798 87106 55800
rect 87130 55798 87186 55800
rect 86890 54764 86946 54766
rect 86970 54764 87026 54766
rect 87050 54764 87106 54766
rect 87130 54764 87186 54766
rect 86890 54712 86916 54764
rect 86916 54712 86946 54764
rect 86970 54712 86980 54764
rect 86980 54712 87026 54764
rect 87050 54712 87096 54764
rect 87096 54712 87106 54764
rect 87130 54712 87160 54764
rect 87160 54712 87186 54764
rect 86890 54710 86946 54712
rect 86970 54710 87026 54712
rect 87050 54710 87106 54712
rect 87130 54710 87186 54712
rect 86890 53676 86946 53678
rect 86970 53676 87026 53678
rect 87050 53676 87106 53678
rect 87130 53676 87186 53678
rect 86890 53624 86916 53676
rect 86916 53624 86946 53676
rect 86970 53624 86980 53676
rect 86980 53624 87026 53676
rect 87050 53624 87096 53676
rect 87096 53624 87106 53676
rect 87130 53624 87160 53676
rect 87160 53624 87186 53676
rect 86890 53622 86946 53624
rect 86970 53622 87026 53624
rect 87050 53622 87106 53624
rect 87130 53622 87186 53624
rect 86890 52588 86946 52590
rect 86970 52588 87026 52590
rect 87050 52588 87106 52590
rect 87130 52588 87186 52590
rect 86890 52536 86916 52588
rect 86916 52536 86946 52588
rect 86970 52536 86980 52588
rect 86980 52536 87026 52588
rect 87050 52536 87096 52588
rect 87096 52536 87106 52588
rect 87130 52536 87160 52588
rect 87160 52536 87186 52588
rect 86890 52534 86946 52536
rect 86970 52534 87026 52536
rect 87050 52534 87106 52536
rect 87130 52534 87186 52536
rect 86890 51500 86946 51502
rect 86970 51500 87026 51502
rect 87050 51500 87106 51502
rect 87130 51500 87186 51502
rect 86890 51448 86916 51500
rect 86916 51448 86946 51500
rect 86970 51448 86980 51500
rect 86980 51448 87026 51500
rect 87050 51448 87096 51500
rect 87096 51448 87106 51500
rect 87130 51448 87160 51500
rect 87160 51448 87186 51500
rect 86890 51446 86946 51448
rect 86970 51446 87026 51448
rect 87050 51446 87106 51448
rect 87130 51446 87186 51448
rect 86890 50412 86946 50414
rect 86970 50412 87026 50414
rect 87050 50412 87106 50414
rect 87130 50412 87186 50414
rect 86890 50360 86916 50412
rect 86916 50360 86946 50412
rect 86970 50360 86980 50412
rect 86980 50360 87026 50412
rect 87050 50360 87096 50412
rect 87096 50360 87106 50412
rect 87130 50360 87160 50412
rect 87160 50360 87186 50412
rect 86890 50358 86946 50360
rect 86970 50358 87026 50360
rect 87050 50358 87106 50360
rect 87130 50358 87186 50360
rect 86890 49324 86946 49326
rect 86970 49324 87026 49326
rect 87050 49324 87106 49326
rect 87130 49324 87186 49326
rect 86890 49272 86916 49324
rect 86916 49272 86946 49324
rect 86970 49272 86980 49324
rect 86980 49272 87026 49324
rect 87050 49272 87096 49324
rect 87096 49272 87106 49324
rect 87130 49272 87160 49324
rect 87160 49272 87186 49324
rect 86890 49270 86946 49272
rect 86970 49270 87026 49272
rect 87050 49270 87106 49272
rect 87130 49270 87186 49272
rect 86890 48236 86946 48238
rect 86970 48236 87026 48238
rect 87050 48236 87106 48238
rect 87130 48236 87186 48238
rect 86890 48184 86916 48236
rect 86916 48184 86946 48236
rect 86970 48184 86980 48236
rect 86980 48184 87026 48236
rect 87050 48184 87096 48236
rect 87096 48184 87106 48236
rect 87130 48184 87160 48236
rect 87160 48184 87186 48236
rect 86890 48182 86946 48184
rect 86970 48182 87026 48184
rect 87050 48182 87106 48184
rect 87130 48182 87186 48184
rect 86890 47148 86946 47150
rect 86970 47148 87026 47150
rect 87050 47148 87106 47150
rect 87130 47148 87186 47150
rect 86890 47096 86916 47148
rect 86916 47096 86946 47148
rect 86970 47096 86980 47148
rect 86980 47096 87026 47148
rect 87050 47096 87096 47148
rect 87096 47096 87106 47148
rect 87130 47096 87160 47148
rect 87160 47096 87186 47148
rect 86890 47094 86946 47096
rect 86970 47094 87026 47096
rect 87050 47094 87106 47096
rect 87130 47094 87186 47096
rect 86890 46060 86946 46062
rect 86970 46060 87026 46062
rect 87050 46060 87106 46062
rect 87130 46060 87186 46062
rect 86890 46008 86916 46060
rect 86916 46008 86946 46060
rect 86970 46008 86980 46060
rect 86980 46008 87026 46060
rect 87050 46008 87096 46060
rect 87096 46008 87106 46060
rect 87130 46008 87160 46060
rect 87160 46008 87186 46060
rect 86890 46006 86946 46008
rect 86970 46006 87026 46008
rect 87050 46006 87106 46008
rect 87130 46006 87186 46008
rect 86890 44972 86946 44974
rect 86970 44972 87026 44974
rect 87050 44972 87106 44974
rect 87130 44972 87186 44974
rect 86890 44920 86916 44972
rect 86916 44920 86946 44972
rect 86970 44920 86980 44972
rect 86980 44920 87026 44972
rect 87050 44920 87096 44972
rect 87096 44920 87106 44972
rect 87130 44920 87160 44972
rect 87160 44920 87186 44972
rect 86890 44918 86946 44920
rect 86970 44918 87026 44920
rect 87050 44918 87106 44920
rect 87130 44918 87186 44920
rect 86890 43884 86946 43886
rect 86970 43884 87026 43886
rect 87050 43884 87106 43886
rect 87130 43884 87186 43886
rect 86890 43832 86916 43884
rect 86916 43832 86946 43884
rect 86970 43832 86980 43884
rect 86980 43832 87026 43884
rect 87050 43832 87096 43884
rect 87096 43832 87106 43884
rect 87130 43832 87160 43884
rect 87160 43832 87186 43884
rect 86890 43830 86946 43832
rect 86970 43830 87026 43832
rect 87050 43830 87106 43832
rect 87130 43830 87186 43832
rect 86890 42796 86946 42798
rect 86970 42796 87026 42798
rect 87050 42796 87106 42798
rect 87130 42796 87186 42798
rect 86890 42744 86916 42796
rect 86916 42744 86946 42796
rect 86970 42744 86980 42796
rect 86980 42744 87026 42796
rect 87050 42744 87096 42796
rect 87096 42744 87106 42796
rect 87130 42744 87160 42796
rect 87160 42744 87186 42796
rect 86890 42742 86946 42744
rect 86970 42742 87026 42744
rect 87050 42742 87106 42744
rect 87130 42742 87186 42744
rect 86890 41708 86946 41710
rect 86970 41708 87026 41710
rect 87050 41708 87106 41710
rect 87130 41708 87186 41710
rect 86890 41656 86916 41708
rect 86916 41656 86946 41708
rect 86970 41656 86980 41708
rect 86980 41656 87026 41708
rect 87050 41656 87096 41708
rect 87096 41656 87106 41708
rect 87130 41656 87160 41708
rect 87160 41656 87186 41708
rect 86890 41654 86946 41656
rect 86970 41654 87026 41656
rect 87050 41654 87106 41656
rect 87130 41654 87186 41656
rect 86890 40620 86946 40622
rect 86970 40620 87026 40622
rect 87050 40620 87106 40622
rect 87130 40620 87186 40622
rect 86890 40568 86916 40620
rect 86916 40568 86946 40620
rect 86970 40568 86980 40620
rect 86980 40568 87026 40620
rect 87050 40568 87096 40620
rect 87096 40568 87106 40620
rect 87130 40568 87160 40620
rect 87160 40568 87186 40620
rect 86890 40566 86946 40568
rect 86970 40566 87026 40568
rect 87050 40566 87106 40568
rect 87130 40566 87186 40568
rect 86890 39532 86946 39534
rect 86970 39532 87026 39534
rect 87050 39532 87106 39534
rect 87130 39532 87186 39534
rect 86890 39480 86916 39532
rect 86916 39480 86946 39532
rect 86970 39480 86980 39532
rect 86980 39480 87026 39532
rect 87050 39480 87096 39532
rect 87096 39480 87106 39532
rect 87130 39480 87160 39532
rect 87160 39480 87186 39532
rect 86890 39478 86946 39480
rect 86970 39478 87026 39480
rect 87050 39478 87106 39480
rect 87130 39478 87186 39480
rect 86890 38444 86946 38446
rect 86970 38444 87026 38446
rect 87050 38444 87106 38446
rect 87130 38444 87186 38446
rect 86890 38392 86916 38444
rect 86916 38392 86946 38444
rect 86970 38392 86980 38444
rect 86980 38392 87026 38444
rect 87050 38392 87096 38444
rect 87096 38392 87106 38444
rect 87130 38392 87160 38444
rect 87160 38392 87186 38444
rect 86890 38390 86946 38392
rect 86970 38390 87026 38392
rect 87050 38390 87106 38392
rect 87130 38390 87186 38392
rect 86890 37356 86946 37358
rect 86970 37356 87026 37358
rect 87050 37356 87106 37358
rect 87130 37356 87186 37358
rect 86890 37304 86916 37356
rect 86916 37304 86946 37356
rect 86970 37304 86980 37356
rect 86980 37304 87026 37356
rect 87050 37304 87096 37356
rect 87096 37304 87106 37356
rect 87130 37304 87160 37356
rect 87160 37304 87186 37356
rect 86890 37302 86946 37304
rect 86970 37302 87026 37304
rect 87050 37302 87106 37304
rect 87130 37302 87186 37304
rect 86890 36268 86946 36270
rect 86970 36268 87026 36270
rect 87050 36268 87106 36270
rect 87130 36268 87186 36270
rect 86890 36216 86916 36268
rect 86916 36216 86946 36268
rect 86970 36216 86980 36268
rect 86980 36216 87026 36268
rect 87050 36216 87096 36268
rect 87096 36216 87106 36268
rect 87130 36216 87160 36268
rect 87160 36216 87186 36268
rect 86890 36214 86946 36216
rect 86970 36214 87026 36216
rect 87050 36214 87106 36216
rect 87130 36214 87186 36216
rect 86890 35180 86946 35182
rect 86970 35180 87026 35182
rect 87050 35180 87106 35182
rect 87130 35180 87186 35182
rect 86890 35128 86916 35180
rect 86916 35128 86946 35180
rect 86970 35128 86980 35180
rect 86980 35128 87026 35180
rect 87050 35128 87096 35180
rect 87096 35128 87106 35180
rect 87130 35128 87160 35180
rect 87160 35128 87186 35180
rect 86890 35126 86946 35128
rect 86970 35126 87026 35128
rect 87050 35126 87106 35128
rect 87130 35126 87186 35128
rect 86890 34092 86946 34094
rect 86970 34092 87026 34094
rect 87050 34092 87106 34094
rect 87130 34092 87186 34094
rect 86890 34040 86916 34092
rect 86916 34040 86946 34092
rect 86970 34040 86980 34092
rect 86980 34040 87026 34092
rect 87050 34040 87096 34092
rect 87096 34040 87106 34092
rect 87130 34040 87160 34092
rect 87160 34040 87186 34092
rect 86890 34038 86946 34040
rect 86970 34038 87026 34040
rect 87050 34038 87106 34040
rect 87130 34038 87186 34040
rect 86890 33004 86946 33006
rect 86970 33004 87026 33006
rect 87050 33004 87106 33006
rect 87130 33004 87186 33006
rect 86890 32952 86916 33004
rect 86916 32952 86946 33004
rect 86970 32952 86980 33004
rect 86980 32952 87026 33004
rect 87050 32952 87096 33004
rect 87096 32952 87106 33004
rect 87130 32952 87160 33004
rect 87160 32952 87186 33004
rect 86890 32950 86946 32952
rect 86970 32950 87026 32952
rect 87050 32950 87106 32952
rect 87130 32950 87186 32952
rect 86890 31916 86946 31918
rect 86970 31916 87026 31918
rect 87050 31916 87106 31918
rect 87130 31916 87186 31918
rect 86890 31864 86916 31916
rect 86916 31864 86946 31916
rect 86970 31864 86980 31916
rect 86980 31864 87026 31916
rect 87050 31864 87096 31916
rect 87096 31864 87106 31916
rect 87130 31864 87160 31916
rect 87160 31864 87186 31916
rect 86890 31862 86946 31864
rect 86970 31862 87026 31864
rect 87050 31862 87106 31864
rect 87130 31862 87186 31864
rect 86890 30828 86946 30830
rect 86970 30828 87026 30830
rect 87050 30828 87106 30830
rect 87130 30828 87186 30830
rect 86890 30776 86916 30828
rect 86916 30776 86946 30828
rect 86970 30776 86980 30828
rect 86980 30776 87026 30828
rect 87050 30776 87096 30828
rect 87096 30776 87106 30828
rect 87130 30776 87160 30828
rect 87160 30776 87186 30828
rect 86890 30774 86946 30776
rect 86970 30774 87026 30776
rect 87050 30774 87106 30776
rect 87130 30774 87186 30776
rect 86890 29740 86946 29742
rect 86970 29740 87026 29742
rect 87050 29740 87106 29742
rect 87130 29740 87186 29742
rect 86890 29688 86916 29740
rect 86916 29688 86946 29740
rect 86970 29688 86980 29740
rect 86980 29688 87026 29740
rect 87050 29688 87096 29740
rect 87096 29688 87106 29740
rect 87130 29688 87160 29740
rect 87160 29688 87186 29740
rect 86890 29686 86946 29688
rect 86970 29686 87026 29688
rect 87050 29686 87106 29688
rect 87130 29686 87186 29688
rect 86890 28652 86946 28654
rect 86970 28652 87026 28654
rect 87050 28652 87106 28654
rect 87130 28652 87186 28654
rect 86890 28600 86916 28652
rect 86916 28600 86946 28652
rect 86970 28600 86980 28652
rect 86980 28600 87026 28652
rect 87050 28600 87096 28652
rect 87096 28600 87106 28652
rect 87130 28600 87160 28652
rect 87160 28600 87186 28652
rect 86890 28598 86946 28600
rect 86970 28598 87026 28600
rect 87050 28598 87106 28600
rect 87130 28598 87186 28600
rect 86890 27564 86946 27566
rect 86970 27564 87026 27566
rect 87050 27564 87106 27566
rect 87130 27564 87186 27566
rect 86890 27512 86916 27564
rect 86916 27512 86946 27564
rect 86970 27512 86980 27564
rect 86980 27512 87026 27564
rect 87050 27512 87096 27564
rect 87096 27512 87106 27564
rect 87130 27512 87160 27564
rect 87160 27512 87186 27564
rect 86890 27510 86946 27512
rect 86970 27510 87026 27512
rect 87050 27510 87106 27512
rect 87130 27510 87186 27512
rect 86890 26476 86946 26478
rect 86970 26476 87026 26478
rect 87050 26476 87106 26478
rect 87130 26476 87186 26478
rect 86890 26424 86916 26476
rect 86916 26424 86946 26476
rect 86970 26424 86980 26476
rect 86980 26424 87026 26476
rect 87050 26424 87096 26476
rect 87096 26424 87106 26476
rect 87130 26424 87160 26476
rect 87160 26424 87186 26476
rect 86890 26422 86946 26424
rect 86970 26422 87026 26424
rect 87050 26422 87106 26424
rect 87130 26422 87186 26424
rect 86890 25388 86946 25390
rect 86970 25388 87026 25390
rect 87050 25388 87106 25390
rect 87130 25388 87186 25390
rect 86890 25336 86916 25388
rect 86916 25336 86946 25388
rect 86970 25336 86980 25388
rect 86980 25336 87026 25388
rect 87050 25336 87096 25388
rect 87096 25336 87106 25388
rect 87130 25336 87160 25388
rect 87160 25336 87186 25388
rect 86890 25334 86946 25336
rect 86970 25334 87026 25336
rect 87050 25334 87106 25336
rect 87130 25334 87186 25336
rect 86890 24300 86946 24302
rect 86970 24300 87026 24302
rect 87050 24300 87106 24302
rect 87130 24300 87186 24302
rect 86890 24248 86916 24300
rect 86916 24248 86946 24300
rect 86970 24248 86980 24300
rect 86980 24248 87026 24300
rect 87050 24248 87096 24300
rect 87096 24248 87106 24300
rect 87130 24248 87160 24300
rect 87160 24248 87186 24300
rect 86890 24246 86946 24248
rect 86970 24246 87026 24248
rect 87050 24246 87106 24248
rect 87130 24246 87186 24248
rect 86890 23212 86946 23214
rect 86970 23212 87026 23214
rect 87050 23212 87106 23214
rect 87130 23212 87186 23214
rect 86890 23160 86916 23212
rect 86916 23160 86946 23212
rect 86970 23160 86980 23212
rect 86980 23160 87026 23212
rect 87050 23160 87096 23212
rect 87096 23160 87106 23212
rect 87130 23160 87160 23212
rect 87160 23160 87186 23212
rect 86890 23158 86946 23160
rect 86970 23158 87026 23160
rect 87050 23158 87106 23160
rect 87130 23158 87186 23160
rect 86890 22124 86946 22126
rect 86970 22124 87026 22126
rect 87050 22124 87106 22126
rect 87130 22124 87186 22126
rect 86890 22072 86916 22124
rect 86916 22072 86946 22124
rect 86970 22072 86980 22124
rect 86980 22072 87026 22124
rect 87050 22072 87096 22124
rect 87096 22072 87106 22124
rect 87130 22072 87160 22124
rect 87160 22072 87186 22124
rect 86890 22070 86946 22072
rect 86970 22070 87026 22072
rect 87050 22070 87106 22072
rect 87130 22070 87186 22072
rect 86890 21036 86946 21038
rect 86970 21036 87026 21038
rect 87050 21036 87106 21038
rect 87130 21036 87186 21038
rect 86890 20984 86916 21036
rect 86916 20984 86946 21036
rect 86970 20984 86980 21036
rect 86980 20984 87026 21036
rect 87050 20984 87096 21036
rect 87096 20984 87106 21036
rect 87130 20984 87160 21036
rect 87160 20984 87186 21036
rect 86890 20982 86946 20984
rect 86970 20982 87026 20984
rect 87050 20982 87106 20984
rect 87130 20982 87186 20984
rect 86890 19948 86946 19950
rect 86970 19948 87026 19950
rect 87050 19948 87106 19950
rect 87130 19948 87186 19950
rect 86890 19896 86916 19948
rect 86916 19896 86946 19948
rect 86970 19896 86980 19948
rect 86980 19896 87026 19948
rect 87050 19896 87096 19948
rect 87096 19896 87106 19948
rect 87130 19896 87160 19948
rect 87160 19896 87186 19948
rect 86890 19894 86946 19896
rect 86970 19894 87026 19896
rect 87050 19894 87106 19896
rect 87130 19894 87186 19896
rect 86890 18860 86946 18862
rect 86970 18860 87026 18862
rect 87050 18860 87106 18862
rect 87130 18860 87186 18862
rect 86890 18808 86916 18860
rect 86916 18808 86946 18860
rect 86970 18808 86980 18860
rect 86980 18808 87026 18860
rect 87050 18808 87096 18860
rect 87096 18808 87106 18860
rect 87130 18808 87160 18860
rect 87160 18808 87186 18860
rect 86890 18806 86946 18808
rect 86970 18806 87026 18808
rect 87050 18806 87106 18808
rect 87130 18806 87186 18808
rect 86890 17772 86946 17774
rect 86970 17772 87026 17774
rect 87050 17772 87106 17774
rect 87130 17772 87186 17774
rect 86890 17720 86916 17772
rect 86916 17720 86946 17772
rect 86970 17720 86980 17772
rect 86980 17720 87026 17772
rect 87050 17720 87096 17772
rect 87096 17720 87106 17772
rect 87130 17720 87160 17772
rect 87160 17720 87186 17772
rect 86890 17718 86946 17720
rect 86970 17718 87026 17720
rect 87050 17718 87106 17720
rect 87130 17718 87186 17720
rect 86890 16684 86946 16686
rect 86970 16684 87026 16686
rect 87050 16684 87106 16686
rect 87130 16684 87186 16686
rect 86890 16632 86916 16684
rect 86916 16632 86946 16684
rect 86970 16632 86980 16684
rect 86980 16632 87026 16684
rect 87050 16632 87096 16684
rect 87096 16632 87106 16684
rect 87130 16632 87160 16684
rect 87160 16632 87186 16684
rect 86890 16630 86946 16632
rect 86970 16630 87026 16632
rect 87050 16630 87106 16632
rect 87130 16630 87186 16632
rect 86890 15596 86946 15598
rect 86970 15596 87026 15598
rect 87050 15596 87106 15598
rect 87130 15596 87186 15598
rect 86890 15544 86916 15596
rect 86916 15544 86946 15596
rect 86970 15544 86980 15596
rect 86980 15544 87026 15596
rect 87050 15544 87096 15596
rect 87096 15544 87106 15596
rect 87130 15544 87160 15596
rect 87160 15544 87186 15596
rect 86890 15542 86946 15544
rect 86970 15542 87026 15544
rect 87050 15542 87106 15544
rect 87130 15542 87186 15544
rect 86890 14508 86946 14510
rect 86970 14508 87026 14510
rect 87050 14508 87106 14510
rect 87130 14508 87186 14510
rect 86890 14456 86916 14508
rect 86916 14456 86946 14508
rect 86970 14456 86980 14508
rect 86980 14456 87026 14508
rect 87050 14456 87096 14508
rect 87096 14456 87106 14508
rect 87130 14456 87160 14508
rect 87160 14456 87186 14508
rect 86890 14454 86946 14456
rect 86970 14454 87026 14456
rect 87050 14454 87106 14456
rect 87130 14454 87186 14456
rect 86890 13420 86946 13422
rect 86970 13420 87026 13422
rect 87050 13420 87106 13422
rect 87130 13420 87186 13422
rect 86890 13368 86916 13420
rect 86916 13368 86946 13420
rect 86970 13368 86980 13420
rect 86980 13368 87026 13420
rect 87050 13368 87096 13420
rect 87096 13368 87106 13420
rect 87130 13368 87160 13420
rect 87160 13368 87186 13420
rect 86890 13366 86946 13368
rect 86970 13366 87026 13368
rect 87050 13366 87106 13368
rect 87130 13366 87186 13368
rect 86890 12332 86946 12334
rect 86970 12332 87026 12334
rect 87050 12332 87106 12334
rect 87130 12332 87186 12334
rect 86890 12280 86916 12332
rect 86916 12280 86946 12332
rect 86970 12280 86980 12332
rect 86980 12280 87026 12332
rect 87050 12280 87096 12332
rect 87096 12280 87106 12332
rect 87130 12280 87160 12332
rect 87160 12280 87186 12332
rect 86890 12278 86946 12280
rect 86970 12278 87026 12280
rect 87050 12278 87106 12280
rect 87130 12278 87186 12280
rect 86890 11244 86946 11246
rect 86970 11244 87026 11246
rect 87050 11244 87106 11246
rect 87130 11244 87186 11246
rect 86890 11192 86916 11244
rect 86916 11192 86946 11244
rect 86970 11192 86980 11244
rect 86980 11192 87026 11244
rect 87050 11192 87096 11244
rect 87096 11192 87106 11244
rect 87130 11192 87160 11244
rect 87160 11192 87186 11244
rect 86890 11190 86946 11192
rect 86970 11190 87026 11192
rect 87050 11190 87106 11192
rect 87130 11190 87186 11192
rect 86890 10156 86946 10158
rect 86970 10156 87026 10158
rect 87050 10156 87106 10158
rect 87130 10156 87186 10158
rect 86890 10104 86916 10156
rect 86916 10104 86946 10156
rect 86970 10104 86980 10156
rect 86980 10104 87026 10156
rect 87050 10104 87096 10156
rect 87096 10104 87106 10156
rect 87130 10104 87160 10156
rect 87160 10104 87186 10156
rect 86890 10102 86946 10104
rect 86970 10102 87026 10104
rect 87050 10102 87106 10104
rect 87130 10102 87186 10104
rect 86890 9068 86946 9070
rect 86970 9068 87026 9070
rect 87050 9068 87106 9070
rect 87130 9068 87186 9070
rect 86890 9016 86916 9068
rect 86916 9016 86946 9068
rect 86970 9016 86980 9068
rect 86980 9016 87026 9068
rect 87050 9016 87096 9068
rect 87096 9016 87106 9068
rect 87130 9016 87160 9068
rect 87160 9016 87186 9068
rect 86890 9014 86946 9016
rect 86970 9014 87026 9016
rect 87050 9014 87106 9016
rect 87130 9014 87186 9016
rect 86890 7980 86946 7982
rect 86970 7980 87026 7982
rect 87050 7980 87106 7982
rect 87130 7980 87186 7982
rect 86890 7928 86916 7980
rect 86916 7928 86946 7980
rect 86970 7928 86980 7980
rect 86980 7928 87026 7980
rect 87050 7928 87096 7980
rect 87096 7928 87106 7980
rect 87130 7928 87160 7980
rect 87160 7928 87186 7980
rect 86890 7926 86946 7928
rect 86970 7926 87026 7928
rect 87050 7926 87106 7928
rect 87130 7926 87186 7928
rect 86890 6892 86946 6894
rect 86970 6892 87026 6894
rect 87050 6892 87106 6894
rect 87130 6892 87186 6894
rect 86890 6840 86916 6892
rect 86916 6840 86946 6892
rect 86970 6840 86980 6892
rect 86980 6840 87026 6892
rect 87050 6840 87096 6892
rect 87096 6840 87106 6892
rect 87130 6840 87160 6892
rect 87160 6840 87186 6892
rect 86890 6838 86946 6840
rect 86970 6838 87026 6840
rect 87050 6838 87106 6840
rect 87130 6838 87186 6840
rect 86890 5804 86946 5806
rect 86970 5804 87026 5806
rect 87050 5804 87106 5806
rect 87130 5804 87186 5806
rect 86890 5752 86916 5804
rect 86916 5752 86946 5804
rect 86970 5752 86980 5804
rect 86980 5752 87026 5804
rect 87050 5752 87096 5804
rect 87096 5752 87106 5804
rect 87130 5752 87160 5804
rect 87160 5752 87186 5804
rect 86890 5750 86946 5752
rect 86970 5750 87026 5752
rect 87050 5750 87106 5752
rect 87130 5750 87186 5752
rect 86890 4716 86946 4718
rect 86970 4716 87026 4718
rect 87050 4716 87106 4718
rect 87130 4716 87186 4718
rect 86890 4664 86916 4716
rect 86916 4664 86946 4716
rect 86970 4664 86980 4716
rect 86980 4664 87026 4716
rect 87050 4664 87096 4716
rect 87096 4664 87106 4716
rect 87130 4664 87160 4716
rect 87160 4664 87186 4716
rect 86890 4662 86946 4664
rect 86970 4662 87026 4664
rect 87050 4662 87106 4664
rect 87130 4662 87186 4664
rect 86890 3628 86946 3630
rect 86970 3628 87026 3630
rect 87050 3628 87106 3630
rect 87130 3628 87186 3630
rect 86890 3576 86916 3628
rect 86916 3576 86946 3628
rect 86970 3576 86980 3628
rect 86980 3576 87026 3628
rect 87050 3576 87096 3628
rect 87096 3576 87106 3628
rect 87130 3576 87160 3628
rect 87160 3576 87186 3628
rect 86890 3574 86946 3576
rect 86970 3574 87026 3576
rect 87050 3574 87106 3576
rect 87130 3574 87186 3576
rect 86890 2540 86946 2542
rect 86970 2540 87026 2542
rect 87050 2540 87106 2542
rect 87130 2540 87186 2542
rect 86890 2488 86916 2540
rect 86916 2488 86946 2540
rect 86970 2488 86980 2540
rect 86980 2488 87026 2540
rect 87050 2488 87096 2540
rect 87096 2488 87106 2540
rect 87130 2488 87160 2540
rect 87160 2488 87186 2540
rect 86890 2486 86946 2488
rect 86970 2486 87026 2488
rect 87050 2486 87106 2488
rect 87130 2486 87186 2488
<< metal3 >>
rect 84323 189204 84389 189207
rect 88454 189204 88934 189234
rect 84323 189202 88934 189204
rect 84323 189146 84328 189202
rect 84384 189146 88934 189202
rect 84323 189144 88934 189146
rect 84323 189141 84389 189144
rect 88454 189114 88934 189144
rect 5244 187918 5250 187982
rect 5314 187980 5320 187982
rect 81747 187980 81813 187983
rect 5314 187978 81813 187980
rect 5314 187922 81752 187978
rect 81808 187922 81813 187978
rect 5314 187920 81813 187922
rect 5314 187918 5320 187920
rect 81747 187917 81813 187920
rect 85151 187980 85217 187983
rect 88454 187980 88934 188010
rect 85151 187978 88934 187980
rect 85151 187922 85156 187978
rect 85212 187922 88934 187978
rect 85151 187920 88934 187922
rect 85151 187917 85217 187920
rect 88454 187890 88934 187920
rect 2878 187506 3198 187507
rect 2878 187442 2886 187506
rect 2950 187442 2966 187506
rect 3030 187442 3046 187506
rect 3110 187442 3126 187506
rect 3190 187442 3198 187506
rect 2878 187441 3198 187442
rect 86878 187506 87198 187507
rect 86878 187442 86886 187506
rect 86950 187442 86966 187506
rect 87030 187442 87046 187506
rect 87110 187442 87126 187506
rect 87190 187442 87198 187506
rect 86878 187441 87198 187442
rect 4140 187374 4146 187438
rect 4210 187436 4216 187438
rect 84231 187436 84297 187439
rect 4210 187434 84297 187436
rect 4210 187378 84236 187434
rect 84292 187378 84297 187434
rect 4210 187376 84297 187378
rect 4210 187374 4216 187376
rect 84231 187373 84297 187376
rect 1247 187300 1313 187303
rect 84180 187300 84186 187302
rect 1247 187298 84186 187300
rect 1247 187242 1252 187298
rect 1308 187242 84186 187298
rect 1247 187240 84186 187242
rect 1247 187237 1313 187240
rect 84180 187238 84186 187240
rect 84250 187238 84256 187302
rect 3588 187102 3594 187166
rect 3658 187164 3664 187166
rect 84548 187164 84554 187166
rect 3658 187104 84554 187164
rect 3658 187102 3664 187104
rect 84548 187102 84554 187104
rect 84618 187102 84624 187166
rect 3772 186966 3778 187030
rect 3842 187028 3848 187030
rect 84599 187028 84665 187031
rect 3842 187026 84665 187028
rect 3842 186970 84604 187026
rect 84660 186970 84665 187026
rect 3842 186968 84665 186970
rect 3842 186966 3848 186968
rect 84599 186965 84665 186968
rect 878 186962 1198 186963
rect 878 186898 886 186962
rect 950 186898 966 186962
rect 1030 186898 1046 186962
rect 1110 186898 1126 186962
rect 1190 186898 1198 186962
rect 878 186897 1198 186898
rect 84878 186962 85198 186963
rect 84878 186898 84886 186962
rect 84950 186898 84966 186962
rect 85030 186898 85046 186962
rect 85110 186898 85126 186962
rect 85190 186898 85198 186962
rect 84878 186897 85198 186898
rect 1431 186756 1497 186759
rect 85151 186756 85217 186759
rect 88454 186756 88934 186786
rect 1431 186754 82408 186756
rect 1431 186698 1436 186754
rect 1492 186698 82408 186754
rect 1431 186696 82408 186698
rect 1431 186693 1497 186696
rect 82348 186620 82408 186696
rect 85151 186754 88934 186756
rect 85151 186698 85156 186754
rect 85212 186698 88934 186754
rect 85151 186696 88934 186698
rect 85151 186693 85217 186696
rect 88454 186666 88934 186696
rect 84732 186620 84738 186622
rect 82348 186560 84738 186620
rect 84732 186558 84738 186560
rect 84802 186558 84808 186622
rect 2878 186418 3198 186419
rect 2878 186354 2886 186418
rect 2950 186354 2966 186418
rect 3030 186354 3046 186418
rect 3110 186354 3126 186418
rect 3190 186354 3198 186418
rect 2878 186353 3198 186354
rect 86878 186418 87198 186419
rect 86878 186354 86886 186418
rect 86950 186354 86966 186418
rect 87030 186354 87046 186418
rect 87110 186354 87126 186418
rect 87190 186354 87198 186418
rect 86878 186353 87198 186354
rect 878 185874 1198 185875
rect 878 185810 886 185874
rect 950 185810 966 185874
rect 1030 185810 1046 185874
rect 1110 185810 1126 185874
rect 1190 185810 1198 185874
rect 878 185809 1198 185810
rect 84878 185874 85198 185875
rect 84878 185810 84886 185874
rect 84950 185810 84966 185874
rect 85030 185810 85046 185874
rect 85110 185810 85126 185874
rect 85190 185810 85198 185874
rect 84878 185809 85198 185810
rect 84783 185532 84849 185535
rect 88454 185532 88934 185562
rect 84783 185530 88934 185532
rect 84783 185474 84788 185530
rect 84844 185474 88934 185530
rect 84783 185472 88934 185474
rect 84783 185469 84849 185472
rect 88454 185442 88934 185472
rect 2878 185330 3198 185331
rect 2878 185266 2886 185330
rect 2950 185266 2966 185330
rect 3030 185266 3046 185330
rect 3110 185266 3126 185330
rect 3190 185266 3198 185330
rect 2878 185265 3198 185266
rect 86878 185330 87198 185331
rect 86878 185266 86886 185330
rect 86950 185266 86966 185330
rect 87030 185266 87046 185330
rect 87110 185266 87126 185330
rect 87190 185266 87198 185330
rect 86878 185265 87198 185266
rect 878 184786 1198 184787
rect 878 184722 886 184786
rect 950 184722 966 184786
rect 1030 184722 1046 184786
rect 1110 184722 1126 184786
rect 1190 184722 1198 184786
rect 878 184721 1198 184722
rect 84878 184786 85198 184787
rect 84878 184722 84886 184786
rect 84950 184722 84966 184786
rect 85030 184722 85046 184786
rect 85110 184722 85126 184786
rect 85190 184722 85198 184786
rect 84878 184721 85198 184722
rect 84732 184382 84738 184446
rect 84802 184444 84808 184446
rect 84802 184384 87376 184444
rect 84802 184382 84808 184384
rect 87316 184308 87376 184384
rect 88454 184308 88934 184338
rect 87316 184248 88934 184308
rect 2878 184242 3198 184243
rect 2878 184178 2886 184242
rect 2950 184178 2966 184242
rect 3030 184178 3046 184242
rect 3110 184178 3126 184242
rect 3190 184178 3198 184242
rect 2878 184177 3198 184178
rect 86878 184242 87198 184243
rect 86878 184178 86886 184242
rect 86950 184178 86966 184242
rect 87030 184178 87046 184242
rect 87110 184178 87126 184242
rect 87190 184178 87198 184242
rect 88454 184218 88934 184248
rect 86878 184177 87198 184178
rect 878 183698 1198 183699
rect 878 183634 886 183698
rect 950 183634 966 183698
rect 1030 183634 1046 183698
rect 1110 183634 1126 183698
rect 1190 183634 1198 183698
rect 878 183633 1198 183634
rect 84878 183698 85198 183699
rect 84878 183634 84886 183698
rect 84950 183634 84966 183698
rect 85030 183634 85046 183698
rect 85110 183634 85126 183698
rect 85190 183634 85198 183698
rect 84878 183633 85198 183634
rect 84548 183294 84554 183358
rect 84618 183356 84624 183358
rect 84618 183296 87376 183356
rect 84618 183294 84624 183296
rect 2878 183154 3198 183155
rect 2878 183090 2886 183154
rect 2950 183090 2966 183154
rect 3030 183090 3046 183154
rect 3110 183090 3126 183154
rect 3190 183090 3198 183154
rect 2878 183089 3198 183090
rect 86878 183154 87198 183155
rect 86878 183090 86886 183154
rect 86950 183090 86966 183154
rect 87030 183090 87046 183154
rect 87110 183090 87126 183154
rect 87190 183090 87198 183154
rect 86878 183089 87198 183090
rect 87316 183084 87376 183296
rect 88454 183084 88934 183114
rect 87316 183024 88934 183084
rect 88454 182994 88934 183024
rect 3915 182812 3981 182815
rect 3915 182810 5128 182812
rect 3915 182754 3920 182810
rect 3976 182754 5128 182810
rect 3915 182752 5128 182754
rect 3915 182749 3981 182752
rect 878 182610 1198 182611
rect 878 182546 886 182610
rect 950 182546 966 182610
rect 1030 182546 1046 182610
rect 1110 182546 1126 182610
rect 1190 182546 1198 182610
rect 878 182545 1198 182546
rect 84878 182610 85198 182611
rect 84878 182546 84886 182610
rect 84950 182546 84966 182610
rect 85030 182546 85046 182610
rect 85110 182546 85126 182610
rect 85190 182546 85198 182610
rect 84878 182545 85198 182546
rect 84231 182404 84297 182407
rect 84231 182402 84432 182404
rect 84231 182346 84236 182402
rect 84292 182346 84432 182402
rect 84231 182344 84432 182346
rect 84231 182341 84297 182344
rect 84372 182132 84432 182344
rect 84548 182206 84554 182270
rect 84618 182268 84624 182270
rect 84618 182208 87560 182268
rect 84618 182206 84624 182208
rect 84372 182072 84616 182132
rect 2878 182066 3198 182067
rect 2878 182002 2886 182066
rect 2950 182002 2966 182066
rect 3030 182002 3046 182066
rect 3110 182002 3126 182066
rect 3190 182002 3198 182066
rect 2878 182001 3198 182002
rect 84556 181999 84616 182072
rect 86878 182066 87198 182067
rect 86878 182002 86886 182066
rect 86950 182002 86966 182066
rect 87030 182002 87046 182066
rect 87110 182002 87126 182066
rect 87190 182002 87198 182066
rect 86878 182001 87198 182002
rect 84556 181994 84665 181999
rect 84556 181938 84604 181994
rect 84660 181938 84665 181994
rect 84556 181936 84665 181938
rect 87500 181996 87560 182208
rect 88454 181996 88934 182026
rect 87500 181936 88934 181996
rect 84599 181933 84665 181936
rect 88454 181906 88934 181936
rect 3547 181724 3613 181727
rect 3547 181722 5128 181724
rect 3547 181666 3552 181722
rect 3608 181666 5128 181722
rect 3547 181664 5128 181666
rect 3547 181661 3613 181664
rect 5068 181661 5128 181664
rect 878 181522 1198 181523
rect 878 181458 886 181522
rect 950 181458 966 181522
rect 1030 181458 1046 181522
rect 1110 181458 1126 181522
rect 1190 181458 1198 181522
rect 878 181457 1198 181458
rect 84878 181522 85198 181523
rect 84878 181458 84886 181522
rect 84950 181458 84966 181522
rect 85030 181458 85046 181522
rect 85110 181458 85126 181522
rect 85190 181458 85198 181522
rect 84878 181457 85198 181458
rect 2878 180978 3198 180979
rect 2878 180914 2886 180978
rect 2950 180914 2966 180978
rect 3030 180914 3046 180978
rect 3110 180914 3126 180978
rect 3190 180914 3198 180978
rect 2878 180913 3198 180914
rect 86878 180978 87198 180979
rect 86878 180914 86886 180978
rect 86950 180914 86966 180978
rect 87030 180914 87046 180978
rect 87110 180914 87126 180978
rect 87190 180914 87198 180978
rect 86878 180913 87198 180914
rect 83955 180772 84021 180775
rect 88454 180772 88934 180802
rect 83955 180770 88934 180772
rect 83955 180714 83960 180770
rect 84016 180714 88934 180770
rect 83955 180712 88934 180714
rect 83955 180709 84021 180712
rect 88454 180682 88934 180712
rect 878 180434 1198 180435
rect 878 180370 886 180434
rect 950 180370 966 180434
rect 1030 180370 1046 180434
rect 1110 180370 1126 180434
rect 1190 180370 1198 180434
rect 878 180369 1198 180370
rect 84878 180434 85198 180435
rect 84878 180370 84886 180434
rect 84950 180370 84966 180434
rect 85030 180370 85046 180434
rect 85110 180370 85126 180434
rect 85190 180370 85198 180434
rect 84878 180369 85198 180370
rect 3547 179956 3613 179959
rect 3823 179956 3889 179959
rect 5068 179956 5128 179961
rect 3547 179954 5128 179956
rect 3547 179898 3552 179954
rect 3608 179898 3828 179954
rect 3884 179898 5128 179954
rect 3547 179896 5128 179898
rect 3547 179893 3613 179896
rect 3823 179893 3889 179896
rect 2878 179890 3198 179891
rect 2878 179826 2886 179890
rect 2950 179826 2966 179890
rect 3030 179826 3046 179890
rect 3110 179826 3126 179890
rect 3190 179826 3198 179890
rect 2878 179825 3198 179826
rect 86878 179890 87198 179891
rect 86878 179826 86886 179890
rect 86950 179826 86966 179890
rect 87030 179826 87046 179890
rect 87110 179826 87126 179890
rect 87190 179826 87198 179890
rect 86878 179825 87198 179826
rect 84139 179548 84205 179551
rect 88454 179548 88934 179578
rect 84139 179546 88934 179548
rect 84139 179490 84144 179546
rect 84200 179490 88934 179546
rect 84139 179488 88934 179490
rect 84139 179485 84205 179488
rect 88454 179458 88934 179488
rect 878 179346 1198 179347
rect 878 179282 886 179346
rect 950 179282 966 179346
rect 1030 179282 1046 179346
rect 1110 179282 1126 179346
rect 1190 179282 1198 179346
rect 878 179281 1198 179282
rect 84878 179346 85198 179347
rect 84878 179282 84886 179346
rect 84950 179282 84966 179346
rect 85030 179282 85046 179346
rect 85110 179282 85126 179346
rect 85190 179282 85198 179346
rect 84878 179281 85198 179282
rect 4007 178868 4073 178871
rect 4007 178866 5128 178868
rect 4007 178810 4012 178866
rect 4068 178810 5128 178866
rect 4007 178808 5128 178810
rect 4007 178805 4073 178808
rect 2878 178802 3198 178803
rect 2878 178738 2886 178802
rect 2950 178738 2966 178802
rect 3030 178738 3046 178802
rect 3110 178738 3126 178802
rect 3190 178738 3198 178802
rect 2878 178737 3198 178738
rect 86878 178802 87198 178803
rect 86878 178738 86886 178802
rect 86950 178738 86966 178802
rect 87030 178738 87046 178802
rect 87110 178738 87126 178802
rect 87190 178738 87198 178802
rect 86878 178737 87198 178738
rect 84599 178596 84665 178599
rect 84599 178594 85352 178596
rect 84599 178538 84604 178594
rect 84660 178538 85352 178594
rect 84599 178536 85352 178538
rect 84599 178533 84665 178536
rect 85292 178324 85352 178536
rect 88454 178324 88934 178354
rect 85292 178264 88934 178324
rect 878 178258 1198 178259
rect 878 178194 886 178258
rect 950 178194 966 178258
rect 1030 178194 1046 178258
rect 1110 178194 1126 178258
rect 1190 178194 1198 178258
rect 878 178193 1198 178194
rect 84878 178258 85198 178259
rect 84878 178194 84886 178258
rect 84950 178194 84966 178258
rect 85030 178194 85046 178258
rect 85110 178194 85126 178258
rect 85190 178194 85198 178258
rect 88454 178234 88934 178264
rect 84878 178193 85198 178194
rect 2878 177714 3198 177715
rect 2878 177650 2886 177714
rect 2950 177650 2966 177714
rect 3030 177650 3046 177714
rect 3110 177650 3126 177714
rect 3190 177650 3198 177714
rect 2878 177649 3198 177650
rect 86878 177714 87198 177715
rect 86878 177650 86886 177714
rect 86950 177650 86966 177714
rect 87030 177650 87046 177714
rect 87110 177650 87126 177714
rect 87190 177650 87198 177714
rect 86878 177649 87198 177650
rect 878 177170 1198 177171
rect 878 177106 886 177170
rect 950 177106 966 177170
rect 1030 177106 1046 177170
rect 1110 177106 1126 177170
rect 1190 177106 1198 177170
rect 84878 177170 85198 177171
rect 878 177105 1198 177106
rect 3639 176828 3705 176831
rect 5068 176828 5128 177133
rect 84878 177106 84886 177170
rect 84950 177106 84966 177170
rect 85030 177106 85046 177170
rect 85110 177106 85126 177170
rect 85190 177106 85198 177170
rect 84878 177105 85198 177106
rect 88454 177100 88934 177130
rect 85292 177040 88934 177100
rect 3639 176826 5128 176828
rect 3639 176770 3644 176826
rect 3700 176770 5128 176826
rect 3639 176768 5128 176770
rect 83771 176828 83837 176831
rect 85292 176828 85352 177040
rect 88454 177010 88934 177040
rect 83771 176826 85352 176828
rect 83771 176770 83776 176826
rect 83832 176770 85352 176826
rect 83771 176768 85352 176770
rect 3639 176765 3705 176768
rect 83771 176765 83837 176768
rect 2878 176626 3198 176627
rect 2878 176562 2886 176626
rect 2950 176562 2966 176626
rect 3030 176562 3046 176626
rect 3110 176562 3126 176626
rect 3190 176562 3198 176626
rect 2878 176561 3198 176562
rect 86878 176626 87198 176627
rect 86878 176562 86886 176626
rect 86950 176562 86966 176626
rect 87030 176562 87046 176626
rect 87110 176562 87126 176626
rect 87190 176562 87198 176626
rect 86878 176561 87198 176562
rect 878 176082 1198 176083
rect 878 176018 886 176082
rect 950 176018 966 176082
rect 1030 176018 1046 176082
rect 1110 176018 1126 176082
rect 1190 176018 1198 176082
rect 878 176017 1198 176018
rect 84878 176082 85198 176083
rect 84878 176018 84886 176082
rect 84950 176018 84966 176082
rect 85030 176018 85046 176082
rect 85110 176018 85126 176082
rect 85190 176018 85198 176082
rect 84878 176017 85198 176018
rect 3271 175740 3337 175743
rect 5068 175740 5128 176005
rect 83863 175876 83929 175879
rect 88454 175876 88934 175906
rect 83863 175874 88934 175876
rect 83863 175818 83868 175874
rect 83924 175818 88934 175874
rect 83863 175816 88934 175818
rect 83863 175813 83929 175816
rect 88454 175786 88934 175816
rect 3271 175738 5128 175740
rect 3271 175682 3276 175738
rect 3332 175682 5128 175738
rect 3271 175680 5128 175682
rect 3271 175677 3337 175680
rect 2878 175538 3198 175539
rect 2878 175474 2886 175538
rect 2950 175474 2966 175538
rect 3030 175474 3046 175538
rect 3110 175474 3126 175538
rect 3190 175474 3198 175538
rect 2878 175473 3198 175474
rect 86878 175538 87198 175539
rect 86878 175474 86886 175538
rect 86950 175474 86966 175538
rect 87030 175474 87046 175538
rect 87110 175474 87126 175538
rect 87190 175474 87198 175538
rect 86878 175473 87198 175474
rect 878 174994 1198 174995
rect 878 174930 886 174994
rect 950 174930 966 174994
rect 1030 174930 1046 174994
rect 1110 174930 1126 174994
rect 1190 174930 1198 174994
rect 878 174929 1198 174930
rect 84878 174994 85198 174995
rect 84878 174930 84886 174994
rect 84950 174930 84966 174994
rect 85030 174930 85046 174994
rect 85110 174930 85126 174994
rect 85190 174930 85198 174994
rect 84878 174929 85198 174930
rect 84139 174788 84205 174791
rect 88454 174788 88934 174818
rect 84139 174786 88934 174788
rect 84139 174730 84144 174786
rect 84200 174730 88934 174786
rect 84139 174728 88934 174730
rect 84139 174725 84205 174728
rect 88454 174698 88934 174728
rect 2878 174450 3198 174451
rect 2878 174386 2886 174450
rect 2950 174386 2966 174450
rect 3030 174386 3046 174450
rect 3110 174386 3126 174450
rect 3190 174386 3198 174450
rect 2878 174385 3198 174386
rect 86878 174450 87198 174451
rect 86878 174386 86886 174450
rect 86950 174386 86966 174450
rect 87030 174386 87046 174450
rect 87110 174386 87126 174450
rect 87190 174386 87198 174450
rect 86878 174385 87198 174386
rect 3639 174108 3705 174111
rect 5068 174108 5128 174305
rect 3639 174106 5128 174108
rect 3639 174050 3644 174106
rect 3700 174050 5128 174106
rect 3639 174048 5128 174050
rect 3639 174045 3705 174048
rect 878 173906 1198 173907
rect 878 173842 886 173906
rect 950 173842 966 173906
rect 1030 173842 1046 173906
rect 1110 173842 1126 173906
rect 1190 173842 1198 173906
rect 878 173841 1198 173842
rect 84878 173906 85198 173907
rect 84878 173842 84886 173906
rect 84950 173842 84966 173906
rect 85030 173842 85046 173906
rect 85110 173842 85126 173906
rect 85190 173842 85198 173906
rect 84878 173841 85198 173842
rect 84047 173564 84113 173567
rect 88454 173564 88934 173594
rect 84047 173562 88934 173564
rect 84047 173506 84052 173562
rect 84108 173506 88934 173562
rect 84047 173504 88934 173506
rect 84047 173501 84113 173504
rect 88454 173474 88934 173504
rect 2878 173362 3198 173363
rect 2878 173298 2886 173362
rect 2950 173298 2966 173362
rect 3030 173298 3046 173362
rect 3110 173298 3126 173362
rect 3190 173298 3198 173362
rect 2878 173297 3198 173298
rect 86878 173362 87198 173363
rect 86878 173298 86886 173362
rect 86950 173298 86966 173362
rect 87030 173298 87046 173362
rect 87110 173298 87126 173362
rect 87190 173298 87198 173362
rect 86878 173297 87198 173298
rect 878 172818 1198 172819
rect 878 172754 886 172818
rect 950 172754 966 172818
rect 1030 172754 1046 172818
rect 1110 172754 1126 172818
rect 1190 172754 1198 172818
rect 878 172753 1198 172754
rect 84878 172818 85198 172819
rect 84878 172754 84886 172818
rect 84950 172754 84966 172818
rect 85030 172754 85046 172818
rect 85110 172754 85126 172818
rect 85190 172754 85198 172818
rect 84878 172753 85198 172754
rect 88454 172340 88934 172370
rect 87316 172280 88934 172340
rect 2878 172274 3198 172275
rect 2878 172210 2886 172274
rect 2950 172210 2966 172274
rect 3030 172210 3046 172274
rect 3110 172210 3126 172274
rect 3190 172210 3198 172274
rect 2878 172209 3198 172210
rect 86878 172274 87198 172275
rect 86878 172210 86886 172274
rect 86950 172210 86966 172274
rect 87030 172210 87046 172274
rect 87110 172210 87126 172274
rect 87190 172210 87198 172274
rect 86878 172209 87198 172210
rect 84732 172006 84738 172070
rect 84802 172068 84808 172070
rect 87316 172068 87376 172280
rect 88454 172250 88934 172280
rect 84802 172008 87376 172068
rect 84802 172006 84808 172008
rect 878 171730 1198 171731
rect 878 171666 886 171730
rect 950 171666 966 171730
rect 1030 171666 1046 171730
rect 1110 171666 1126 171730
rect 1190 171666 1198 171730
rect 878 171665 1198 171666
rect 84878 171730 85198 171731
rect 84878 171666 84886 171730
rect 84950 171666 84966 171730
rect 85030 171666 85046 171730
rect 85110 171666 85126 171730
rect 85190 171666 85198 171730
rect 84878 171665 85198 171666
rect 2878 171186 3198 171187
rect 2878 171122 2886 171186
rect 2950 171122 2966 171186
rect 3030 171122 3046 171186
rect 3110 171122 3126 171186
rect 3190 171122 3198 171186
rect 2878 171121 3198 171122
rect 86878 171186 87198 171187
rect 86878 171122 86886 171186
rect 86950 171122 86966 171186
rect 87030 171122 87046 171186
rect 87110 171122 87126 171186
rect 87190 171122 87198 171186
rect 86878 171121 87198 171122
rect 1891 171116 1957 171119
rect 2259 171116 2325 171119
rect 88454 171116 88934 171146
rect 1891 171114 2325 171116
rect 1891 171058 1896 171114
rect 1952 171058 2264 171114
rect 2320 171058 2325 171114
rect 1891 171056 2325 171058
rect 1891 171053 1957 171056
rect 2259 171053 2325 171056
rect 87316 171056 88934 171116
rect 84783 170980 84849 170983
rect 87316 170980 87376 171056
rect 88454 171026 88934 171056
rect 84783 170978 87376 170980
rect 84783 170922 84788 170978
rect 84844 170922 87376 170978
rect 84783 170920 87376 170922
rect 84783 170917 84849 170920
rect 878 170642 1198 170643
rect 878 170578 886 170642
rect 950 170578 966 170642
rect 1030 170578 1046 170642
rect 1110 170578 1126 170642
rect 1190 170578 1198 170642
rect 878 170577 1198 170578
rect 84878 170642 85198 170643
rect 84878 170578 84886 170642
rect 84950 170578 84966 170642
rect 85030 170578 85046 170642
rect 85110 170578 85126 170642
rect 85190 170578 85198 170642
rect 84878 170577 85198 170578
rect 2878 170098 3198 170099
rect 2878 170034 2886 170098
rect 2950 170034 2966 170098
rect 3030 170034 3046 170098
rect 3110 170034 3126 170098
rect 3190 170034 3198 170098
rect 2878 170033 3198 170034
rect 86878 170098 87198 170099
rect 86878 170034 86886 170098
rect 86950 170034 86966 170098
rect 87030 170034 87046 170098
rect 87110 170034 87126 170098
rect 87190 170034 87198 170098
rect 86878 170033 87198 170034
rect 83812 169830 83818 169894
rect 83882 169892 83888 169894
rect 88454 169892 88934 169922
rect 83882 169832 88934 169892
rect 83882 169830 83888 169832
rect 88454 169802 88934 169832
rect 878 169554 1198 169555
rect 878 169490 886 169554
rect 950 169490 966 169554
rect 1030 169490 1046 169554
rect 1110 169490 1126 169554
rect 1190 169490 1198 169554
rect 878 169489 1198 169490
rect 84878 169554 85198 169555
rect 84878 169490 84886 169554
rect 84950 169490 84966 169554
rect 85030 169490 85046 169554
rect 85110 169490 85126 169554
rect 85190 169490 85198 169554
rect 84878 169489 85198 169490
rect 2878 169010 3198 169011
rect 2878 168946 2886 169010
rect 2950 168946 2966 169010
rect 3030 168946 3046 169010
rect 3110 168946 3126 169010
rect 3190 168946 3198 169010
rect 2878 168945 3198 168946
rect 86878 169010 87198 169011
rect 86878 168946 86886 169010
rect 86950 168946 86966 169010
rect 87030 168946 87046 169010
rect 87110 168946 87126 169010
rect 87190 168946 87198 169010
rect 86878 168945 87198 168946
rect 83628 168606 83634 168670
rect 83698 168668 83704 168670
rect 88454 168668 88934 168698
rect 83698 168608 88934 168668
rect 83698 168606 83704 168608
rect 88454 168578 88934 168608
rect 878 168466 1198 168467
rect 878 168402 886 168466
rect 950 168402 966 168466
rect 1030 168402 1046 168466
rect 1110 168402 1126 168466
rect 1190 168402 1198 168466
rect 878 168401 1198 168402
rect 84878 168466 85198 168467
rect 84878 168402 84886 168466
rect 84950 168402 84966 168466
rect 85030 168402 85046 168466
rect 85110 168402 85126 168466
rect 85190 168402 85198 168466
rect 84878 168401 85198 168402
rect 2878 167922 3198 167923
rect 2878 167858 2886 167922
rect 2950 167858 2966 167922
rect 3030 167858 3046 167922
rect 3110 167858 3126 167922
rect 3190 167858 3198 167922
rect 2878 167857 3198 167858
rect 86878 167922 87198 167923
rect 86878 167858 86886 167922
rect 86950 167858 86966 167922
rect 87030 167858 87046 167922
rect 87110 167858 87126 167922
rect 87190 167858 87198 167922
rect 86878 167857 87198 167858
rect 84180 167518 84186 167582
rect 84250 167580 84256 167582
rect 88454 167580 88934 167610
rect 84250 167520 88934 167580
rect 84250 167518 84256 167520
rect 88454 167490 88934 167520
rect 878 167378 1198 167379
rect 878 167314 886 167378
rect 950 167314 966 167378
rect 1030 167314 1046 167378
rect 1110 167314 1126 167378
rect 1190 167314 1198 167378
rect 878 167313 1198 167314
rect 84878 167378 85198 167379
rect 84878 167314 84886 167378
rect 84950 167314 84966 167378
rect 85030 167314 85046 167378
rect 85110 167314 85126 167378
rect 85190 167314 85198 167378
rect 84878 167313 85198 167314
rect 2878 166834 3198 166835
rect 2878 166770 2886 166834
rect 2950 166770 2966 166834
rect 3030 166770 3046 166834
rect 3110 166770 3126 166834
rect 3190 166770 3198 166834
rect 2878 166769 3198 166770
rect 86878 166834 87198 166835
rect 86878 166770 86886 166834
rect 86950 166770 86966 166834
rect 87030 166770 87046 166834
rect 87110 166770 87126 166834
rect 87190 166770 87198 166834
rect 86878 166769 87198 166770
rect 88454 166356 88934 166386
rect 85292 166296 88934 166356
rect 878 166290 1198 166291
rect 878 166226 886 166290
rect 950 166226 966 166290
rect 1030 166226 1046 166290
rect 1110 166226 1126 166290
rect 1190 166226 1198 166290
rect 878 166225 1198 166226
rect 84878 166290 85198 166291
rect 84878 166226 84886 166290
rect 84950 166226 84966 166290
rect 85030 166226 85046 166290
rect 85110 166226 85126 166290
rect 85190 166226 85198 166290
rect 84878 166225 85198 166226
rect 83444 166022 83450 166086
rect 83514 166084 83520 166086
rect 85292 166084 85352 166296
rect 88454 166266 88934 166296
rect 83514 166024 85352 166084
rect 83514 166022 83520 166024
rect 2878 165746 3198 165747
rect 2878 165682 2886 165746
rect 2950 165682 2966 165746
rect 3030 165682 3046 165746
rect 3110 165682 3126 165746
rect 3190 165682 3198 165746
rect 2878 165681 3198 165682
rect 86878 165746 87198 165747
rect 86878 165682 86886 165746
rect 86950 165682 86966 165746
rect 87030 165682 87046 165746
rect 87110 165682 87126 165746
rect 87190 165682 87198 165746
rect 86878 165681 87198 165682
rect 83311 165404 83377 165407
rect 83311 165402 85352 165404
rect 83311 165346 83316 165402
rect 83372 165346 85352 165402
rect 83311 165344 85352 165346
rect 83311 165341 83377 165344
rect 878 165202 1198 165203
rect 878 165138 886 165202
rect 950 165138 966 165202
rect 1030 165138 1046 165202
rect 1110 165138 1126 165202
rect 1190 165138 1198 165202
rect 878 165137 1198 165138
rect 84878 165202 85198 165203
rect 84878 165138 84886 165202
rect 84950 165138 84966 165202
rect 85030 165138 85046 165202
rect 85110 165138 85126 165202
rect 85190 165138 85198 165202
rect 84878 165137 85198 165138
rect 85292 165132 85352 165344
rect 88454 165132 88934 165162
rect 85292 165072 88934 165132
rect 88454 165042 88934 165072
rect 84415 164998 84481 164999
rect 84364 164996 84370 164998
rect 84324 164936 84370 164996
rect 84434 164994 84481 164998
rect 84476 164938 84481 164994
rect 84364 164934 84370 164936
rect 84434 164934 84481 164938
rect 84415 164933 84481 164934
rect 84599 164862 84665 164863
rect 84548 164860 84554 164862
rect 84508 164800 84554 164860
rect 84618 164858 84665 164862
rect 84660 164802 84665 164858
rect 84548 164798 84554 164800
rect 84618 164798 84665 164802
rect 84599 164797 84665 164798
rect 2878 164658 3198 164659
rect 2878 164594 2886 164658
rect 2950 164594 2966 164658
rect 3030 164594 3046 164658
rect 3110 164594 3126 164658
rect 3190 164594 3198 164658
rect 2878 164593 3198 164594
rect 86878 164658 87198 164659
rect 86878 164594 86886 164658
rect 86950 164594 86966 164658
rect 87030 164594 87046 164658
rect 87110 164594 87126 164658
rect 87190 164594 87198 164658
rect 86878 164593 87198 164594
rect 84231 164452 84297 164455
rect 84364 164452 84370 164454
rect 84231 164450 84370 164452
rect 84231 164394 84236 164450
rect 84292 164394 84370 164450
rect 84231 164392 84370 164394
rect 84231 164389 84297 164392
rect 84364 164390 84370 164392
rect 84434 164390 84440 164454
rect 84415 164316 84481 164319
rect 84548 164316 84554 164318
rect 84415 164314 84554 164316
rect 84415 164258 84420 164314
rect 84476 164258 84554 164314
rect 84415 164256 84554 164258
rect 84415 164253 84481 164256
rect 84548 164254 84554 164256
rect 84618 164254 84624 164318
rect 878 164114 1198 164115
rect 878 164050 886 164114
rect 950 164050 966 164114
rect 1030 164050 1046 164114
rect 1110 164050 1126 164114
rect 1190 164050 1198 164114
rect 878 164049 1198 164050
rect 84878 164114 85198 164115
rect 84878 164050 84886 164114
rect 84950 164050 84966 164114
rect 85030 164050 85046 164114
rect 85110 164050 85126 164114
rect 85190 164050 85198 164114
rect 84878 164049 85198 164050
rect 85151 163908 85217 163911
rect 88454 163908 88934 163938
rect 85151 163906 88934 163908
rect 85151 163850 85156 163906
rect 85212 163850 88934 163906
rect 85151 163848 88934 163850
rect 85151 163845 85217 163848
rect 88454 163818 88934 163848
rect 2878 163570 3198 163571
rect 2878 163506 2886 163570
rect 2950 163506 2966 163570
rect 3030 163506 3046 163570
rect 3110 163506 3126 163570
rect 3190 163506 3198 163570
rect 2878 163505 3198 163506
rect 86878 163570 87198 163571
rect 86878 163506 86886 163570
rect 86950 163506 86966 163570
rect 87030 163506 87046 163570
rect 87110 163506 87126 163570
rect 87190 163506 87198 163570
rect 86878 163505 87198 163506
rect 878 163026 1198 163027
rect 878 162962 886 163026
rect 950 162962 966 163026
rect 1030 162962 1046 163026
rect 1110 162962 1126 163026
rect 1190 162962 1198 163026
rect 878 162961 1198 162962
rect 84878 163026 85198 163027
rect 84878 162962 84886 163026
rect 84950 162962 84966 163026
rect 85030 162962 85046 163026
rect 85110 162962 85126 163026
rect 85190 162962 85198 163026
rect 84878 162961 85198 162962
rect 84323 162684 84389 162687
rect 88454 162684 88934 162714
rect 84323 162682 88934 162684
rect 84323 162626 84328 162682
rect 84384 162626 88934 162682
rect 84323 162624 88934 162626
rect 84323 162621 84389 162624
rect 88454 162594 88934 162624
rect 2878 162482 3198 162483
rect 2878 162418 2886 162482
rect 2950 162418 2966 162482
rect 3030 162418 3046 162482
rect 3110 162418 3126 162482
rect 3190 162418 3198 162482
rect 2878 162417 3198 162418
rect 86878 162482 87198 162483
rect 86878 162418 86886 162482
rect 86950 162418 86966 162482
rect 87030 162418 87046 162482
rect 87110 162418 87126 162482
rect 87190 162418 87198 162482
rect 86878 162417 87198 162418
rect 878 161938 1198 161939
rect 878 161874 886 161938
rect 950 161874 966 161938
rect 1030 161874 1046 161938
rect 1110 161874 1126 161938
rect 1190 161874 1198 161938
rect 878 161873 1198 161874
rect 84878 161938 85198 161939
rect 84878 161874 84886 161938
rect 84950 161874 84966 161938
rect 85030 161874 85046 161938
rect 85110 161874 85126 161938
rect 85190 161874 85198 161938
rect 84878 161873 85198 161874
rect 85151 161596 85217 161599
rect 85151 161594 87376 161596
rect 85151 161538 85156 161594
rect 85212 161538 87376 161594
rect 85151 161536 87376 161538
rect 85151 161533 85217 161536
rect 87316 161460 87376 161536
rect 88454 161460 88934 161490
rect 87316 161400 88934 161460
rect 2878 161394 3198 161395
rect 2878 161330 2886 161394
rect 2950 161330 2966 161394
rect 3030 161330 3046 161394
rect 3110 161330 3126 161394
rect 3190 161330 3198 161394
rect 2878 161329 3198 161330
rect 86878 161394 87198 161395
rect 86878 161330 86886 161394
rect 86950 161330 86966 161394
rect 87030 161330 87046 161394
rect 87110 161330 87126 161394
rect 87190 161330 87198 161394
rect 88454 161370 88934 161400
rect 86878 161329 87198 161330
rect 878 160850 1198 160851
rect 878 160786 886 160850
rect 950 160786 966 160850
rect 1030 160786 1046 160850
rect 1110 160786 1126 160850
rect 1190 160786 1198 160850
rect 878 160785 1198 160786
rect 84878 160850 85198 160851
rect 84878 160786 84886 160850
rect 84950 160786 84966 160850
rect 85030 160786 85046 160850
rect 85110 160786 85126 160850
rect 85190 160786 85198 160850
rect 84878 160785 85198 160786
rect 84599 160508 84665 160511
rect 84599 160506 87376 160508
rect 84599 160450 84604 160506
rect 84660 160450 87376 160506
rect 84599 160448 87376 160450
rect 84599 160445 84665 160448
rect 2878 160306 3198 160307
rect 2878 160242 2886 160306
rect 2950 160242 2966 160306
rect 3030 160242 3046 160306
rect 3110 160242 3126 160306
rect 3190 160242 3198 160306
rect 2878 160241 3198 160242
rect 86878 160306 87198 160307
rect 86878 160242 86886 160306
rect 86950 160242 86966 160306
rect 87030 160242 87046 160306
rect 87110 160242 87126 160306
rect 87190 160242 87198 160306
rect 86878 160241 87198 160242
rect 87316 160236 87376 160448
rect 88454 160236 88934 160266
rect 87316 160176 88934 160236
rect 88454 160146 88934 160176
rect 878 159762 1198 159763
rect 878 159698 886 159762
rect 950 159698 966 159762
rect 1030 159698 1046 159762
rect 1110 159698 1126 159762
rect 1190 159698 1198 159762
rect 878 159697 1198 159698
rect 84878 159762 85198 159763
rect 84878 159698 84886 159762
rect 84950 159698 84966 159762
rect 85030 159698 85046 159762
rect 85110 159698 85126 159762
rect 85190 159698 85198 159762
rect 84878 159697 85198 159698
rect 84323 159420 84389 159423
rect 84323 159418 87376 159420
rect 84323 159362 84328 159418
rect 84384 159362 87376 159418
rect 84323 159360 87376 159362
rect 84323 159357 84389 159360
rect 2878 159218 3198 159219
rect 2878 159154 2886 159218
rect 2950 159154 2966 159218
rect 3030 159154 3046 159218
rect 3110 159154 3126 159218
rect 3190 159154 3198 159218
rect 2878 159153 3198 159154
rect 86878 159218 87198 159219
rect 86878 159154 86886 159218
rect 86950 159154 86966 159218
rect 87030 159154 87046 159218
rect 87110 159154 87126 159218
rect 87190 159154 87198 159218
rect 86878 159153 87198 159154
rect 87316 159148 87376 159360
rect 88454 159148 88934 159178
rect 87316 159088 88934 159148
rect 88454 159058 88934 159088
rect 878 158674 1198 158675
rect 878 158610 886 158674
rect 950 158610 966 158674
rect 1030 158610 1046 158674
rect 1110 158610 1126 158674
rect 1190 158610 1198 158674
rect 878 158609 1198 158610
rect 84878 158674 85198 158675
rect 84878 158610 84886 158674
rect 84950 158610 84966 158674
rect 85030 158610 85046 158674
rect 85110 158610 85126 158674
rect 85190 158610 85198 158674
rect 84878 158609 85198 158610
rect 2878 158130 3198 158131
rect 2878 158066 2886 158130
rect 2950 158066 2966 158130
rect 3030 158066 3046 158130
rect 3110 158066 3126 158130
rect 3190 158066 3198 158130
rect 2878 158065 3198 158066
rect 86878 158130 87198 158131
rect 86878 158066 86886 158130
rect 86950 158066 86966 158130
rect 87030 158066 87046 158130
rect 87110 158066 87126 158130
rect 87190 158066 87198 158130
rect 86878 158065 87198 158066
rect 83955 157924 84021 157927
rect 88454 157924 88934 157954
rect 83955 157922 88934 157924
rect 83955 157866 83960 157922
rect 84016 157866 88934 157922
rect 83955 157864 88934 157866
rect 83955 157861 84021 157864
rect 88454 157834 88934 157864
rect 878 157586 1198 157587
rect 878 157522 886 157586
rect 950 157522 966 157586
rect 1030 157522 1046 157586
rect 1110 157522 1126 157586
rect 1190 157522 1198 157586
rect 878 157521 1198 157522
rect 84878 157586 85198 157587
rect 84878 157522 84886 157586
rect 84950 157522 84966 157586
rect 85030 157522 85046 157586
rect 85110 157522 85126 157586
rect 85190 157522 85198 157586
rect 84878 157521 85198 157522
rect 2878 157042 3198 157043
rect 2878 156978 2886 157042
rect 2950 156978 2966 157042
rect 3030 156978 3046 157042
rect 3110 156978 3126 157042
rect 3190 156978 3198 157042
rect 2878 156977 3198 156978
rect 86878 157042 87198 157043
rect 86878 156978 86886 157042
rect 86950 156978 86966 157042
rect 87030 156978 87046 157042
rect 87110 156978 87126 157042
rect 87190 156978 87198 157042
rect 86878 156977 87198 156978
rect 85059 156700 85125 156703
rect 88454 156700 88934 156730
rect 85059 156698 88934 156700
rect 85059 156642 85064 156698
rect 85120 156642 88934 156698
rect 85059 156640 88934 156642
rect 85059 156637 85125 156640
rect 88454 156610 88934 156640
rect 878 156498 1198 156499
rect 878 156434 886 156498
rect 950 156434 966 156498
rect 1030 156434 1046 156498
rect 1110 156434 1126 156498
rect 1190 156434 1198 156498
rect 878 156433 1198 156434
rect 84878 156498 85198 156499
rect 84878 156434 84886 156498
rect 84950 156434 84966 156498
rect 85030 156434 85046 156498
rect 85110 156434 85126 156498
rect 85190 156434 85198 156498
rect 84878 156433 85198 156434
rect 2878 155954 3198 155955
rect 2878 155890 2886 155954
rect 2950 155890 2966 155954
rect 3030 155890 3046 155954
rect 3110 155890 3126 155954
rect 3190 155890 3198 155954
rect 2878 155889 3198 155890
rect 86878 155954 87198 155955
rect 86878 155890 86886 155954
rect 86950 155890 86966 155954
rect 87030 155890 87046 155954
rect 87110 155890 87126 155954
rect 87190 155890 87198 155954
rect 86878 155889 87198 155890
rect 84415 155612 84481 155615
rect 84415 155610 85536 155612
rect 84415 155554 84420 155610
rect 84476 155554 85536 155610
rect 84415 155552 85536 155554
rect 84415 155549 84481 155552
rect 85476 155476 85536 155552
rect 88454 155476 88934 155506
rect 85476 155416 88934 155476
rect 878 155410 1198 155411
rect 878 155346 886 155410
rect 950 155346 966 155410
rect 1030 155346 1046 155410
rect 1110 155346 1126 155410
rect 1190 155346 1198 155410
rect 878 155345 1198 155346
rect 84878 155410 85198 155411
rect 84878 155346 84886 155410
rect 84950 155346 84966 155410
rect 85030 155346 85046 155410
rect 85110 155346 85126 155410
rect 85190 155346 85198 155410
rect 88454 155386 88934 155416
rect 84878 155345 85198 155346
rect 2878 154866 3198 154867
rect 2878 154802 2886 154866
rect 2950 154802 2966 154866
rect 3030 154802 3046 154866
rect 3110 154802 3126 154866
rect 3190 154802 3198 154866
rect 2878 154801 3198 154802
rect 86878 154866 87198 154867
rect 86878 154802 86886 154866
rect 86950 154802 86966 154866
rect 87030 154802 87046 154866
rect 87110 154802 87126 154866
rect 87190 154802 87198 154866
rect 86878 154801 87198 154802
rect 878 154322 1198 154323
rect 878 154258 886 154322
rect 950 154258 966 154322
rect 1030 154258 1046 154322
rect 1110 154258 1126 154322
rect 1190 154258 1198 154322
rect 878 154257 1198 154258
rect 84878 154322 85198 154323
rect 84878 154258 84886 154322
rect 84950 154258 84966 154322
rect 85030 154258 85046 154322
rect 85110 154258 85126 154322
rect 85190 154258 85198 154322
rect 84878 154257 85198 154258
rect 85335 154252 85401 154255
rect 88454 154252 88934 154282
rect 85335 154250 88934 154252
rect 85335 154194 85340 154250
rect 85396 154194 88934 154250
rect 85335 154192 88934 154194
rect 85335 154189 85401 154192
rect 88454 154162 88934 154192
rect 2878 153778 3198 153779
rect 2878 153714 2886 153778
rect 2950 153714 2966 153778
rect 3030 153714 3046 153778
rect 3110 153714 3126 153778
rect 3190 153714 3198 153778
rect 2878 153713 3198 153714
rect 86878 153778 87198 153779
rect 86878 153714 86886 153778
rect 86950 153714 86966 153778
rect 87030 153714 87046 153778
rect 87110 153714 87126 153778
rect 87190 153714 87198 153778
rect 86878 153713 87198 153714
rect 878 153234 1198 153235
rect 878 153170 886 153234
rect 950 153170 966 153234
rect 1030 153170 1046 153234
rect 1110 153170 1126 153234
rect 1190 153170 1198 153234
rect 878 153169 1198 153170
rect 84878 153234 85198 153235
rect 84878 153170 84886 153234
rect 84950 153170 84966 153234
rect 85030 153170 85046 153234
rect 85110 153170 85126 153234
rect 85190 153170 85198 153234
rect 84878 153169 85198 153170
rect 84507 153028 84573 153031
rect 88454 153028 88934 153058
rect 84507 153026 88934 153028
rect 84507 152970 84512 153026
rect 84568 152970 88934 153026
rect 84507 152968 88934 152970
rect 84507 152965 84573 152968
rect 88454 152938 88934 152968
rect 2878 152690 3198 152691
rect 2878 152626 2886 152690
rect 2950 152626 2966 152690
rect 3030 152626 3046 152690
rect 3110 152626 3126 152690
rect 3190 152626 3198 152690
rect 2878 152625 3198 152626
rect 86878 152690 87198 152691
rect 86878 152626 86886 152690
rect 86950 152626 86966 152690
rect 87030 152626 87046 152690
rect 87110 152626 87126 152690
rect 87190 152626 87198 152690
rect 86878 152625 87198 152626
rect 878 152146 1198 152147
rect 878 152082 886 152146
rect 950 152082 966 152146
rect 1030 152082 1046 152146
rect 1110 152082 1126 152146
rect 1190 152082 1198 152146
rect 878 152081 1198 152082
rect 84878 152146 85198 152147
rect 84878 152082 84886 152146
rect 84950 152082 84966 152146
rect 85030 152082 85046 152146
rect 85110 152082 85126 152146
rect 85190 152082 85198 152146
rect 84878 152081 85198 152082
rect 84691 151940 84757 151943
rect 88454 151940 88934 151970
rect 84691 151938 88934 151940
rect 84691 151882 84696 151938
rect 84752 151882 88934 151938
rect 84691 151880 88934 151882
rect 84691 151877 84757 151880
rect 88454 151850 88934 151880
rect 5571 151806 5637 151807
rect 5571 151804 5618 151806
rect 5526 151802 5618 151804
rect 5526 151746 5576 151802
rect 5526 151744 5618 151746
rect 5571 151742 5618 151744
rect 5682 151742 5688 151806
rect 82340 151742 82346 151806
rect 82410 151804 82416 151806
rect 82483 151804 82549 151807
rect 82410 151802 82549 151804
rect 82410 151746 82488 151802
rect 82544 151746 82549 151802
rect 82410 151744 82549 151746
rect 82410 151742 82416 151744
rect 5571 151741 5637 151742
rect 82483 151741 82549 151744
rect 2878 151602 3198 151603
rect 2878 151538 2886 151602
rect 2950 151538 2966 151602
rect 3030 151538 3046 151602
rect 3110 151538 3126 151602
rect 3190 151538 3198 151602
rect 2878 151537 3198 151538
rect 86878 151602 87198 151603
rect 86878 151538 86886 151602
rect 86950 151538 86966 151602
rect 87030 151538 87046 151602
rect 87110 151538 87126 151602
rect 87190 151538 87198 151602
rect 86878 151537 87198 151538
rect 878 151058 1198 151059
rect 878 150994 886 151058
rect 950 150994 966 151058
rect 1030 150994 1046 151058
rect 1110 150994 1126 151058
rect 1190 150994 1198 151058
rect 878 150993 1198 150994
rect 84878 151058 85198 151059
rect 84878 150994 84886 151058
rect 84950 150994 84966 151058
rect 85030 150994 85046 151058
rect 85110 150994 85126 151058
rect 85190 150994 85198 151058
rect 84878 150993 85198 150994
rect 83219 150716 83285 150719
rect 88454 150716 88934 150746
rect 83219 150714 88934 150716
rect 83219 150658 83224 150714
rect 83280 150658 88934 150714
rect 83219 150656 88934 150658
rect 83219 150653 83285 150656
rect 88454 150626 88934 150656
rect 2878 150514 3198 150515
rect 2878 150450 2886 150514
rect 2950 150450 2966 150514
rect 3030 150450 3046 150514
rect 3110 150450 3126 150514
rect 3190 150450 3198 150514
rect 2878 150449 3198 150450
rect 86878 150514 87198 150515
rect 86878 150450 86886 150514
rect 86950 150450 86966 150514
rect 87030 150450 87046 150514
rect 87110 150450 87126 150514
rect 87190 150450 87198 150514
rect 86878 150449 87198 150450
rect 878 149970 1198 149971
rect 878 149906 886 149970
rect 950 149906 966 149970
rect 1030 149906 1046 149970
rect 1110 149906 1126 149970
rect 1190 149906 1198 149970
rect 878 149905 1198 149906
rect 84878 149970 85198 149971
rect 84878 149906 84886 149970
rect 84950 149906 84966 149970
rect 85030 149906 85046 149970
rect 85110 149906 85126 149970
rect 85190 149906 85198 149970
rect 84878 149905 85198 149906
rect 83955 149628 84021 149631
rect 83955 149626 87560 149628
rect 83955 149570 83960 149626
rect 84016 149570 87560 149626
rect 83955 149568 87560 149570
rect 83955 149565 84021 149568
rect 87500 149492 87560 149568
rect 88454 149492 88934 149522
rect 87500 149432 88934 149492
rect 2878 149426 3198 149427
rect 2878 149362 2886 149426
rect 2950 149362 2966 149426
rect 3030 149362 3046 149426
rect 3110 149362 3126 149426
rect 3190 149362 3198 149426
rect 2878 149361 3198 149362
rect 86878 149426 87198 149427
rect 86878 149362 86886 149426
rect 86950 149362 86966 149426
rect 87030 149362 87046 149426
rect 87110 149362 87126 149426
rect 87190 149362 87198 149426
rect 88454 149402 88934 149432
rect 86878 149361 87198 149362
rect 878 148882 1198 148883
rect 878 148818 886 148882
rect 950 148818 966 148882
rect 1030 148818 1046 148882
rect 1110 148818 1126 148882
rect 1190 148818 1198 148882
rect 878 148817 1198 148818
rect 84878 148882 85198 148883
rect 84878 148818 84886 148882
rect 84950 148818 84966 148882
rect 85030 148818 85046 148882
rect 85110 148818 85126 148882
rect 85190 148818 85198 148882
rect 84878 148817 85198 148818
rect 83955 148540 84021 148543
rect 83955 148538 87560 148540
rect 83955 148482 83960 148538
rect 84016 148482 87560 148538
rect 83955 148480 87560 148482
rect 83955 148477 84021 148480
rect 2878 148338 3198 148339
rect 2878 148274 2886 148338
rect 2950 148274 2966 148338
rect 3030 148274 3046 148338
rect 3110 148274 3126 148338
rect 3190 148274 3198 148338
rect 2878 148273 3198 148274
rect 86878 148338 87198 148339
rect 86878 148274 86886 148338
rect 86950 148274 86966 148338
rect 87030 148274 87046 148338
rect 87110 148274 87126 148338
rect 87190 148274 87198 148338
rect 86878 148273 87198 148274
rect 87500 148268 87560 148480
rect 88454 148268 88934 148298
rect 87500 148208 88934 148268
rect 88454 148178 88934 148208
rect 878 147794 1198 147795
rect 878 147730 886 147794
rect 950 147730 966 147794
rect 1030 147730 1046 147794
rect 1110 147730 1126 147794
rect 1190 147730 1198 147794
rect 878 147729 1198 147730
rect 84878 147794 85198 147795
rect 84878 147730 84886 147794
rect 84950 147730 84966 147794
rect 85030 147730 85046 147794
rect 85110 147730 85126 147794
rect 85190 147730 85198 147794
rect 84878 147729 85198 147730
rect 2878 147250 3198 147251
rect 2878 147186 2886 147250
rect 2950 147186 2966 147250
rect 3030 147186 3046 147250
rect 3110 147186 3126 147250
rect 3190 147186 3198 147250
rect 2878 147185 3198 147186
rect 86878 147250 87198 147251
rect 86878 147186 86886 147250
rect 86950 147186 86966 147250
rect 87030 147186 87046 147250
rect 87110 147186 87126 147250
rect 87190 147186 87198 147250
rect 86878 147185 87198 147186
rect 83955 147044 84021 147047
rect 88454 147044 88934 147074
rect 83955 147042 88934 147044
rect 83955 146986 83960 147042
rect 84016 146986 88934 147042
rect 83955 146984 88934 146986
rect 83955 146981 84021 146984
rect 88454 146954 88934 146984
rect 3731 146772 3797 146775
rect 4007 146772 4073 146775
rect 3731 146770 4073 146772
rect 3731 146714 3736 146770
rect 3792 146714 4012 146770
rect 4068 146714 4073 146770
rect 3731 146712 4073 146714
rect 3731 146709 3797 146712
rect 4007 146709 4073 146712
rect 878 146706 1198 146707
rect 878 146642 886 146706
rect 950 146642 966 146706
rect 1030 146642 1046 146706
rect 1110 146642 1126 146706
rect 1190 146642 1198 146706
rect 878 146641 1198 146642
rect 84878 146706 85198 146707
rect 84878 146642 84886 146706
rect 84950 146642 84966 146706
rect 85030 146642 85046 146706
rect 85110 146642 85126 146706
rect 85190 146642 85198 146706
rect 84878 146641 85198 146642
rect 2878 146162 3198 146163
rect 2878 146098 2886 146162
rect 2950 146098 2966 146162
rect 3030 146098 3046 146162
rect 3110 146098 3126 146162
rect 3190 146098 3198 146162
rect 2878 146097 3198 146098
rect 86878 146162 87198 146163
rect 86878 146098 86886 146162
rect 86950 146098 86966 146162
rect 87030 146098 87046 146162
rect 87110 146098 87126 146162
rect 87190 146098 87198 146162
rect 86878 146097 87198 146098
rect 83955 145820 84021 145823
rect 88454 145820 88934 145850
rect 83955 145818 88934 145820
rect 83955 145762 83960 145818
rect 84016 145762 88934 145818
rect 83955 145760 88934 145762
rect 83955 145757 84021 145760
rect 88454 145730 88934 145760
rect 878 145618 1198 145619
rect 878 145554 886 145618
rect 950 145554 966 145618
rect 1030 145554 1046 145618
rect 1110 145554 1126 145618
rect 1190 145554 1198 145618
rect 878 145553 1198 145554
rect 84878 145618 85198 145619
rect 84878 145554 84886 145618
rect 84950 145554 84966 145618
rect 85030 145554 85046 145618
rect 85110 145554 85126 145618
rect 85190 145554 85198 145618
rect 84878 145553 85198 145554
rect 2878 145074 3198 145075
rect 2878 145010 2886 145074
rect 2950 145010 2966 145074
rect 3030 145010 3046 145074
rect 3110 145010 3126 145074
rect 3190 145010 3198 145074
rect 2878 145009 3198 145010
rect 86878 145074 87198 145075
rect 86878 145010 86886 145074
rect 86950 145010 86966 145074
rect 87030 145010 87046 145074
rect 87110 145010 87126 145074
rect 87190 145010 87198 145074
rect 86878 145009 87198 145010
rect 83955 144732 84021 144735
rect 88454 144732 88934 144762
rect 83955 144730 88934 144732
rect 83955 144674 83960 144730
rect 84016 144674 88934 144730
rect 83955 144672 88934 144674
rect 83955 144669 84021 144672
rect 88454 144642 88934 144672
rect 878 144530 1198 144531
rect 878 144466 886 144530
rect 950 144466 966 144530
rect 1030 144466 1046 144530
rect 1110 144466 1126 144530
rect 1190 144466 1198 144530
rect 878 144465 1198 144466
rect 84878 144530 85198 144531
rect 84878 144466 84886 144530
rect 84950 144466 84966 144530
rect 85030 144466 85046 144530
rect 85110 144466 85126 144530
rect 85190 144466 85198 144530
rect 84878 144465 85198 144466
rect 2878 143986 3198 143987
rect 2878 143922 2886 143986
rect 2950 143922 2966 143986
rect 3030 143922 3046 143986
rect 3110 143922 3126 143986
rect 3190 143922 3198 143986
rect 2878 143921 3198 143922
rect 86878 143986 87198 143987
rect 86878 143922 86886 143986
rect 86950 143922 86966 143986
rect 87030 143922 87046 143986
rect 87110 143922 87126 143986
rect 87190 143922 87198 143986
rect 86878 143921 87198 143922
rect 84231 143780 84297 143783
rect 84231 143778 85352 143780
rect 84231 143722 84236 143778
rect 84292 143722 85352 143778
rect 84231 143720 85352 143722
rect 84231 143717 84297 143720
rect 85292 143508 85352 143720
rect 88454 143508 88934 143538
rect 85292 143448 88934 143508
rect 878 143442 1198 143443
rect 878 143378 886 143442
rect 950 143378 966 143442
rect 1030 143378 1046 143442
rect 1110 143378 1126 143442
rect 1190 143378 1198 143442
rect 878 143377 1198 143378
rect 84878 143442 85198 143443
rect 84878 143378 84886 143442
rect 84950 143378 84966 143442
rect 85030 143378 85046 143442
rect 85110 143378 85126 143442
rect 85190 143378 85198 143442
rect 88454 143418 88934 143448
rect 84878 143377 85198 143378
rect 2878 142898 3198 142899
rect 2878 142834 2886 142898
rect 2950 142834 2966 142898
rect 3030 142834 3046 142898
rect 3110 142834 3126 142898
rect 3190 142834 3198 142898
rect 2878 142833 3198 142834
rect 86878 142898 87198 142899
rect 86878 142834 86886 142898
rect 86950 142834 86966 142898
rect 87030 142834 87046 142898
rect 87110 142834 87126 142898
rect 87190 142834 87198 142898
rect 86878 142833 87198 142834
rect 878 142354 1198 142355
rect 878 142290 886 142354
rect 950 142290 966 142354
rect 1030 142290 1046 142354
rect 1110 142290 1126 142354
rect 1190 142290 1198 142354
rect 878 142289 1198 142290
rect 84878 142354 85198 142355
rect 84878 142290 84886 142354
rect 84950 142290 84966 142354
rect 85030 142290 85046 142354
rect 85110 142290 85126 142354
rect 85190 142290 85198 142354
rect 84878 142289 85198 142290
rect 88454 142284 88934 142314
rect 85292 142224 88934 142284
rect 84507 142148 84573 142151
rect 85292 142148 85352 142224
rect 88454 142194 88934 142224
rect 84507 142146 85352 142148
rect 84507 142090 84512 142146
rect 84568 142090 85352 142146
rect 84507 142088 85352 142090
rect 84507 142085 84573 142088
rect 2878 141810 3198 141811
rect 2878 141746 2886 141810
rect 2950 141746 2966 141810
rect 3030 141746 3046 141810
rect 3110 141746 3126 141810
rect 3190 141746 3198 141810
rect 2878 141745 3198 141746
rect 86878 141810 87198 141811
rect 86878 141746 86886 141810
rect 86950 141746 86966 141810
rect 87030 141746 87046 141810
rect 87110 141746 87126 141810
rect 87190 141746 87198 141810
rect 86878 141745 87198 141746
rect 878 141266 1198 141267
rect 878 141202 886 141266
rect 950 141202 966 141266
rect 1030 141202 1046 141266
rect 1110 141202 1126 141266
rect 1190 141202 1198 141266
rect 878 141201 1198 141202
rect 84878 141266 85198 141267
rect 84878 141202 84886 141266
rect 84950 141202 84966 141266
rect 85030 141202 85046 141266
rect 85110 141202 85126 141266
rect 85190 141202 85198 141266
rect 84878 141201 85198 141202
rect 82340 140998 82346 141062
rect 82410 141060 82416 141062
rect 88454 141060 88934 141090
rect 82410 141000 88934 141060
rect 82410 140998 82416 141000
rect 88454 140970 88934 141000
rect 2878 140722 3198 140723
rect 2878 140658 2886 140722
rect 2950 140658 2966 140722
rect 3030 140658 3046 140722
rect 3110 140658 3126 140722
rect 3190 140658 3198 140722
rect 2878 140657 3198 140658
rect 86878 140722 87198 140723
rect 86878 140658 86886 140722
rect 86950 140658 86966 140722
rect 87030 140658 87046 140722
rect 87110 140658 87126 140722
rect 87190 140658 87198 140722
rect 86878 140657 87198 140658
rect 878 140178 1198 140179
rect 878 140114 886 140178
rect 950 140114 966 140178
rect 1030 140114 1046 140178
rect 1110 140114 1126 140178
rect 1190 140114 1198 140178
rect 878 140113 1198 140114
rect 84878 140178 85198 140179
rect 84878 140114 84886 140178
rect 84950 140114 84966 140178
rect 85030 140114 85046 140178
rect 85110 140114 85126 140178
rect 85190 140114 85198 140178
rect 84878 140113 85198 140114
rect 84599 139836 84665 139839
rect 88454 139836 88934 139866
rect 84599 139834 88934 139836
rect 84599 139778 84604 139834
rect 84660 139778 88934 139834
rect 84599 139776 88934 139778
rect 84599 139773 84665 139776
rect 88454 139746 88934 139776
rect 2878 139634 3198 139635
rect 2878 139570 2886 139634
rect 2950 139570 2966 139634
rect 3030 139570 3046 139634
rect 3110 139570 3126 139634
rect 3190 139570 3198 139634
rect 2878 139569 3198 139570
rect 86878 139634 87198 139635
rect 86878 139570 86886 139634
rect 86950 139570 86966 139634
rect 87030 139570 87046 139634
rect 87110 139570 87126 139634
rect 87190 139570 87198 139634
rect 86878 139569 87198 139570
rect 878 139090 1198 139091
rect 878 139026 886 139090
rect 950 139026 966 139090
rect 1030 139026 1046 139090
rect 1110 139026 1126 139090
rect 1190 139026 1198 139090
rect 878 139025 1198 139026
rect 84878 139090 85198 139091
rect 84878 139026 84886 139090
rect 84950 139026 84966 139090
rect 85030 139026 85046 139090
rect 85110 139026 85126 139090
rect 85190 139026 85198 139090
rect 84878 139025 85198 139026
rect 88454 138612 88934 138642
rect 87500 138552 88934 138612
rect 2878 138546 3198 138547
rect 2878 138482 2886 138546
rect 2950 138482 2966 138546
rect 3030 138482 3046 138546
rect 3110 138482 3126 138546
rect 3190 138482 3198 138546
rect 2878 138481 3198 138482
rect 86878 138546 87198 138547
rect 86878 138482 86886 138546
rect 86950 138482 86966 138546
rect 87030 138482 87046 138546
rect 87110 138482 87126 138546
rect 87190 138482 87198 138546
rect 86878 138481 87198 138482
rect 84231 138340 84297 138343
rect 87500 138340 87560 138552
rect 88454 138522 88934 138552
rect 84231 138338 87560 138340
rect 84231 138282 84236 138338
rect 84292 138282 87560 138338
rect 84231 138280 87560 138282
rect 84231 138277 84297 138280
rect 878 138002 1198 138003
rect 878 137938 886 138002
rect 950 137938 966 138002
rect 1030 137938 1046 138002
rect 1110 137938 1126 138002
rect 1190 137938 1198 138002
rect 878 137937 1198 137938
rect 84878 138002 85198 138003
rect 84878 137938 84886 138002
rect 84950 137938 84966 138002
rect 85030 137938 85046 138002
rect 85110 137938 85126 138002
rect 85190 137938 85198 138002
rect 84878 137937 85198 137938
rect 2878 137458 3198 137459
rect 2878 137394 2886 137458
rect 2950 137394 2966 137458
rect 3030 137394 3046 137458
rect 3110 137394 3126 137458
rect 3190 137394 3198 137458
rect 2878 137393 3198 137394
rect 86878 137458 87198 137459
rect 86878 137394 86886 137458
rect 86950 137394 86966 137458
rect 87030 137394 87046 137458
rect 87110 137394 87126 137458
rect 87190 137394 87198 137458
rect 86878 137393 87198 137394
rect 88454 137388 88934 137418
rect 87500 137328 88934 137388
rect 85795 137252 85861 137255
rect 87500 137252 87560 137328
rect 88454 137298 88934 137328
rect 85795 137250 87560 137252
rect 85795 137194 85800 137250
rect 85856 137194 87560 137250
rect 85795 137192 87560 137194
rect 85795 137189 85861 137192
rect 878 136914 1198 136915
rect 878 136850 886 136914
rect 950 136850 966 136914
rect 1030 136850 1046 136914
rect 1110 136850 1126 136914
rect 1190 136850 1198 136914
rect 878 136849 1198 136850
rect 84878 136914 85198 136915
rect 84878 136850 84886 136914
rect 84950 136850 84966 136914
rect 85030 136850 85046 136914
rect 85110 136850 85126 136914
rect 85190 136850 85198 136914
rect 84878 136849 85198 136850
rect 2878 136370 3198 136371
rect 2878 136306 2886 136370
rect 2950 136306 2966 136370
rect 3030 136306 3046 136370
rect 3110 136306 3126 136370
rect 3190 136306 3198 136370
rect 2878 136305 3198 136306
rect 86878 136370 87198 136371
rect 86878 136306 86886 136370
rect 86950 136306 86966 136370
rect 87030 136306 87046 136370
rect 87110 136306 87126 136370
rect 87190 136306 87198 136370
rect 86878 136305 87198 136306
rect 88454 136300 88934 136330
rect 87500 136240 88934 136300
rect 83311 136164 83377 136167
rect 87500 136164 87560 136240
rect 88454 136210 88934 136240
rect 83311 136162 87560 136164
rect 83311 136106 83316 136162
rect 83372 136106 87560 136162
rect 83311 136104 87560 136106
rect 83311 136101 83377 136104
rect 878 135826 1198 135827
rect 878 135762 886 135826
rect 950 135762 966 135826
rect 1030 135762 1046 135826
rect 1110 135762 1126 135826
rect 1190 135762 1198 135826
rect 878 135761 1198 135762
rect 84878 135826 85198 135827
rect 84878 135762 84886 135826
rect 84950 135762 84966 135826
rect 85030 135762 85046 135826
rect 85110 135762 85126 135826
rect 85190 135762 85198 135826
rect 84878 135761 85198 135762
rect 2878 135282 3198 135283
rect 2878 135218 2886 135282
rect 2950 135218 2966 135282
rect 3030 135218 3046 135282
rect 3110 135218 3126 135282
rect 3190 135218 3198 135282
rect 2878 135217 3198 135218
rect 86878 135282 87198 135283
rect 86878 135218 86886 135282
rect 86950 135218 86966 135282
rect 87030 135218 87046 135282
rect 87110 135218 87126 135282
rect 87190 135218 87198 135282
rect 86878 135217 87198 135218
rect 84691 135076 84757 135079
rect 88454 135076 88934 135106
rect 84691 135074 88934 135076
rect 84691 135018 84696 135074
rect 84752 135018 88934 135074
rect 84691 135016 88934 135018
rect 84691 135013 84757 135016
rect 88454 134986 88934 135016
rect 878 134738 1198 134739
rect 878 134674 886 134738
rect 950 134674 966 134738
rect 1030 134674 1046 134738
rect 1110 134674 1126 134738
rect 1190 134674 1198 134738
rect 878 134673 1198 134674
rect 84878 134738 85198 134739
rect 84878 134674 84886 134738
rect 84950 134674 84966 134738
rect 85030 134674 85046 134738
rect 85110 134674 85126 134738
rect 85190 134674 85198 134738
rect 84878 134673 85198 134674
rect 2878 134194 3198 134195
rect 2878 134130 2886 134194
rect 2950 134130 2966 134194
rect 3030 134130 3046 134194
rect 3110 134130 3126 134194
rect 3190 134130 3198 134194
rect 2878 134129 3198 134130
rect 86878 134194 87198 134195
rect 86878 134130 86886 134194
rect 86950 134130 86966 134194
rect 87030 134130 87046 134194
rect 87110 134130 87126 134194
rect 87190 134130 87198 134194
rect 86878 134129 87198 134130
rect 84415 133852 84481 133855
rect 88454 133852 88934 133882
rect 84415 133850 88934 133852
rect 84415 133794 84420 133850
rect 84476 133794 88934 133850
rect 84415 133792 88934 133794
rect 84415 133789 84481 133792
rect 88454 133762 88934 133792
rect 878 133650 1198 133651
rect 878 133586 886 133650
rect 950 133586 966 133650
rect 1030 133586 1046 133650
rect 1110 133586 1126 133650
rect 1190 133586 1198 133650
rect 878 133585 1198 133586
rect 84878 133650 85198 133651
rect 84878 133586 84886 133650
rect 84950 133586 84966 133650
rect 85030 133586 85046 133650
rect 85110 133586 85126 133650
rect 85190 133586 85198 133650
rect 84878 133585 85198 133586
rect 2878 133106 3198 133107
rect 2878 133042 2886 133106
rect 2950 133042 2966 133106
rect 3030 133042 3046 133106
rect 3110 133042 3126 133106
rect 3190 133042 3198 133106
rect 2878 133041 3198 133042
rect 86878 133106 87198 133107
rect 86878 133042 86886 133106
rect 86950 133042 86966 133106
rect 87030 133042 87046 133106
rect 87110 133042 87126 133106
rect 87190 133042 87198 133106
rect 86878 133041 87198 133042
rect 84323 132900 84389 132903
rect 84323 132898 85352 132900
rect 84323 132842 84328 132898
rect 84384 132842 85352 132898
rect 84323 132840 85352 132842
rect 84323 132837 84389 132840
rect 85292 132628 85352 132840
rect 88454 132628 88934 132658
rect 85292 132568 88934 132628
rect 878 132562 1198 132563
rect 878 132498 886 132562
rect 950 132498 966 132562
rect 1030 132498 1046 132562
rect 1110 132498 1126 132562
rect 1190 132498 1198 132562
rect 878 132497 1198 132498
rect 84878 132562 85198 132563
rect 84878 132498 84886 132562
rect 84950 132498 84966 132562
rect 85030 132498 85046 132562
rect 85110 132498 85126 132562
rect 85190 132498 85198 132562
rect 88454 132538 88934 132568
rect 84878 132497 85198 132498
rect 2878 132018 3198 132019
rect 2878 131954 2886 132018
rect 2950 131954 2966 132018
rect 3030 131954 3046 132018
rect 3110 131954 3126 132018
rect 3190 131954 3198 132018
rect 2878 131953 3198 131954
rect 86878 132018 87198 132019
rect 86878 131954 86886 132018
rect 86950 131954 86966 132018
rect 87030 131954 87046 132018
rect 87110 131954 87126 132018
rect 87190 131954 87198 132018
rect 86878 131953 87198 131954
rect 84231 131812 84297 131815
rect 84231 131810 85352 131812
rect 84231 131754 84236 131810
rect 84292 131754 85352 131810
rect 84231 131752 85352 131754
rect 84231 131749 84297 131752
rect 878 131474 1198 131475
rect 878 131410 886 131474
rect 950 131410 966 131474
rect 1030 131410 1046 131474
rect 1110 131410 1126 131474
rect 1190 131410 1198 131474
rect 878 131409 1198 131410
rect 84878 131474 85198 131475
rect 84878 131410 84886 131474
rect 84950 131410 84966 131474
rect 85030 131410 85046 131474
rect 85110 131410 85126 131474
rect 85190 131410 85198 131474
rect 84878 131409 85198 131410
rect 85292 131404 85352 131752
rect 88454 131404 88934 131434
rect 85292 131344 88934 131404
rect 88454 131314 88934 131344
rect 2878 130930 3198 130931
rect 2878 130866 2886 130930
rect 2950 130866 2966 130930
rect 3030 130866 3046 130930
rect 3110 130866 3126 130930
rect 3190 130866 3198 130930
rect 2878 130865 3198 130866
rect 86878 130930 87198 130931
rect 86878 130866 86886 130930
rect 86950 130866 86966 130930
rect 87030 130866 87046 130930
rect 87110 130866 87126 130930
rect 87190 130866 87198 130930
rect 86878 130865 87198 130866
rect 878 130386 1198 130387
rect 878 130322 886 130386
rect 950 130322 966 130386
rect 1030 130322 1046 130386
rect 1110 130322 1126 130386
rect 1190 130322 1198 130386
rect 878 130321 1198 130322
rect 84878 130386 85198 130387
rect 84878 130322 84886 130386
rect 84950 130322 84966 130386
rect 85030 130322 85046 130386
rect 85110 130322 85126 130386
rect 85190 130322 85198 130386
rect 84878 130321 85198 130322
rect 83587 130180 83653 130183
rect 88454 130180 88934 130210
rect 83587 130178 88934 130180
rect 83587 130122 83592 130178
rect 83648 130122 88934 130178
rect 83587 130120 88934 130122
rect 83587 130117 83653 130120
rect 88454 130090 88934 130120
rect 2878 129842 3198 129843
rect 2878 129778 2886 129842
rect 2950 129778 2966 129842
rect 3030 129778 3046 129842
rect 3110 129778 3126 129842
rect 3190 129778 3198 129842
rect 2878 129777 3198 129778
rect 86878 129842 87198 129843
rect 86878 129778 86886 129842
rect 86950 129778 86966 129842
rect 87030 129778 87046 129842
rect 87110 129778 87126 129842
rect 87190 129778 87198 129842
rect 86878 129777 87198 129778
rect 878 129298 1198 129299
rect 878 129234 886 129298
rect 950 129234 966 129298
rect 1030 129234 1046 129298
rect 1110 129234 1126 129298
rect 1190 129234 1198 129298
rect 878 129233 1198 129234
rect 84878 129298 85198 129299
rect 84878 129234 84886 129298
rect 84950 129234 84966 129298
rect 85030 129234 85046 129298
rect 85110 129234 85126 129298
rect 85190 129234 85198 129298
rect 84878 129233 85198 129234
rect 85887 129092 85953 129095
rect 88454 129092 88934 129122
rect 85887 129090 88934 129092
rect 85887 129034 85892 129090
rect 85948 129034 88934 129090
rect 85887 129032 88934 129034
rect 85887 129029 85953 129032
rect 88454 129002 88934 129032
rect 2878 128754 3198 128755
rect 2878 128690 2886 128754
rect 2950 128690 2966 128754
rect 3030 128690 3046 128754
rect 3110 128690 3126 128754
rect 3190 128690 3198 128754
rect 2878 128689 3198 128690
rect 86878 128754 87198 128755
rect 86878 128690 86886 128754
rect 86950 128690 86966 128754
rect 87030 128690 87046 128754
rect 87110 128690 87126 128754
rect 87190 128690 87198 128754
rect 86878 128689 87198 128690
rect 878 128210 1198 128211
rect 878 128146 886 128210
rect 950 128146 966 128210
rect 1030 128146 1046 128210
rect 1110 128146 1126 128210
rect 1190 128146 1198 128210
rect 878 128145 1198 128146
rect 84878 128210 85198 128211
rect 84878 128146 84886 128210
rect 84950 128146 84966 128210
rect 85030 128146 85046 128210
rect 85110 128146 85126 128210
rect 85190 128146 85198 128210
rect 84878 128145 85198 128146
rect 84507 127868 84573 127871
rect 88454 127868 88934 127898
rect 84507 127866 88934 127868
rect 84507 127810 84512 127866
rect 84568 127810 88934 127866
rect 84507 127808 88934 127810
rect 84507 127805 84573 127808
rect 88454 127778 88934 127808
rect 2878 127666 3198 127667
rect 2878 127602 2886 127666
rect 2950 127602 2966 127666
rect 3030 127602 3046 127666
rect 3110 127602 3126 127666
rect 3190 127602 3198 127666
rect 2878 127601 3198 127602
rect 86878 127666 87198 127667
rect 86878 127602 86886 127666
rect 86950 127602 86966 127666
rect 87030 127602 87046 127666
rect 87110 127602 87126 127666
rect 87190 127602 87198 127666
rect 86878 127601 87198 127602
rect 878 127122 1198 127123
rect 878 127058 886 127122
rect 950 127058 966 127122
rect 1030 127058 1046 127122
rect 1110 127058 1126 127122
rect 1190 127058 1198 127122
rect 878 127057 1198 127058
rect 84878 127122 85198 127123
rect 84878 127058 84886 127122
rect 84950 127058 84966 127122
rect 85030 127058 85046 127122
rect 85110 127058 85126 127122
rect 85190 127058 85198 127122
rect 84878 127057 85198 127058
rect 88454 126644 88934 126674
rect 87500 126584 88934 126644
rect 2878 126578 3198 126579
rect 2878 126514 2886 126578
rect 2950 126514 2966 126578
rect 3030 126514 3046 126578
rect 3110 126514 3126 126578
rect 3190 126514 3198 126578
rect 2878 126513 3198 126514
rect 86878 126578 87198 126579
rect 86878 126514 86886 126578
rect 86950 126514 86966 126578
rect 87030 126514 87046 126578
rect 87110 126514 87126 126578
rect 87190 126514 87198 126578
rect 86878 126513 87198 126514
rect 85979 126372 86045 126375
rect 87500 126372 87560 126584
rect 88454 126554 88934 126584
rect 85979 126370 87560 126372
rect 85979 126314 85984 126370
rect 86040 126314 87560 126370
rect 85979 126312 87560 126314
rect 85979 126309 86045 126312
rect 878 126034 1198 126035
rect 878 125970 886 126034
rect 950 125970 966 126034
rect 1030 125970 1046 126034
rect 1110 125970 1126 126034
rect 1190 125970 1198 126034
rect 878 125969 1198 125970
rect 84878 126034 85198 126035
rect 84878 125970 84886 126034
rect 84950 125970 84966 126034
rect 85030 125970 85046 126034
rect 85110 125970 85126 126034
rect 85190 125970 85198 126034
rect 84878 125969 85198 125970
rect 2878 125490 3198 125491
rect 2878 125426 2886 125490
rect 2950 125426 2966 125490
rect 3030 125426 3046 125490
rect 3110 125426 3126 125490
rect 3190 125426 3198 125490
rect 2878 125425 3198 125426
rect 86878 125490 87198 125491
rect 86878 125426 86886 125490
rect 86950 125426 86966 125490
rect 87030 125426 87046 125490
rect 87110 125426 87126 125490
rect 87190 125426 87198 125490
rect 86878 125425 87198 125426
rect 88454 125420 88934 125450
rect 87500 125360 88934 125420
rect 84231 125284 84297 125287
rect 87500 125284 87560 125360
rect 88454 125330 88934 125360
rect 84231 125282 87560 125284
rect 84231 125226 84236 125282
rect 84292 125226 87560 125282
rect 84231 125224 87560 125226
rect 84231 125221 84297 125224
rect 878 124946 1198 124947
rect 878 124882 886 124946
rect 950 124882 966 124946
rect 1030 124882 1046 124946
rect 1110 124882 1126 124946
rect 1190 124882 1198 124946
rect 878 124881 1198 124882
rect 84878 124946 85198 124947
rect 84878 124882 84886 124946
rect 84950 124882 84966 124946
rect 85030 124882 85046 124946
rect 85110 124882 85126 124946
rect 85190 124882 85198 124946
rect 84878 124881 85198 124882
rect 2167 124740 2233 124743
rect 2300 124740 2306 124742
rect 2167 124738 2306 124740
rect 2167 124682 2172 124738
rect 2228 124682 2306 124738
rect 2167 124680 2306 124682
rect 2167 124677 2233 124680
rect 2300 124678 2306 124680
rect 2370 124678 2376 124742
rect 2878 124402 3198 124403
rect 2878 124338 2886 124402
rect 2950 124338 2966 124402
rect 3030 124338 3046 124402
rect 3110 124338 3126 124402
rect 3190 124338 3198 124402
rect 2878 124337 3198 124338
rect 86878 124402 87198 124403
rect 86878 124338 86886 124402
rect 86950 124338 86966 124402
rect 87030 124338 87046 124402
rect 87110 124338 87126 124402
rect 87190 124338 87198 124402
rect 86878 124337 87198 124338
rect 84415 124196 84481 124199
rect 88454 124196 88934 124226
rect 84415 124194 88934 124196
rect 84415 124138 84420 124194
rect 84476 124138 88934 124194
rect 84415 124136 88934 124138
rect 84415 124133 84481 124136
rect 88454 124106 88934 124136
rect 878 123858 1198 123859
rect 878 123794 886 123858
rect 950 123794 966 123858
rect 1030 123794 1046 123858
rect 1110 123794 1126 123858
rect 1190 123794 1198 123858
rect 878 123793 1198 123794
rect 84878 123858 85198 123859
rect 84878 123794 84886 123858
rect 84950 123794 84966 123858
rect 85030 123794 85046 123858
rect 85110 123794 85126 123858
rect 85190 123794 85198 123858
rect 84878 123793 85198 123794
rect 2878 123314 3198 123315
rect 2878 123250 2886 123314
rect 2950 123250 2966 123314
rect 3030 123250 3046 123314
rect 3110 123250 3126 123314
rect 3190 123250 3198 123314
rect 2878 123249 3198 123250
rect 86878 123314 87198 123315
rect 86878 123250 86886 123314
rect 86950 123250 86966 123314
rect 87030 123250 87046 123314
rect 87110 123250 87126 123314
rect 87190 123250 87198 123314
rect 86878 123249 87198 123250
rect 84415 122972 84481 122975
rect 88454 122972 88934 123002
rect 84415 122970 88934 122972
rect 84415 122914 84420 122970
rect 84476 122914 88934 122970
rect 84415 122912 88934 122914
rect 84415 122909 84481 122912
rect 88454 122882 88934 122912
rect 878 122770 1198 122771
rect 878 122706 886 122770
rect 950 122706 966 122770
rect 1030 122706 1046 122770
rect 1110 122706 1126 122770
rect 1190 122706 1198 122770
rect 878 122705 1198 122706
rect 84878 122770 85198 122771
rect 84878 122706 84886 122770
rect 84950 122706 84966 122770
rect 85030 122706 85046 122770
rect 85110 122706 85126 122770
rect 85190 122706 85198 122770
rect 84878 122705 85198 122706
rect 2878 122226 3198 122227
rect 2878 122162 2886 122226
rect 2950 122162 2966 122226
rect 3030 122162 3046 122226
rect 3110 122162 3126 122226
rect 3190 122162 3198 122226
rect 2878 122161 3198 122162
rect 86878 122226 87198 122227
rect 86878 122162 86886 122226
rect 86950 122162 86966 122226
rect 87030 122162 87046 122226
rect 87110 122162 87126 122226
rect 87190 122162 87198 122226
rect 86878 122161 87198 122162
rect 83955 121884 84021 121887
rect 88454 121884 88934 121914
rect 83955 121882 88934 121884
rect 83955 121826 83960 121882
rect 84016 121826 88934 121882
rect 83955 121824 88934 121826
rect 83955 121821 84021 121824
rect 88454 121794 88934 121824
rect 878 121682 1198 121683
rect 878 121618 886 121682
rect 950 121618 966 121682
rect 1030 121618 1046 121682
rect 1110 121618 1126 121682
rect 1190 121618 1198 121682
rect 878 121617 1198 121618
rect 84878 121682 85198 121683
rect 84878 121618 84886 121682
rect 84950 121618 84966 121682
rect 85030 121618 85046 121682
rect 85110 121618 85126 121682
rect 85190 121618 85198 121682
rect 84878 121617 85198 121618
rect 2878 121138 3198 121139
rect 2878 121074 2886 121138
rect 2950 121074 2966 121138
rect 3030 121074 3046 121138
rect 3110 121074 3126 121138
rect 3190 121074 3198 121138
rect 2878 121073 3198 121074
rect 86878 121138 87198 121139
rect 86878 121074 86886 121138
rect 86950 121074 86966 121138
rect 87030 121074 87046 121138
rect 87110 121074 87126 121138
rect 87190 121074 87198 121138
rect 86878 121073 87198 121074
rect 88454 120660 88934 120690
rect 85292 120600 88934 120660
rect 878 120594 1198 120595
rect 878 120530 886 120594
rect 950 120530 966 120594
rect 1030 120530 1046 120594
rect 1110 120530 1126 120594
rect 1190 120530 1198 120594
rect 878 120529 1198 120530
rect 84878 120594 85198 120595
rect 84878 120530 84886 120594
rect 84950 120530 84966 120594
rect 85030 120530 85046 120594
rect 85110 120530 85126 120594
rect 85190 120530 85198 120594
rect 84878 120529 85198 120530
rect 84231 120252 84297 120255
rect 85292 120252 85352 120600
rect 88454 120570 88934 120600
rect 84231 120250 85352 120252
rect 84231 120194 84236 120250
rect 84292 120194 85352 120250
rect 84231 120192 85352 120194
rect 84231 120189 84297 120192
rect 2878 120050 3198 120051
rect 2878 119986 2886 120050
rect 2950 119986 2966 120050
rect 3030 119986 3046 120050
rect 3110 119986 3126 120050
rect 3190 119986 3198 120050
rect 2878 119985 3198 119986
rect 86878 120050 87198 120051
rect 86878 119986 86886 120050
rect 86950 119986 86966 120050
rect 87030 119986 87046 120050
rect 87110 119986 87126 120050
rect 87190 119986 87198 120050
rect 86878 119985 87198 119986
rect 878 119506 1198 119507
rect 878 119442 886 119506
rect 950 119442 966 119506
rect 1030 119442 1046 119506
rect 1110 119442 1126 119506
rect 1190 119442 1198 119506
rect 878 119441 1198 119442
rect 84878 119506 85198 119507
rect 84878 119442 84886 119506
rect 84950 119442 84966 119506
rect 85030 119442 85046 119506
rect 85110 119442 85126 119506
rect 85190 119442 85198 119506
rect 84878 119441 85198 119442
rect 85335 119436 85401 119439
rect 88454 119436 88934 119466
rect 85335 119434 88934 119436
rect 85335 119378 85340 119434
rect 85396 119378 88934 119434
rect 85335 119376 88934 119378
rect 85335 119373 85401 119376
rect 88454 119346 88934 119376
rect 2878 118962 3198 118963
rect 2878 118898 2886 118962
rect 2950 118898 2966 118962
rect 3030 118898 3046 118962
rect 3110 118898 3126 118962
rect 3190 118898 3198 118962
rect 2878 118897 3198 118898
rect 86878 118962 87198 118963
rect 86878 118898 86886 118962
rect 86950 118898 86966 118962
rect 87030 118898 87046 118962
rect 87110 118898 87126 118962
rect 87190 118898 87198 118962
rect 86878 118897 87198 118898
rect 878 118418 1198 118419
rect 878 118354 886 118418
rect 950 118354 966 118418
rect 1030 118354 1046 118418
rect 1110 118354 1126 118418
rect 1190 118354 1198 118418
rect 878 118353 1198 118354
rect 84878 118418 85198 118419
rect 84878 118354 84886 118418
rect 84950 118354 84966 118418
rect 85030 118354 85046 118418
rect 85110 118354 85126 118418
rect 85190 118354 85198 118418
rect 84878 118353 85198 118354
rect 84323 118212 84389 118215
rect 88454 118212 88934 118242
rect 84323 118210 88934 118212
rect 84323 118154 84328 118210
rect 84384 118154 88934 118210
rect 84323 118152 88934 118154
rect 84323 118149 84389 118152
rect 88454 118122 88934 118152
rect 2878 117874 3198 117875
rect 2878 117810 2886 117874
rect 2950 117810 2966 117874
rect 3030 117810 3046 117874
rect 3110 117810 3126 117874
rect 3190 117810 3198 117874
rect 2878 117809 3198 117810
rect 86878 117874 87198 117875
rect 86878 117810 86886 117874
rect 86950 117810 86966 117874
rect 87030 117810 87046 117874
rect 87110 117810 87126 117874
rect 87190 117810 87198 117874
rect 86878 117809 87198 117810
rect 878 117330 1198 117331
rect 878 117266 886 117330
rect 950 117266 966 117330
rect 1030 117266 1046 117330
rect 1110 117266 1126 117330
rect 1190 117266 1198 117330
rect 878 117265 1198 117266
rect 84878 117330 85198 117331
rect 84878 117266 84886 117330
rect 84950 117266 84966 117330
rect 85030 117266 85046 117330
rect 85110 117266 85126 117330
rect 85190 117266 85198 117330
rect 84878 117265 85198 117266
rect 84231 116988 84297 116991
rect 88454 116988 88934 117018
rect 84231 116986 88934 116988
rect 84231 116930 84236 116986
rect 84292 116930 88934 116986
rect 84231 116928 88934 116930
rect 84231 116925 84297 116928
rect 88454 116898 88934 116928
rect 2878 116786 3198 116787
rect 2878 116722 2886 116786
rect 2950 116722 2966 116786
rect 3030 116722 3046 116786
rect 3110 116722 3126 116786
rect 3190 116722 3198 116786
rect 2878 116721 3198 116722
rect 86878 116786 87198 116787
rect 86878 116722 86886 116786
rect 86950 116722 86966 116786
rect 87030 116722 87046 116786
rect 87110 116722 87126 116786
rect 87190 116722 87198 116786
rect 86878 116721 87198 116722
rect 4283 116444 4349 116447
rect 5068 116444 5128 116457
rect 4283 116442 5128 116444
rect 4283 116386 4288 116442
rect 4344 116386 5128 116442
rect 4283 116384 5128 116386
rect 4283 116381 4349 116384
rect 878 116242 1198 116243
rect 878 116178 886 116242
rect 950 116178 966 116242
rect 1030 116178 1046 116242
rect 1110 116178 1126 116242
rect 1190 116178 1198 116242
rect 878 116177 1198 116178
rect 84878 116242 85198 116243
rect 84878 116178 84886 116242
rect 84950 116178 84966 116242
rect 85030 116178 85046 116242
rect 85110 116178 85126 116242
rect 85190 116178 85198 116242
rect 84878 116177 85198 116178
rect 83955 115900 84021 115903
rect 83955 115898 87560 115900
rect 83955 115842 83960 115898
rect 84016 115842 87560 115898
rect 83955 115840 87560 115842
rect 83955 115837 84021 115840
rect 87500 115764 87560 115840
rect 88454 115764 88934 115794
rect 87500 115704 88934 115764
rect 2878 115698 3198 115699
rect 2878 115634 2886 115698
rect 2950 115634 2966 115698
rect 3030 115634 3046 115698
rect 3110 115634 3126 115698
rect 3190 115634 3198 115698
rect 2878 115633 3198 115634
rect 86878 115698 87198 115699
rect 86878 115634 86886 115698
rect 86950 115634 86966 115698
rect 87030 115634 87046 115698
rect 87110 115634 87126 115698
rect 87190 115634 87198 115698
rect 88454 115674 88934 115704
rect 86878 115633 87198 115634
rect 878 115154 1198 115155
rect 878 115090 886 115154
rect 950 115090 966 115154
rect 1030 115090 1046 115154
rect 1110 115090 1126 115154
rect 1190 115090 1198 115154
rect 878 115089 1198 115090
rect 84878 115154 85198 115155
rect 84878 115090 84886 115154
rect 84950 115090 84966 115154
rect 85030 115090 85046 115154
rect 85110 115090 85126 115154
rect 85190 115090 85198 115154
rect 84878 115089 85198 115090
rect 3455 114812 3521 114815
rect 84323 114812 84389 114815
rect 3455 114810 5128 114812
rect 3455 114754 3460 114810
rect 3516 114754 5128 114810
rect 3455 114752 5128 114754
rect 84323 114810 87560 114812
rect 84323 114754 84328 114810
rect 84384 114754 87560 114810
rect 84323 114752 87560 114754
rect 3455 114749 3521 114752
rect 84323 114749 84389 114752
rect 2878 114610 3198 114611
rect 2878 114546 2886 114610
rect 2950 114546 2966 114610
rect 3030 114546 3046 114610
rect 3110 114546 3126 114610
rect 3190 114546 3198 114610
rect 2878 114545 3198 114546
rect 86878 114610 87198 114611
rect 86878 114546 86886 114610
rect 86950 114546 86966 114610
rect 87030 114546 87046 114610
rect 87110 114546 87126 114610
rect 87190 114546 87198 114610
rect 86878 114545 87198 114546
rect 87500 114540 87560 114752
rect 88454 114540 88934 114570
rect 87500 114480 88934 114540
rect 88454 114450 88934 114480
rect 878 114066 1198 114067
rect 878 114002 886 114066
rect 950 114002 966 114066
rect 1030 114002 1046 114066
rect 1110 114002 1126 114066
rect 1190 114002 1198 114066
rect 878 114001 1198 114002
rect 84878 114066 85198 114067
rect 84878 114002 84886 114066
rect 84950 114002 84966 114066
rect 85030 114002 85046 114066
rect 85110 114002 85126 114066
rect 85190 114002 85198 114066
rect 84878 114001 85198 114002
rect 2878 113522 3198 113523
rect 2878 113458 2886 113522
rect 2950 113458 2966 113522
rect 3030 113458 3046 113522
rect 3110 113458 3126 113522
rect 3190 113458 3198 113522
rect 2878 113457 3198 113458
rect 86878 113522 87198 113523
rect 86878 113458 86886 113522
rect 86950 113458 86966 113522
rect 87030 113458 87046 113522
rect 87110 113458 87126 113522
rect 87190 113458 87198 113522
rect 86878 113457 87198 113458
rect 88454 113452 88934 113482
rect 87500 113392 88934 113452
rect 84323 113316 84389 113319
rect 87500 113316 87560 113392
rect 88454 113362 88934 113392
rect 84323 113314 87560 113316
rect 84323 113258 84328 113314
rect 84384 113258 87560 113314
rect 84323 113256 87560 113258
rect 84323 113253 84389 113256
rect 878 112978 1198 112979
rect 878 112914 886 112978
rect 950 112914 966 112978
rect 1030 112914 1046 112978
rect 1110 112914 1126 112978
rect 1190 112914 1198 112978
rect 878 112913 1198 112914
rect 84878 112978 85198 112979
rect 84878 112914 84886 112978
rect 84950 112914 84966 112978
rect 85030 112914 85046 112978
rect 85110 112914 85126 112978
rect 85190 112914 85198 112978
rect 84878 112913 85198 112914
rect 2878 112434 3198 112435
rect 2878 112370 2886 112434
rect 2950 112370 2966 112434
rect 3030 112370 3046 112434
rect 3110 112370 3126 112434
rect 3190 112370 3198 112434
rect 2878 112369 3198 112370
rect 86878 112434 87198 112435
rect 86878 112370 86886 112434
rect 86950 112370 86966 112434
rect 87030 112370 87046 112434
rect 87110 112370 87126 112434
rect 87190 112370 87198 112434
rect 86878 112369 87198 112370
rect 84875 112228 84941 112231
rect 88454 112228 88934 112258
rect 84875 112226 88934 112228
rect 84875 112170 84880 112226
rect 84936 112170 88934 112226
rect 84875 112168 88934 112170
rect 84875 112165 84941 112168
rect 88454 112138 88934 112168
rect 878 111890 1198 111891
rect 878 111826 886 111890
rect 950 111826 966 111890
rect 1030 111826 1046 111890
rect 1110 111826 1126 111890
rect 1190 111826 1198 111890
rect 878 111825 1198 111826
rect 84878 111890 85198 111891
rect 84878 111826 84886 111890
rect 84950 111826 84966 111890
rect 85030 111826 85046 111890
rect 85110 111826 85126 111890
rect 85190 111826 85198 111890
rect 84878 111825 85198 111826
rect 2878 111346 3198 111347
rect 2878 111282 2886 111346
rect 2950 111282 2966 111346
rect 3030 111282 3046 111346
rect 3110 111282 3126 111346
rect 3190 111282 3198 111346
rect 2878 111281 3198 111282
rect 86878 111346 87198 111347
rect 86878 111282 86886 111346
rect 86950 111282 86966 111346
rect 87030 111282 87046 111346
rect 87110 111282 87126 111346
rect 87190 111282 87198 111346
rect 86878 111281 87198 111282
rect 86071 111004 86137 111007
rect 88454 111004 88934 111034
rect 86071 111002 88934 111004
rect 86071 110946 86076 111002
rect 86132 110946 88934 111002
rect 86071 110944 88934 110946
rect 86071 110941 86137 110944
rect 88454 110914 88934 110944
rect 878 110802 1198 110803
rect 878 110738 886 110802
rect 950 110738 966 110802
rect 1030 110738 1046 110802
rect 1110 110738 1126 110802
rect 1190 110738 1198 110802
rect 878 110737 1198 110738
rect 84878 110802 85198 110803
rect 84878 110738 84886 110802
rect 84950 110738 84966 110802
rect 85030 110738 85046 110802
rect 85110 110738 85126 110802
rect 85190 110738 85198 110802
rect 84878 110737 85198 110738
rect 2878 110258 3198 110259
rect 2878 110194 2886 110258
rect 2950 110194 2966 110258
rect 3030 110194 3046 110258
rect 3110 110194 3126 110258
rect 3190 110194 3198 110258
rect 2878 110193 3198 110194
rect 86878 110258 87198 110259
rect 86878 110194 86886 110258
rect 86950 110194 86966 110258
rect 87030 110194 87046 110258
rect 87110 110194 87126 110258
rect 87190 110194 87198 110258
rect 86878 110193 87198 110194
rect 88454 109780 88934 109810
rect 85292 109720 88934 109780
rect 878 109714 1198 109715
rect 878 109650 886 109714
rect 950 109650 966 109714
rect 1030 109650 1046 109714
rect 1110 109650 1126 109714
rect 1190 109650 1198 109714
rect 878 109649 1198 109650
rect 84878 109714 85198 109715
rect 84878 109650 84886 109714
rect 84950 109650 84966 109714
rect 85030 109650 85046 109714
rect 85110 109650 85126 109714
rect 85190 109650 85198 109714
rect 84878 109649 85198 109650
rect 83955 109372 84021 109375
rect 85292 109372 85352 109720
rect 88454 109690 88934 109720
rect 83955 109370 85352 109372
rect 83955 109314 83960 109370
rect 84016 109314 85352 109370
rect 83955 109312 85352 109314
rect 83955 109309 84021 109312
rect 2878 109170 3198 109171
rect 2878 109106 2886 109170
rect 2950 109106 2966 109170
rect 3030 109106 3046 109170
rect 3110 109106 3126 109170
rect 3190 109106 3198 109170
rect 2878 109105 3198 109106
rect 86878 109170 87198 109171
rect 86878 109106 86886 109170
rect 86950 109106 86966 109170
rect 87030 109106 87046 109170
rect 87110 109106 87126 109170
rect 87190 109106 87198 109170
rect 86878 109105 87198 109106
rect 878 108626 1198 108627
rect 878 108562 886 108626
rect 950 108562 966 108626
rect 1030 108562 1046 108626
rect 1110 108562 1126 108626
rect 1190 108562 1198 108626
rect 878 108561 1198 108562
rect 84878 108626 85198 108627
rect 84878 108562 84886 108626
rect 84950 108562 84966 108626
rect 85030 108562 85046 108626
rect 85110 108562 85126 108626
rect 85190 108562 85198 108626
rect 84878 108561 85198 108562
rect 88454 108556 88934 108586
rect 85292 108496 88934 108556
rect 83955 108284 84021 108287
rect 85292 108284 85352 108496
rect 88454 108466 88934 108496
rect 83955 108282 85352 108284
rect 83955 108226 83960 108282
rect 84016 108226 85352 108282
rect 83955 108224 85352 108226
rect 83955 108221 84021 108224
rect 2167 108148 2233 108151
rect 2300 108148 2306 108150
rect 2167 108146 2306 108148
rect 2167 108090 2172 108146
rect 2228 108090 2306 108146
rect 2167 108088 2306 108090
rect 2167 108085 2233 108088
rect 2300 108086 2306 108088
rect 2370 108086 2376 108150
rect 2878 108082 3198 108083
rect 2878 108018 2886 108082
rect 2950 108018 2966 108082
rect 3030 108018 3046 108082
rect 3110 108018 3126 108082
rect 3190 108018 3198 108082
rect 2878 108017 3198 108018
rect 86878 108082 87198 108083
rect 86878 108018 86886 108082
rect 86950 108018 86966 108082
rect 87030 108018 87046 108082
rect 87110 108018 87126 108082
rect 87190 108018 87198 108082
rect 86878 108017 87198 108018
rect 878 107538 1198 107539
rect 878 107474 886 107538
rect 950 107474 966 107538
rect 1030 107474 1046 107538
rect 1110 107474 1126 107538
rect 1190 107474 1198 107538
rect 878 107473 1198 107474
rect 84878 107538 85198 107539
rect 84878 107474 84886 107538
rect 84950 107474 84966 107538
rect 85030 107474 85046 107538
rect 85110 107474 85126 107538
rect 85190 107474 85198 107538
rect 84878 107473 85198 107474
rect 83955 107332 84021 107335
rect 88454 107332 88934 107362
rect 83955 107330 88934 107332
rect 83955 107274 83960 107330
rect 84016 107274 88934 107330
rect 83955 107272 88934 107274
rect 83955 107269 84021 107272
rect 88454 107242 88934 107272
rect 2878 106994 3198 106995
rect 2878 106930 2886 106994
rect 2950 106930 2966 106994
rect 3030 106930 3046 106994
rect 3110 106930 3126 106994
rect 3190 106930 3198 106994
rect 2878 106929 3198 106930
rect 86878 106994 87198 106995
rect 86878 106930 86886 106994
rect 86950 106930 86966 106994
rect 87030 106930 87046 106994
rect 87110 106930 87126 106994
rect 87190 106930 87198 106994
rect 86878 106929 87198 106930
rect 878 106450 1198 106451
rect 878 106386 886 106450
rect 950 106386 966 106450
rect 1030 106386 1046 106450
rect 1110 106386 1126 106450
rect 1190 106386 1198 106450
rect 878 106385 1198 106386
rect 84878 106450 85198 106451
rect 84878 106386 84886 106450
rect 84950 106386 84966 106450
rect 85030 106386 85046 106450
rect 85110 106386 85126 106450
rect 85190 106386 85198 106450
rect 84878 106385 85198 106386
rect 84231 106244 84297 106247
rect 88454 106244 88934 106274
rect 84231 106242 88934 106244
rect 84231 106186 84236 106242
rect 84292 106186 88934 106242
rect 84231 106184 88934 106186
rect 84231 106181 84297 106184
rect 88454 106154 88934 106184
rect 2878 105906 3198 105907
rect 2878 105842 2886 105906
rect 2950 105842 2966 105906
rect 3030 105842 3046 105906
rect 3110 105842 3126 105906
rect 3190 105842 3198 105906
rect 2878 105841 3198 105842
rect 86878 105906 87198 105907
rect 86878 105842 86886 105906
rect 86950 105842 86966 105906
rect 87030 105842 87046 105906
rect 87110 105842 87126 105906
rect 87190 105842 87198 105906
rect 86878 105841 87198 105842
rect 878 105362 1198 105363
rect 878 105298 886 105362
rect 950 105298 966 105362
rect 1030 105298 1046 105362
rect 1110 105298 1126 105362
rect 1190 105298 1198 105362
rect 878 105297 1198 105298
rect 84878 105362 85198 105363
rect 84878 105298 84886 105362
rect 84950 105298 84966 105362
rect 85030 105298 85046 105362
rect 85110 105298 85126 105362
rect 85190 105298 85198 105362
rect 84878 105297 85198 105298
rect 86163 105020 86229 105023
rect 88454 105020 88934 105050
rect 86163 105018 88934 105020
rect 86163 104962 86168 105018
rect 86224 104962 88934 105018
rect 86163 104960 88934 104962
rect 86163 104957 86229 104960
rect 88454 104930 88934 104960
rect 2878 104818 3198 104819
rect 2878 104754 2886 104818
rect 2950 104754 2966 104818
rect 3030 104754 3046 104818
rect 3110 104754 3126 104818
rect 3190 104754 3198 104818
rect 2878 104753 3198 104754
rect 86878 104818 87198 104819
rect 86878 104754 86886 104818
rect 86950 104754 86966 104818
rect 87030 104754 87046 104818
rect 87110 104754 87126 104818
rect 87190 104754 87198 104818
rect 86878 104753 87198 104754
rect 878 104274 1198 104275
rect 878 104210 886 104274
rect 950 104210 966 104274
rect 1030 104210 1046 104274
rect 1110 104210 1126 104274
rect 1190 104210 1198 104274
rect 878 104209 1198 104210
rect 84878 104274 85198 104275
rect 84878 104210 84886 104274
rect 84950 104210 84966 104274
rect 85030 104210 85046 104274
rect 85110 104210 85126 104274
rect 85190 104210 85198 104274
rect 84878 104209 85198 104210
rect 88454 103796 88934 103826
rect 87500 103736 88934 103796
rect 2878 103730 3198 103731
rect 2878 103666 2886 103730
rect 2950 103666 2966 103730
rect 3030 103666 3046 103730
rect 3110 103666 3126 103730
rect 3190 103666 3198 103730
rect 2878 103665 3198 103666
rect 86878 103730 87198 103731
rect 86878 103666 86886 103730
rect 86950 103666 86966 103730
rect 87030 103666 87046 103730
rect 87110 103666 87126 103730
rect 87190 103666 87198 103730
rect 86878 103665 87198 103666
rect 86255 103524 86321 103527
rect 87500 103524 87560 103736
rect 88454 103706 88934 103736
rect 86255 103522 87560 103524
rect 86255 103466 86260 103522
rect 86316 103466 87560 103522
rect 86255 103464 87560 103466
rect 86255 103461 86321 103464
rect 878 103186 1198 103187
rect 878 103122 886 103186
rect 950 103122 966 103186
rect 1030 103122 1046 103186
rect 1110 103122 1126 103186
rect 1190 103122 1198 103186
rect 878 103121 1198 103122
rect 84878 103186 85198 103187
rect 84878 103122 84886 103186
rect 84950 103122 84966 103186
rect 85030 103122 85046 103186
rect 85110 103122 85126 103186
rect 85190 103122 85198 103186
rect 84878 103121 85198 103122
rect 2878 102642 3198 102643
rect 2878 102578 2886 102642
rect 2950 102578 2966 102642
rect 3030 102578 3046 102642
rect 3110 102578 3126 102642
rect 3190 102578 3198 102642
rect 2878 102577 3198 102578
rect 86878 102642 87198 102643
rect 86878 102578 86886 102642
rect 86950 102578 86966 102642
rect 87030 102578 87046 102642
rect 87110 102578 87126 102642
rect 87190 102578 87198 102642
rect 86878 102577 87198 102578
rect 88454 102572 88934 102602
rect 87500 102512 88934 102572
rect 84139 102436 84205 102439
rect 87500 102436 87560 102512
rect 88454 102482 88934 102512
rect 84139 102434 87560 102436
rect 84139 102378 84144 102434
rect 84200 102378 87560 102434
rect 84139 102376 87560 102378
rect 84139 102373 84205 102376
rect 878 102098 1198 102099
rect 878 102034 886 102098
rect 950 102034 966 102098
rect 1030 102034 1046 102098
rect 1110 102034 1126 102098
rect 1190 102034 1198 102098
rect 878 102033 1198 102034
rect 84878 102098 85198 102099
rect 84878 102034 84886 102098
rect 84950 102034 84966 102098
rect 85030 102034 85046 102098
rect 85110 102034 85126 102098
rect 85190 102034 85198 102098
rect 84878 102033 85198 102034
rect 2878 101554 3198 101555
rect 2878 101490 2886 101554
rect 2950 101490 2966 101554
rect 3030 101490 3046 101554
rect 3110 101490 3126 101554
rect 3190 101490 3198 101554
rect 2878 101489 3198 101490
rect 86878 101554 87198 101555
rect 86878 101490 86886 101554
rect 86950 101490 86966 101554
rect 87030 101490 87046 101554
rect 87110 101490 87126 101554
rect 87190 101490 87198 101554
rect 86878 101489 87198 101490
rect 85703 101348 85769 101351
rect 88454 101348 88934 101378
rect 85703 101346 88934 101348
rect 85703 101290 85708 101346
rect 85764 101290 88934 101346
rect 85703 101288 88934 101290
rect 85703 101285 85769 101288
rect 88454 101258 88934 101288
rect 878 101010 1198 101011
rect 878 100946 886 101010
rect 950 100946 966 101010
rect 1030 100946 1046 101010
rect 1110 100946 1126 101010
rect 1190 100946 1198 101010
rect 878 100945 1198 100946
rect 84878 101010 85198 101011
rect 84878 100946 84886 101010
rect 84950 100946 84966 101010
rect 85030 100946 85046 101010
rect 85110 100946 85126 101010
rect 85190 100946 85198 101010
rect 84878 100945 85198 100946
rect 2878 100466 3198 100467
rect 2878 100402 2886 100466
rect 2950 100402 2966 100466
rect 3030 100402 3046 100466
rect 3110 100402 3126 100466
rect 3190 100402 3198 100466
rect 2878 100401 3198 100402
rect 86878 100466 87198 100467
rect 86878 100402 86886 100466
rect 86950 100402 86966 100466
rect 87030 100402 87046 100466
rect 87110 100402 87126 100466
rect 87190 100402 87198 100466
rect 86878 100401 87198 100402
rect 84691 100124 84757 100127
rect 88454 100124 88934 100154
rect 84691 100122 88934 100124
rect 84691 100066 84696 100122
rect 84752 100066 88934 100122
rect 84691 100064 88934 100066
rect 84691 100061 84757 100064
rect 88454 100034 88934 100064
rect 878 99922 1198 99923
rect 878 99858 886 99922
rect 950 99858 966 99922
rect 1030 99858 1046 99922
rect 1110 99858 1126 99922
rect 1190 99858 1198 99922
rect 878 99857 1198 99858
rect 84878 99922 85198 99923
rect 84878 99858 84886 99922
rect 84950 99858 84966 99922
rect 85030 99858 85046 99922
rect 85110 99858 85126 99922
rect 85190 99858 85198 99922
rect 84878 99857 85198 99858
rect 2878 99378 3198 99379
rect 2878 99314 2886 99378
rect 2950 99314 2966 99378
rect 3030 99314 3046 99378
rect 3110 99314 3126 99378
rect 3190 99314 3198 99378
rect 2878 99313 3198 99314
rect 86878 99378 87198 99379
rect 86878 99314 86886 99378
rect 86950 99314 86966 99378
rect 87030 99314 87046 99378
rect 87110 99314 87126 99378
rect 87190 99314 87198 99378
rect 86878 99313 87198 99314
rect 84599 99036 84665 99039
rect 88454 99036 88934 99066
rect 84599 99034 88934 99036
rect 84599 98978 84604 99034
rect 84660 98978 88934 99034
rect 84599 98976 88934 98978
rect 84599 98973 84665 98976
rect 88454 98946 88934 98976
rect 878 98834 1198 98835
rect 878 98770 886 98834
rect 950 98770 966 98834
rect 1030 98770 1046 98834
rect 1110 98770 1126 98834
rect 1190 98770 1198 98834
rect 878 98769 1198 98770
rect 84878 98834 85198 98835
rect 84878 98770 84886 98834
rect 84950 98770 84966 98834
rect 85030 98770 85046 98834
rect 85110 98770 85126 98834
rect 85190 98770 85198 98834
rect 84878 98769 85198 98770
rect 4099 98356 4165 98359
rect 4324 98356 4330 98358
rect 4099 98354 4330 98356
rect 4099 98298 4104 98354
rect 4160 98298 4330 98354
rect 4099 98296 4330 98298
rect 4099 98293 4165 98296
rect 4324 98294 4330 98296
rect 4394 98356 4400 98358
rect 4467 98356 4533 98359
rect 4394 98354 4533 98356
rect 4394 98298 4472 98354
rect 4528 98298 4533 98354
rect 4394 98296 4533 98298
rect 4394 98294 4400 98296
rect 4467 98293 4533 98296
rect 2878 98290 3198 98291
rect 2878 98226 2886 98290
rect 2950 98226 2966 98290
rect 3030 98226 3046 98290
rect 3110 98226 3126 98290
rect 3190 98226 3198 98290
rect 2878 98225 3198 98226
rect 86878 98290 87198 98291
rect 86878 98226 86886 98290
rect 86950 98226 86966 98290
rect 87030 98226 87046 98290
rect 87110 98226 87126 98290
rect 87190 98226 87198 98290
rect 86878 98225 87198 98226
rect 3772 98158 3778 98222
rect 3842 98220 3848 98222
rect 4099 98220 4165 98223
rect 3842 98218 4165 98220
rect 3842 98162 4104 98218
rect 4160 98162 4165 98218
rect 3842 98160 4165 98162
rect 3842 98158 3848 98160
rect 4099 98157 4165 98160
rect 84323 97948 84389 97951
rect 84323 97946 85352 97948
rect 84323 97890 84328 97946
rect 84384 97890 85352 97946
rect 84323 97888 85352 97890
rect 84323 97885 84389 97888
rect 85292 97812 85352 97888
rect 88454 97812 88934 97842
rect 85292 97752 88934 97812
rect 878 97746 1198 97747
rect 878 97682 886 97746
rect 950 97682 966 97746
rect 1030 97682 1046 97746
rect 1110 97682 1126 97746
rect 1190 97682 1198 97746
rect 878 97681 1198 97682
rect 84878 97746 85198 97747
rect 84878 97682 84886 97746
rect 84950 97682 84966 97746
rect 85030 97682 85046 97746
rect 85110 97682 85126 97746
rect 85190 97682 85198 97746
rect 88454 97722 88934 97752
rect 84878 97681 85198 97682
rect 83628 97614 83634 97678
rect 83698 97676 83704 97678
rect 83771 97676 83837 97679
rect 83698 97674 83837 97676
rect 83698 97618 83776 97674
rect 83832 97618 83837 97674
rect 83698 97616 83837 97618
rect 83698 97614 83704 97616
rect 83771 97613 83837 97616
rect 2878 97202 3198 97203
rect 2878 97138 2886 97202
rect 2950 97138 2966 97202
rect 3030 97138 3046 97202
rect 3110 97138 3126 97202
rect 3190 97138 3198 97202
rect 2878 97137 3198 97138
rect 86878 97202 87198 97203
rect 86878 97138 86886 97202
rect 86950 97138 86966 97202
rect 87030 97138 87046 97202
rect 87110 97138 87126 97202
rect 87190 97138 87198 97202
rect 86878 97137 87198 97138
rect 83771 97132 83837 97135
rect 84139 97134 84205 97135
rect 84139 97132 84186 97134
rect 45364 97130 83837 97132
rect 45364 97074 83776 97130
rect 83832 97074 83837 97130
rect 45364 97072 83837 97074
rect 84094 97130 84186 97132
rect 84094 97074 84144 97130
rect 84094 97072 84186 97074
rect 2535 96996 2601 96999
rect 39100 96996 39106 96998
rect 2535 96994 39106 96996
rect 2535 96938 2540 96994
rect 2596 96938 39106 96994
rect 2535 96936 39106 96938
rect 2535 96933 2601 96936
rect 39100 96934 39106 96936
rect 39170 96934 39176 96998
rect 14587 96862 14653 96863
rect 14587 96860 14634 96862
rect 14542 96858 14634 96860
rect 14542 96802 14592 96858
rect 14542 96800 14634 96802
rect 14587 96798 14634 96800
rect 14698 96798 14704 96862
rect 28479 96860 28545 96863
rect 45364 96862 45424 97072
rect 83771 97069 83837 97072
rect 84139 97070 84186 97072
rect 84250 97070 84256 97134
rect 84139 97069 84205 97070
rect 48719 96996 48785 96999
rect 55527 96996 55593 96999
rect 48719 96994 55593 96996
rect 48719 96938 48724 96994
rect 48780 96938 55532 96994
rect 55588 96938 55593 96994
rect 48719 96936 55593 96938
rect 48719 96933 48785 96936
rect 55527 96933 55593 96936
rect 77975 96996 78041 96999
rect 82340 96996 82346 96998
rect 77975 96994 82346 96996
rect 77975 96938 77980 96994
rect 78036 96938 82346 96994
rect 77975 96936 82346 96938
rect 77975 96933 78041 96936
rect 82340 96934 82346 96936
rect 82410 96934 82416 96998
rect 33396 96860 33402 96862
rect 28479 96858 33402 96860
rect 28479 96802 28484 96858
rect 28540 96802 33402 96858
rect 28479 96800 33402 96802
rect 14587 96797 14653 96798
rect 28479 96797 28545 96800
rect 33396 96798 33402 96800
rect 33466 96798 33472 96862
rect 45356 96798 45362 96862
rect 45426 96798 45432 96862
rect 46603 96860 46669 96863
rect 51019 96860 51085 96863
rect 83495 96862 83561 96863
rect 83444 96860 83450 96862
rect 46603 96858 50464 96860
rect 46603 96802 46608 96858
rect 46664 96802 50464 96858
rect 46603 96800 50464 96802
rect 46603 96797 46669 96800
rect 2995 96724 3061 96727
rect 3404 96724 3410 96726
rect 2995 96722 3410 96724
rect 2995 96666 3000 96722
rect 3056 96666 3410 96722
rect 2995 96664 3410 96666
rect 2995 96661 3061 96664
rect 3404 96662 3410 96664
rect 3474 96662 3480 96726
rect 5203 96724 5269 96727
rect 15732 96724 15738 96726
rect 5203 96722 15738 96724
rect 5203 96666 5208 96722
rect 5264 96666 15738 96722
rect 5203 96664 15738 96666
rect 5203 96661 5269 96664
rect 15732 96662 15738 96664
rect 15802 96662 15808 96726
rect 21988 96662 21994 96726
rect 22058 96724 22064 96726
rect 22131 96724 22197 96727
rect 25259 96726 25325 96727
rect 28939 96726 29005 96727
rect 29951 96726 30017 96727
rect 35011 96726 35077 96727
rect 25259 96724 25306 96726
rect 22058 96722 22197 96724
rect 22058 96666 22136 96722
rect 22192 96666 22197 96722
rect 22058 96664 22197 96666
rect 25214 96722 25306 96724
rect 25214 96666 25264 96722
rect 25214 96664 25306 96666
rect 22058 96662 22064 96664
rect 22131 96661 22197 96664
rect 25259 96662 25306 96664
rect 25370 96662 25376 96726
rect 28939 96724 28986 96726
rect 28894 96722 28986 96724
rect 28894 96666 28944 96722
rect 28894 96664 28986 96666
rect 28939 96662 28986 96664
rect 29050 96662 29056 96726
rect 29951 96724 29977 96726
rect 29885 96722 29977 96724
rect 29885 96666 29956 96722
rect 29885 96664 29977 96666
rect 29951 96662 29977 96664
rect 30041 96662 30047 96726
rect 34963 96662 34969 96726
rect 35033 96724 35077 96726
rect 36851 96726 36917 96727
rect 36851 96724 36898 96726
rect 35033 96722 35125 96724
rect 35072 96666 35125 96722
rect 35033 96664 35125 96666
rect 36806 96722 36898 96724
rect 36806 96666 36856 96722
rect 36806 96664 36898 96666
rect 35033 96662 35077 96664
rect 25259 96661 25325 96662
rect 28939 96661 29005 96662
rect 29951 96661 30017 96662
rect 35011 96661 35077 96662
rect 36851 96662 36898 96664
rect 36962 96662 36968 96726
rect 37035 96724 37101 96727
rect 37035 96722 42112 96724
rect 37035 96666 37040 96722
rect 37096 96666 42112 96722
rect 37035 96664 42112 96666
rect 36851 96661 36917 96662
rect 37035 96661 37101 96664
rect 878 96658 1198 96659
rect 878 96594 886 96658
rect 950 96594 966 96658
rect 1030 96594 1046 96658
rect 1110 96594 1126 96658
rect 1190 96594 1198 96658
rect 878 96593 1198 96594
rect 5244 96588 5250 96590
rect 4516 96528 5250 96588
rect 4099 96452 4165 96455
rect 4516 96454 4576 96528
rect 5244 96526 5250 96528
rect 5314 96588 5320 96590
rect 15691 96588 15757 96591
rect 5314 96586 15757 96588
rect 5314 96530 15696 96586
rect 15752 96530 15757 96586
rect 5314 96528 15757 96530
rect 5314 96526 5320 96528
rect 15691 96525 15757 96528
rect 24707 96588 24773 96591
rect 42052 96588 42112 96664
rect 44252 96662 44258 96726
rect 44322 96724 44328 96726
rect 48719 96724 48785 96727
rect 48903 96726 48969 96727
rect 50191 96726 50257 96727
rect 44322 96722 48785 96724
rect 44322 96666 48724 96722
rect 48780 96666 48785 96722
rect 44322 96664 48785 96666
rect 44322 96662 44328 96664
rect 48719 96661 48785 96664
rect 48852 96662 48858 96726
rect 48922 96724 48969 96726
rect 48922 96722 49014 96724
rect 48964 96666 49014 96722
rect 48922 96664 49014 96666
rect 48922 96662 48969 96664
rect 50140 96662 50146 96726
rect 50210 96724 50257 96726
rect 50404 96724 50464 96800
rect 51019 96858 83450 96860
rect 83514 96860 83561 96862
rect 83771 96860 83837 96863
rect 83514 96858 83837 96860
rect 51019 96802 51024 96858
rect 51080 96802 83450 96858
rect 83556 96802 83776 96858
rect 83832 96802 83837 96858
rect 51019 96800 83450 96802
rect 51019 96797 51085 96800
rect 83444 96798 83450 96800
rect 83514 96800 83837 96802
rect 83514 96798 83561 96800
rect 83495 96797 83561 96798
rect 83771 96797 83837 96800
rect 84732 96798 84738 96862
rect 84802 96860 84808 96862
rect 85335 96860 85401 96863
rect 84802 96858 85401 96860
rect 84802 96802 85340 96858
rect 85396 96802 85401 96858
rect 84802 96800 85401 96802
rect 84802 96798 84808 96800
rect 85335 96797 85401 96800
rect 64543 96724 64609 96727
rect 50210 96722 50302 96724
rect 50252 96666 50302 96722
rect 50210 96664 50302 96666
rect 50404 96722 64609 96724
rect 50404 96666 64548 96722
rect 64604 96666 64609 96722
rect 50404 96664 64609 96666
rect 50210 96662 50257 96664
rect 48903 96661 48969 96662
rect 50191 96661 50257 96662
rect 64543 96661 64609 96664
rect 66567 96724 66633 96727
rect 73467 96724 73533 96727
rect 66567 96722 73533 96724
rect 66567 96666 66572 96722
rect 66628 96666 73472 96722
rect 73528 96666 73533 96722
rect 66567 96664 73533 96666
rect 66567 96661 66633 96664
rect 73467 96661 73533 96664
rect 81471 96724 81537 96727
rect 82156 96724 82162 96726
rect 81471 96722 82162 96724
rect 81471 96666 81476 96722
rect 81532 96666 82162 96722
rect 81471 96664 82162 96666
rect 81471 96661 81537 96664
rect 82156 96662 82162 96664
rect 82226 96662 82232 96726
rect 84139 96724 84205 96727
rect 82532 96722 84205 96724
rect 82532 96666 84144 96722
rect 84200 96666 84205 96722
rect 82532 96664 84205 96666
rect 46603 96588 46669 96591
rect 24707 96586 24816 96588
rect 24707 96530 24712 96586
rect 24768 96530 24816 96586
rect 24707 96525 24816 96530
rect 42052 96586 46669 96588
rect 42052 96530 46608 96586
rect 46664 96530 46669 96586
rect 42052 96528 46669 96530
rect 46603 96525 46669 96528
rect 64911 96588 64977 96591
rect 77975 96588 78041 96591
rect 82532 96590 82592 96664
rect 84139 96661 84205 96664
rect 84878 96658 85198 96659
rect 84878 96594 84886 96658
rect 84950 96594 84966 96658
rect 85030 96594 85046 96658
rect 85110 96594 85126 96658
rect 85190 96594 85198 96658
rect 84878 96593 85198 96594
rect 82524 96588 82530 96590
rect 64911 96586 78041 96588
rect 64911 96530 64916 96586
rect 64972 96530 77980 96586
rect 78036 96530 78041 96586
rect 64911 96528 78041 96530
rect 64911 96525 64977 96528
rect 77975 96525 78041 96528
rect 82348 96528 82530 96588
rect 4508 96452 4514 96454
rect 4099 96450 4514 96452
rect 4099 96394 4104 96450
rect 4160 96394 4514 96450
rect 4099 96392 4514 96394
rect 4099 96389 4165 96392
rect 4508 96390 4514 96392
rect 4578 96390 4584 96454
rect 24756 96452 24816 96525
rect 24708 96392 24816 96452
rect 33631 96452 33697 96455
rect 34692 96452 34936 96486
rect 40388 96452 40394 96454
rect 33631 96450 40394 96452
rect 33631 96394 33636 96450
rect 33692 96426 40394 96450
rect 33692 96394 34752 96426
rect 33631 96392 34752 96394
rect 34876 96392 40394 96426
rect 3179 96316 3245 96319
rect 3772 96316 3778 96318
rect 3179 96314 3778 96316
rect 3179 96258 3184 96314
rect 3240 96258 3778 96314
rect 3179 96256 3778 96258
rect 3179 96253 3245 96256
rect 3772 96254 3778 96256
rect 3842 96316 3848 96318
rect 4191 96316 4257 96319
rect 3842 96314 4257 96316
rect 3842 96258 4196 96314
rect 4252 96258 4257 96314
rect 3842 96256 4257 96258
rect 24708 96316 24768 96392
rect 33631 96389 33697 96392
rect 40388 96390 40394 96392
rect 40458 96390 40464 96454
rect 55527 96452 55593 96455
rect 62059 96452 62125 96455
rect 55527 96450 62125 96452
rect 55527 96394 55532 96450
rect 55588 96394 62064 96450
rect 62120 96394 62125 96450
rect 55527 96392 62125 96394
rect 55527 96389 55593 96392
rect 62059 96389 62125 96392
rect 73559 96452 73625 96455
rect 82348 96452 82408 96528
rect 82524 96526 82530 96528
rect 82594 96526 82600 96590
rect 85427 96588 85493 96591
rect 88454 96588 88934 96618
rect 85427 96586 88934 96588
rect 85427 96530 85432 96586
rect 85488 96530 88934 96586
rect 85427 96528 88934 96530
rect 85427 96525 85493 96528
rect 88454 96498 88934 96528
rect 73559 96450 82408 96452
rect 73559 96394 73564 96450
rect 73620 96394 82408 96450
rect 73559 96392 82408 96394
rect 73559 96389 73625 96392
rect 24983 96316 25049 96319
rect 83587 96316 83653 96319
rect 83771 96318 83837 96319
rect 83771 96316 83818 96318
rect 24708 96314 25049 96316
rect 24708 96258 24988 96314
rect 25044 96258 25049 96314
rect 24708 96256 25049 96258
rect 3842 96254 3848 96256
rect 4191 96253 4257 96256
rect 24983 96253 25049 96256
rect 47020 96314 83818 96316
rect 47020 96258 83592 96314
rect 83648 96258 83776 96314
rect 47020 96256 83818 96258
rect 38139 96182 38205 96183
rect 47020 96182 47080 96256
rect 83587 96253 83653 96256
rect 83771 96254 83818 96256
rect 83882 96254 83888 96318
rect 83771 96253 83837 96254
rect 47615 96182 47681 96183
rect 38139 96180 38186 96182
rect 38094 96178 38186 96180
rect 38094 96122 38144 96178
rect 38094 96120 38186 96122
rect 38139 96118 38186 96120
rect 38250 96118 38256 96182
rect 47012 96118 47018 96182
rect 47082 96118 47088 96182
rect 47564 96118 47570 96182
rect 47634 96180 47681 96182
rect 62427 96180 62493 96183
rect 82483 96180 82549 96183
rect 47634 96178 47726 96180
rect 47676 96122 47726 96178
rect 47634 96120 47726 96122
rect 62427 96178 82549 96180
rect 62427 96122 62432 96178
rect 62488 96122 82488 96178
rect 82544 96122 82549 96178
rect 62427 96120 82549 96122
rect 47634 96118 47681 96120
rect 38139 96117 38205 96118
rect 47615 96117 47681 96118
rect 62427 96117 62493 96120
rect 82483 96117 82549 96120
rect 2878 96114 3198 96115
rect 2878 96050 2886 96114
rect 2950 96050 2966 96114
rect 3030 96050 3046 96114
rect 3110 96050 3126 96114
rect 3190 96050 3198 96114
rect 2878 96049 3198 96050
rect 86878 96114 87198 96115
rect 86878 96050 86886 96114
rect 86950 96050 86966 96114
rect 87030 96050 87046 96114
rect 87110 96050 87126 96114
rect 87190 96050 87198 96114
rect 86878 96049 87198 96050
rect 18359 96044 18425 96047
rect 23419 96046 23485 96047
rect 18492 96044 18498 96046
rect 18359 96042 18498 96044
rect 18359 95986 18364 96042
rect 18420 95986 18498 96042
rect 18359 95984 18498 95986
rect 18359 95981 18425 95984
rect 18492 95982 18498 95984
rect 18562 95982 18568 96046
rect 23408 95982 23414 96046
rect 23478 96044 23485 96046
rect 23478 96042 23570 96044
rect 23480 95986 23570 96042
rect 23478 95984 23570 95986
rect 23478 95982 23485 95984
rect 32660 95982 32666 96046
rect 32730 96044 32736 96046
rect 81839 96044 81905 96047
rect 32730 96042 81905 96044
rect 32730 95986 81844 96042
rect 81900 95986 81905 96042
rect 32730 95984 81905 95986
rect 32730 95982 32736 95984
rect 23419 95981 23485 95982
rect 81839 95981 81905 95984
rect 14035 95910 14101 95911
rect 14035 95908 14070 95910
rect 13978 95906 14070 95908
rect 13978 95850 14040 95906
rect 13978 95848 14070 95850
rect 14035 95846 14070 95848
rect 14134 95846 14140 95910
rect 16979 95908 17045 95911
rect 23971 95910 24037 95911
rect 17568 95908 17574 95910
rect 16979 95906 17574 95908
rect 16979 95850 16984 95906
rect 17040 95850 17574 95906
rect 16979 95848 17574 95850
rect 14035 95845 14101 95846
rect 16979 95845 17045 95848
rect 17568 95846 17574 95848
rect 17638 95846 17644 95910
rect 23971 95908 24018 95910
rect 23926 95906 24018 95908
rect 23926 95850 23976 95906
rect 23926 95848 24018 95850
rect 23971 95846 24018 95848
rect 24082 95846 24088 95910
rect 31740 95846 31746 95910
rect 31810 95908 31816 95910
rect 81655 95908 81721 95911
rect 31810 95906 81721 95908
rect 31810 95850 81660 95906
rect 81716 95850 81721 95906
rect 31810 95848 81721 95850
rect 31810 95846 31816 95848
rect 23971 95845 24037 95846
rect 81655 95845 81721 95848
rect 19831 95774 19897 95775
rect 19780 95772 19786 95774
rect 19740 95712 19786 95772
rect 19850 95770 19897 95774
rect 19892 95714 19897 95770
rect 19780 95710 19786 95712
rect 19850 95710 19897 95714
rect 29348 95710 29354 95774
rect 29418 95772 29424 95774
rect 80091 95772 80157 95775
rect 29418 95770 80157 95772
rect 29418 95714 80096 95770
rect 80152 95714 80157 95770
rect 29418 95712 80157 95714
rect 29418 95710 29424 95712
rect 19831 95709 19897 95710
rect 80091 95709 80157 95712
rect 27191 95638 27257 95639
rect 51479 95638 51545 95639
rect 27140 95574 27146 95638
rect 27210 95636 27257 95638
rect 27210 95634 27302 95636
rect 27252 95578 27302 95634
rect 27210 95576 27302 95578
rect 27210 95574 27257 95576
rect 51428 95574 51434 95638
rect 51498 95636 51545 95638
rect 51498 95634 51590 95636
rect 51540 95578 51590 95634
rect 51498 95576 51590 95578
rect 51498 95574 51545 95576
rect 27191 95573 27257 95574
rect 51479 95573 51545 95574
rect 878 95570 1198 95571
rect 878 95506 886 95570
rect 950 95506 966 95570
rect 1030 95506 1046 95570
rect 1110 95506 1126 95570
rect 1190 95506 1198 95570
rect 878 95505 1198 95506
rect 84878 95570 85198 95571
rect 84878 95506 84886 95570
rect 84950 95506 84966 95570
rect 85030 95506 85046 95570
rect 85110 95506 85126 95570
rect 85190 95506 85198 95570
rect 84878 95505 85198 95506
rect 16979 95500 17045 95503
rect 84507 95500 84573 95503
rect 16979 95498 84573 95500
rect 16979 95442 16984 95498
rect 17040 95442 84512 95498
rect 84568 95442 84573 95498
rect 16979 95440 84573 95442
rect 16979 95437 17045 95440
rect 84507 95437 84573 95440
rect 20751 95364 20817 95367
rect 83219 95364 83285 95367
rect 20751 95362 83285 95364
rect 20751 95306 20756 95362
rect 20812 95306 83224 95362
rect 83280 95306 83285 95362
rect 20751 95304 83285 95306
rect 20751 95301 20817 95304
rect 83219 95301 83285 95304
rect 85151 95364 85217 95367
rect 88454 95364 88934 95394
rect 85151 95362 88934 95364
rect 85151 95306 85156 95362
rect 85212 95306 88934 95362
rect 85151 95304 88934 95306
rect 85151 95301 85217 95304
rect 88454 95274 88934 95304
rect 24431 95230 24497 95231
rect 25719 95230 25785 95231
rect 26639 95230 26705 95231
rect 24380 95228 24386 95230
rect 24340 95168 24386 95228
rect 24450 95226 24497 95230
rect 25668 95228 25674 95230
rect 24492 95170 24497 95226
rect 24380 95166 24386 95168
rect 24450 95166 24497 95170
rect 25628 95168 25674 95228
rect 25738 95226 25785 95230
rect 26588 95228 26594 95230
rect 25780 95170 25785 95226
rect 25668 95166 25674 95168
rect 25738 95166 25785 95170
rect 26548 95168 26594 95228
rect 26658 95226 26705 95230
rect 26700 95170 26705 95226
rect 26588 95166 26594 95168
rect 26658 95166 26705 95170
rect 34316 95166 34322 95230
rect 34386 95228 34392 95230
rect 34459 95228 34525 95231
rect 35655 95230 35721 95231
rect 36207 95230 36273 95231
rect 37495 95230 37561 95231
rect 38599 95230 38665 95231
rect 35604 95228 35610 95230
rect 34386 95226 34525 95228
rect 34386 95170 34464 95226
rect 34520 95170 34525 95226
rect 34386 95168 34525 95170
rect 35564 95168 35610 95228
rect 35674 95226 35721 95230
rect 36156 95228 36162 95230
rect 35716 95170 35721 95226
rect 34386 95166 34392 95168
rect 24431 95165 24497 95166
rect 25719 95165 25785 95166
rect 26639 95165 26705 95166
rect 34459 95165 34525 95168
rect 35604 95166 35610 95168
rect 35674 95166 35721 95170
rect 36116 95168 36162 95228
rect 36226 95226 36273 95230
rect 37444 95228 37450 95230
rect 36268 95170 36273 95226
rect 36156 95166 36162 95168
rect 36226 95166 36273 95170
rect 37404 95168 37450 95228
rect 37514 95226 37561 95230
rect 38548 95228 38554 95230
rect 37556 95170 37561 95226
rect 37444 95166 37450 95168
rect 37514 95166 37561 95170
rect 38508 95168 38554 95228
rect 38618 95226 38665 95230
rect 38660 95170 38665 95226
rect 38548 95166 38554 95168
rect 38618 95166 38665 95170
rect 35655 95165 35721 95166
rect 36207 95165 36273 95166
rect 37495 95165 37561 95166
rect 38599 95165 38665 95166
rect 41819 95230 41885 95231
rect 43751 95230 43817 95231
rect 44487 95230 44553 95231
rect 46511 95230 46577 95231
rect 47799 95230 47865 95231
rect 48719 95230 48785 95231
rect 50191 95230 50257 95231
rect 41819 95226 41866 95230
rect 41930 95228 41936 95230
rect 43700 95228 43706 95230
rect 41819 95170 41824 95226
rect 41819 95166 41866 95170
rect 41930 95168 41976 95228
rect 43660 95168 43706 95228
rect 43770 95226 43817 95230
rect 44436 95228 44442 95230
rect 43812 95170 43817 95226
rect 41930 95166 41936 95168
rect 43700 95166 43706 95168
rect 43770 95166 43817 95170
rect 44396 95168 44442 95228
rect 44506 95226 44553 95230
rect 46460 95228 46466 95230
rect 44548 95170 44553 95226
rect 44436 95166 44442 95168
rect 44506 95166 44553 95170
rect 46420 95168 46466 95228
rect 46530 95226 46577 95230
rect 47748 95228 47754 95230
rect 46572 95170 46577 95226
rect 46460 95166 46466 95168
rect 46530 95166 46577 95170
rect 47708 95168 47754 95228
rect 47818 95226 47865 95230
rect 48668 95228 48674 95230
rect 47860 95170 47865 95226
rect 47748 95166 47754 95168
rect 47818 95166 47865 95170
rect 48628 95168 48674 95228
rect 48738 95226 48785 95230
rect 50140 95228 50146 95230
rect 48780 95170 48785 95226
rect 48668 95166 48674 95168
rect 48738 95166 48785 95170
rect 50100 95168 50146 95228
rect 50210 95226 50257 95230
rect 50252 95170 50257 95226
rect 50140 95166 50146 95168
rect 50210 95166 50257 95170
rect 51428 95166 51434 95230
rect 51498 95228 51504 95230
rect 51571 95228 51637 95231
rect 56631 95230 56697 95231
rect 57919 95230 57985 95231
rect 59391 95230 59457 95231
rect 61783 95230 61849 95231
rect 56580 95228 56586 95230
rect 51498 95226 51637 95228
rect 51498 95170 51576 95226
rect 51632 95170 51637 95226
rect 51498 95168 51637 95170
rect 56540 95168 56586 95228
rect 56650 95226 56697 95230
rect 57868 95228 57874 95230
rect 56692 95170 56697 95226
rect 51498 95166 51504 95168
rect 41819 95165 41885 95166
rect 43751 95165 43817 95166
rect 44487 95165 44553 95166
rect 46511 95165 46577 95166
rect 47799 95165 47865 95166
rect 48719 95165 48785 95166
rect 50191 95165 50257 95166
rect 51571 95165 51637 95168
rect 56580 95166 56586 95168
rect 56650 95166 56697 95170
rect 57828 95168 57874 95228
rect 57938 95226 57985 95230
rect 59340 95228 59346 95230
rect 57980 95170 57985 95226
rect 57868 95166 57874 95168
rect 57938 95166 57985 95170
rect 59300 95168 59346 95228
rect 59410 95226 59457 95230
rect 61732 95228 61738 95230
rect 59452 95170 59457 95226
rect 59340 95166 59346 95168
rect 59410 95166 59457 95170
rect 61692 95168 61738 95228
rect 61802 95226 61849 95230
rect 61844 95170 61849 95226
rect 61732 95166 61738 95168
rect 61802 95166 61849 95170
rect 62652 95166 62658 95230
rect 62722 95228 62728 95230
rect 62795 95228 62861 95231
rect 62722 95226 62861 95228
rect 62722 95170 62800 95226
rect 62856 95170 62861 95226
rect 62722 95168 62861 95170
rect 62722 95166 62728 95168
rect 56631 95165 56697 95166
rect 57919 95165 57985 95166
rect 59391 95165 59457 95166
rect 61783 95165 61849 95166
rect 62795 95165 62861 95168
rect 4283 95094 4349 95095
rect 8147 95094 8213 95095
rect 4283 95090 4330 95094
rect 4394 95092 4400 95094
rect 4283 95034 4288 95090
rect 4283 95030 4330 95034
rect 4394 95032 4440 95092
rect 8147 95090 8194 95094
rect 8258 95092 8264 95094
rect 11827 95092 11893 95095
rect 12236 95092 12242 95094
rect 8147 95034 8152 95090
rect 4394 95030 4400 95032
rect 8147 95030 8194 95034
rect 8258 95032 8304 95092
rect 11827 95090 12242 95092
rect 11827 95034 11832 95090
rect 11888 95034 12242 95090
rect 11827 95032 12242 95034
rect 8258 95030 8264 95032
rect 4283 95029 4349 95030
rect 8147 95029 8213 95030
rect 11827 95029 11893 95032
rect 12236 95030 12242 95032
rect 12306 95030 12312 95094
rect 31147 95092 31213 95095
rect 36299 95094 36365 95095
rect 31372 95092 31378 95094
rect 31147 95090 31378 95092
rect 31147 95034 31152 95090
rect 31208 95034 31378 95090
rect 31147 95032 31378 95034
rect 31147 95029 31213 95032
rect 31372 95030 31378 95032
rect 31442 95030 31448 95094
rect 36299 95092 36346 95094
rect 36254 95090 36346 95092
rect 36254 95034 36304 95090
rect 36254 95032 36346 95034
rect 36299 95030 36346 95032
rect 36410 95030 36416 95094
rect 36708 95030 36714 95094
rect 36778 95092 36784 95094
rect 37311 95092 37377 95095
rect 38783 95094 38849 95095
rect 36778 95090 37377 95092
rect 36778 95034 37316 95090
rect 37372 95034 37377 95090
rect 36778 95032 37377 95034
rect 36778 95030 36784 95032
rect 36299 95029 36365 95030
rect 37311 95029 37377 95032
rect 38732 95030 38738 95094
rect 38802 95092 38849 95094
rect 38802 95090 38894 95092
rect 38844 95034 38894 95090
rect 38802 95032 38894 95034
rect 38802 95030 38849 95032
rect 43332 95030 43338 95094
rect 43402 95092 43408 95094
rect 43935 95092 44001 95095
rect 43402 95090 44001 95092
rect 43402 95034 43940 95090
rect 43996 95034 44001 95090
rect 43402 95032 44001 95034
rect 43402 95030 43408 95032
rect 38783 95029 38849 95030
rect 43935 95029 44001 95032
rect 47932 95030 47938 95094
rect 48002 95092 48008 95094
rect 49087 95092 49153 95095
rect 50375 95094 50441 95095
rect 54239 95094 54305 95095
rect 48002 95090 49153 95092
rect 48002 95034 49092 95090
rect 49148 95034 49153 95090
rect 48002 95032 49153 95034
rect 48002 95030 48008 95032
rect 49087 95029 49153 95032
rect 50324 95030 50330 95094
rect 50394 95092 50441 95094
rect 50394 95090 50486 95092
rect 50436 95034 50486 95090
rect 50394 95032 50486 95034
rect 50394 95030 50441 95032
rect 54188 95030 54194 95094
rect 54258 95092 54305 95094
rect 58103 95092 58169 95095
rect 66475 95092 66541 95095
rect 54258 95090 54350 95092
rect 54300 95034 54350 95090
rect 54258 95032 54350 95034
rect 58103 95090 66541 95092
rect 58103 95034 58108 95090
rect 58164 95034 66480 95090
rect 66536 95034 66541 95090
rect 58103 95032 66541 95034
rect 54258 95030 54305 95032
rect 50375 95029 50441 95030
rect 54239 95029 54305 95030
rect 58103 95029 58169 95032
rect 66475 95029 66541 95032
rect 2878 95026 3198 95027
rect 2878 94962 2886 95026
rect 2950 94962 2966 95026
rect 3030 94962 3046 95026
rect 3110 94962 3126 95026
rect 3190 94962 3198 95026
rect 2878 94961 3198 94962
rect 86878 95026 87198 95027
rect 86878 94962 86886 95026
rect 86950 94962 86966 95026
rect 87030 94962 87046 95026
rect 87110 94962 87126 95026
rect 87190 94962 87198 95026
rect 86878 94961 87198 94962
rect 11091 94956 11157 94959
rect 11316 94956 11322 94958
rect 11091 94954 11322 94956
rect 11091 94898 11096 94954
rect 11152 94898 11322 94954
rect 11091 94896 11322 94898
rect 11091 94893 11157 94896
rect 11316 94894 11322 94896
rect 11386 94894 11392 94958
rect 22724 94894 22730 94958
rect 22794 94956 22800 94958
rect 23327 94956 23393 94959
rect 22794 94954 23393 94956
rect 22794 94898 23332 94954
rect 23388 94898 23393 94954
rect 22794 94896 23393 94898
rect 22794 94894 22800 94896
rect 23327 94893 23393 94896
rect 25300 94894 25306 94958
rect 25370 94956 25376 94958
rect 25903 94956 25969 94959
rect 25370 94954 25969 94956
rect 25370 94898 25908 94954
rect 25964 94898 25969 94954
rect 25370 94896 25969 94898
rect 25370 94894 25376 94896
rect 25903 94893 25969 94896
rect 35011 94956 35077 94959
rect 80091 94956 80157 94959
rect 35011 94954 80157 94956
rect 35011 94898 35016 94954
rect 35072 94898 80096 94954
rect 80152 94898 80157 94954
rect 35011 94896 80157 94898
rect 35011 94893 35077 94896
rect 80091 94893 80157 94896
rect 18175 94822 18241 94823
rect 18124 94758 18130 94822
rect 18194 94820 18241 94822
rect 19831 94820 19897 94823
rect 19964 94820 19970 94822
rect 18194 94818 18286 94820
rect 18236 94762 18286 94818
rect 18194 94760 18286 94762
rect 19831 94818 19970 94820
rect 19831 94762 19836 94818
rect 19892 94762 19970 94818
rect 19831 94760 19970 94762
rect 18194 94758 18241 94760
rect 18175 94757 18241 94758
rect 19831 94757 19897 94760
rect 19964 94758 19970 94760
rect 20034 94758 20040 94822
rect 20843 94820 20909 94823
rect 21436 94820 21442 94822
rect 20843 94818 21442 94820
rect 20843 94762 20848 94818
rect 20904 94762 21442 94818
rect 20843 94760 21442 94762
rect 20843 94757 20909 94760
rect 21436 94758 21442 94760
rect 21506 94758 21512 94822
rect 25995 94820 26061 94823
rect 26404 94820 26410 94822
rect 25995 94818 26410 94820
rect 25995 94762 26000 94818
rect 26056 94762 26410 94818
rect 25995 94760 26410 94762
rect 25995 94757 26061 94760
rect 26404 94758 26410 94760
rect 26474 94758 26480 94822
rect 49772 94758 49778 94822
rect 49842 94820 49848 94822
rect 50283 94820 50349 94823
rect 49842 94818 50349 94820
rect 49842 94762 50288 94818
rect 50344 94762 50349 94818
rect 49842 94760 50349 94762
rect 49842 94758 49848 94760
rect 50283 94757 50349 94760
rect 52348 94758 52354 94822
rect 52418 94820 52424 94822
rect 54147 94820 54213 94823
rect 85887 94820 85953 94823
rect 52418 94760 54072 94820
rect 52418 94758 52424 94760
rect 27283 94684 27349 94687
rect 32435 94686 32501 94687
rect 27508 94684 27514 94686
rect 27283 94682 27514 94684
rect 27283 94626 27288 94682
rect 27344 94626 27514 94682
rect 27283 94624 27514 94626
rect 27283 94621 27349 94624
rect 27508 94622 27514 94624
rect 27578 94622 27584 94686
rect 32435 94684 32482 94686
rect 32390 94682 32482 94684
rect 32390 94626 32440 94682
rect 32390 94624 32482 94626
rect 32435 94622 32482 94624
rect 32546 94622 32552 94686
rect 48484 94622 48490 94686
rect 48554 94684 48560 94686
rect 49087 94684 49153 94687
rect 48554 94682 49153 94684
rect 48554 94626 49092 94682
rect 49148 94626 49153 94682
rect 48554 94624 49153 94626
rect 48554 94622 48560 94624
rect 32435 94621 32501 94622
rect 49087 94621 49153 94624
rect 52716 94622 52722 94686
rect 52786 94684 52792 94686
rect 52951 94684 53017 94687
rect 52786 94682 53017 94684
rect 52786 94626 52956 94682
rect 53012 94626 53017 94682
rect 52786 94624 53017 94626
rect 54012 94684 54072 94760
rect 54147 94818 85953 94820
rect 54147 94762 54152 94818
rect 54208 94762 85892 94818
rect 85948 94762 85953 94818
rect 54147 94760 85953 94762
rect 54147 94757 54213 94760
rect 85887 94757 85953 94760
rect 82667 94684 82733 94687
rect 83812 94684 83818 94686
rect 54012 94682 83818 94684
rect 54012 94626 82672 94682
rect 82728 94626 83818 94682
rect 54012 94624 83818 94626
rect 52786 94622 52792 94624
rect 52951 94621 53017 94624
rect 82667 94621 82733 94624
rect 83812 94622 83818 94624
rect 83882 94622 83888 94686
rect 40071 94550 40137 94551
rect 40020 94486 40026 94550
rect 40090 94548 40137 94550
rect 41451 94550 41517 94551
rect 42647 94550 42713 94551
rect 41451 94548 41498 94550
rect 40090 94546 40182 94548
rect 40132 94490 40182 94546
rect 40090 94488 40182 94490
rect 41406 94546 41498 94548
rect 41406 94490 41456 94546
rect 41406 94488 41498 94490
rect 40090 94486 40137 94488
rect 40071 94485 40137 94486
rect 41451 94486 41498 94488
rect 41562 94486 41568 94550
rect 42596 94486 42602 94550
rect 42666 94548 42713 94550
rect 42666 94546 42758 94548
rect 42708 94490 42758 94546
rect 42666 94488 42758 94490
rect 42666 94486 42713 94488
rect 53820 94486 53826 94550
rect 53890 94548 53896 94550
rect 68499 94548 68565 94551
rect 53890 94546 68565 94548
rect 53890 94490 68504 94546
rect 68560 94490 68565 94546
rect 53890 94488 68565 94490
rect 53890 94486 53896 94488
rect 41451 94485 41517 94486
rect 42647 94485 42713 94486
rect 68499 94485 68565 94488
rect 70983 94548 71049 94551
rect 83219 94548 83285 94551
rect 84139 94548 84205 94551
rect 70983 94546 84205 94548
rect 70983 94490 70988 94546
rect 71044 94490 83224 94546
rect 83280 94490 84144 94546
rect 84200 94490 84205 94546
rect 70983 94488 84205 94490
rect 70983 94485 71049 94488
rect 83219 94485 83285 94488
rect 84139 94485 84205 94488
rect 878 94482 1198 94483
rect 878 94418 886 94482
rect 950 94418 966 94482
rect 1030 94418 1046 94482
rect 1110 94418 1126 94482
rect 1190 94418 1198 94482
rect 878 94417 1198 94418
rect 84878 94482 85198 94483
rect 84878 94418 84886 94482
rect 84950 94418 84966 94482
rect 85030 94418 85046 94482
rect 85110 94418 85126 94482
rect 85190 94418 85198 94482
rect 84878 94417 85198 94418
rect 18267 94412 18333 94415
rect 29767 94414 29833 94415
rect 18676 94412 18682 94414
rect 18267 94410 18682 94412
rect 18267 94354 18272 94410
rect 18328 94354 18682 94410
rect 18267 94352 18682 94354
rect 18267 94349 18333 94352
rect 18676 94350 18682 94352
rect 18746 94350 18752 94414
rect 29716 94350 29722 94414
rect 29786 94412 29833 94414
rect 41267 94414 41333 94415
rect 41727 94414 41793 94415
rect 43935 94414 44001 94415
rect 41267 94412 41314 94414
rect 29786 94410 29878 94412
rect 29828 94354 29878 94410
rect 29786 94352 29878 94354
rect 41222 94410 41314 94412
rect 41222 94354 41272 94410
rect 41222 94352 41314 94354
rect 29786 94350 29833 94352
rect 29767 94349 29833 94350
rect 41267 94350 41314 94352
rect 41378 94350 41384 94414
rect 41676 94412 41682 94414
rect 41636 94352 41682 94412
rect 41746 94410 41793 94414
rect 41788 94354 41793 94410
rect 41676 94350 41682 94352
rect 41746 94350 41793 94354
rect 43884 94350 43890 94414
rect 43954 94412 44001 94414
rect 43954 94410 44046 94412
rect 43996 94354 44046 94410
rect 43954 94352 44046 94354
rect 43954 94350 44001 94352
rect 44620 94350 44626 94414
rect 44690 94412 44696 94414
rect 45223 94412 45289 94415
rect 51663 94414 51729 94415
rect 44690 94410 45289 94412
rect 44690 94354 45228 94410
rect 45284 94354 45289 94410
rect 44690 94352 45289 94354
rect 44690 94350 44696 94352
rect 41267 94349 41333 94350
rect 41727 94349 41793 94350
rect 43935 94349 44001 94350
rect 45223 94349 45289 94352
rect 51612 94350 51618 94414
rect 51682 94412 51729 94414
rect 56355 94412 56421 94415
rect 66475 94412 66541 94415
rect 51682 94410 51774 94412
rect 51724 94354 51774 94410
rect 51682 94352 51774 94354
rect 56355 94410 66541 94412
rect 56355 94354 56360 94410
rect 56416 94354 66480 94410
rect 66536 94354 66541 94410
rect 56355 94352 66541 94354
rect 51682 94350 51729 94352
rect 51663 94349 51729 94350
rect 56355 94349 56421 94352
rect 66475 94349 66541 94352
rect 69828 94350 69834 94414
rect 69898 94350 69904 94414
rect 70983 94412 71049 94415
rect 81747 94412 81813 94415
rect 70983 94410 81813 94412
rect 70983 94354 70988 94410
rect 71044 94354 81752 94410
rect 81808 94354 81813 94410
rect 70983 94352 81813 94354
rect 21804 94214 21810 94278
rect 21874 94276 21880 94278
rect 56907 94276 56973 94279
rect 21874 94274 56973 94276
rect 21874 94218 56912 94274
rect 56968 94218 56973 94274
rect 21874 94216 56973 94218
rect 21874 94214 21880 94216
rect 56907 94213 56973 94216
rect 61967 94276 62033 94279
rect 69836 94276 69896 94350
rect 70983 94349 71049 94352
rect 81747 94349 81813 94352
rect 61967 94274 69896 94276
rect 61967 94218 61972 94274
rect 62028 94218 69896 94274
rect 61967 94216 69896 94218
rect 61967 94213 62033 94216
rect 23828 94078 23834 94142
rect 23898 94140 23904 94142
rect 24615 94140 24681 94143
rect 23898 94138 24681 94140
rect 23898 94082 24620 94138
rect 24676 94082 24681 94138
rect 23898 94080 24681 94082
rect 23898 94078 23904 94080
rect 24615 94077 24681 94080
rect 28244 94078 28250 94142
rect 28314 94140 28320 94142
rect 28387 94140 28453 94143
rect 28314 94138 28453 94140
rect 28314 94082 28392 94138
rect 28448 94082 28453 94138
rect 28314 94080 28453 94082
rect 28314 94078 28320 94080
rect 28387 94077 28453 94080
rect 42647 94140 42713 94143
rect 84783 94140 84849 94143
rect 88454 94140 88934 94170
rect 42647 94138 84064 94140
rect 42647 94082 42652 94138
rect 42708 94082 84064 94138
rect 42647 94080 84064 94082
rect 42647 94077 42713 94080
rect 30636 93942 30642 94006
rect 30706 94004 30712 94006
rect 31055 94004 31121 94007
rect 30706 94002 31121 94004
rect 30706 93946 31060 94002
rect 31116 93946 31121 94002
rect 30706 93944 31121 93946
rect 30706 93942 30712 93944
rect 31055 93941 31121 93944
rect 45724 93942 45730 94006
rect 45794 94004 45800 94006
rect 46143 94004 46209 94007
rect 45794 94002 46209 94004
rect 45794 93946 46148 94002
rect 46204 93946 46209 94002
rect 45794 93944 46209 93946
rect 45794 93942 45800 93944
rect 46143 93941 46209 93944
rect 52900 93942 52906 94006
rect 52970 94004 52976 94006
rect 54147 94004 54213 94007
rect 82708 94004 82714 94006
rect 52970 94002 54213 94004
rect 52970 93946 54152 94002
rect 54208 93946 54213 94002
rect 52970 93944 54213 93946
rect 52970 93942 52976 93944
rect 54147 93941 54213 93944
rect 73746 93944 82714 94004
rect 2878 93938 3198 93939
rect 2878 93874 2886 93938
rect 2950 93874 2966 93938
rect 3030 93874 3046 93938
rect 3110 93874 3126 93938
rect 3190 93874 3198 93938
rect 2878 93873 3198 93874
rect 30687 93870 30753 93871
rect 32343 93870 32409 93871
rect 30636 93868 30642 93870
rect 30596 93808 30642 93868
rect 30706 93866 30753 93870
rect 30748 93810 30753 93866
rect 30636 93806 30642 93808
rect 30706 93806 30753 93810
rect 32292 93806 32298 93870
rect 32362 93868 32409 93870
rect 32362 93866 32454 93868
rect 32404 93810 32454 93866
rect 32362 93808 32454 93810
rect 32362 93806 32409 93808
rect 33396 93806 33402 93870
rect 33466 93868 33472 93870
rect 33631 93868 33697 93871
rect 33466 93866 33697 93868
rect 33466 93810 33636 93866
rect 33692 93810 33697 93866
rect 33466 93808 33697 93810
rect 33466 93806 33472 93808
rect 30687 93805 30753 93806
rect 32343 93805 32409 93806
rect 33631 93805 33697 93808
rect 34684 93806 34690 93870
rect 34754 93868 34760 93870
rect 34919 93868 34985 93871
rect 34754 93866 34985 93868
rect 34754 93810 34924 93866
rect 34980 93810 34985 93866
rect 34754 93808 34985 93810
rect 34754 93806 34760 93808
rect 34919 93805 34985 93808
rect 35788 93806 35794 93870
rect 35858 93868 35864 93870
rect 36207 93868 36273 93871
rect 35858 93866 36273 93868
rect 35858 93810 36212 93866
rect 36268 93810 36273 93866
rect 35858 93808 36273 93810
rect 35858 93806 35864 93808
rect 36207 93805 36273 93808
rect 37996 93806 38002 93870
rect 38066 93868 38072 93870
rect 38875 93868 38941 93871
rect 38066 93866 38941 93868
rect 38066 93810 38880 93866
rect 38936 93810 38941 93866
rect 38066 93808 38941 93810
rect 38066 93806 38072 93808
rect 38875 93805 38941 93808
rect 39955 93806 39961 93870
rect 40025 93868 40031 93870
rect 42739 93868 42805 93871
rect 53687 93870 53753 93871
rect 40025 93866 42805 93868
rect 40025 93810 42744 93866
rect 42800 93810 42805 93866
rect 40025 93808 42805 93810
rect 40025 93806 40031 93808
rect 42739 93805 42805 93808
rect 53683 93806 53689 93870
rect 53753 93868 53759 93870
rect 53753 93808 53844 93868
rect 53753 93806 53759 93808
rect 69828 93806 69834 93870
rect 69898 93868 69904 93870
rect 73746 93868 73806 93944
rect 82708 93942 82714 93944
rect 82778 94004 82784 94006
rect 83863 94004 83929 94007
rect 82778 94002 83929 94004
rect 82778 93946 83868 94002
rect 83924 93946 83929 94002
rect 82778 93944 83929 93946
rect 84004 94004 84064 94080
rect 84783 94138 88934 94140
rect 84783 94082 84788 94138
rect 84844 94082 88934 94138
rect 84783 94080 88934 94082
rect 84783 94077 84849 94080
rect 88454 94050 88934 94080
rect 86163 94004 86229 94007
rect 84004 94002 86229 94004
rect 84004 93946 86168 94002
rect 86224 93946 86229 94002
rect 84004 93944 86229 93946
rect 82778 93942 82784 93944
rect 83863 93941 83929 93944
rect 86163 93941 86229 93944
rect 86878 93938 87198 93939
rect 86878 93874 86886 93938
rect 86950 93874 86966 93938
rect 87030 93874 87046 93938
rect 87110 93874 87126 93938
rect 87190 93874 87198 93938
rect 86878 93873 87198 93874
rect 69898 93808 73806 93868
rect 78435 93870 78501 93871
rect 78435 93866 78482 93870
rect 78546 93868 78552 93870
rect 78435 93810 78440 93866
rect 69898 93806 69904 93808
rect 78435 93806 78482 93810
rect 78546 93808 78592 93868
rect 78546 93806 78552 93808
rect 53687 93805 53753 93806
rect 78435 93805 78501 93806
rect 36299 93732 36365 93735
rect 81839 93732 81905 93735
rect 36299 93730 81905 93732
rect 36299 93674 36304 93730
rect 36360 93674 81844 93730
rect 81900 93674 81905 93730
rect 36299 93672 81905 93674
rect 36299 93669 36365 93672
rect 81839 93669 81905 93672
rect 27475 93534 27481 93598
rect 27545 93596 27551 93598
rect 38047 93596 38113 93599
rect 27545 93594 38113 93596
rect 27545 93538 38052 93594
rect 38108 93538 38113 93594
rect 27545 93536 38113 93538
rect 27545 93534 27551 93536
rect 38047 93533 38113 93536
rect 38231 93596 38297 93599
rect 81655 93596 81721 93599
rect 38231 93594 81721 93596
rect 38231 93538 38236 93594
rect 38292 93538 81660 93594
rect 81716 93538 81721 93594
rect 38231 93536 81721 93538
rect 38231 93533 38297 93536
rect 81655 93533 81721 93536
rect 29675 93460 29741 93463
rect 82483 93460 82549 93463
rect 29675 93458 82549 93460
rect 29675 93402 29680 93458
rect 29736 93402 82488 93458
rect 82544 93402 82549 93458
rect 29675 93400 82549 93402
rect 29675 93397 29741 93400
rect 82483 93397 82549 93400
rect 878 93394 1198 93395
rect 878 93330 886 93394
rect 950 93330 966 93394
rect 1030 93330 1046 93394
rect 1110 93330 1126 93394
rect 1190 93330 1198 93394
rect 878 93329 1198 93330
rect 84878 93394 85198 93395
rect 84878 93330 84886 93394
rect 84950 93330 84966 93394
rect 85030 93330 85046 93394
rect 85110 93330 85126 93394
rect 85190 93330 85198 93394
rect 84878 93329 85198 93330
rect 27191 93324 27257 93327
rect 82115 93324 82181 93327
rect 27191 93322 82181 93324
rect 27191 93266 27196 93322
rect 27252 93266 82120 93322
rect 82176 93266 82181 93322
rect 27191 93264 82181 93266
rect 27191 93261 27257 93264
rect 82115 93261 82181 93264
rect 25852 93126 25858 93190
rect 25922 93188 25928 93190
rect 81379 93188 81445 93191
rect 25922 93186 81445 93188
rect 25922 93130 81384 93186
rect 81440 93130 81445 93186
rect 25922 93128 81445 93130
rect 25922 93126 25928 93128
rect 81379 93125 81445 93128
rect 48811 93052 48877 93055
rect 82299 93052 82365 93055
rect 48811 93050 82365 93052
rect 48811 92994 48816 93050
rect 48872 92994 82304 93050
rect 82360 92994 82365 93050
rect 48811 92992 82365 92994
rect 48811 92989 48877 92992
rect 82299 92989 82365 92992
rect 85151 93052 85217 93055
rect 85151 93050 87376 93052
rect 85151 92994 85156 93050
rect 85212 92994 87376 93050
rect 85151 92992 87376 92994
rect 85151 92989 85217 92992
rect 87316 92916 87376 92992
rect 88454 92916 88934 92946
rect 87316 92856 88934 92916
rect 2878 92850 3198 92851
rect 2878 92786 2886 92850
rect 2950 92786 2966 92850
rect 3030 92786 3046 92850
rect 3110 92786 3126 92850
rect 3190 92786 3198 92850
rect 2878 92785 3198 92786
rect 86878 92850 87198 92851
rect 86878 92786 86886 92850
rect 86950 92786 86966 92850
rect 87030 92786 87046 92850
rect 87110 92786 87126 92850
rect 87190 92786 87198 92850
rect 88454 92826 88934 92856
rect 86878 92785 87198 92786
rect 56907 92780 56973 92783
rect 80091 92780 80157 92783
rect 56907 92778 80157 92780
rect 56907 92722 56912 92778
rect 56968 92722 80096 92778
rect 80152 92722 80157 92778
rect 56907 92720 80157 92722
rect 56907 92717 56973 92720
rect 80091 92717 80157 92720
rect 55343 92646 55409 92647
rect 60495 92646 60561 92647
rect 73743 92646 73809 92647
rect 55292 92582 55298 92646
rect 55362 92644 55409 92646
rect 60444 92644 60450 92646
rect 55362 92642 55454 92644
rect 55404 92586 55454 92642
rect 55362 92584 55454 92586
rect 60404 92584 60450 92644
rect 60514 92642 60561 92646
rect 73692 92644 73698 92646
rect 60556 92586 60561 92642
rect 55362 92582 55409 92584
rect 60444 92582 60450 92584
rect 60514 92582 60561 92586
rect 73652 92584 73698 92644
rect 73762 92642 73809 92646
rect 73804 92586 73809 92642
rect 73692 92582 73698 92584
rect 73762 92582 73809 92586
rect 55343 92581 55409 92582
rect 60495 92581 60561 92582
rect 73743 92581 73809 92582
rect 878 92306 1198 92307
rect 878 92242 886 92306
rect 950 92242 966 92306
rect 1030 92242 1046 92306
rect 1110 92242 1126 92306
rect 1190 92242 1198 92306
rect 878 92241 1198 92242
rect 84878 92306 85198 92307
rect 84878 92242 84886 92306
rect 84950 92242 84966 92306
rect 85030 92242 85046 92306
rect 85110 92242 85126 92306
rect 85190 92242 85198 92306
rect 84878 92241 85198 92242
rect 85151 91964 85217 91967
rect 85151 91962 87376 91964
rect 85151 91906 85156 91962
rect 85212 91906 87376 91962
rect 85151 91904 87376 91906
rect 85151 91901 85217 91904
rect 82164 91828 82224 91838
rect 83955 91828 84021 91831
rect 82164 91826 84021 91828
rect 82164 91770 83960 91826
rect 84016 91770 84021 91826
rect 82164 91768 84021 91770
rect 83955 91765 84021 91768
rect 2878 91762 3198 91763
rect 2878 91698 2886 91762
rect 2950 91698 2966 91762
rect 3030 91698 3046 91762
rect 3110 91698 3126 91762
rect 3190 91698 3198 91762
rect 2878 91697 3198 91698
rect 86878 91762 87198 91763
rect 86878 91698 86886 91762
rect 86950 91698 86966 91762
rect 87030 91698 87046 91762
rect 87110 91698 87126 91762
rect 87190 91698 87198 91762
rect 86878 91697 87198 91698
rect 87316 91692 87376 91904
rect 88454 91692 88934 91722
rect 87316 91632 88934 91692
rect 88454 91602 88934 91632
rect 878 91218 1198 91219
rect 878 91154 886 91218
rect 950 91154 966 91218
rect 1030 91154 1046 91218
rect 1110 91154 1126 91218
rect 1190 91154 1198 91218
rect 878 91153 1198 91154
rect 84878 91218 85198 91219
rect 84878 91154 84886 91218
rect 84950 91154 84966 91218
rect 85030 91154 85046 91218
rect 85110 91154 85126 91218
rect 85190 91154 85198 91218
rect 84878 91153 85198 91154
rect 84047 90876 84113 90879
rect 84047 90874 87376 90876
rect 84047 90818 84052 90874
rect 84108 90818 87376 90874
rect 84047 90816 87376 90818
rect 84047 90813 84113 90816
rect 2878 90674 3198 90675
rect 2878 90610 2886 90674
rect 2950 90610 2966 90674
rect 3030 90610 3046 90674
rect 3110 90610 3126 90674
rect 3190 90610 3198 90674
rect 2878 90609 3198 90610
rect 86878 90674 87198 90675
rect 86878 90610 86886 90674
rect 86950 90610 86966 90674
rect 87030 90610 87046 90674
rect 87110 90610 87126 90674
rect 87190 90610 87198 90674
rect 86878 90609 87198 90610
rect 87316 90604 87376 90816
rect 88454 90604 88934 90634
rect 87316 90544 88934 90604
rect 88454 90514 88934 90544
rect 878 90130 1198 90131
rect 878 90066 886 90130
rect 950 90066 966 90130
rect 1030 90066 1046 90130
rect 1110 90066 1126 90130
rect 1190 90066 1198 90130
rect 878 90065 1198 90066
rect 84878 90130 85198 90131
rect 84878 90066 84886 90130
rect 84950 90066 84966 90130
rect 85030 90066 85046 90130
rect 85110 90066 85126 90130
rect 85190 90066 85198 90130
rect 84878 90065 85198 90066
rect 2878 89586 3198 89587
rect 2878 89522 2886 89586
rect 2950 89522 2966 89586
rect 3030 89522 3046 89586
rect 3110 89522 3126 89586
rect 3190 89522 3198 89586
rect 2878 89521 3198 89522
rect 86878 89586 87198 89587
rect 86878 89522 86886 89586
rect 86950 89522 86966 89586
rect 87030 89522 87046 89586
rect 87110 89522 87126 89586
rect 87190 89522 87198 89586
rect 86878 89521 87198 89522
rect 84139 89380 84205 89383
rect 88454 89380 88934 89410
rect 84139 89378 88934 89380
rect 84139 89322 84144 89378
rect 84200 89322 88934 89378
rect 84139 89320 88934 89322
rect 84139 89317 84205 89320
rect 88454 89290 88934 89320
rect 878 89042 1198 89043
rect 878 88978 886 89042
rect 950 88978 966 89042
rect 1030 88978 1046 89042
rect 1110 88978 1126 89042
rect 1190 88978 1198 89042
rect 878 88977 1198 88978
rect 84878 89042 85198 89043
rect 84878 88978 84886 89042
rect 84950 88978 84966 89042
rect 85030 88978 85046 89042
rect 85110 88978 85126 89042
rect 85190 88978 85198 89042
rect 84878 88977 85198 88978
rect 3731 88836 3797 88839
rect 3731 88834 3840 88836
rect 3731 88778 3736 88834
rect 3792 88778 3840 88834
rect 3731 88773 3840 88778
rect 3780 88564 3840 88773
rect 3915 88564 3981 88567
rect 3780 88562 3981 88564
rect 3780 88506 3920 88562
rect 3976 88506 3981 88562
rect 3780 88504 3981 88506
rect 3915 88501 3981 88504
rect 4099 88564 4165 88567
rect 5436 88564 5496 88742
rect 4099 88562 5496 88564
rect 4099 88506 4104 88562
rect 4160 88506 5496 88562
rect 4099 88504 5496 88506
rect 4099 88501 4165 88504
rect 2878 88498 3198 88499
rect 2878 88434 2886 88498
rect 2950 88434 2966 88498
rect 3030 88434 3046 88498
rect 3110 88434 3126 88498
rect 3190 88434 3198 88498
rect 2878 88433 3198 88434
rect 86878 88498 87198 88499
rect 86878 88434 86886 88498
rect 86950 88434 86966 88498
rect 87030 88434 87046 88498
rect 87110 88434 87126 88498
rect 87190 88434 87198 88498
rect 86878 88433 87198 88434
rect 84415 88156 84481 88159
rect 88454 88156 88934 88186
rect 84415 88154 88934 88156
rect 84415 88098 84420 88154
rect 84476 88098 88934 88154
rect 84415 88096 88934 88098
rect 84415 88093 84481 88096
rect 88454 88066 88934 88096
rect 878 87954 1198 87955
rect 878 87890 886 87954
rect 950 87890 966 87954
rect 1030 87890 1046 87954
rect 1110 87890 1126 87954
rect 1190 87890 1198 87954
rect 878 87889 1198 87890
rect 84878 87954 85198 87955
rect 84878 87890 84886 87954
rect 84950 87890 84966 87954
rect 85030 87890 85046 87954
rect 85110 87890 85126 87954
rect 85190 87890 85198 87954
rect 84878 87889 85198 87890
rect 3731 87612 3797 87615
rect 5068 87612 5128 87614
rect 3731 87610 5128 87612
rect 3731 87554 3736 87610
rect 3792 87554 5128 87610
rect 3731 87552 5128 87554
rect 3731 87549 3797 87552
rect 2878 87410 3198 87411
rect 2878 87346 2886 87410
rect 2950 87346 2966 87410
rect 3030 87346 3046 87410
rect 3110 87346 3126 87410
rect 3190 87346 3198 87410
rect 2878 87345 3198 87346
rect 86878 87410 87198 87411
rect 86878 87346 86886 87410
rect 86950 87346 86966 87410
rect 87030 87346 87046 87410
rect 87110 87346 87126 87410
rect 87190 87346 87198 87410
rect 86878 87345 87198 87346
rect 84691 87068 84757 87071
rect 84691 87066 85352 87068
rect 84691 87010 84696 87066
rect 84752 87010 85352 87066
rect 84691 87008 85352 87010
rect 84691 87005 84757 87008
rect 85292 86932 85352 87008
rect 88454 86932 88934 86962
rect 85292 86872 88934 86932
rect 878 86866 1198 86867
rect 878 86802 886 86866
rect 950 86802 966 86866
rect 1030 86802 1046 86866
rect 1110 86802 1126 86866
rect 1190 86802 1198 86866
rect 878 86801 1198 86802
rect 84878 86866 85198 86867
rect 84878 86802 84886 86866
rect 84950 86802 84966 86866
rect 85030 86802 85046 86866
rect 85110 86802 85126 86866
rect 85190 86802 85198 86866
rect 88454 86842 88934 86872
rect 84878 86801 85198 86802
rect 2878 86322 3198 86323
rect 2878 86258 2886 86322
rect 2950 86258 2966 86322
rect 3030 86258 3046 86322
rect 3110 86258 3126 86322
rect 3190 86258 3198 86322
rect 2878 86257 3198 86258
rect 86878 86322 87198 86323
rect 86878 86258 86886 86322
rect 86950 86258 86966 86322
rect 87030 86258 87046 86322
rect 87110 86258 87126 86322
rect 87190 86258 87198 86322
rect 86878 86257 87198 86258
rect 4191 85980 4257 85983
rect 84323 85980 84389 85983
rect 4191 85978 5128 85980
rect 4191 85922 4196 85978
rect 4252 85922 5128 85978
rect 4191 85920 5128 85922
rect 4191 85917 4257 85920
rect 5068 85914 5128 85920
rect 84323 85978 85720 85980
rect 84323 85922 84328 85978
rect 84384 85922 85720 85978
rect 84323 85920 85720 85922
rect 84323 85917 84389 85920
rect 878 85778 1198 85779
rect 878 85714 886 85778
rect 950 85714 966 85778
rect 1030 85714 1046 85778
rect 1110 85714 1126 85778
rect 1190 85714 1198 85778
rect 878 85713 1198 85714
rect 84878 85778 85198 85779
rect 84878 85714 84886 85778
rect 84950 85714 84966 85778
rect 85030 85714 85046 85778
rect 85110 85714 85126 85778
rect 85190 85714 85198 85778
rect 84878 85713 85198 85714
rect 85660 85708 85720 85920
rect 88454 85708 88934 85738
rect 85660 85648 88934 85708
rect 88454 85618 88934 85648
rect 2878 85234 3198 85235
rect 2878 85170 2886 85234
rect 2950 85170 2966 85234
rect 3030 85170 3046 85234
rect 3110 85170 3126 85234
rect 3190 85170 3198 85234
rect 2878 85169 3198 85170
rect 86878 85234 87198 85235
rect 86878 85170 86886 85234
rect 86950 85170 86966 85234
rect 87030 85170 87046 85234
rect 87110 85170 87126 85234
rect 87190 85170 87198 85234
rect 86878 85169 87198 85170
rect 4007 84756 4073 84759
rect 5068 84756 5128 84786
rect 4007 84754 5128 84756
rect 4007 84698 4012 84754
rect 4068 84698 5128 84754
rect 4007 84696 5128 84698
rect 4007 84693 4073 84696
rect 878 84690 1198 84691
rect 878 84626 886 84690
rect 950 84626 966 84690
rect 1030 84626 1046 84690
rect 1110 84626 1126 84690
rect 1190 84626 1198 84690
rect 878 84625 1198 84626
rect 84878 84690 85198 84691
rect 84878 84626 84886 84690
rect 84950 84626 84966 84690
rect 85030 84626 85046 84690
rect 85110 84626 85126 84690
rect 85190 84626 85198 84690
rect 84878 84625 85198 84626
rect 84231 84484 84297 84487
rect 88454 84484 88934 84514
rect 84231 84482 88934 84484
rect 84231 84426 84236 84482
rect 84292 84426 88934 84482
rect 84231 84424 88934 84426
rect 84231 84421 84297 84424
rect 88454 84394 88934 84424
rect 2878 84146 3198 84147
rect 2878 84082 2886 84146
rect 2950 84082 2966 84146
rect 3030 84082 3046 84146
rect 3110 84082 3126 84146
rect 3190 84082 3198 84146
rect 2878 84081 3198 84082
rect 86878 84146 87198 84147
rect 86878 84082 86886 84146
rect 86950 84082 86966 84146
rect 87030 84082 87046 84146
rect 87110 84082 87126 84146
rect 87190 84082 87198 84146
rect 86878 84081 87198 84082
rect 4692 83606 4698 83670
rect 4762 83606 4768 83670
rect 878 83602 1198 83603
rect 878 83538 886 83602
rect 950 83538 966 83602
rect 1030 83538 1046 83602
rect 1110 83538 1126 83602
rect 1190 83538 1198 83602
rect 878 83537 1198 83538
rect 4700 83398 4760 83606
rect 84878 83602 85198 83603
rect 84878 83538 84886 83602
rect 84950 83538 84966 83602
rect 85030 83538 85046 83602
rect 85110 83538 85126 83602
rect 85190 83538 85198 83602
rect 84878 83537 85198 83538
rect 4692 83334 4698 83398
rect 4762 83334 4768 83398
rect 84507 83396 84573 83399
rect 88454 83396 88934 83426
rect 84507 83394 88934 83396
rect 84507 83338 84512 83394
rect 84568 83338 88934 83394
rect 84507 83336 88934 83338
rect 84507 83333 84573 83336
rect 88454 83306 88934 83336
rect 3547 83124 3613 83127
rect 3547 83122 5128 83124
rect 3547 83066 3552 83122
rect 3608 83066 5128 83122
rect 3547 83064 5128 83066
rect 3547 83061 3613 83064
rect 2878 83058 3198 83059
rect 2878 82994 2886 83058
rect 2950 82994 2966 83058
rect 3030 82994 3046 83058
rect 3110 82994 3126 83058
rect 3190 82994 3198 83058
rect 2878 82993 3198 82994
rect 86878 83058 87198 83059
rect 86878 82994 86886 83058
rect 86950 82994 86966 83058
rect 87030 82994 87046 83058
rect 87110 82994 87126 83058
rect 87190 82994 87198 83058
rect 86878 82993 87198 82994
rect 878 82514 1198 82515
rect 878 82450 886 82514
rect 950 82450 966 82514
rect 1030 82450 1046 82514
rect 1110 82450 1126 82514
rect 1190 82450 1198 82514
rect 878 82449 1198 82450
rect 84878 82514 85198 82515
rect 84878 82450 84886 82514
rect 84950 82450 84966 82514
rect 85030 82450 85046 82514
rect 85110 82450 85126 82514
rect 85190 82450 85198 82514
rect 84878 82449 85198 82450
rect 84415 82172 84481 82175
rect 88454 82172 88934 82202
rect 84415 82170 88934 82172
rect 84415 82114 84420 82170
rect 84476 82114 88934 82170
rect 84415 82112 88934 82114
rect 84415 82109 84481 82112
rect 88454 82082 88934 82112
rect 3271 82036 3337 82039
rect 3271 82034 5128 82036
rect 3271 81978 3276 82034
rect 3332 81978 5128 82034
rect 3271 81976 5128 81978
rect 3271 81973 3337 81976
rect 2878 81970 3198 81971
rect 2878 81906 2886 81970
rect 2950 81906 2966 81970
rect 3030 81906 3046 81970
rect 3110 81906 3126 81970
rect 3190 81906 3198 81970
rect 5068 81958 5128 81976
rect 86878 81970 87198 81971
rect 2878 81905 3198 81906
rect 86878 81906 86886 81970
rect 86950 81906 86966 81970
rect 87030 81906 87046 81970
rect 87110 81906 87126 81970
rect 87190 81906 87198 81970
rect 86878 81905 87198 81906
rect 878 81426 1198 81427
rect 878 81362 886 81426
rect 950 81362 966 81426
rect 1030 81362 1046 81426
rect 1110 81362 1126 81426
rect 1190 81362 1198 81426
rect 878 81361 1198 81362
rect 84878 81426 85198 81427
rect 84878 81362 84886 81426
rect 84950 81362 84966 81426
rect 85030 81362 85046 81426
rect 85110 81362 85126 81426
rect 85190 81362 85198 81426
rect 84878 81361 85198 81362
rect 88454 80948 88934 80978
rect 87316 80888 88934 80948
rect 2878 80882 3198 80883
rect 2878 80818 2886 80882
rect 2950 80818 2966 80882
rect 3030 80818 3046 80882
rect 3110 80818 3126 80882
rect 3190 80818 3198 80882
rect 2878 80817 3198 80818
rect 86878 80882 87198 80883
rect 86878 80818 86886 80882
rect 86950 80818 86966 80882
rect 87030 80818 87046 80882
rect 87110 80818 87126 80882
rect 87190 80818 87198 80882
rect 86878 80817 87198 80818
rect 84783 80676 84849 80679
rect 87316 80676 87376 80888
rect 88454 80858 88934 80888
rect 84783 80674 87376 80676
rect 84783 80618 84788 80674
rect 84844 80618 87376 80674
rect 84783 80616 87376 80618
rect 84783 80613 84849 80616
rect 878 80338 1198 80339
rect 878 80274 886 80338
rect 950 80274 966 80338
rect 1030 80274 1046 80338
rect 1110 80274 1126 80338
rect 1190 80274 1198 80338
rect 878 80273 1198 80274
rect 84878 80338 85198 80339
rect 84878 80274 84886 80338
rect 84950 80274 84966 80338
rect 85030 80274 85046 80338
rect 85110 80274 85126 80338
rect 85190 80274 85198 80338
rect 84878 80273 85198 80274
rect 3639 79996 3705 79999
rect 5068 79996 5128 80258
rect 3639 79994 5128 79996
rect 3639 79938 3644 79994
rect 3700 79938 5128 79994
rect 3639 79936 5128 79938
rect 84599 79996 84665 79999
rect 84599 79994 87376 79996
rect 84599 79938 84604 79994
rect 84660 79938 87376 79994
rect 84599 79936 87376 79938
rect 3639 79933 3705 79936
rect 84599 79933 84665 79936
rect 2878 79794 3198 79795
rect 2878 79730 2886 79794
rect 2950 79730 2966 79794
rect 3030 79730 3046 79794
rect 3110 79730 3126 79794
rect 3190 79730 3198 79794
rect 2878 79729 3198 79730
rect 86878 79794 87198 79795
rect 86878 79730 86886 79794
rect 86950 79730 86966 79794
rect 87030 79730 87046 79794
rect 87110 79730 87126 79794
rect 87190 79730 87198 79794
rect 86878 79729 87198 79730
rect 87316 79724 87376 79936
rect 88454 79724 88934 79754
rect 87316 79664 88934 79724
rect 88454 79634 88934 79664
rect 878 79250 1198 79251
rect 878 79186 886 79250
rect 950 79186 966 79250
rect 1030 79186 1046 79250
rect 1110 79186 1126 79250
rect 1190 79186 1198 79250
rect 878 79185 1198 79186
rect 84878 79250 85198 79251
rect 84878 79186 84886 79250
rect 84950 79186 84966 79250
rect 85030 79186 85046 79250
rect 85110 79186 85126 79250
rect 85190 79186 85198 79250
rect 84878 79185 85198 79186
rect 2878 78706 3198 78707
rect 2878 78642 2886 78706
rect 2950 78642 2966 78706
rect 3030 78642 3046 78706
rect 3110 78642 3126 78706
rect 3190 78642 3198 78706
rect 2878 78641 3198 78642
rect 86878 78706 87198 78707
rect 86878 78642 86886 78706
rect 86950 78642 86966 78706
rect 87030 78642 87046 78706
rect 87110 78642 87126 78706
rect 87190 78642 87198 78706
rect 86878 78641 87198 78642
rect 84231 78500 84297 78503
rect 88454 78500 88934 78530
rect 84231 78498 88934 78500
rect 84231 78442 84236 78498
rect 84292 78442 88934 78498
rect 84231 78440 88934 78442
rect 84231 78437 84297 78440
rect 88454 78410 88934 78440
rect 878 78162 1198 78163
rect 878 78098 886 78162
rect 950 78098 966 78162
rect 1030 78098 1046 78162
rect 1110 78098 1126 78162
rect 1190 78098 1198 78162
rect 878 78097 1198 78098
rect 84878 78162 85198 78163
rect 84878 78098 84886 78162
rect 84950 78098 84966 78162
rect 85030 78098 85046 78162
rect 85110 78098 85126 78162
rect 85190 78098 85198 78162
rect 84878 78097 85198 78098
rect 2878 77618 3198 77619
rect 2878 77554 2886 77618
rect 2950 77554 2966 77618
rect 3030 77554 3046 77618
rect 3110 77554 3126 77618
rect 3190 77554 3198 77618
rect 2878 77553 3198 77554
rect 86878 77618 87198 77619
rect 86878 77554 86886 77618
rect 86950 77554 86966 77618
rect 87030 77554 87046 77618
rect 87110 77554 87126 77618
rect 87190 77554 87198 77618
rect 86878 77553 87198 77554
rect 84139 77276 84205 77279
rect 88454 77276 88934 77306
rect 84139 77274 88934 77276
rect 84139 77218 84144 77274
rect 84200 77218 88934 77274
rect 84139 77216 88934 77218
rect 84139 77213 84205 77216
rect 88454 77186 88934 77216
rect 878 77074 1198 77075
rect 878 77010 886 77074
rect 950 77010 966 77074
rect 1030 77010 1046 77074
rect 1110 77010 1126 77074
rect 1190 77010 1198 77074
rect 878 77009 1198 77010
rect 84878 77074 85198 77075
rect 84878 77010 84886 77074
rect 84950 77010 84966 77074
rect 85030 77010 85046 77074
rect 85110 77010 85126 77074
rect 85190 77010 85198 77074
rect 84878 77009 85198 77010
rect 2878 76530 3198 76531
rect 2878 76466 2886 76530
rect 2950 76466 2966 76530
rect 3030 76466 3046 76530
rect 3110 76466 3126 76530
rect 3190 76466 3198 76530
rect 2878 76465 3198 76466
rect 86878 76530 87198 76531
rect 86878 76466 86886 76530
rect 86950 76466 86966 76530
rect 87030 76466 87046 76530
rect 87110 76466 87126 76530
rect 87190 76466 87198 76530
rect 86878 76465 87198 76466
rect 83311 76188 83377 76191
rect 88454 76188 88934 76218
rect 83311 76186 88934 76188
rect 83311 76130 83316 76186
rect 83372 76130 88934 76186
rect 83311 76128 88934 76130
rect 83311 76125 83377 76128
rect 88454 76098 88934 76128
rect 878 75986 1198 75987
rect 878 75922 886 75986
rect 950 75922 966 75986
rect 1030 75922 1046 75986
rect 1110 75922 1126 75986
rect 1190 75922 1198 75986
rect 878 75921 1198 75922
rect 84878 75986 85198 75987
rect 84878 75922 84886 75986
rect 84950 75922 84966 75986
rect 85030 75922 85046 75986
rect 85110 75922 85126 75986
rect 85190 75922 85198 75986
rect 84878 75921 85198 75922
rect 2878 75442 3198 75443
rect 2878 75378 2886 75442
rect 2950 75378 2966 75442
rect 3030 75378 3046 75442
rect 3110 75378 3126 75442
rect 3190 75378 3198 75442
rect 2878 75377 3198 75378
rect 86878 75442 87198 75443
rect 86878 75378 86886 75442
rect 86950 75378 86966 75442
rect 87030 75378 87046 75442
rect 87110 75378 87126 75442
rect 87190 75378 87198 75442
rect 86878 75377 87198 75378
rect 84783 75100 84849 75103
rect 84783 75098 85352 75100
rect 84783 75042 84788 75098
rect 84844 75042 85352 75098
rect 84783 75040 85352 75042
rect 84783 75037 84849 75040
rect 85292 74964 85352 75040
rect 88454 74964 88934 74994
rect 85292 74904 88934 74964
rect 878 74898 1198 74899
rect 878 74834 886 74898
rect 950 74834 966 74898
rect 1030 74834 1046 74898
rect 1110 74834 1126 74898
rect 1190 74834 1198 74898
rect 878 74833 1198 74834
rect 84878 74898 85198 74899
rect 84878 74834 84886 74898
rect 84950 74834 84966 74898
rect 85030 74834 85046 74898
rect 85110 74834 85126 74898
rect 85190 74834 85198 74898
rect 88454 74874 88934 74904
rect 84878 74833 85198 74834
rect 4692 74692 4698 74694
rect 4516 74632 4698 74692
rect 4516 74422 4576 74632
rect 4692 74630 4698 74632
rect 4762 74630 4768 74694
rect 4508 74358 4514 74422
rect 4578 74358 4584 74422
rect 2878 74354 3198 74355
rect 2878 74290 2886 74354
rect 2950 74290 2966 74354
rect 3030 74290 3046 74354
rect 3110 74290 3126 74354
rect 3190 74290 3198 74354
rect 2878 74289 3198 74290
rect 86878 74354 87198 74355
rect 86878 74290 86886 74354
rect 86950 74290 86966 74354
rect 87030 74290 87046 74354
rect 87110 74290 87126 74354
rect 87190 74290 87198 74354
rect 86878 74289 87198 74290
rect 84875 74012 84941 74015
rect 84875 74010 85352 74012
rect 84875 73954 84880 74010
rect 84936 73954 85352 74010
rect 84875 73952 85352 73954
rect 84875 73949 84941 73952
rect 878 73810 1198 73811
rect 878 73746 886 73810
rect 950 73746 966 73810
rect 1030 73746 1046 73810
rect 1110 73746 1126 73810
rect 1190 73746 1198 73810
rect 878 73745 1198 73746
rect 84878 73810 85198 73811
rect 84878 73746 84886 73810
rect 84950 73746 84966 73810
rect 85030 73746 85046 73810
rect 85110 73746 85126 73810
rect 85190 73746 85198 73810
rect 84878 73745 85198 73746
rect 85292 73740 85352 73952
rect 88454 73740 88934 73770
rect 85292 73680 88934 73740
rect 88454 73650 88934 73680
rect 2878 73266 3198 73267
rect 2878 73202 2886 73266
rect 2950 73202 2966 73266
rect 3030 73202 3046 73266
rect 3110 73202 3126 73266
rect 3190 73202 3198 73266
rect 2878 73201 3198 73202
rect 86878 73266 87198 73267
rect 86878 73202 86886 73266
rect 86950 73202 86966 73266
rect 87030 73202 87046 73266
rect 87110 73202 87126 73266
rect 87190 73202 87198 73266
rect 86878 73201 87198 73202
rect 878 72722 1198 72723
rect 878 72658 886 72722
rect 950 72658 966 72722
rect 1030 72658 1046 72722
rect 1110 72658 1126 72722
rect 1190 72658 1198 72722
rect 878 72657 1198 72658
rect 84878 72722 85198 72723
rect 84878 72658 84886 72722
rect 84950 72658 84966 72722
rect 85030 72658 85046 72722
rect 85110 72658 85126 72722
rect 85190 72658 85198 72722
rect 84878 72657 85198 72658
rect 84691 72516 84757 72519
rect 88454 72516 88934 72546
rect 84691 72514 88934 72516
rect 84691 72458 84696 72514
rect 84752 72458 88934 72514
rect 84691 72456 88934 72458
rect 84691 72453 84757 72456
rect 88454 72426 88934 72456
rect 2878 72178 3198 72179
rect 2878 72114 2886 72178
rect 2950 72114 2966 72178
rect 3030 72114 3046 72178
rect 3110 72114 3126 72178
rect 3190 72114 3198 72178
rect 2878 72113 3198 72114
rect 86878 72178 87198 72179
rect 86878 72114 86886 72178
rect 86950 72114 86966 72178
rect 87030 72114 87046 72178
rect 87110 72114 87126 72178
rect 87190 72114 87198 72178
rect 86878 72113 87198 72114
rect 878 71634 1198 71635
rect 878 71570 886 71634
rect 950 71570 966 71634
rect 1030 71570 1046 71634
rect 1110 71570 1126 71634
rect 1190 71570 1198 71634
rect 878 71569 1198 71570
rect 84878 71634 85198 71635
rect 84878 71570 84886 71634
rect 84950 71570 84966 71634
rect 85030 71570 85046 71634
rect 85110 71570 85126 71634
rect 85190 71570 85198 71634
rect 84878 71569 85198 71570
rect 84599 71292 84665 71295
rect 88454 71292 88934 71322
rect 84599 71290 88934 71292
rect 84599 71234 84604 71290
rect 84660 71234 88934 71290
rect 84599 71232 88934 71234
rect 84599 71229 84665 71232
rect 88454 71202 88934 71232
rect 2878 71090 3198 71091
rect 2878 71026 2886 71090
rect 2950 71026 2966 71090
rect 3030 71026 3046 71090
rect 3110 71026 3126 71090
rect 3190 71026 3198 71090
rect 2878 71025 3198 71026
rect 86878 71090 87198 71091
rect 86878 71026 86886 71090
rect 86950 71026 86966 71090
rect 87030 71026 87046 71090
rect 87110 71026 87126 71090
rect 87190 71026 87198 71090
rect 86878 71025 87198 71026
rect 878 70546 1198 70547
rect 878 70482 886 70546
rect 950 70482 966 70546
rect 1030 70482 1046 70546
rect 1110 70482 1126 70546
rect 1190 70482 1198 70546
rect 878 70481 1198 70482
rect 84878 70546 85198 70547
rect 84878 70482 84886 70546
rect 84950 70482 84966 70546
rect 85030 70482 85046 70546
rect 85110 70482 85126 70546
rect 85190 70482 85198 70546
rect 84878 70481 85198 70482
rect 84323 70204 84389 70207
rect 84323 70202 87376 70204
rect 84323 70146 84328 70202
rect 84384 70146 87376 70202
rect 84323 70144 87376 70146
rect 84323 70141 84389 70144
rect 87316 70068 87376 70144
rect 88454 70068 88934 70098
rect 87316 70008 88934 70068
rect 2878 70002 3198 70003
rect 2878 69938 2886 70002
rect 2950 69938 2966 70002
rect 3030 69938 3046 70002
rect 3110 69938 3126 70002
rect 3190 69938 3198 70002
rect 2878 69937 3198 69938
rect 86878 70002 87198 70003
rect 86878 69938 86886 70002
rect 86950 69938 86966 70002
rect 87030 69938 87046 70002
rect 87110 69938 87126 70002
rect 87190 69938 87198 70002
rect 88454 69978 88934 70008
rect 86878 69937 87198 69938
rect 878 69458 1198 69459
rect 878 69394 886 69458
rect 950 69394 966 69458
rect 1030 69394 1046 69458
rect 1110 69394 1126 69458
rect 1190 69394 1198 69458
rect 878 69393 1198 69394
rect 84878 69458 85198 69459
rect 84878 69394 84886 69458
rect 84950 69394 84966 69458
rect 85030 69394 85046 69458
rect 85110 69394 85126 69458
rect 85190 69394 85198 69458
rect 84878 69393 85198 69394
rect 84415 69116 84481 69119
rect 84415 69114 87376 69116
rect 84415 69058 84420 69114
rect 84476 69058 87376 69114
rect 84415 69056 87376 69058
rect 84415 69053 84481 69056
rect 2878 68914 3198 68915
rect 2878 68850 2886 68914
rect 2950 68850 2966 68914
rect 3030 68850 3046 68914
rect 3110 68850 3126 68914
rect 3190 68850 3198 68914
rect 2878 68849 3198 68850
rect 86878 68914 87198 68915
rect 86878 68850 86886 68914
rect 86950 68850 86966 68914
rect 87030 68850 87046 68914
rect 87110 68850 87126 68914
rect 87190 68850 87198 68914
rect 86878 68849 87198 68850
rect 87316 68844 87376 69056
rect 88454 68844 88934 68874
rect 87316 68784 88934 68844
rect 88454 68754 88934 68784
rect 878 68370 1198 68371
rect 878 68306 886 68370
rect 950 68306 966 68370
rect 1030 68306 1046 68370
rect 1110 68306 1126 68370
rect 1190 68306 1198 68370
rect 878 68305 1198 68306
rect 84878 68370 85198 68371
rect 84878 68306 84886 68370
rect 84950 68306 84966 68370
rect 85030 68306 85046 68370
rect 85110 68306 85126 68370
rect 85190 68306 85198 68370
rect 84878 68305 85198 68306
rect 84783 68028 84849 68031
rect 84783 68026 87376 68028
rect 84783 67970 84788 68026
rect 84844 67970 87376 68026
rect 84783 67968 87376 67970
rect 84783 67965 84849 67968
rect 2878 67826 3198 67827
rect 2878 67762 2886 67826
rect 2950 67762 2966 67826
rect 3030 67762 3046 67826
rect 3110 67762 3126 67826
rect 3190 67762 3198 67826
rect 2878 67761 3198 67762
rect 86878 67826 87198 67827
rect 86878 67762 86886 67826
rect 86950 67762 86966 67826
rect 87030 67762 87046 67826
rect 87110 67762 87126 67826
rect 87190 67762 87198 67826
rect 86878 67761 87198 67762
rect 87316 67756 87376 67968
rect 88454 67756 88934 67786
rect 87316 67696 88934 67756
rect 88454 67666 88934 67696
rect 878 67282 1198 67283
rect 878 67218 886 67282
rect 950 67218 966 67282
rect 1030 67218 1046 67282
rect 1110 67218 1126 67282
rect 1190 67218 1198 67282
rect 878 67217 1198 67218
rect 84878 67282 85198 67283
rect 84878 67218 84886 67282
rect 84950 67218 84966 67282
rect 85030 67218 85046 67282
rect 85110 67218 85126 67282
rect 85190 67218 85198 67282
rect 84878 67217 85198 67218
rect 2878 66738 3198 66739
rect 2878 66674 2886 66738
rect 2950 66674 2966 66738
rect 3030 66674 3046 66738
rect 3110 66674 3126 66738
rect 3190 66674 3198 66738
rect 2878 66673 3198 66674
rect 86878 66738 87198 66739
rect 86878 66674 86886 66738
rect 86950 66674 86966 66738
rect 87030 66674 87046 66738
rect 87110 66674 87126 66738
rect 87190 66674 87198 66738
rect 86878 66673 87198 66674
rect 85151 66532 85217 66535
rect 88454 66532 88934 66562
rect 85151 66530 88934 66532
rect 85151 66474 85156 66530
rect 85212 66474 88934 66530
rect 85151 66472 88934 66474
rect 85151 66469 85217 66472
rect 88454 66442 88934 66472
rect 878 66194 1198 66195
rect 878 66130 886 66194
rect 950 66130 966 66194
rect 1030 66130 1046 66194
rect 1110 66130 1126 66194
rect 1190 66130 1198 66194
rect 878 66129 1198 66130
rect 84878 66194 85198 66195
rect 84878 66130 84886 66194
rect 84950 66130 84966 66194
rect 85030 66130 85046 66194
rect 85110 66130 85126 66194
rect 85190 66130 85198 66194
rect 84878 66129 85198 66130
rect 2878 65650 3198 65651
rect 2878 65586 2886 65650
rect 2950 65586 2966 65650
rect 3030 65586 3046 65650
rect 3110 65586 3126 65650
rect 3190 65586 3198 65650
rect 2878 65585 3198 65586
rect 86878 65650 87198 65651
rect 86878 65586 86886 65650
rect 86950 65586 86966 65650
rect 87030 65586 87046 65650
rect 87110 65586 87126 65650
rect 87190 65586 87198 65650
rect 86878 65585 87198 65586
rect 4508 65518 4514 65582
rect 4578 65518 4584 65582
rect 4516 65308 4576 65518
rect 4692 65308 4698 65310
rect 4516 65248 4698 65308
rect 4692 65246 4698 65248
rect 4762 65246 4768 65310
rect 84599 65308 84665 65311
rect 88454 65308 88934 65338
rect 84599 65306 88934 65308
rect 84599 65250 84604 65306
rect 84660 65250 88934 65306
rect 84599 65248 88934 65250
rect 84599 65245 84665 65248
rect 88454 65218 88934 65248
rect 878 65106 1198 65107
rect 878 65042 886 65106
rect 950 65042 966 65106
rect 1030 65042 1046 65106
rect 1110 65042 1126 65106
rect 1190 65042 1198 65106
rect 878 65041 1198 65042
rect 84878 65106 85198 65107
rect 84878 65042 84886 65106
rect 84950 65042 84966 65106
rect 85030 65042 85046 65106
rect 85110 65042 85126 65106
rect 85190 65042 85198 65106
rect 84878 65041 85198 65042
rect 2878 64562 3198 64563
rect 2878 64498 2886 64562
rect 2950 64498 2966 64562
rect 3030 64498 3046 64562
rect 3110 64498 3126 64562
rect 3190 64498 3198 64562
rect 2878 64497 3198 64498
rect 86878 64562 87198 64563
rect 86878 64498 86886 64562
rect 86950 64498 86966 64562
rect 87030 64498 87046 64562
rect 87110 64498 87126 64562
rect 87190 64498 87198 64562
rect 86878 64497 87198 64498
rect 88454 64084 88934 64114
rect 85844 64024 88934 64084
rect 878 64018 1198 64019
rect 878 63954 886 64018
rect 950 63954 966 64018
rect 1030 63954 1046 64018
rect 1110 63954 1126 64018
rect 1190 63954 1198 64018
rect 878 63953 1198 63954
rect 84878 64018 85198 64019
rect 84878 63954 84886 64018
rect 84950 63954 84966 64018
rect 85030 63954 85046 64018
rect 85110 63954 85126 64018
rect 85190 63954 85198 64018
rect 84878 63953 85198 63954
rect 84691 63812 84757 63815
rect 85844 63812 85904 64024
rect 88454 63994 88934 64024
rect 84691 63810 85904 63812
rect 84691 63754 84696 63810
rect 84752 63754 85904 63810
rect 84691 63752 85904 63754
rect 84691 63749 84757 63752
rect 2878 63474 3198 63475
rect 2878 63410 2886 63474
rect 2950 63410 2966 63474
rect 3030 63410 3046 63474
rect 3110 63410 3126 63474
rect 3190 63410 3198 63474
rect 2878 63409 3198 63410
rect 86878 63474 87198 63475
rect 86878 63410 86886 63474
rect 86950 63410 86966 63474
rect 87030 63410 87046 63474
rect 87110 63410 87126 63474
rect 87190 63410 87198 63474
rect 86878 63409 87198 63410
rect 3823 63132 3889 63135
rect 83127 63132 83193 63135
rect 3780 63130 3889 63132
rect 3780 63074 3828 63130
rect 3884 63074 3889 63130
rect 3780 63069 3889 63074
rect 83084 63130 83193 63132
rect 83084 63074 83132 63130
rect 83188 63074 83193 63130
rect 83084 63069 83193 63074
rect 3780 62999 3840 63069
rect 3731 62994 3840 62999
rect 3731 62938 3736 62994
rect 3792 62938 3840 62994
rect 3731 62936 3840 62938
rect 83084 62999 83144 63069
rect 83084 62994 83193 62999
rect 83084 62938 83132 62994
rect 83188 62938 83193 62994
rect 83084 62936 83193 62938
rect 3731 62933 3797 62936
rect 83127 62933 83193 62936
rect 878 62930 1198 62931
rect 878 62866 886 62930
rect 950 62866 966 62930
rect 1030 62866 1046 62930
rect 1110 62866 1126 62930
rect 1190 62866 1198 62930
rect 878 62865 1198 62866
rect 84878 62930 85198 62931
rect 84878 62866 84886 62930
rect 84950 62866 84966 62930
rect 85030 62866 85046 62930
rect 85110 62866 85126 62930
rect 85190 62866 85198 62930
rect 84878 62865 85198 62866
rect 88454 62860 88934 62890
rect 85292 62800 88934 62860
rect 84783 62724 84849 62727
rect 85292 62724 85352 62800
rect 88454 62770 88934 62800
rect 84783 62722 85352 62724
rect 84783 62666 84788 62722
rect 84844 62666 85352 62722
rect 84783 62664 85352 62666
rect 84783 62661 84849 62664
rect 2878 62386 3198 62387
rect 2878 62322 2886 62386
rect 2950 62322 2966 62386
rect 3030 62322 3046 62386
rect 3110 62322 3126 62386
rect 3190 62322 3198 62386
rect 2878 62321 3198 62322
rect 86878 62386 87198 62387
rect 86878 62322 86886 62386
rect 86950 62322 86966 62386
rect 87030 62322 87046 62386
rect 87110 62322 87126 62386
rect 87190 62322 87198 62386
rect 86878 62321 87198 62322
rect 878 61842 1198 61843
rect 878 61778 886 61842
rect 950 61778 966 61842
rect 1030 61778 1046 61842
rect 1110 61778 1126 61842
rect 1190 61778 1198 61842
rect 878 61777 1198 61778
rect 84878 61842 85198 61843
rect 84878 61778 84886 61842
rect 84950 61778 84966 61842
rect 85030 61778 85046 61842
rect 85110 61778 85126 61842
rect 85190 61778 85198 61842
rect 84878 61777 85198 61778
rect 83311 61636 83377 61639
rect 88454 61636 88934 61666
rect 83311 61634 88934 61636
rect 83311 61578 83316 61634
rect 83372 61578 88934 61634
rect 83311 61576 88934 61578
rect 83311 61573 83377 61576
rect 88454 61546 88934 61576
rect 2878 61298 3198 61299
rect 2878 61234 2886 61298
rect 2950 61234 2966 61298
rect 3030 61234 3046 61298
rect 3110 61234 3126 61298
rect 3190 61234 3198 61298
rect 2878 61233 3198 61234
rect 86878 61298 87198 61299
rect 86878 61234 86886 61298
rect 86950 61234 86966 61298
rect 87030 61234 87046 61298
rect 87110 61234 87126 61298
rect 87190 61234 87198 61298
rect 86878 61233 87198 61234
rect 878 60754 1198 60755
rect 878 60690 886 60754
rect 950 60690 966 60754
rect 1030 60690 1046 60754
rect 1110 60690 1126 60754
rect 1190 60690 1198 60754
rect 878 60689 1198 60690
rect 84878 60754 85198 60755
rect 84878 60690 84886 60754
rect 84950 60690 84966 60754
rect 85030 60690 85046 60754
rect 85110 60690 85126 60754
rect 85190 60690 85198 60754
rect 84878 60689 85198 60690
rect 84047 60548 84113 60551
rect 88454 60548 88934 60578
rect 84047 60546 88934 60548
rect 84047 60490 84052 60546
rect 84108 60490 88934 60546
rect 84047 60488 88934 60490
rect 84047 60485 84113 60488
rect 88454 60458 88934 60488
rect 2878 60210 3198 60211
rect 2878 60146 2886 60210
rect 2950 60146 2966 60210
rect 3030 60146 3046 60210
rect 3110 60146 3126 60210
rect 3190 60146 3198 60210
rect 2878 60145 3198 60146
rect 86878 60210 87198 60211
rect 86878 60146 86886 60210
rect 86950 60146 86966 60210
rect 87030 60146 87046 60210
rect 87110 60146 87126 60210
rect 87190 60146 87198 60210
rect 86878 60145 87198 60146
rect 878 59666 1198 59667
rect 878 59602 886 59666
rect 950 59602 966 59666
rect 1030 59602 1046 59666
rect 1110 59602 1126 59666
rect 1190 59602 1198 59666
rect 878 59601 1198 59602
rect 84878 59666 85198 59667
rect 84878 59602 84886 59666
rect 84950 59602 84966 59666
rect 85030 59602 85046 59666
rect 85110 59602 85126 59666
rect 85190 59602 85198 59666
rect 84878 59601 85198 59602
rect 83260 59262 83266 59326
rect 83330 59324 83336 59326
rect 88454 59324 88934 59354
rect 83330 59264 88934 59324
rect 83330 59262 83336 59264
rect 88454 59234 88934 59264
rect 2878 59122 3198 59123
rect 2878 59058 2886 59122
rect 2950 59058 2966 59122
rect 3030 59058 3046 59122
rect 3110 59058 3126 59122
rect 3190 59058 3198 59122
rect 2878 59057 3198 59058
rect 86878 59122 87198 59123
rect 86878 59058 86886 59122
rect 86950 59058 86966 59122
rect 87030 59058 87046 59122
rect 87110 59058 87126 59122
rect 87190 59058 87198 59122
rect 86878 59057 87198 59058
rect 878 58578 1198 58579
rect 878 58514 886 58578
rect 950 58514 966 58578
rect 1030 58514 1046 58578
rect 1110 58514 1126 58578
rect 1190 58514 1198 58578
rect 878 58513 1198 58514
rect 84878 58578 85198 58579
rect 84878 58514 84886 58578
rect 84950 58514 84966 58578
rect 85030 58514 85046 58578
rect 85110 58514 85126 58578
rect 85190 58514 85198 58578
rect 84878 58513 85198 58514
rect 88454 58100 88934 58130
rect 87316 58040 88934 58100
rect 2878 58034 3198 58035
rect 2878 57970 2886 58034
rect 2950 57970 2966 58034
rect 3030 57970 3046 58034
rect 3110 57970 3126 58034
rect 3190 57970 3198 58034
rect 2878 57969 3198 57970
rect 86878 58034 87198 58035
rect 86878 57970 86886 58034
rect 86950 57970 86966 58034
rect 87030 57970 87046 58034
rect 87110 57970 87126 58034
rect 87190 57970 87198 58034
rect 86878 57969 87198 57970
rect 84548 57766 84554 57830
rect 84618 57828 84624 57830
rect 87316 57828 87376 58040
rect 88454 58010 88934 58040
rect 84618 57768 87376 57828
rect 84618 57766 84624 57768
rect 878 57490 1198 57491
rect 878 57426 886 57490
rect 950 57426 966 57490
rect 1030 57426 1046 57490
rect 1110 57426 1126 57490
rect 1190 57426 1198 57490
rect 878 57425 1198 57426
rect 84878 57490 85198 57491
rect 84878 57426 84886 57490
rect 84950 57426 84966 57490
rect 85030 57426 85046 57490
rect 85110 57426 85126 57490
rect 85190 57426 85198 57490
rect 84878 57425 85198 57426
rect 2878 56946 3198 56947
rect 2878 56882 2886 56946
rect 2950 56882 2966 56946
rect 3030 56882 3046 56946
rect 3110 56882 3126 56946
rect 3190 56882 3198 56946
rect 2878 56881 3198 56882
rect 86878 56946 87198 56947
rect 86878 56882 86886 56946
rect 86950 56882 86966 56946
rect 87030 56882 87046 56946
rect 87110 56882 87126 56946
rect 87190 56882 87198 56946
rect 86878 56881 87198 56882
rect 88454 56876 88934 56906
rect 87316 56816 88934 56876
rect 84783 56740 84849 56743
rect 87316 56740 87376 56816
rect 88454 56786 88934 56816
rect 84783 56738 87376 56740
rect 84783 56682 84788 56738
rect 84844 56682 87376 56738
rect 84783 56680 87376 56682
rect 84783 56677 84849 56680
rect 878 56402 1198 56403
rect 878 56338 886 56402
rect 950 56338 966 56402
rect 1030 56338 1046 56402
rect 1110 56338 1126 56402
rect 1190 56338 1198 56402
rect 878 56337 1198 56338
rect 84878 56402 85198 56403
rect 84878 56338 84886 56402
rect 84950 56338 84966 56402
rect 85030 56338 85046 56402
rect 85110 56338 85126 56402
rect 85190 56338 85198 56402
rect 84878 56337 85198 56338
rect 2878 55858 3198 55859
rect 2878 55794 2886 55858
rect 2950 55794 2966 55858
rect 3030 55794 3046 55858
rect 3110 55794 3126 55858
rect 3190 55794 3198 55858
rect 2878 55793 3198 55794
rect 86878 55858 87198 55859
rect 86878 55794 86886 55858
rect 86950 55794 86966 55858
rect 87030 55794 87046 55858
rect 87110 55794 87126 55858
rect 87190 55794 87198 55858
rect 86878 55793 87198 55794
rect 84415 55652 84481 55655
rect 88454 55652 88934 55682
rect 84415 55650 88934 55652
rect 84415 55594 84420 55650
rect 84476 55594 88934 55650
rect 84415 55592 88934 55594
rect 84415 55589 84481 55592
rect 88454 55562 88934 55592
rect 878 55314 1198 55315
rect 878 55250 886 55314
rect 950 55250 966 55314
rect 1030 55250 1046 55314
rect 1110 55250 1126 55314
rect 1190 55250 1198 55314
rect 878 55249 1198 55250
rect 84878 55314 85198 55315
rect 84878 55250 84886 55314
rect 84950 55250 84966 55314
rect 85030 55250 85046 55314
rect 85110 55250 85126 55314
rect 85190 55250 85198 55314
rect 84878 55249 85198 55250
rect 83444 55182 83450 55246
rect 83514 55244 83520 55246
rect 84047 55244 84113 55247
rect 83514 55242 84113 55244
rect 83514 55186 84052 55242
rect 84108 55186 84113 55242
rect 83514 55184 84113 55186
rect 83514 55182 83520 55184
rect 84047 55181 84113 55184
rect 2878 54770 3198 54771
rect 2878 54706 2886 54770
rect 2950 54706 2966 54770
rect 3030 54706 3046 54770
rect 3110 54706 3126 54770
rect 3190 54706 3198 54770
rect 2878 54705 3198 54706
rect 86878 54770 87198 54771
rect 86878 54706 86886 54770
rect 86950 54706 86966 54770
rect 87030 54706 87046 54770
rect 87110 54706 87126 54770
rect 87190 54706 87198 54770
rect 86878 54705 87198 54706
rect 84507 54428 84573 54431
rect 88454 54428 88934 54458
rect 84507 54426 88934 54428
rect 84507 54370 84512 54426
rect 84568 54370 88934 54426
rect 84507 54368 88934 54370
rect 84507 54365 84573 54368
rect 88454 54338 88934 54368
rect 878 54226 1198 54227
rect 878 54162 886 54226
rect 950 54162 966 54226
rect 1030 54162 1046 54226
rect 1110 54162 1126 54226
rect 1190 54162 1198 54226
rect 878 54161 1198 54162
rect 84878 54226 85198 54227
rect 84878 54162 84886 54226
rect 84950 54162 84966 54226
rect 85030 54162 85046 54226
rect 85110 54162 85126 54226
rect 85190 54162 85198 54226
rect 84878 54161 85198 54162
rect 2878 53682 3198 53683
rect 2878 53618 2886 53682
rect 2950 53618 2966 53682
rect 3030 53618 3046 53682
rect 3110 53618 3126 53682
rect 3190 53618 3198 53682
rect 2878 53617 3198 53618
rect 86878 53682 87198 53683
rect 86878 53618 86886 53682
rect 86950 53618 86966 53682
rect 87030 53618 87046 53682
rect 87110 53618 87126 53682
rect 87190 53618 87198 53682
rect 86878 53617 87198 53618
rect 83403 53340 83469 53343
rect 88454 53340 88934 53370
rect 83403 53338 88934 53340
rect 83403 53282 83408 53338
rect 83464 53282 88934 53338
rect 83403 53280 88934 53282
rect 83403 53277 83469 53280
rect 88454 53250 88934 53280
rect 878 53138 1198 53139
rect 878 53074 886 53138
rect 950 53074 966 53138
rect 1030 53074 1046 53138
rect 1110 53074 1126 53138
rect 1190 53074 1198 53138
rect 878 53073 1198 53074
rect 84878 53138 85198 53139
rect 84878 53074 84886 53138
rect 84950 53074 84966 53138
rect 85030 53074 85046 53138
rect 85110 53074 85126 53138
rect 85190 53074 85198 53138
rect 84878 53073 85198 53074
rect 2878 52594 3198 52595
rect 2878 52530 2886 52594
rect 2950 52530 2966 52594
rect 3030 52530 3046 52594
rect 3110 52530 3126 52594
rect 3190 52530 3198 52594
rect 2878 52529 3198 52530
rect 86878 52594 87198 52595
rect 86878 52530 86886 52594
rect 86950 52530 86966 52594
rect 87030 52530 87046 52594
rect 87110 52530 87126 52594
rect 87190 52530 87198 52594
rect 86878 52529 87198 52530
rect 88454 52116 88934 52146
rect 85292 52056 88934 52116
rect 878 52050 1198 52051
rect 878 51986 886 52050
rect 950 51986 966 52050
rect 1030 51986 1046 52050
rect 1110 51986 1126 52050
rect 1190 51986 1198 52050
rect 878 51985 1198 51986
rect 84878 52050 85198 52051
rect 84878 51986 84886 52050
rect 84950 51986 84966 52050
rect 85030 51986 85046 52050
rect 85110 51986 85126 52050
rect 85190 51986 85198 52050
rect 84878 51985 85198 51986
rect 83587 51844 83653 51847
rect 85292 51844 85352 52056
rect 88454 52026 88934 52056
rect 83587 51842 85352 51844
rect 83587 51786 83592 51842
rect 83648 51786 85352 51842
rect 83587 51784 85352 51786
rect 83587 51781 83653 51784
rect 2878 51506 3198 51507
rect 2878 51442 2886 51506
rect 2950 51442 2966 51506
rect 3030 51442 3046 51506
rect 3110 51442 3126 51506
rect 3190 51442 3198 51506
rect 2878 51441 3198 51442
rect 86878 51506 87198 51507
rect 86878 51442 86886 51506
rect 86950 51442 86966 51506
rect 87030 51442 87046 51506
rect 87110 51442 87126 51506
rect 87190 51442 87198 51506
rect 86878 51441 87198 51442
rect 878 50962 1198 50963
rect 878 50898 886 50962
rect 950 50898 966 50962
rect 1030 50898 1046 50962
rect 1110 50898 1126 50962
rect 1190 50898 1198 50962
rect 878 50897 1198 50898
rect 84878 50962 85198 50963
rect 84878 50898 84886 50962
rect 84950 50898 84966 50962
rect 85030 50898 85046 50962
rect 85110 50898 85126 50962
rect 85190 50898 85198 50962
rect 84878 50897 85198 50898
rect 88454 50892 88934 50922
rect 85292 50832 88934 50892
rect 85151 50756 85217 50759
rect 85292 50756 85352 50832
rect 88454 50802 88934 50832
rect 85151 50754 85352 50756
rect 85151 50698 85156 50754
rect 85212 50698 85352 50754
rect 85151 50696 85352 50698
rect 85151 50693 85217 50696
rect 2878 50418 3198 50419
rect 2878 50354 2886 50418
rect 2950 50354 2966 50418
rect 3030 50354 3046 50418
rect 3110 50354 3126 50418
rect 3190 50354 3198 50418
rect 2878 50353 3198 50354
rect 86878 50418 87198 50419
rect 86878 50354 86886 50418
rect 86950 50354 86966 50418
rect 87030 50354 87046 50418
rect 87110 50354 87126 50418
rect 87190 50354 87198 50418
rect 86878 50353 87198 50354
rect 878 49874 1198 49875
rect 878 49810 886 49874
rect 950 49810 966 49874
rect 1030 49810 1046 49874
rect 1110 49810 1126 49874
rect 1190 49810 1198 49874
rect 878 49809 1198 49810
rect 84878 49874 85198 49875
rect 84878 49810 84886 49874
rect 84950 49810 84966 49874
rect 85030 49810 85046 49874
rect 85110 49810 85126 49874
rect 85190 49810 85198 49874
rect 84878 49809 85198 49810
rect 84783 49668 84849 49671
rect 88454 49668 88934 49698
rect 84783 49666 88934 49668
rect 84783 49610 84788 49666
rect 84844 49610 88934 49666
rect 84783 49608 88934 49610
rect 84783 49605 84849 49608
rect 88454 49578 88934 49608
rect 2878 49330 3198 49331
rect 2878 49266 2886 49330
rect 2950 49266 2966 49330
rect 3030 49266 3046 49330
rect 3110 49266 3126 49330
rect 3190 49266 3198 49330
rect 2878 49265 3198 49266
rect 86878 49330 87198 49331
rect 86878 49266 86886 49330
rect 86950 49266 86966 49330
rect 87030 49266 87046 49330
rect 87110 49266 87126 49330
rect 87190 49266 87198 49330
rect 86878 49265 87198 49266
rect 878 48786 1198 48787
rect 878 48722 886 48786
rect 950 48722 966 48786
rect 1030 48722 1046 48786
rect 1110 48722 1126 48786
rect 1190 48722 1198 48786
rect 878 48721 1198 48722
rect 84878 48786 85198 48787
rect 84878 48722 84886 48786
rect 84950 48722 84966 48786
rect 85030 48722 85046 48786
rect 85110 48722 85126 48786
rect 85190 48722 85198 48786
rect 84878 48721 85198 48722
rect 85795 48444 85861 48447
rect 88454 48444 88934 48474
rect 85795 48442 88934 48444
rect 85795 48386 85800 48442
rect 85856 48386 88934 48442
rect 85795 48384 88934 48386
rect 85795 48381 85861 48384
rect 88454 48354 88934 48384
rect 2878 48242 3198 48243
rect 2878 48178 2886 48242
rect 2950 48178 2966 48242
rect 3030 48178 3046 48242
rect 3110 48178 3126 48242
rect 3190 48178 3198 48242
rect 2878 48177 3198 48178
rect 86878 48242 87198 48243
rect 86878 48178 86886 48242
rect 86950 48178 86966 48242
rect 87030 48178 87046 48242
rect 87110 48178 87126 48242
rect 87190 48178 87198 48242
rect 86878 48177 87198 48178
rect 878 47698 1198 47699
rect 878 47634 886 47698
rect 950 47634 966 47698
rect 1030 47634 1046 47698
rect 1110 47634 1126 47698
rect 1190 47634 1198 47698
rect 878 47633 1198 47634
rect 84878 47698 85198 47699
rect 84878 47634 84886 47698
rect 84950 47634 84966 47698
rect 85030 47634 85046 47698
rect 85110 47634 85126 47698
rect 85190 47634 85198 47698
rect 84878 47633 85198 47634
rect 88454 47220 88934 47250
rect 87316 47160 88934 47220
rect 2878 47154 3198 47155
rect 2878 47090 2886 47154
rect 2950 47090 2966 47154
rect 3030 47090 3046 47154
rect 3110 47090 3126 47154
rect 3190 47090 3198 47154
rect 2878 47089 3198 47090
rect 86878 47154 87198 47155
rect 86878 47090 86886 47154
rect 86950 47090 86966 47154
rect 87030 47090 87046 47154
rect 87110 47090 87126 47154
rect 87190 47090 87198 47154
rect 86878 47089 87198 47090
rect 83863 46948 83929 46951
rect 87316 46948 87376 47160
rect 88454 47130 88934 47160
rect 83863 46946 87376 46948
rect 83863 46890 83868 46946
rect 83924 46890 87376 46946
rect 83863 46888 87376 46890
rect 83863 46885 83929 46888
rect 878 46610 1198 46611
rect 878 46546 886 46610
rect 950 46546 966 46610
rect 1030 46546 1046 46610
rect 1110 46546 1126 46610
rect 1190 46546 1198 46610
rect 878 46545 1198 46546
rect 84878 46610 85198 46611
rect 84878 46546 84886 46610
rect 84950 46546 84966 46610
rect 85030 46546 85046 46610
rect 85110 46546 85126 46610
rect 85190 46546 85198 46610
rect 84878 46545 85198 46546
rect 2878 46066 3198 46067
rect 2878 46002 2886 46066
rect 2950 46002 2966 46066
rect 3030 46002 3046 46066
rect 3110 46002 3126 46066
rect 3190 46002 3198 46066
rect 2878 46001 3198 46002
rect 86878 46066 87198 46067
rect 86878 46002 86886 46066
rect 86950 46002 86966 46066
rect 87030 46002 87046 46066
rect 87110 46002 87126 46066
rect 87190 46002 87198 46066
rect 86878 46001 87198 46002
rect 88454 45996 88934 46026
rect 87316 45936 88934 45996
rect 85887 45860 85953 45863
rect 87316 45860 87376 45936
rect 88454 45906 88934 45936
rect 85887 45858 87376 45860
rect 85887 45802 85892 45858
rect 85948 45802 87376 45858
rect 85887 45800 87376 45802
rect 85887 45797 85953 45800
rect 878 45522 1198 45523
rect 878 45458 886 45522
rect 950 45458 966 45522
rect 1030 45458 1046 45522
rect 1110 45458 1126 45522
rect 1190 45458 1198 45522
rect 878 45457 1198 45458
rect 84878 45522 85198 45523
rect 84878 45458 84886 45522
rect 84950 45458 84966 45522
rect 85030 45458 85046 45522
rect 85110 45458 85126 45522
rect 85190 45458 85198 45522
rect 84878 45457 85198 45458
rect 84323 45180 84389 45183
rect 84323 45178 87376 45180
rect 84323 45122 84328 45178
rect 84384 45122 87376 45178
rect 84323 45120 87376 45122
rect 84323 45117 84389 45120
rect 2878 44978 3198 44979
rect 2878 44914 2886 44978
rect 2950 44914 2966 44978
rect 3030 44914 3046 44978
rect 3110 44914 3126 44978
rect 3190 44914 3198 44978
rect 2878 44913 3198 44914
rect 86878 44978 87198 44979
rect 86878 44914 86886 44978
rect 86950 44914 86966 44978
rect 87030 44914 87046 44978
rect 87110 44914 87126 44978
rect 87190 44914 87198 44978
rect 86878 44913 87198 44914
rect 87316 44908 87376 45120
rect 88454 44908 88934 44938
rect 87316 44848 88934 44908
rect 88454 44818 88934 44848
rect 878 44434 1198 44435
rect 878 44370 886 44434
rect 950 44370 966 44434
rect 1030 44370 1046 44434
rect 1110 44370 1126 44434
rect 1190 44370 1198 44434
rect 878 44369 1198 44370
rect 84878 44434 85198 44435
rect 84878 44370 84886 44434
rect 84950 44370 84966 44434
rect 85030 44370 85046 44434
rect 85110 44370 85126 44434
rect 85190 44370 85198 44434
rect 84878 44369 85198 44370
rect 2878 43890 3198 43891
rect 2878 43826 2886 43890
rect 2950 43826 2966 43890
rect 3030 43826 3046 43890
rect 3110 43826 3126 43890
rect 3190 43826 3198 43890
rect 2878 43825 3198 43826
rect 86878 43890 87198 43891
rect 86878 43826 86886 43890
rect 86950 43826 86966 43890
rect 87030 43826 87046 43890
rect 87110 43826 87126 43890
rect 87190 43826 87198 43890
rect 86878 43825 87198 43826
rect 82851 43684 82917 43687
rect 83035 43684 83101 43687
rect 82851 43682 83101 43684
rect 82851 43626 82856 43682
rect 82912 43626 83040 43682
rect 83096 43626 83101 43682
rect 82851 43624 83101 43626
rect 82851 43621 82917 43624
rect 83035 43621 83101 43624
rect 85151 43684 85217 43687
rect 88454 43684 88934 43714
rect 85151 43682 88934 43684
rect 85151 43626 85156 43682
rect 85212 43626 88934 43682
rect 85151 43624 88934 43626
rect 85151 43621 85217 43624
rect 88454 43594 88934 43624
rect 878 43346 1198 43347
rect 878 43282 886 43346
rect 950 43282 966 43346
rect 1030 43282 1046 43346
rect 1110 43282 1126 43346
rect 1190 43282 1198 43346
rect 878 43281 1198 43282
rect 84878 43346 85198 43347
rect 84878 43282 84886 43346
rect 84950 43282 84966 43346
rect 85030 43282 85046 43346
rect 85110 43282 85126 43346
rect 85190 43282 85198 43346
rect 84878 43281 85198 43282
rect 2878 42802 3198 42803
rect 2878 42738 2886 42802
rect 2950 42738 2966 42802
rect 3030 42738 3046 42802
rect 3110 42738 3126 42802
rect 3190 42738 3198 42802
rect 2878 42737 3198 42738
rect 86878 42802 87198 42803
rect 86878 42738 86886 42802
rect 86950 42738 86966 42802
rect 87030 42738 87046 42802
rect 87110 42738 87126 42802
rect 87190 42738 87198 42802
rect 86878 42737 87198 42738
rect 84139 42460 84205 42463
rect 88454 42460 88934 42490
rect 84139 42458 88934 42460
rect 84139 42402 84144 42458
rect 84200 42402 88934 42458
rect 84139 42400 88934 42402
rect 84139 42397 84205 42400
rect 88454 42370 88934 42400
rect 878 42258 1198 42259
rect 878 42194 886 42258
rect 950 42194 966 42258
rect 1030 42194 1046 42258
rect 1110 42194 1126 42258
rect 1190 42194 1198 42258
rect 878 42193 1198 42194
rect 84878 42258 85198 42259
rect 84878 42194 84886 42258
rect 84950 42194 84966 42258
rect 85030 42194 85046 42258
rect 85110 42194 85126 42258
rect 85190 42194 85198 42258
rect 84878 42193 85198 42194
rect 2878 41714 3198 41715
rect 2878 41650 2886 41714
rect 2950 41650 2966 41714
rect 3030 41650 3046 41714
rect 3110 41650 3126 41714
rect 3190 41650 3198 41714
rect 2878 41649 3198 41650
rect 86878 41714 87198 41715
rect 86878 41650 86886 41714
rect 86950 41650 86966 41714
rect 87030 41650 87046 41714
rect 87110 41650 87126 41714
rect 87190 41650 87198 41714
rect 86878 41649 87198 41650
rect 84231 41372 84297 41375
rect 84231 41370 85352 41372
rect 84231 41314 84236 41370
rect 84292 41314 85352 41370
rect 84231 41312 85352 41314
rect 84231 41309 84297 41312
rect 85292 41236 85352 41312
rect 88454 41236 88934 41266
rect 85292 41176 88934 41236
rect 878 41170 1198 41171
rect 878 41106 886 41170
rect 950 41106 966 41170
rect 1030 41106 1046 41170
rect 1110 41106 1126 41170
rect 1190 41106 1198 41170
rect 878 41105 1198 41106
rect 84878 41170 85198 41171
rect 84878 41106 84886 41170
rect 84950 41106 84966 41170
rect 85030 41106 85046 41170
rect 85110 41106 85126 41170
rect 85190 41106 85198 41170
rect 88454 41146 88934 41176
rect 84878 41105 85198 41106
rect 2878 40626 3198 40627
rect 2878 40562 2886 40626
rect 2950 40562 2966 40626
rect 3030 40562 3046 40626
rect 3110 40562 3126 40626
rect 3190 40562 3198 40626
rect 2878 40561 3198 40562
rect 86878 40626 87198 40627
rect 86878 40562 86886 40626
rect 86950 40562 86966 40626
rect 87030 40562 87046 40626
rect 87110 40562 87126 40626
rect 87190 40562 87198 40626
rect 86878 40561 87198 40562
rect 878 40082 1198 40083
rect 878 40018 886 40082
rect 950 40018 966 40082
rect 1030 40018 1046 40082
rect 1110 40018 1126 40082
rect 1190 40018 1198 40082
rect 878 40017 1198 40018
rect 84878 40082 85198 40083
rect 84878 40018 84886 40082
rect 84950 40018 84966 40082
rect 85030 40018 85046 40082
rect 85110 40018 85126 40082
rect 85190 40018 85198 40082
rect 84878 40017 85198 40018
rect 88454 40012 88934 40042
rect 85292 39952 88934 40012
rect 84783 39876 84849 39879
rect 85292 39876 85352 39952
rect 88454 39922 88934 39952
rect 84783 39874 85352 39876
rect 84783 39818 84788 39874
rect 84844 39818 85352 39874
rect 84783 39816 85352 39818
rect 84783 39813 84849 39816
rect 2878 39538 3198 39539
rect 2878 39474 2886 39538
rect 2950 39474 2966 39538
rect 3030 39474 3046 39538
rect 3110 39474 3126 39538
rect 3190 39474 3198 39538
rect 2878 39473 3198 39474
rect 86878 39538 87198 39539
rect 86878 39474 86886 39538
rect 86950 39474 86966 39538
rect 87030 39474 87046 39538
rect 87110 39474 87126 39538
rect 87190 39474 87198 39538
rect 86878 39473 87198 39474
rect 878 38994 1198 38995
rect 878 38930 886 38994
rect 950 38930 966 38994
rect 1030 38930 1046 38994
rect 1110 38930 1126 38994
rect 1190 38930 1198 38994
rect 878 38929 1198 38930
rect 84878 38994 85198 38995
rect 84878 38930 84886 38994
rect 84950 38930 84966 38994
rect 85030 38930 85046 38994
rect 85110 38930 85126 38994
rect 85190 38930 85198 38994
rect 84878 38929 85198 38930
rect 83127 38788 83193 38791
rect 88454 38788 88934 38818
rect 83127 38786 88934 38788
rect 83127 38730 83132 38786
rect 83188 38730 88934 38786
rect 83127 38728 88934 38730
rect 83127 38725 83193 38728
rect 88454 38698 88934 38728
rect 2878 38450 3198 38451
rect 2878 38386 2886 38450
rect 2950 38386 2966 38450
rect 3030 38386 3046 38450
rect 3110 38386 3126 38450
rect 3190 38386 3198 38450
rect 2878 38385 3198 38386
rect 86878 38450 87198 38451
rect 86878 38386 86886 38450
rect 86950 38386 86966 38450
rect 87030 38386 87046 38450
rect 87110 38386 87126 38450
rect 87190 38386 87198 38450
rect 86878 38385 87198 38386
rect 878 37906 1198 37907
rect 878 37842 886 37906
rect 950 37842 966 37906
rect 1030 37842 1046 37906
rect 1110 37842 1126 37906
rect 1190 37842 1198 37906
rect 878 37841 1198 37842
rect 84878 37906 85198 37907
rect 84878 37842 84886 37906
rect 84950 37842 84966 37906
rect 85030 37842 85046 37906
rect 85110 37842 85126 37906
rect 85190 37842 85198 37906
rect 84878 37841 85198 37842
rect 83035 37700 83101 37703
rect 88454 37700 88934 37730
rect 83035 37698 88934 37700
rect 83035 37642 83040 37698
rect 83096 37642 88934 37698
rect 83035 37640 88934 37642
rect 83035 37637 83101 37640
rect 88454 37610 88934 37640
rect 2878 37362 3198 37363
rect 2878 37298 2886 37362
rect 2950 37298 2966 37362
rect 3030 37298 3046 37362
rect 3110 37298 3126 37362
rect 3190 37298 3198 37362
rect 2878 37297 3198 37298
rect 86878 37362 87198 37363
rect 86878 37298 86886 37362
rect 86950 37298 86966 37362
rect 87030 37298 87046 37362
rect 87110 37298 87126 37362
rect 87190 37298 87198 37362
rect 86878 37297 87198 37298
rect 878 36818 1198 36819
rect 878 36754 886 36818
rect 950 36754 966 36818
rect 1030 36754 1046 36818
rect 1110 36754 1126 36818
rect 1190 36754 1198 36818
rect 878 36753 1198 36754
rect 84878 36818 85198 36819
rect 84878 36754 84886 36818
rect 84950 36754 84966 36818
rect 85030 36754 85046 36818
rect 85110 36754 85126 36818
rect 85190 36754 85198 36818
rect 84878 36753 85198 36754
rect 84783 36476 84849 36479
rect 88454 36476 88934 36506
rect 84783 36474 88934 36476
rect 84783 36418 84788 36474
rect 84844 36418 88934 36474
rect 84783 36416 88934 36418
rect 84783 36413 84849 36416
rect 88454 36386 88934 36416
rect 2878 36274 3198 36275
rect 2878 36210 2886 36274
rect 2950 36210 2966 36274
rect 3030 36210 3046 36274
rect 3110 36210 3126 36274
rect 3190 36210 3198 36274
rect 2878 36209 3198 36210
rect 86878 36274 87198 36275
rect 86878 36210 86886 36274
rect 86950 36210 86966 36274
rect 87030 36210 87046 36274
rect 87110 36210 87126 36274
rect 87190 36210 87198 36274
rect 86878 36209 87198 36210
rect 878 35730 1198 35731
rect 878 35666 886 35730
rect 950 35666 966 35730
rect 1030 35666 1046 35730
rect 1110 35666 1126 35730
rect 1190 35666 1198 35730
rect 878 35665 1198 35666
rect 84878 35730 85198 35731
rect 84878 35666 84886 35730
rect 84950 35666 84966 35730
rect 85030 35666 85046 35730
rect 85110 35666 85126 35730
rect 85190 35666 85198 35730
rect 84878 35665 85198 35666
rect 88454 35252 88934 35282
rect 87316 35192 88934 35252
rect 2878 35186 3198 35187
rect 2878 35122 2886 35186
rect 2950 35122 2966 35186
rect 3030 35122 3046 35186
rect 3110 35122 3126 35186
rect 3190 35122 3198 35186
rect 2878 35121 3198 35122
rect 86878 35186 87198 35187
rect 86878 35122 86886 35186
rect 86950 35122 86966 35186
rect 87030 35122 87046 35186
rect 87110 35122 87126 35186
rect 87190 35122 87198 35186
rect 86878 35121 87198 35122
rect 84732 34918 84738 34982
rect 84802 34980 84808 34982
rect 87316 34980 87376 35192
rect 88454 35162 88934 35192
rect 84802 34920 87376 34980
rect 84802 34918 84808 34920
rect 878 34642 1198 34643
rect 878 34578 886 34642
rect 950 34578 966 34642
rect 1030 34578 1046 34642
rect 1110 34578 1126 34642
rect 1190 34578 1198 34642
rect 878 34577 1198 34578
rect 84878 34642 85198 34643
rect 84878 34578 84886 34642
rect 84950 34578 84966 34642
rect 85030 34578 85046 34642
rect 85110 34578 85126 34642
rect 85190 34578 85198 34642
rect 84878 34577 85198 34578
rect 3271 34572 3337 34575
rect 3915 34572 3981 34575
rect 3271 34570 3981 34572
rect 3271 34514 3276 34570
rect 3332 34514 3920 34570
rect 3976 34514 3981 34570
rect 3271 34512 3981 34514
rect 3271 34509 3337 34512
rect 3915 34509 3981 34512
rect 2878 34098 3198 34099
rect 2878 34034 2886 34098
rect 2950 34034 2966 34098
rect 3030 34034 3046 34098
rect 3110 34034 3126 34098
rect 3190 34034 3198 34098
rect 2878 34033 3198 34034
rect 86878 34098 87198 34099
rect 86878 34034 86886 34098
rect 86950 34034 86966 34098
rect 87030 34034 87046 34098
rect 87110 34034 87126 34098
rect 87190 34034 87198 34098
rect 86878 34033 87198 34034
rect 88454 34028 88934 34058
rect 87316 33968 88934 34028
rect 83628 33830 83634 33894
rect 83698 33892 83704 33894
rect 87316 33892 87376 33968
rect 88454 33938 88934 33968
rect 83698 33832 87376 33892
rect 83698 33830 83704 33832
rect 878 33554 1198 33555
rect 878 33490 886 33554
rect 950 33490 966 33554
rect 1030 33490 1046 33554
rect 1110 33490 1126 33554
rect 1190 33490 1198 33554
rect 878 33489 1198 33490
rect 84878 33554 85198 33555
rect 84878 33490 84886 33554
rect 84950 33490 84966 33554
rect 85030 33490 85046 33554
rect 85110 33490 85126 33554
rect 85190 33490 85198 33554
rect 84878 33489 85198 33490
rect 2878 33010 3198 33011
rect 2878 32946 2886 33010
rect 2950 32946 2966 33010
rect 3030 32946 3046 33010
rect 3110 32946 3126 33010
rect 3190 32946 3198 33010
rect 2878 32945 3198 32946
rect 86878 33010 87198 33011
rect 86878 32946 86886 33010
rect 86950 32946 86966 33010
rect 87030 32946 87046 33010
rect 87110 32946 87126 33010
rect 87190 32946 87198 33010
rect 86878 32945 87198 32946
rect 84364 32742 84370 32806
rect 84434 32804 84440 32806
rect 88454 32804 88934 32834
rect 84434 32744 88934 32804
rect 84434 32742 84440 32744
rect 88454 32714 88934 32744
rect 878 32466 1198 32467
rect 878 32402 886 32466
rect 950 32402 966 32466
rect 1030 32402 1046 32466
rect 1110 32402 1126 32466
rect 1190 32402 1198 32466
rect 878 32401 1198 32402
rect 84878 32466 85198 32467
rect 84878 32402 84886 32466
rect 84950 32402 84966 32466
rect 85030 32402 85046 32466
rect 85110 32402 85126 32466
rect 85190 32402 85198 32466
rect 84878 32401 85198 32402
rect 2878 31922 3198 31923
rect 2878 31858 2886 31922
rect 2950 31858 2966 31922
rect 3030 31858 3046 31922
rect 3110 31858 3126 31922
rect 3190 31858 3198 31922
rect 2878 31857 3198 31858
rect 86878 31922 87198 31923
rect 86878 31858 86886 31922
rect 86950 31858 86966 31922
rect 87030 31858 87046 31922
rect 87110 31858 87126 31922
rect 87190 31858 87198 31922
rect 86878 31857 87198 31858
rect 84139 31580 84205 31583
rect 88454 31580 88934 31610
rect 84139 31578 88934 31580
rect 82164 31444 82224 31567
rect 84139 31522 84144 31578
rect 84200 31522 88934 31578
rect 84139 31520 88934 31522
rect 84139 31517 84205 31520
rect 88454 31490 88934 31520
rect 84047 31444 84113 31447
rect 82164 31442 84113 31444
rect 82164 31386 84052 31442
rect 84108 31386 84113 31442
rect 82164 31384 84113 31386
rect 84047 31381 84113 31384
rect 878 31378 1198 31379
rect 878 31314 886 31378
rect 950 31314 966 31378
rect 1030 31314 1046 31378
rect 1110 31314 1126 31378
rect 1190 31314 1198 31378
rect 878 31313 1198 31314
rect 84878 31378 85198 31379
rect 84878 31314 84886 31378
rect 84950 31314 84966 31378
rect 85030 31314 85046 31378
rect 85110 31314 85126 31378
rect 85190 31314 85198 31378
rect 84878 31313 85198 31314
rect 2878 30834 3198 30835
rect 2878 30770 2886 30834
rect 2950 30770 2966 30834
rect 3030 30770 3046 30834
rect 3110 30770 3126 30834
rect 3190 30770 3198 30834
rect 2878 30769 3198 30770
rect 86878 30834 87198 30835
rect 86878 30770 86886 30834
rect 86950 30770 86966 30834
rect 87030 30770 87046 30834
rect 87110 30770 87126 30834
rect 87190 30770 87198 30834
rect 86878 30769 87198 30770
rect 83679 30492 83745 30495
rect 88454 30492 88934 30522
rect 83679 30490 88934 30492
rect 83679 30434 83684 30490
rect 83740 30434 88934 30490
rect 83679 30432 88934 30434
rect 83679 30429 83745 30432
rect 88454 30402 88934 30432
rect 878 30290 1198 30291
rect 878 30226 886 30290
rect 950 30226 966 30290
rect 1030 30226 1046 30290
rect 1110 30226 1126 30290
rect 1190 30226 1198 30290
rect 878 30225 1198 30226
rect 84878 30290 85198 30291
rect 84878 30226 84886 30290
rect 84950 30226 84966 30290
rect 85030 30226 85046 30290
rect 85110 30226 85126 30290
rect 85190 30226 85198 30290
rect 84878 30225 85198 30226
rect 84047 29948 84113 29951
rect 82164 29946 84113 29948
rect 82164 29890 84052 29946
rect 84108 29890 84113 29946
rect 82164 29888 84113 29890
rect 82164 29867 82224 29888
rect 84047 29885 84113 29888
rect 2878 29746 3198 29747
rect 2878 29682 2886 29746
rect 2950 29682 2966 29746
rect 3030 29682 3046 29746
rect 3110 29682 3126 29746
rect 3190 29682 3198 29746
rect 2878 29681 3198 29682
rect 86878 29746 87198 29747
rect 86878 29682 86886 29746
rect 86950 29682 86966 29746
rect 87030 29682 87046 29746
rect 87110 29682 87126 29746
rect 87190 29682 87198 29746
rect 86878 29681 87198 29682
rect 5612 29478 5618 29542
rect 5682 29540 5688 29542
rect 5755 29540 5821 29543
rect 5682 29538 5821 29540
rect 5682 29482 5760 29538
rect 5816 29482 5821 29538
rect 5682 29480 5821 29482
rect 5682 29478 5688 29480
rect 5755 29477 5821 29480
rect 84691 29404 84757 29407
rect 85468 29404 85474 29406
rect 84691 29402 85474 29404
rect 84691 29346 84696 29402
rect 84752 29346 85474 29402
rect 84691 29344 85474 29346
rect 84691 29341 84757 29344
rect 85468 29342 85474 29344
rect 85538 29342 85544 29406
rect 88454 29268 88934 29298
rect 85292 29208 88934 29268
rect 878 29202 1198 29203
rect 878 29138 886 29202
rect 950 29138 966 29202
rect 1030 29138 1046 29202
rect 1110 29138 1126 29202
rect 1190 29138 1198 29202
rect 878 29137 1198 29138
rect 84878 29202 85198 29203
rect 84878 29138 84886 29202
rect 84950 29138 84966 29202
rect 85030 29138 85046 29202
rect 85110 29138 85126 29202
rect 85190 29138 85198 29202
rect 84878 29137 85198 29138
rect 84691 28996 84757 28999
rect 85292 28996 85352 29208
rect 88454 29178 88934 29208
rect 84691 28994 85352 28996
rect 84691 28938 84696 28994
rect 84752 28938 85352 28994
rect 84691 28936 85352 28938
rect 84691 28933 84757 28936
rect 82164 28724 82224 28739
rect 84139 28724 84205 28727
rect 82164 28722 84205 28724
rect 82164 28666 84144 28722
rect 84200 28666 84205 28722
rect 82164 28664 84205 28666
rect 84139 28661 84205 28664
rect 2878 28658 3198 28659
rect 2878 28594 2886 28658
rect 2950 28594 2966 28658
rect 3030 28594 3046 28658
rect 3110 28594 3126 28658
rect 3190 28594 3198 28658
rect 2878 28593 3198 28594
rect 86878 28658 87198 28659
rect 86878 28594 86886 28658
rect 86950 28594 86966 28658
rect 87030 28594 87046 28658
rect 87110 28594 87126 28658
rect 87190 28594 87198 28658
rect 86878 28593 87198 28594
rect 84599 28316 84665 28319
rect 85468 28316 85474 28318
rect 84599 28314 85474 28316
rect 84599 28258 84604 28314
rect 84660 28258 85474 28314
rect 84599 28256 85474 28258
rect 84599 28253 84665 28256
rect 85468 28254 85474 28256
rect 85538 28254 85544 28318
rect 82667 28180 82733 28183
rect 83495 28180 83561 28183
rect 82667 28178 83561 28180
rect 82667 28122 82672 28178
rect 82728 28122 83500 28178
rect 83556 28122 83561 28178
rect 82667 28120 83561 28122
rect 82667 28117 82733 28120
rect 83495 28117 83561 28120
rect 878 28114 1198 28115
rect 878 28050 886 28114
rect 950 28050 966 28114
rect 1030 28050 1046 28114
rect 1110 28050 1126 28114
rect 1190 28050 1198 28114
rect 878 28049 1198 28050
rect 84878 28114 85198 28115
rect 84878 28050 84886 28114
rect 84950 28050 84966 28114
rect 85030 28050 85046 28114
rect 85110 28050 85126 28114
rect 85190 28050 85198 28114
rect 84878 28049 85198 28050
rect 5295 28044 5361 28047
rect 5612 28044 5618 28046
rect 5295 28042 5618 28044
rect 5295 27986 5300 28042
rect 5356 27986 5618 28042
rect 5295 27984 5618 27986
rect 5295 27981 5361 27984
rect 5612 27982 5618 27984
rect 5682 27982 5688 28046
rect 88454 28044 88934 28074
rect 85292 27984 88934 28044
rect 83219 27908 83285 27911
rect 85292 27908 85352 27984
rect 88454 27954 88934 27984
rect 83219 27906 85352 27908
rect 83219 27850 83224 27906
rect 83280 27850 85352 27906
rect 83219 27848 85352 27850
rect 83219 27845 83285 27848
rect 2878 27570 3198 27571
rect 2878 27506 2886 27570
rect 2950 27506 2966 27570
rect 3030 27506 3046 27570
rect 3110 27506 3126 27570
rect 3190 27506 3198 27570
rect 2878 27505 3198 27506
rect 86878 27570 87198 27571
rect 86878 27506 86886 27570
rect 86950 27506 86966 27570
rect 87030 27506 87046 27570
rect 87110 27506 87126 27570
rect 87190 27506 87198 27570
rect 86878 27505 87198 27506
rect 84231 27092 84297 27095
rect 82164 27090 84297 27092
rect 82164 27034 84236 27090
rect 84292 27034 84297 27090
rect 82164 27032 84297 27034
rect 84231 27029 84297 27032
rect 878 27026 1198 27027
rect 878 26962 886 27026
rect 950 26962 966 27026
rect 1030 26962 1046 27026
rect 1110 26962 1126 27026
rect 1190 26962 1198 27026
rect 878 26961 1198 26962
rect 84878 27026 85198 27027
rect 84878 26962 84886 27026
rect 84950 26962 84966 27026
rect 85030 26962 85046 27026
rect 85110 26962 85126 27026
rect 85190 26962 85198 27026
rect 84878 26961 85198 26962
rect 84323 26820 84389 26823
rect 88454 26820 88934 26850
rect 84323 26818 88934 26820
rect 84323 26762 84328 26818
rect 84384 26762 88934 26818
rect 84323 26760 88934 26762
rect 84323 26757 84389 26760
rect 88454 26730 88934 26760
rect 2878 26482 3198 26483
rect 2878 26418 2886 26482
rect 2950 26418 2966 26482
rect 3030 26418 3046 26482
rect 3110 26418 3126 26482
rect 3190 26418 3198 26482
rect 2878 26417 3198 26418
rect 86878 26482 87198 26483
rect 86878 26418 86886 26482
rect 86950 26418 86966 26482
rect 87030 26418 87046 26482
rect 87110 26418 87126 26482
rect 87190 26418 87198 26482
rect 86878 26417 87198 26418
rect 878 25938 1198 25939
rect 878 25874 886 25938
rect 950 25874 966 25938
rect 1030 25874 1046 25938
rect 1110 25874 1126 25938
rect 1190 25874 1198 25938
rect 84878 25938 85198 25939
rect 878 25873 1198 25874
rect 81796 25732 81856 25911
rect 84878 25874 84886 25938
rect 84950 25874 84966 25938
rect 85030 25874 85046 25938
rect 85110 25874 85126 25938
rect 85190 25874 85198 25938
rect 84878 25873 85198 25874
rect 83495 25732 83561 25735
rect 81796 25730 83561 25732
rect 81796 25674 83500 25730
rect 83556 25674 83561 25730
rect 81796 25672 83561 25674
rect 83495 25669 83561 25672
rect 3363 25596 3429 25599
rect 3915 25596 3981 25599
rect 3363 25594 3981 25596
rect 3363 25538 3368 25594
rect 3424 25538 3920 25594
rect 3976 25538 3981 25594
rect 3363 25536 3981 25538
rect 3363 25533 3429 25536
rect 3915 25533 3981 25536
rect 84875 25596 84941 25599
rect 88454 25596 88934 25626
rect 84875 25594 88934 25596
rect 84875 25538 84880 25594
rect 84936 25538 88934 25594
rect 84875 25536 88934 25538
rect 84875 25533 84941 25536
rect 88454 25506 88934 25536
rect 2878 25394 3198 25395
rect 2878 25330 2886 25394
rect 2950 25330 2966 25394
rect 3030 25330 3046 25394
rect 3110 25330 3126 25394
rect 3190 25330 3198 25394
rect 2878 25329 3198 25330
rect 86878 25394 87198 25395
rect 86878 25330 86886 25394
rect 86950 25330 86966 25394
rect 87030 25330 87046 25394
rect 87110 25330 87126 25394
rect 87190 25330 87198 25394
rect 86878 25329 87198 25330
rect 878 24850 1198 24851
rect 878 24786 886 24850
rect 950 24786 966 24850
rect 1030 24786 1046 24850
rect 1110 24786 1126 24850
rect 1190 24786 1198 24850
rect 878 24785 1198 24786
rect 84878 24850 85198 24851
rect 84878 24786 84886 24850
rect 84950 24786 84966 24850
rect 85030 24786 85046 24850
rect 85110 24786 85126 24850
rect 85190 24786 85198 24850
rect 84878 24785 85198 24786
rect 82340 24446 82346 24510
rect 82410 24508 82416 24510
rect 84599 24508 84665 24511
rect 82410 24448 82960 24508
rect 82410 24446 82416 24448
rect 82667 24372 82733 24375
rect 82532 24370 82733 24372
rect 82532 24314 82672 24370
rect 82728 24314 82733 24370
rect 82532 24312 82733 24314
rect 2878 24306 3198 24307
rect 2878 24242 2886 24306
rect 2950 24242 2966 24306
rect 3030 24242 3046 24306
rect 3110 24242 3126 24306
rect 3190 24242 3198 24306
rect 2878 24241 3198 24242
rect 82532 24236 82592 24312
rect 82667 24309 82733 24312
rect 82667 24236 82733 24239
rect 82532 24234 82733 24236
rect 82164 23964 82224 24211
rect 82532 24178 82672 24234
rect 82728 24178 82733 24234
rect 82532 24176 82733 24178
rect 82667 24173 82733 24176
rect 82340 24038 82346 24102
rect 82410 24100 82416 24102
rect 82900 24100 82960 24448
rect 84599 24506 87376 24508
rect 84599 24450 84604 24506
rect 84660 24450 87376 24506
rect 84599 24448 87376 24450
rect 84599 24445 84665 24448
rect 87316 24372 87376 24448
rect 88454 24372 88934 24402
rect 87316 24312 88934 24372
rect 86878 24306 87198 24307
rect 86878 24242 86886 24306
rect 86950 24242 86966 24306
rect 87030 24242 87046 24306
rect 87110 24242 87126 24306
rect 87190 24242 87198 24306
rect 88454 24282 88934 24312
rect 86878 24241 87198 24242
rect 83996 24174 84002 24238
rect 84066 24236 84072 24238
rect 84691 24236 84757 24239
rect 84066 24234 84757 24236
rect 84066 24178 84696 24234
rect 84752 24178 84757 24234
rect 84066 24176 84757 24178
rect 84066 24174 84072 24176
rect 84691 24173 84757 24176
rect 82410 24040 82960 24100
rect 82410 24038 82416 24040
rect 84231 23964 84297 23967
rect 82164 23962 84297 23964
rect 82164 23906 84236 23962
rect 84292 23906 84297 23962
rect 82164 23904 84297 23906
rect 84231 23901 84297 23904
rect 878 23762 1198 23763
rect 878 23698 886 23762
rect 950 23698 966 23762
rect 1030 23698 1046 23762
rect 1110 23698 1126 23762
rect 1190 23698 1198 23762
rect 878 23697 1198 23698
rect 84878 23762 85198 23763
rect 84878 23698 84886 23762
rect 84950 23698 84966 23762
rect 85030 23698 85046 23762
rect 85110 23698 85126 23762
rect 85190 23698 85198 23762
rect 84878 23697 85198 23698
rect 83955 23420 84021 23423
rect 83955 23418 87376 23420
rect 83955 23362 83960 23418
rect 84016 23362 87376 23418
rect 83955 23360 87376 23362
rect 83955 23357 84021 23360
rect 2878 23218 3198 23219
rect 2878 23154 2886 23218
rect 2950 23154 2966 23218
rect 3030 23154 3046 23218
rect 3110 23154 3126 23218
rect 3190 23154 3198 23218
rect 2878 23153 3198 23154
rect 86878 23218 87198 23219
rect 86878 23154 86886 23218
rect 86950 23154 86966 23218
rect 87030 23154 87046 23218
rect 87110 23154 87126 23218
rect 87190 23154 87198 23218
rect 86878 23153 87198 23154
rect 83955 23148 84021 23151
rect 82164 23146 84021 23148
rect 82164 23090 83960 23146
rect 84016 23090 84021 23146
rect 82164 23088 84021 23090
rect 87316 23148 87376 23360
rect 88454 23148 88934 23178
rect 87316 23088 88934 23148
rect 82164 23083 82224 23088
rect 83955 23085 84021 23088
rect 88454 23058 88934 23088
rect 3823 22876 3889 22879
rect 4140 22876 4146 22878
rect 3823 22874 4146 22876
rect 3823 22818 3828 22874
rect 3884 22818 4146 22874
rect 3823 22816 4146 22818
rect 3823 22813 3889 22816
rect 4140 22814 4146 22816
rect 4210 22876 4216 22878
rect 4210 22816 5128 22876
rect 4210 22814 4216 22816
rect 878 22674 1198 22675
rect 878 22610 886 22674
rect 950 22610 966 22674
rect 1030 22610 1046 22674
rect 1110 22610 1126 22674
rect 1190 22610 1198 22674
rect 878 22609 1198 22610
rect 5068 22410 5128 22816
rect 84878 22674 85198 22675
rect 84878 22610 84886 22674
rect 84950 22610 84966 22674
rect 85030 22610 85046 22674
rect 85110 22610 85126 22674
rect 85190 22610 85198 22674
rect 84878 22609 85198 22610
rect 2878 22130 3198 22131
rect 2878 22066 2886 22130
rect 2950 22066 2966 22130
rect 3030 22066 3046 22130
rect 3110 22066 3126 22130
rect 3190 22066 3198 22130
rect 2878 22065 3198 22066
rect 86878 22130 87198 22131
rect 86878 22066 86886 22130
rect 86950 22066 86966 22130
rect 87030 22066 87046 22130
rect 87110 22066 87126 22130
rect 87190 22066 87198 22130
rect 86878 22065 87198 22066
rect 88454 22060 88934 22090
rect 87316 22000 88934 22060
rect 84180 21862 84186 21926
rect 84250 21924 84256 21926
rect 87316 21924 87376 22000
rect 88454 21970 88934 22000
rect 84250 21864 87376 21924
rect 84250 21862 84256 21864
rect 878 21586 1198 21587
rect 878 21522 886 21586
rect 950 21522 966 21586
rect 1030 21522 1046 21586
rect 1110 21522 1126 21586
rect 1190 21522 1198 21586
rect 878 21521 1198 21522
rect 84878 21586 85198 21587
rect 84878 21522 84886 21586
rect 84950 21522 84966 21586
rect 85030 21522 85046 21586
rect 85110 21522 85126 21586
rect 85190 21522 85198 21586
rect 84878 21521 85198 21522
rect 2878 21042 3198 21043
rect 2878 20978 2886 21042
rect 2950 20978 2966 21042
rect 3030 20978 3046 21042
rect 3110 20978 3126 21042
rect 3190 20978 3198 21042
rect 2878 20977 3198 20978
rect 86878 21042 87198 21043
rect 86878 20978 86886 21042
rect 86950 20978 86966 21042
rect 87030 20978 87046 21042
rect 87110 20978 87126 21042
rect 87190 20978 87198 21042
rect 86878 20977 87198 20978
rect 84415 20836 84481 20839
rect 88454 20836 88934 20866
rect 84415 20834 88934 20836
rect 84415 20778 84420 20834
rect 84476 20778 88934 20834
rect 84415 20776 88934 20778
rect 84415 20773 84481 20776
rect 88454 20746 88934 20776
rect 4283 20564 4349 20567
rect 5068 20564 5128 20710
rect 4283 20562 5128 20564
rect 4283 20506 4288 20562
rect 4344 20506 5128 20562
rect 4283 20504 5128 20506
rect 4283 20501 4349 20504
rect 878 20498 1198 20499
rect 878 20434 886 20498
rect 950 20434 966 20498
rect 1030 20434 1046 20498
rect 1110 20434 1126 20498
rect 1190 20434 1198 20498
rect 878 20433 1198 20434
rect 84878 20498 85198 20499
rect 84878 20434 84886 20498
rect 84950 20434 84966 20498
rect 85030 20434 85046 20498
rect 85110 20434 85126 20498
rect 85190 20434 85198 20498
rect 84878 20433 85198 20434
rect 2878 19954 3198 19955
rect 2878 19890 2886 19954
rect 2950 19890 2966 19954
rect 3030 19890 3046 19954
rect 3110 19890 3126 19954
rect 3190 19890 3198 19954
rect 2878 19889 3198 19890
rect 86878 19954 87198 19955
rect 86878 19890 86886 19954
rect 86950 19890 86966 19954
rect 87030 19890 87046 19954
rect 87110 19890 87126 19954
rect 87190 19890 87198 19954
rect 86878 19889 87198 19890
rect 83996 19550 84002 19614
rect 84066 19612 84072 19614
rect 84231 19612 84297 19615
rect 84066 19610 84297 19612
rect 84066 19554 84236 19610
rect 84292 19554 84297 19610
rect 84066 19552 84297 19554
rect 84066 19550 84072 19552
rect 84231 19549 84297 19552
rect 85519 19612 85585 19615
rect 88454 19612 88934 19642
rect 85519 19610 88934 19612
rect 85519 19554 85524 19610
rect 85580 19554 88934 19610
rect 85519 19552 88934 19554
rect 85519 19549 85585 19552
rect 88454 19522 88934 19552
rect 878 19410 1198 19411
rect 878 19346 886 19410
rect 950 19346 966 19410
rect 1030 19346 1046 19410
rect 1110 19346 1126 19410
rect 1190 19346 1198 19410
rect 878 19345 1198 19346
rect 84878 19410 85198 19411
rect 84878 19346 84886 19410
rect 84950 19346 84966 19410
rect 85030 19346 85046 19410
rect 85110 19346 85126 19410
rect 85190 19346 85198 19410
rect 84878 19345 85198 19346
rect 2878 18866 3198 18867
rect 2878 18802 2886 18866
rect 2950 18802 2966 18866
rect 3030 18802 3046 18866
rect 3110 18802 3126 18866
rect 3190 18802 3198 18866
rect 2878 18801 3198 18802
rect 86878 18866 87198 18867
rect 86878 18802 86886 18866
rect 86950 18802 86966 18866
rect 87030 18802 87046 18866
rect 87110 18802 87126 18866
rect 87190 18802 87198 18866
rect 86878 18801 87198 18802
rect 83955 18524 84021 18527
rect 83955 18522 85352 18524
rect 83955 18466 83960 18522
rect 84016 18466 85352 18522
rect 83955 18464 85352 18466
rect 83955 18461 84021 18464
rect 85292 18388 85352 18464
rect 88454 18388 88934 18418
rect 85292 18328 88934 18388
rect 878 18322 1198 18323
rect 878 18258 886 18322
rect 950 18258 966 18322
rect 1030 18258 1046 18322
rect 1110 18258 1126 18322
rect 1190 18258 1198 18322
rect 878 18257 1198 18258
rect 84878 18322 85198 18323
rect 84878 18258 84886 18322
rect 84950 18258 84966 18322
rect 85030 18258 85046 18322
rect 85110 18258 85126 18322
rect 85190 18258 85198 18322
rect 88454 18298 88934 18328
rect 84878 18257 85198 18258
rect 82483 17844 82549 17847
rect 82759 17844 82825 17847
rect 82483 17842 82825 17844
rect 82483 17786 82488 17842
rect 82544 17786 82764 17842
rect 82820 17786 82825 17842
rect 82483 17784 82825 17786
rect 82483 17781 82549 17784
rect 82759 17781 82825 17784
rect 83495 17844 83561 17847
rect 83863 17844 83929 17847
rect 83495 17842 83929 17844
rect 83495 17786 83500 17842
rect 83556 17786 83868 17842
rect 83924 17786 83929 17842
rect 83495 17784 83929 17786
rect 83495 17781 83561 17784
rect 83863 17781 83929 17784
rect 2878 17778 3198 17779
rect 2878 17714 2886 17778
rect 2950 17714 2966 17778
rect 3030 17714 3046 17778
rect 3110 17714 3126 17778
rect 3190 17714 3198 17778
rect 2878 17713 3198 17714
rect 86878 17778 87198 17779
rect 86878 17714 86886 17778
rect 86950 17714 86966 17778
rect 87030 17714 87046 17778
rect 87110 17714 87126 17778
rect 87190 17714 87198 17778
rect 86878 17713 87198 17714
rect 84139 17436 84205 17439
rect 84139 17434 85720 17436
rect 84139 17378 84144 17434
rect 84200 17378 85720 17434
rect 84139 17376 85720 17378
rect 84139 17373 84205 17376
rect 878 17234 1198 17235
rect 878 17170 886 17234
rect 950 17170 966 17234
rect 1030 17170 1046 17234
rect 1110 17170 1126 17234
rect 1190 17170 1198 17234
rect 878 17169 1198 17170
rect 84878 17234 85198 17235
rect 84878 17170 84886 17234
rect 84950 17170 84966 17234
rect 85030 17170 85046 17234
rect 85110 17170 85126 17234
rect 85190 17170 85198 17234
rect 84878 17169 85198 17170
rect 85660 17164 85720 17376
rect 88454 17164 88934 17194
rect 85660 17104 88934 17164
rect 88454 17074 88934 17104
rect 3455 17028 3521 17031
rect 3455 17026 3840 17028
rect 3455 16970 3460 17026
rect 3516 16970 3840 17026
rect 3455 16968 3840 16970
rect 3455 16965 3521 16968
rect 2878 16690 3198 16691
rect 2878 16626 2886 16690
rect 2950 16626 2966 16690
rect 3030 16626 3046 16690
rect 3110 16626 3126 16690
rect 3190 16626 3198 16690
rect 2878 16625 3198 16626
rect 3455 16620 3521 16623
rect 3780 16620 3840 16968
rect 86878 16690 87198 16691
rect 86878 16626 86886 16690
rect 86950 16626 86966 16690
rect 87030 16626 87046 16690
rect 87110 16626 87126 16690
rect 87190 16626 87198 16690
rect 86878 16625 87198 16626
rect 3455 16618 3840 16620
rect 3455 16562 3460 16618
rect 3516 16562 3840 16618
rect 3455 16560 3840 16562
rect 3455 16557 3521 16560
rect 84875 16348 84941 16351
rect 84875 16346 85352 16348
rect 84875 16290 84880 16346
rect 84936 16290 85352 16346
rect 84875 16288 85352 16290
rect 84875 16285 84941 16288
rect 878 16146 1198 16147
rect 878 16082 886 16146
rect 950 16082 966 16146
rect 1030 16082 1046 16146
rect 1110 16082 1126 16146
rect 1190 16082 1198 16146
rect 878 16081 1198 16082
rect 84878 16146 85198 16147
rect 84878 16082 84886 16146
rect 84950 16082 84966 16146
rect 85030 16082 85046 16146
rect 85110 16082 85126 16146
rect 85190 16082 85198 16146
rect 84878 16081 85198 16082
rect 85292 15940 85352 16288
rect 88454 15940 88934 15970
rect 85292 15880 88934 15940
rect 88454 15850 88934 15880
rect 2878 15602 3198 15603
rect 2878 15538 2886 15602
rect 2950 15538 2966 15602
rect 3030 15538 3046 15602
rect 3110 15538 3126 15602
rect 3190 15538 3198 15602
rect 2878 15537 3198 15538
rect 86878 15602 87198 15603
rect 86878 15538 86886 15602
rect 86950 15538 86966 15602
rect 87030 15538 87046 15602
rect 87110 15538 87126 15602
rect 87190 15538 87198 15602
rect 86878 15537 87198 15538
rect 82340 15470 82346 15534
rect 82410 15532 82416 15534
rect 82892 15532 82898 15534
rect 82410 15472 82898 15532
rect 82410 15470 82416 15472
rect 82892 15470 82898 15472
rect 82962 15470 82968 15534
rect 82340 15334 82346 15398
rect 82410 15396 82416 15398
rect 82667 15396 82733 15399
rect 82410 15394 82733 15396
rect 82410 15338 82672 15394
rect 82728 15338 82733 15394
rect 82410 15336 82733 15338
rect 82410 15334 82416 15336
rect 82667 15333 82733 15336
rect 878 15058 1198 15059
rect 878 14994 886 15058
rect 950 14994 966 15058
rect 1030 14994 1046 15058
rect 1110 14994 1126 15058
rect 1190 14994 1198 15058
rect 878 14993 1198 14994
rect 84878 15058 85198 15059
rect 84878 14994 84886 15058
rect 84950 14994 84966 15058
rect 85030 14994 85046 15058
rect 85110 14994 85126 15058
rect 85190 14994 85198 15058
rect 84878 14993 85198 14994
rect 84231 14852 84297 14855
rect 88454 14852 88934 14882
rect 84231 14850 88934 14852
rect 84231 14794 84236 14850
rect 84292 14794 88934 14850
rect 84231 14792 88934 14794
rect 84231 14789 84297 14792
rect 88454 14762 88934 14792
rect 2878 14514 3198 14515
rect 2878 14450 2886 14514
rect 2950 14450 2966 14514
rect 3030 14450 3046 14514
rect 3110 14450 3126 14514
rect 3190 14450 3198 14514
rect 2878 14449 3198 14450
rect 86878 14514 87198 14515
rect 86878 14450 86886 14514
rect 86950 14450 86966 14514
rect 87030 14450 87046 14514
rect 87110 14450 87126 14514
rect 87190 14450 87198 14514
rect 86878 14449 87198 14450
rect 878 13970 1198 13971
rect 878 13906 886 13970
rect 950 13906 966 13970
rect 1030 13906 1046 13970
rect 1110 13906 1126 13970
rect 1190 13906 1198 13970
rect 878 13905 1198 13906
rect 84878 13970 85198 13971
rect 84878 13906 84886 13970
rect 84950 13906 84966 13970
rect 85030 13906 85046 13970
rect 85110 13906 85126 13970
rect 85190 13906 85198 13970
rect 84878 13905 85198 13906
rect 84047 13628 84113 13631
rect 88454 13628 88934 13658
rect 84047 13626 88934 13628
rect 84047 13570 84052 13626
rect 84108 13570 88934 13626
rect 84047 13568 88934 13570
rect 84047 13565 84113 13568
rect 88454 13538 88934 13568
rect 2878 13426 3198 13427
rect 2878 13362 2886 13426
rect 2950 13362 2966 13426
rect 3030 13362 3046 13426
rect 3110 13362 3126 13426
rect 3190 13362 3198 13426
rect 2878 13361 3198 13362
rect 86878 13426 87198 13427
rect 86878 13362 86886 13426
rect 86950 13362 86966 13426
rect 87030 13362 87046 13426
rect 87110 13362 87126 13426
rect 87190 13362 87198 13426
rect 86878 13361 87198 13362
rect 878 12882 1198 12883
rect 878 12818 886 12882
rect 950 12818 966 12882
rect 1030 12818 1046 12882
rect 1110 12818 1126 12882
rect 1190 12818 1198 12882
rect 878 12817 1198 12818
rect 84878 12882 85198 12883
rect 84878 12818 84886 12882
rect 84950 12818 84966 12882
rect 85030 12818 85046 12882
rect 85110 12818 85126 12882
rect 85190 12818 85198 12882
rect 84878 12817 85198 12818
rect 83955 12540 84021 12543
rect 83955 12538 87376 12540
rect 83955 12482 83960 12538
rect 84016 12482 87376 12538
rect 83955 12480 87376 12482
rect 83955 12477 84021 12480
rect 87316 12404 87376 12480
rect 88454 12404 88934 12434
rect 87316 12344 88934 12404
rect 2878 12338 3198 12339
rect 2878 12274 2886 12338
rect 2950 12274 2966 12338
rect 3030 12274 3046 12338
rect 3110 12274 3126 12338
rect 3190 12274 3198 12338
rect 2878 12273 3198 12274
rect 86878 12338 87198 12339
rect 86878 12274 86886 12338
rect 86950 12274 86966 12338
rect 87030 12274 87046 12338
rect 87110 12274 87126 12338
rect 87190 12274 87198 12338
rect 88454 12314 88934 12344
rect 86878 12273 87198 12274
rect 878 11794 1198 11795
rect 878 11730 886 11794
rect 950 11730 966 11794
rect 1030 11730 1046 11794
rect 1110 11730 1126 11794
rect 1190 11730 1198 11794
rect 878 11729 1198 11730
rect 84878 11794 85198 11795
rect 84878 11730 84886 11794
rect 84950 11730 84966 11794
rect 85030 11730 85046 11794
rect 85110 11730 85126 11794
rect 85190 11730 85198 11794
rect 84878 11729 85198 11730
rect 2878 11250 3198 11251
rect 2878 11186 2886 11250
rect 2950 11186 2966 11250
rect 3030 11186 3046 11250
rect 3110 11186 3126 11250
rect 3190 11186 3198 11250
rect 2878 11185 3198 11186
rect 86878 11250 87198 11251
rect 86878 11186 86886 11250
rect 86950 11186 86966 11250
rect 87030 11186 87046 11250
rect 87110 11186 87126 11250
rect 87190 11186 87198 11250
rect 86878 11185 87198 11186
rect 88454 11180 88934 11210
rect 87316 11120 88934 11180
rect 85979 11044 86045 11047
rect 87316 11044 87376 11120
rect 88454 11090 88934 11120
rect 85979 11042 87376 11044
rect 85979 10986 85984 11042
rect 86040 10986 87376 11042
rect 85979 10984 87376 10986
rect 85979 10981 86045 10984
rect 878 10706 1198 10707
rect 878 10642 886 10706
rect 950 10642 966 10706
rect 1030 10642 1046 10706
rect 1110 10642 1126 10706
rect 1190 10642 1198 10706
rect 878 10641 1198 10642
rect 84878 10706 85198 10707
rect 84878 10642 84886 10706
rect 84950 10642 84966 10706
rect 85030 10642 85046 10706
rect 85110 10642 85126 10706
rect 85190 10642 85198 10706
rect 84878 10641 85198 10642
rect 2878 10162 3198 10163
rect 2878 10098 2886 10162
rect 2950 10098 2966 10162
rect 3030 10098 3046 10162
rect 3110 10098 3126 10162
rect 3190 10098 3198 10162
rect 2878 10097 3198 10098
rect 86878 10162 87198 10163
rect 86878 10098 86886 10162
rect 86950 10098 86966 10162
rect 87030 10098 87046 10162
rect 87110 10098 87126 10162
rect 87190 10098 87198 10162
rect 86878 10097 87198 10098
rect 84139 9956 84205 9959
rect 88454 9956 88934 9986
rect 84139 9954 88934 9956
rect 84139 9898 84144 9954
rect 84200 9898 88934 9954
rect 84139 9896 88934 9898
rect 84139 9893 84205 9896
rect 88454 9866 88934 9896
rect 878 9618 1198 9619
rect 878 9554 886 9618
rect 950 9554 966 9618
rect 1030 9554 1046 9618
rect 1110 9554 1126 9618
rect 1190 9554 1198 9618
rect 878 9553 1198 9554
rect 84878 9618 85198 9619
rect 84878 9554 84886 9618
rect 84950 9554 84966 9618
rect 85030 9554 85046 9618
rect 85110 9554 85126 9618
rect 85190 9554 85198 9618
rect 84878 9553 85198 9554
rect 2878 9074 3198 9075
rect 2878 9010 2886 9074
rect 2950 9010 2966 9074
rect 3030 9010 3046 9074
rect 3110 9010 3126 9074
rect 3190 9010 3198 9074
rect 2878 9009 3198 9010
rect 86878 9074 87198 9075
rect 86878 9010 86886 9074
rect 86950 9010 86966 9074
rect 87030 9010 87046 9074
rect 87110 9010 87126 9074
rect 87190 9010 87198 9074
rect 86878 9009 87198 9010
rect 82575 8868 82641 8871
rect 82759 8868 82825 8871
rect 82575 8866 82825 8868
rect 82575 8810 82580 8866
rect 82636 8810 82764 8866
rect 82820 8810 82825 8866
rect 82575 8808 82825 8810
rect 82575 8805 82641 8808
rect 82759 8805 82825 8808
rect 83495 8868 83561 8871
rect 83495 8866 83834 8868
rect 83495 8810 83500 8866
rect 83556 8810 83834 8866
rect 83495 8808 83834 8810
rect 83495 8805 83561 8808
rect 82483 8596 82549 8599
rect 83774 8596 83834 8808
rect 83955 8732 84021 8735
rect 88454 8732 88934 8762
rect 83955 8730 88934 8732
rect 83955 8674 83960 8730
rect 84016 8674 88934 8730
rect 83955 8672 88934 8674
rect 83955 8669 84021 8672
rect 88454 8642 88934 8672
rect 82483 8594 83834 8596
rect 82483 8538 82488 8594
rect 82544 8538 83834 8594
rect 82483 8536 83834 8538
rect 82483 8533 82549 8536
rect 878 8530 1198 8531
rect 878 8466 886 8530
rect 950 8466 966 8530
rect 1030 8466 1046 8530
rect 1110 8466 1126 8530
rect 1190 8466 1198 8530
rect 878 8465 1198 8466
rect 84878 8530 85198 8531
rect 84878 8466 84886 8530
rect 84950 8466 84966 8530
rect 85030 8466 85046 8530
rect 85110 8466 85126 8530
rect 85190 8466 85198 8530
rect 84878 8465 85198 8466
rect 2878 7986 3198 7987
rect 2878 7922 2886 7986
rect 2950 7922 2966 7986
rect 3030 7922 3046 7986
rect 3110 7922 3126 7986
rect 3190 7922 3198 7986
rect 2878 7921 3198 7922
rect 86878 7986 87198 7987
rect 86878 7922 86886 7986
rect 86950 7922 86966 7986
rect 87030 7922 87046 7986
rect 87110 7922 87126 7986
rect 87190 7922 87198 7986
rect 86878 7921 87198 7922
rect 85059 7644 85125 7647
rect 88454 7644 88934 7674
rect 85059 7642 88934 7644
rect 85059 7586 85064 7642
rect 85120 7586 88934 7642
rect 85059 7584 88934 7586
rect 85059 7581 85125 7584
rect 88454 7554 88934 7584
rect 878 7442 1198 7443
rect 878 7378 886 7442
rect 950 7378 966 7442
rect 1030 7378 1046 7442
rect 1110 7378 1126 7442
rect 1190 7378 1198 7442
rect 878 7377 1198 7378
rect 84878 7442 85198 7443
rect 84878 7378 84886 7442
rect 84950 7378 84966 7442
rect 85030 7378 85046 7442
rect 85110 7378 85126 7442
rect 85190 7378 85198 7442
rect 84878 7377 85198 7378
rect 2878 6898 3198 6899
rect 2878 6834 2886 6898
rect 2950 6834 2966 6898
rect 3030 6834 3046 6898
rect 3110 6834 3126 6898
rect 3190 6834 3198 6898
rect 2878 6833 3198 6834
rect 86878 6898 87198 6899
rect 86878 6834 86886 6898
rect 86950 6834 86966 6898
rect 87030 6834 87046 6898
rect 87110 6834 87126 6898
rect 87190 6834 87198 6898
rect 86878 6833 87198 6834
rect 84507 6556 84573 6559
rect 84507 6554 85352 6556
rect 84507 6498 84512 6554
rect 84568 6498 85352 6554
rect 84507 6496 85352 6498
rect 84507 6493 84573 6496
rect 85292 6420 85352 6496
rect 88454 6420 88934 6450
rect 85292 6360 88934 6420
rect 878 6354 1198 6355
rect 878 6290 886 6354
rect 950 6290 966 6354
rect 1030 6290 1046 6354
rect 1110 6290 1126 6354
rect 1190 6290 1198 6354
rect 878 6289 1198 6290
rect 84878 6354 85198 6355
rect 84878 6290 84886 6354
rect 84950 6290 84966 6354
rect 85030 6290 85046 6354
rect 85110 6290 85126 6354
rect 85190 6290 85198 6354
rect 88454 6330 88934 6360
rect 84878 6289 85198 6290
rect 82340 6086 82346 6150
rect 82410 6148 82416 6150
rect 82667 6148 82733 6151
rect 82410 6146 82733 6148
rect 82410 6090 82672 6146
rect 82728 6090 82733 6146
rect 82410 6088 82733 6090
rect 82410 6086 82416 6088
rect 82667 6085 82733 6088
rect 2878 5810 3198 5811
rect 2878 5746 2886 5810
rect 2950 5746 2966 5810
rect 3030 5746 3046 5810
rect 3110 5746 3126 5810
rect 3190 5746 3198 5810
rect 2878 5745 3198 5746
rect 86878 5810 87198 5811
rect 86878 5746 86886 5810
rect 86950 5746 86966 5810
rect 87030 5746 87046 5810
rect 87110 5746 87126 5810
rect 87190 5746 87198 5810
rect 86878 5745 87198 5746
rect 878 5266 1198 5267
rect 878 5202 886 5266
rect 950 5202 966 5266
rect 1030 5202 1046 5266
rect 1110 5202 1126 5266
rect 1190 5202 1198 5266
rect 878 5201 1198 5202
rect 84878 5266 85198 5267
rect 84878 5202 84886 5266
rect 84950 5202 84966 5266
rect 85030 5202 85046 5266
rect 85110 5202 85126 5266
rect 85190 5202 85198 5266
rect 84878 5201 85198 5202
rect 3639 5198 3705 5199
rect 3588 5134 3594 5198
rect 3658 5196 3705 5198
rect 88454 5196 88934 5226
rect 3658 5194 3750 5196
rect 3700 5138 3750 5194
rect 3658 5136 3750 5138
rect 85292 5136 88934 5196
rect 3658 5134 3705 5136
rect 3639 5133 3705 5134
rect 84139 5060 84205 5063
rect 85292 5060 85352 5136
rect 88454 5106 88934 5136
rect 84139 5058 85352 5060
rect 84139 5002 84144 5058
rect 84200 5002 85352 5058
rect 84139 5000 85352 5002
rect 84139 4997 84205 5000
rect 2878 4722 3198 4723
rect 2878 4658 2886 4722
rect 2950 4658 2966 4722
rect 3030 4658 3046 4722
rect 3110 4658 3126 4722
rect 3190 4658 3198 4722
rect 2878 4657 3198 4658
rect 86878 4722 87198 4723
rect 86878 4658 86886 4722
rect 86950 4658 86966 4722
rect 87030 4658 87046 4722
rect 87110 4658 87126 4722
rect 87190 4658 87198 4722
rect 86878 4657 87198 4658
rect 4140 4590 4146 4654
rect 4210 4652 4216 4654
rect 4375 4652 4441 4655
rect 4508 4652 4514 4654
rect 4210 4650 4514 4652
rect 4210 4594 4380 4650
rect 4436 4594 4514 4650
rect 4210 4592 4514 4594
rect 4210 4590 4216 4592
rect 4375 4589 4441 4592
rect 4508 4590 4514 4592
rect 4578 4590 4584 4654
rect 2903 4244 2969 4247
rect 4140 4244 4146 4246
rect 2903 4242 4146 4244
rect 2903 4186 2908 4242
rect 2964 4186 4146 4242
rect 2903 4184 4146 4186
rect 2903 4181 2969 4184
rect 4140 4182 4146 4184
rect 4210 4182 4216 4246
rect 878 4178 1198 4179
rect 878 4114 886 4178
rect 950 4114 966 4178
rect 1030 4114 1046 4178
rect 1110 4114 1126 4178
rect 1190 4114 1198 4178
rect 878 4113 1198 4114
rect 84878 4178 85198 4179
rect 84878 4114 84886 4178
rect 84950 4114 84966 4178
rect 85030 4114 85046 4178
rect 85110 4114 85126 4178
rect 85190 4114 85198 4178
rect 84878 4113 85198 4114
rect 83771 4110 83837 4111
rect 83771 4108 83818 4110
rect 83726 4106 83818 4108
rect 83726 4050 83776 4106
rect 83726 4048 83818 4050
rect 83771 4046 83818 4048
rect 83882 4046 83888 4110
rect 83771 4045 83837 4046
rect 84047 3972 84113 3975
rect 88454 3972 88934 4002
rect 84047 3970 88934 3972
rect 84047 3914 84052 3970
rect 84108 3914 88934 3970
rect 84047 3912 88934 3914
rect 84047 3909 84113 3912
rect 88454 3882 88934 3912
rect 82759 3836 82825 3839
rect 82892 3836 82898 3838
rect 82759 3834 82898 3836
rect 82759 3778 82764 3834
rect 82820 3778 82898 3834
rect 82759 3776 82898 3778
rect 82759 3773 82825 3776
rect 82892 3774 82898 3776
rect 82962 3774 82968 3838
rect 2878 3634 3198 3635
rect 2878 3570 2886 3634
rect 2950 3570 2966 3634
rect 3030 3570 3046 3634
rect 3110 3570 3126 3634
rect 3190 3570 3198 3634
rect 2878 3569 3198 3570
rect 86878 3634 87198 3635
rect 86878 3570 86886 3634
rect 86950 3570 86966 3634
rect 87030 3570 87046 3634
rect 87110 3570 87126 3634
rect 87190 3570 87198 3634
rect 86878 3569 87198 3570
rect 3271 3564 3337 3567
rect 3404 3564 3410 3566
rect 3271 3562 3410 3564
rect 3271 3506 3276 3562
rect 3332 3506 3410 3562
rect 3271 3504 3410 3506
rect 3271 3501 3337 3504
rect 3404 3502 3410 3504
rect 3474 3502 3480 3566
rect 1799 3292 1865 3295
rect 4375 3292 4441 3295
rect 1799 3290 4441 3292
rect 1799 3234 1804 3290
rect 1860 3234 4380 3290
rect 4436 3234 4441 3290
rect 1799 3232 4441 3234
rect 1799 3229 1865 3232
rect 4375 3229 4441 3232
rect 81471 3292 81537 3295
rect 84548 3292 84554 3294
rect 81471 3290 84554 3292
rect 81471 3234 81476 3290
rect 81532 3234 84554 3290
rect 81471 3232 84554 3234
rect 81471 3229 81537 3232
rect 84548 3230 84554 3232
rect 84618 3230 84624 3294
rect 2995 3156 3061 3159
rect 3772 3156 3778 3158
rect 2995 3154 3778 3156
rect 2995 3098 3000 3154
rect 3056 3098 3778 3154
rect 2995 3096 3778 3098
rect 2995 3093 3061 3096
rect 3772 3094 3778 3096
rect 3842 3094 3848 3158
rect 81379 3156 81445 3159
rect 84364 3156 84370 3158
rect 81379 3154 84370 3156
rect 81379 3098 81384 3154
rect 81440 3098 84370 3154
rect 81379 3096 84370 3098
rect 81379 3093 81445 3096
rect 84364 3094 84370 3096
rect 84434 3094 84440 3158
rect 878 3090 1198 3091
rect 878 3026 886 3090
rect 950 3026 966 3090
rect 1030 3026 1046 3090
rect 1110 3026 1126 3090
rect 1190 3026 1198 3090
rect 878 3025 1198 3026
rect 84878 3090 85198 3091
rect 84878 3026 84886 3090
rect 84950 3026 84966 3090
rect 85030 3026 85046 3090
rect 85110 3026 85126 3090
rect 85190 3026 85198 3090
rect 84878 3025 85198 3026
rect 2443 3020 2509 3023
rect 39100 3020 39106 3022
rect 2443 3018 39106 3020
rect 2443 2962 2448 3018
rect 2504 2962 39106 3018
rect 2443 2960 39106 2962
rect 2443 2957 2509 2960
rect 39100 2958 39106 2960
rect 39170 2958 39176 3022
rect 42964 2958 42970 3022
rect 43034 3020 43040 3022
rect 82667 3020 82733 3023
rect 43034 3018 82733 3020
rect 43034 2962 82672 3018
rect 82728 2962 82733 3018
rect 43034 2960 82733 2962
rect 43034 2958 43040 2960
rect 82667 2957 82733 2960
rect 1339 2884 1405 2887
rect 19739 2886 19805 2887
rect 13524 2884 13530 2886
rect 1339 2882 13530 2884
rect 1339 2826 1344 2882
rect 1400 2826 13530 2882
rect 1339 2824 13530 2826
rect 1339 2821 1405 2824
rect 13524 2822 13530 2824
rect 13594 2822 13600 2886
rect 19739 2884 19786 2886
rect 19694 2882 19786 2884
rect 19694 2826 19744 2882
rect 19694 2824 19786 2826
rect 19739 2822 19786 2824
rect 19850 2822 19856 2886
rect 21988 2822 21994 2886
rect 22058 2884 22064 2886
rect 22131 2884 22197 2887
rect 23971 2886 24037 2887
rect 25075 2886 25141 2887
rect 27467 2886 27533 2887
rect 31055 2886 31121 2887
rect 33723 2886 33789 2887
rect 36943 2886 37009 2887
rect 23971 2884 24018 2886
rect 22058 2882 22197 2884
rect 22058 2826 22136 2882
rect 22192 2826 22197 2882
rect 22058 2824 22197 2826
rect 23926 2882 24018 2884
rect 23926 2826 23976 2882
rect 23926 2824 24018 2826
rect 22058 2822 22064 2824
rect 19739 2821 19805 2822
rect 22131 2821 22197 2824
rect 23971 2822 24018 2824
rect 24082 2822 24088 2886
rect 25075 2884 25122 2886
rect 25030 2882 25122 2884
rect 25030 2826 25080 2882
rect 25030 2824 25122 2826
rect 25075 2822 25122 2824
rect 25186 2822 25192 2886
rect 27467 2884 27514 2886
rect 27422 2882 27514 2884
rect 27422 2826 27472 2882
rect 27422 2824 27514 2826
rect 27467 2822 27514 2824
rect 27578 2822 27584 2886
rect 31050 2884 31056 2886
rect 30964 2824 31056 2884
rect 31050 2822 31056 2824
rect 31120 2822 31126 2886
rect 33718 2884 33724 2886
rect 33632 2824 33724 2884
rect 33718 2822 33724 2824
rect 33788 2822 33794 2886
rect 36892 2822 36898 2886
rect 36962 2884 37009 2886
rect 38783 2884 38849 2887
rect 41359 2886 41425 2887
rect 38916 2884 38922 2886
rect 36962 2882 37054 2884
rect 37004 2826 37054 2882
rect 36962 2824 37054 2826
rect 38783 2882 38922 2884
rect 38783 2826 38788 2882
rect 38844 2826 38922 2882
rect 38783 2824 38922 2826
rect 36962 2822 37009 2824
rect 23971 2821 24037 2822
rect 25075 2821 25141 2822
rect 27467 2821 27533 2822
rect 31055 2821 31121 2822
rect 33723 2821 33789 2822
rect 36943 2821 37009 2822
rect 38783 2821 38849 2824
rect 38916 2822 38922 2824
rect 38986 2822 38992 2886
rect 41308 2822 41314 2886
rect 41378 2884 41425 2886
rect 41378 2882 41470 2884
rect 41420 2826 41470 2882
rect 41378 2824 41470 2826
rect 41378 2822 41425 2824
rect 44252 2822 44258 2886
rect 44322 2884 44328 2886
rect 82524 2884 82530 2886
rect 44322 2824 82530 2884
rect 44322 2822 44328 2824
rect 82524 2822 82530 2824
rect 82594 2884 82600 2886
rect 83771 2884 83837 2887
rect 82594 2882 83837 2884
rect 82594 2826 83776 2882
rect 83832 2826 83837 2882
rect 82594 2824 83837 2826
rect 82594 2822 82600 2824
rect 41359 2821 41425 2822
rect 83771 2821 83837 2824
rect 2719 2748 2785 2751
rect 4375 2748 4441 2751
rect 37076 2748 37082 2750
rect 2719 2746 4162 2748
rect 2719 2690 2724 2746
rect 2780 2690 4162 2746
rect 2719 2688 4162 2690
rect 2719 2685 2785 2688
rect 4102 2612 4162 2688
rect 4375 2746 37082 2748
rect 4375 2690 4380 2746
rect 4436 2690 37082 2746
rect 4375 2688 37082 2690
rect 4375 2685 4441 2688
rect 37076 2686 37082 2688
rect 37146 2686 37152 2750
rect 45356 2686 45362 2750
rect 45426 2748 45432 2750
rect 78067 2748 78133 2751
rect 45426 2746 78133 2748
rect 45426 2690 78072 2746
rect 78128 2690 78133 2746
rect 45426 2688 78133 2690
rect 45426 2686 45432 2688
rect 78067 2685 78133 2688
rect 81287 2748 81353 2751
rect 88454 2748 88934 2778
rect 81287 2746 88934 2748
rect 81287 2690 81292 2746
rect 81348 2690 88934 2746
rect 81287 2688 88934 2690
rect 81287 2685 81353 2688
rect 88454 2658 88934 2688
rect 4743 2612 4809 2615
rect 19463 2612 19529 2615
rect 24615 2612 24681 2615
rect 50191 2614 50257 2615
rect 53687 2614 53753 2615
rect 4102 2610 19529 2612
rect 4102 2554 4748 2610
rect 4804 2554 19468 2610
rect 19524 2554 19529 2610
rect 4102 2552 19529 2554
rect 4743 2549 4809 2552
rect 19463 2549 19529 2552
rect 24584 2610 24681 2612
rect 24584 2554 24620 2610
rect 24676 2554 24681 2610
rect 24584 2549 24681 2554
rect 48852 2550 48858 2614
rect 48922 2550 48928 2614
rect 50140 2612 50146 2614
rect 50100 2552 50146 2612
rect 50210 2610 50257 2614
rect 53636 2612 53642 2614
rect 50252 2554 50257 2610
rect 50140 2550 50146 2552
rect 50210 2550 50257 2554
rect 53596 2552 53642 2612
rect 53706 2610 53753 2614
rect 83495 2612 83561 2615
rect 84231 2612 84297 2615
rect 53748 2554 53753 2610
rect 53636 2550 53642 2552
rect 53706 2550 53753 2554
rect 2878 2546 3198 2547
rect 2878 2482 2886 2546
rect 2950 2482 2966 2546
rect 3030 2482 3046 2546
rect 3110 2482 3126 2546
rect 3190 2482 3198 2546
rect 2878 2481 3198 2482
rect 7871 2476 7937 2479
rect 24584 2476 24644 2549
rect 25995 2476 26061 2479
rect 7871 2474 12304 2476
rect 7871 2418 7876 2474
rect 7932 2418 12304 2474
rect 7871 2416 12304 2418
rect 24584 2474 26061 2476
rect 24584 2418 26000 2474
rect 26056 2418 26061 2474
rect 24584 2416 26061 2418
rect 48860 2476 48920 2550
rect 50191 2549 50257 2550
rect 53687 2549 53753 2550
rect 55668 2552 68608 2612
rect 55668 2476 55728 2552
rect 48860 2416 55728 2476
rect 7871 2413 7937 2416
rect 12244 2340 12304 2416
rect 25995 2413 26061 2416
rect 18267 2342 18333 2343
rect 18267 2340 18314 2342
rect 12244 2280 18146 2340
rect 18222 2338 18314 2340
rect 18222 2282 18272 2338
rect 18222 2280 18314 2282
rect 18086 2204 18146 2280
rect 18267 2278 18314 2280
rect 18378 2278 18384 2342
rect 28387 2340 28453 2343
rect 54239 2342 54305 2343
rect 34868 2340 34874 2342
rect 26044 2280 26610 2340
rect 18267 2277 18333 2278
rect 19371 2204 19437 2207
rect 18086 2202 19437 2204
rect 18086 2146 19376 2202
rect 19432 2146 19437 2202
rect 18086 2144 19437 2146
rect 19371 2141 19437 2144
rect 19555 2204 19621 2207
rect 26044 2204 26104 2280
rect 26363 2206 26429 2207
rect 26363 2204 26410 2206
rect 19555 2202 26104 2204
rect 19555 2146 19560 2202
rect 19616 2146 26104 2202
rect 19555 2144 26104 2146
rect 26318 2202 26410 2204
rect 26318 2146 26368 2202
rect 26318 2144 26410 2146
rect 19555 2141 19621 2144
rect 26363 2142 26410 2144
rect 26474 2142 26480 2206
rect 26550 2204 26610 2280
rect 28387 2338 34874 2340
rect 28387 2282 28392 2338
rect 28448 2282 34874 2338
rect 28387 2280 34874 2282
rect 28387 2277 28453 2280
rect 34868 2278 34874 2280
rect 34938 2278 34944 2342
rect 54188 2278 54194 2342
rect 54258 2340 54305 2342
rect 68548 2340 68608 2552
rect 77380 2610 83561 2612
rect 77380 2554 83500 2610
rect 83556 2554 83561 2610
rect 77380 2552 83561 2554
rect 77380 2340 77440 2552
rect 83495 2549 83561 2552
rect 83820 2610 84297 2612
rect 83820 2554 84236 2610
rect 84292 2554 84297 2610
rect 83820 2552 84297 2554
rect 78067 2476 78133 2479
rect 83820 2476 83880 2552
rect 84231 2549 84297 2552
rect 86878 2546 87198 2547
rect 86878 2482 86886 2546
rect 86950 2482 86966 2546
rect 87030 2482 87046 2546
rect 87110 2482 87126 2546
rect 87190 2482 87198 2546
rect 86878 2481 87198 2482
rect 78067 2474 83880 2476
rect 78067 2418 78072 2474
rect 78128 2418 83880 2474
rect 78067 2416 83880 2418
rect 83955 2478 84021 2479
rect 83955 2474 84002 2478
rect 84066 2476 84072 2478
rect 83955 2418 83960 2474
rect 78067 2413 78133 2416
rect 83955 2414 84002 2418
rect 84066 2416 84112 2476
rect 84066 2414 84072 2416
rect 83955 2413 84021 2414
rect 54258 2338 54350 2340
rect 54300 2282 54350 2338
rect 54258 2280 54350 2282
rect 68548 2280 77440 2340
rect 54258 2278 54305 2280
rect 82708 2278 82714 2342
rect 82778 2340 82784 2342
rect 83495 2340 83561 2343
rect 82778 2338 83561 2340
rect 82778 2282 83500 2338
rect 83556 2282 83561 2338
rect 82778 2280 83561 2282
rect 82778 2278 82784 2280
rect 54239 2277 54305 2278
rect 83495 2277 83561 2280
rect 35011 2204 35077 2207
rect 41819 2206 41885 2207
rect 45223 2206 45289 2207
rect 46695 2206 46761 2207
rect 41819 2204 41866 2206
rect 26550 2202 35077 2204
rect 26550 2146 35016 2202
rect 35072 2146 35077 2202
rect 26550 2144 35077 2146
rect 41774 2202 41866 2204
rect 41774 2146 41824 2202
rect 41774 2144 41866 2146
rect 26363 2141 26429 2142
rect 35011 2141 35077 2144
rect 41819 2142 41866 2144
rect 41930 2142 41936 2206
rect 45172 2204 45178 2206
rect 45132 2144 45178 2204
rect 45242 2202 45289 2206
rect 45284 2146 45289 2202
rect 45172 2142 45178 2144
rect 45242 2142 45289 2146
rect 46644 2142 46650 2206
rect 46714 2204 46761 2206
rect 46714 2202 46806 2204
rect 46756 2146 46806 2202
rect 46714 2144 46806 2146
rect 46714 2142 46761 2144
rect 47564 2142 47570 2206
rect 47634 2204 47640 2206
rect 47891 2204 47957 2207
rect 49823 2206 49889 2207
rect 47634 2202 47957 2204
rect 47634 2146 47896 2202
rect 47952 2146 47957 2202
rect 47634 2144 47957 2146
rect 47634 2142 47640 2144
rect 41819 2141 41885 2142
rect 45223 2141 45289 2142
rect 46695 2141 46761 2142
rect 47891 2141 47957 2144
rect 49772 2142 49778 2206
rect 49842 2204 49889 2206
rect 50007 2204 50073 2207
rect 83996 2204 84002 2206
rect 49842 2202 49934 2204
rect 49884 2146 49934 2202
rect 49842 2144 49934 2146
rect 50007 2202 84002 2204
rect 50007 2146 50012 2202
rect 50068 2146 84002 2202
rect 50007 2144 84002 2146
rect 49842 2142 49889 2144
rect 49823 2141 49889 2142
rect 50007 2141 50073 2144
rect 83996 2142 84002 2144
rect 84066 2142 84072 2206
rect 4007 2068 4073 2071
rect 84139 2068 84205 2071
rect 4007 2066 84205 2068
rect 4007 2010 4012 2066
rect 4068 2010 84144 2066
rect 84200 2010 84205 2066
rect 4007 2008 84205 2010
rect 4007 2005 4073 2008
rect 84139 2005 84205 2008
rect 878 2002 1198 2003
rect 878 1938 886 2002
rect 950 1938 966 2002
rect 1030 1938 1046 2002
rect 1110 1938 1126 2002
rect 1190 1938 1198 2002
rect 878 1937 1198 1938
rect 84878 2002 85198 2003
rect 84878 1938 84886 2002
rect 84950 1938 84966 2002
rect 85030 1938 85046 2002
rect 85110 1938 85126 2002
rect 85190 1938 85198 2002
rect 84878 1937 85198 1938
rect 4191 1932 4257 1935
rect 84507 1932 84573 1935
rect 4191 1930 84573 1932
rect 4191 1874 4196 1930
rect 4252 1874 84512 1930
rect 84568 1874 84573 1930
rect 4191 1872 84573 1874
rect 4191 1869 4257 1872
rect 84507 1869 84573 1872
rect 3731 1796 3797 1799
rect 82575 1796 82641 1799
rect 3731 1794 82641 1796
rect 3731 1738 3736 1794
rect 3792 1738 82580 1794
rect 82636 1738 82641 1794
rect 3731 1736 82641 1738
rect 3731 1733 3797 1736
rect 82575 1733 82641 1736
rect 8699 1662 8765 1663
rect 22407 1662 22473 1663
rect 24707 1662 24773 1663
rect 29215 1662 29281 1663
rect 36299 1662 36365 1663
rect 8699 1658 8735 1662
rect 8799 1660 8805 1662
rect 22364 1660 22370 1662
rect 8699 1602 8704 1658
rect 8699 1598 8735 1602
rect 8799 1600 8856 1660
rect 22316 1600 22370 1660
rect 22434 1658 22473 1662
rect 24700 1660 24706 1662
rect 22468 1602 22473 1658
rect 8799 1598 8805 1600
rect 22364 1598 22370 1600
rect 22434 1598 22473 1602
rect 24616 1600 24706 1660
rect 24700 1598 24706 1600
rect 24770 1598 24776 1662
rect 29215 1660 29254 1662
rect 29162 1658 29254 1660
rect 29162 1602 29220 1658
rect 29162 1600 29254 1602
rect 29215 1598 29254 1600
rect 29318 1598 29324 1662
rect 36256 1598 36262 1662
rect 36326 1660 36365 1662
rect 36483 1660 36549 1663
rect 80735 1660 80801 1663
rect 84180 1660 84186 1662
rect 36326 1658 36418 1660
rect 36360 1602 36418 1658
rect 36326 1600 36418 1602
rect 36483 1658 80801 1660
rect 36483 1602 36488 1658
rect 36544 1602 80740 1658
rect 80796 1602 80801 1658
rect 36483 1600 80801 1602
rect 36326 1598 36365 1600
rect 8699 1597 8765 1598
rect 22407 1597 22473 1598
rect 24707 1597 24773 1598
rect 29215 1597 29281 1598
rect 36299 1597 36365 1598
rect 36483 1597 36549 1600
rect 80735 1597 80801 1600
rect 80876 1600 84186 1660
rect 3455 1524 3521 1527
rect 80876 1524 80936 1600
rect 84180 1598 84186 1600
rect 84250 1598 84256 1662
rect 3455 1522 80936 1524
rect 3455 1466 3460 1522
rect 3516 1466 80936 1522
rect 3455 1464 80936 1466
rect 83955 1524 84021 1527
rect 88454 1524 88934 1554
rect 83955 1522 88934 1524
rect 83955 1466 83960 1522
rect 84016 1466 88934 1522
rect 83955 1464 88934 1466
rect 3455 1461 3521 1464
rect 83955 1461 84021 1464
rect 88454 1434 88934 1464
rect 33079 1388 33145 1391
rect 36483 1388 36549 1391
rect 42279 1390 42345 1391
rect 42228 1388 42234 1390
rect 33079 1386 36549 1388
rect 33079 1330 33084 1386
rect 33140 1330 36488 1386
rect 36544 1330 36549 1386
rect 33079 1328 36549 1330
rect 42188 1328 42234 1388
rect 42298 1386 42345 1390
rect 42340 1330 42345 1386
rect 33079 1325 33145 1328
rect 36483 1325 36549 1328
rect 42228 1326 42234 1328
rect 42298 1326 42345 1330
rect 42279 1325 42345 1326
rect 42463 1388 42529 1391
rect 50007 1388 50073 1391
rect 51479 1390 51545 1391
rect 42463 1386 50073 1388
rect 42463 1330 42468 1386
rect 42524 1330 50012 1386
rect 50068 1330 50073 1386
rect 42463 1328 50073 1330
rect 42463 1325 42529 1328
rect 50007 1325 50073 1328
rect 51428 1326 51434 1390
rect 51498 1388 51545 1390
rect 80735 1388 80801 1391
rect 84732 1388 84738 1390
rect 51498 1386 51590 1388
rect 51540 1330 51590 1386
rect 51498 1328 51590 1330
rect 80735 1386 84738 1388
rect 80735 1330 80740 1386
rect 80796 1330 84738 1386
rect 80735 1328 84738 1330
rect 51498 1326 51545 1328
rect 51479 1325 51545 1326
rect 80735 1325 80801 1328
rect 84732 1326 84738 1328
rect 84802 1326 84808 1390
rect 27140 1054 27146 1118
rect 27210 1116 27216 1118
rect 83628 1116 83634 1118
rect 27210 1056 83634 1116
rect 27210 1054 27216 1056
rect 83628 1054 83634 1056
rect 83698 1054 83704 1118
rect 11643 982 11709 983
rect 11643 980 11690 982
rect 11598 978 11690 980
rect 11598 922 11648 978
rect 11598 920 11690 922
rect 11643 918 11690 920
rect 11754 918 11760 982
rect 11827 980 11893 983
rect 12236 980 12242 982
rect 11827 978 12242 980
rect 11827 922 11832 978
rect 11888 922 12242 978
rect 11827 920 12242 922
rect 11643 917 11709 918
rect 11827 917 11893 920
rect 12236 918 12242 920
rect 12306 918 12312 982
rect 14403 980 14469 983
rect 15180 980 15186 982
rect 14403 978 15186 980
rect 14403 922 14408 978
rect 14464 922 15186 978
rect 14403 920 15186 922
rect 14403 917 14469 920
rect 15180 918 15186 920
rect 15250 918 15256 982
rect 16979 980 17045 983
rect 17572 980 17578 982
rect 16979 978 17578 980
rect 16979 922 16984 978
rect 17040 922 17578 978
rect 16979 920 17578 922
rect 16979 917 17045 920
rect 17572 918 17578 920
rect 17642 918 17648 982
rect 17756 918 17762 982
rect 17826 980 17832 982
rect 18083 980 18149 983
rect 18911 982 18977 983
rect 18860 980 18866 982
rect 17826 978 18149 980
rect 17826 922 18088 978
rect 18144 922 18149 978
rect 17826 920 18149 922
rect 18820 920 18866 980
rect 18930 978 18977 982
rect 18972 922 18977 978
rect 17826 918 17832 920
rect 18083 917 18149 920
rect 18860 918 18866 920
rect 18930 918 18977 922
rect 18911 917 18977 918
rect 20843 980 20909 983
rect 21303 982 21369 983
rect 21068 980 21074 982
rect 20843 978 21074 980
rect 20843 922 20848 978
rect 20904 922 21074 978
rect 20843 920 21074 922
rect 20843 917 20909 920
rect 21068 918 21074 920
rect 21138 918 21144 982
rect 21252 980 21258 982
rect 21212 920 21258 980
rect 21322 978 21369 982
rect 23419 982 23485 983
rect 24247 982 24313 983
rect 28295 982 28361 983
rect 29399 982 29465 983
rect 31055 982 31121 983
rect 23419 980 23466 982
rect 21364 922 21369 978
rect 21252 918 21258 920
rect 21322 918 21369 922
rect 23374 978 23466 980
rect 23374 922 23424 978
rect 23374 920 23466 922
rect 21303 917 21369 918
rect 23419 918 23466 920
rect 23530 918 23536 982
rect 24196 980 24202 982
rect 24156 920 24202 980
rect 24266 978 24313 982
rect 28244 980 28250 982
rect 24308 922 24313 978
rect 24196 918 24202 920
rect 24266 918 24313 922
rect 28204 920 28250 980
rect 28314 978 28361 982
rect 29348 980 29354 982
rect 28356 922 28361 978
rect 28244 918 28250 920
rect 28314 918 28361 922
rect 29308 920 29354 980
rect 29418 978 29465 982
rect 31004 980 31010 982
rect 29460 922 29465 978
rect 29348 918 29354 920
rect 29418 918 29465 922
rect 30964 920 31010 980
rect 31074 978 31121 982
rect 31116 922 31121 978
rect 31004 918 31010 920
rect 31074 918 31121 922
rect 31740 918 31746 982
rect 31810 980 31816 982
rect 31883 980 31949 983
rect 32895 982 32961 983
rect 34735 982 34801 983
rect 35287 982 35353 983
rect 32844 980 32850 982
rect 31810 978 31949 980
rect 31810 922 31888 978
rect 31944 922 31949 978
rect 31810 920 31949 922
rect 32804 920 32850 980
rect 32914 978 32961 982
rect 34684 980 34690 982
rect 32956 922 32961 978
rect 31810 918 31816 920
rect 23419 917 23485 918
rect 24247 917 24313 918
rect 28295 917 28361 918
rect 29399 917 29465 918
rect 31055 917 31121 918
rect 31883 917 31949 920
rect 32844 918 32850 920
rect 32914 918 32961 922
rect 34644 920 34690 980
rect 34754 978 34801 982
rect 35236 980 35242 982
rect 34796 922 34801 978
rect 34684 918 34690 920
rect 34754 918 34801 922
rect 35196 920 35242 980
rect 35306 978 35353 982
rect 35348 922 35353 978
rect 35236 918 35242 920
rect 35306 918 35353 922
rect 38180 918 38186 982
rect 38250 980 38256 982
rect 38323 980 38389 983
rect 40071 982 40137 983
rect 43935 982 44001 983
rect 40020 980 40026 982
rect 38250 978 38389 980
rect 38250 922 38328 978
rect 38384 922 38389 978
rect 38250 920 38389 922
rect 39980 920 40026 980
rect 40090 978 40137 982
rect 43884 980 43890 982
rect 40132 922 40137 978
rect 38250 918 38256 920
rect 32895 917 32961 918
rect 34735 917 34801 918
rect 35287 917 35353 918
rect 38323 917 38389 920
rect 40020 918 40026 920
rect 40090 918 40137 922
rect 43844 920 43890 980
rect 43954 978 44001 982
rect 43996 922 44001 978
rect 43884 918 43890 920
rect 43954 918 44001 922
rect 45724 918 45730 982
rect 45794 980 45800 982
rect 46143 980 46209 983
rect 45794 978 46209 980
rect 45794 922 46148 978
rect 46204 922 46209 978
rect 45794 920 46209 922
rect 45794 918 45800 920
rect 40071 917 40137 918
rect 43935 917 44001 918
rect 46143 917 46209 920
rect 47932 918 47938 982
rect 48002 980 48008 982
rect 50467 980 50533 983
rect 48002 978 50533 980
rect 48002 922 50472 978
rect 50528 922 50533 978
rect 48002 920 50533 922
rect 48002 918 48008 920
rect 50467 917 50533 920
rect 4508 782 4514 846
rect 4578 844 4584 846
rect 40940 844 40946 846
rect 4578 784 40946 844
rect 4578 782 4584 784
rect 40940 782 40946 784
rect 41010 782 41016 846
rect 48116 782 48122 846
rect 48186 844 48192 846
rect 81747 844 81813 847
rect 48186 842 81813 844
rect 48186 786 81752 842
rect 81808 786 81813 842
rect 48186 784 81813 786
rect 48186 782 48192 784
rect 81747 781 81813 784
rect 20751 710 20817 711
rect 4140 646 4146 710
rect 4210 708 4216 710
rect 15732 708 15738 710
rect 4210 648 15738 708
rect 4210 646 4216 648
rect 15732 646 15738 648
rect 15802 646 15808 710
rect 20700 708 20706 710
rect 20660 648 20706 708
rect 20770 706 20817 710
rect 29859 710 29925 711
rect 29859 708 29906 710
rect 20812 650 20817 706
rect 20700 646 20706 648
rect 20770 646 20817 650
rect 29814 706 29906 708
rect 29814 650 29864 706
rect 29814 648 29906 650
rect 20751 645 20817 646
rect 29859 646 29906 648
rect 29970 646 29976 710
rect 51612 646 51618 710
rect 51682 708 51688 710
rect 83260 708 83266 710
rect 51682 648 83266 708
rect 51682 646 51688 648
rect 83260 646 83266 648
rect 83330 646 83336 710
rect 29859 645 29925 646
rect 32435 574 32501 575
rect 32435 572 32482 574
rect 32390 570 32482 572
rect 32390 514 32440 570
rect 32390 512 32482 514
rect 32435 510 32482 512
rect 32546 510 32552 574
rect 52716 510 52722 574
rect 52786 572 52792 574
rect 82759 572 82825 575
rect 52786 570 82825 572
rect 52786 514 82764 570
rect 82820 514 82825 570
rect 52786 512 82825 514
rect 52786 510 52792 512
rect 32435 509 32501 510
rect 82759 509 82825 512
rect 38047 436 38113 439
rect 38548 436 38554 438
rect 38047 434 38554 436
rect 38047 378 38052 434
rect 38108 378 38554 434
rect 38047 376 38554 378
rect 38047 373 38113 376
rect 38548 374 38554 376
rect 38618 374 38624 438
rect 52900 374 52906 438
rect 52970 436 52976 438
rect 83444 436 83450 438
rect 52970 376 83450 436
rect 52970 374 52976 376
rect 83444 374 83450 376
rect 83514 374 83520 438
rect 83955 436 84021 439
rect 88454 436 88934 466
rect 83955 434 88934 436
rect 83955 378 83960 434
rect 84016 378 88934 434
rect 83955 376 88934 378
rect 83955 373 84021 376
rect 88454 346 88934 376
rect 50324 238 50330 302
rect 50394 300 50400 302
rect 81287 300 81353 303
rect 50394 298 81353 300
rect 50394 242 81292 298
rect 81348 242 81353 298
rect 50394 240 81353 242
rect 50394 238 50400 240
rect 81287 237 81353 240
rect 25852 102 25858 166
rect 25922 164 25928 166
rect 81195 164 81261 167
rect 25922 162 81261 164
rect 25922 106 81200 162
rect 81256 106 81261 162
rect 25922 104 81261 106
rect 25922 102 25928 104
rect 81195 101 81261 104
<< via3 >>
rect 5250 187918 5314 187982
rect 2886 187502 2950 187506
rect 2886 187446 2890 187502
rect 2890 187446 2946 187502
rect 2946 187446 2950 187502
rect 2886 187442 2950 187446
rect 2966 187502 3030 187506
rect 2966 187446 2970 187502
rect 2970 187446 3026 187502
rect 3026 187446 3030 187502
rect 2966 187442 3030 187446
rect 3046 187502 3110 187506
rect 3046 187446 3050 187502
rect 3050 187446 3106 187502
rect 3106 187446 3110 187502
rect 3046 187442 3110 187446
rect 3126 187502 3190 187506
rect 3126 187446 3130 187502
rect 3130 187446 3186 187502
rect 3186 187446 3190 187502
rect 3126 187442 3190 187446
rect 86886 187502 86950 187506
rect 86886 187446 86890 187502
rect 86890 187446 86946 187502
rect 86946 187446 86950 187502
rect 86886 187442 86950 187446
rect 86966 187502 87030 187506
rect 86966 187446 86970 187502
rect 86970 187446 87026 187502
rect 87026 187446 87030 187502
rect 86966 187442 87030 187446
rect 87046 187502 87110 187506
rect 87046 187446 87050 187502
rect 87050 187446 87106 187502
rect 87106 187446 87110 187502
rect 87046 187442 87110 187446
rect 87126 187502 87190 187506
rect 87126 187446 87130 187502
rect 87130 187446 87186 187502
rect 87186 187446 87190 187502
rect 87126 187442 87190 187446
rect 4146 187374 4210 187438
rect 84186 187238 84250 187302
rect 3594 187102 3658 187166
rect 84554 187102 84618 187166
rect 3778 186966 3842 187030
rect 886 186958 950 186962
rect 886 186902 890 186958
rect 890 186902 946 186958
rect 946 186902 950 186958
rect 886 186898 950 186902
rect 966 186958 1030 186962
rect 966 186902 970 186958
rect 970 186902 1026 186958
rect 1026 186902 1030 186958
rect 966 186898 1030 186902
rect 1046 186958 1110 186962
rect 1046 186902 1050 186958
rect 1050 186902 1106 186958
rect 1106 186902 1110 186958
rect 1046 186898 1110 186902
rect 1126 186958 1190 186962
rect 1126 186902 1130 186958
rect 1130 186902 1186 186958
rect 1186 186902 1190 186958
rect 1126 186898 1190 186902
rect 84886 186958 84950 186962
rect 84886 186902 84890 186958
rect 84890 186902 84946 186958
rect 84946 186902 84950 186958
rect 84886 186898 84950 186902
rect 84966 186958 85030 186962
rect 84966 186902 84970 186958
rect 84970 186902 85026 186958
rect 85026 186902 85030 186958
rect 84966 186898 85030 186902
rect 85046 186958 85110 186962
rect 85046 186902 85050 186958
rect 85050 186902 85106 186958
rect 85106 186902 85110 186958
rect 85046 186898 85110 186902
rect 85126 186958 85190 186962
rect 85126 186902 85130 186958
rect 85130 186902 85186 186958
rect 85186 186902 85190 186958
rect 85126 186898 85190 186902
rect 84738 186558 84802 186622
rect 2886 186414 2950 186418
rect 2886 186358 2890 186414
rect 2890 186358 2946 186414
rect 2946 186358 2950 186414
rect 2886 186354 2950 186358
rect 2966 186414 3030 186418
rect 2966 186358 2970 186414
rect 2970 186358 3026 186414
rect 3026 186358 3030 186414
rect 2966 186354 3030 186358
rect 3046 186414 3110 186418
rect 3046 186358 3050 186414
rect 3050 186358 3106 186414
rect 3106 186358 3110 186414
rect 3046 186354 3110 186358
rect 3126 186414 3190 186418
rect 3126 186358 3130 186414
rect 3130 186358 3186 186414
rect 3186 186358 3190 186414
rect 3126 186354 3190 186358
rect 86886 186414 86950 186418
rect 86886 186358 86890 186414
rect 86890 186358 86946 186414
rect 86946 186358 86950 186414
rect 86886 186354 86950 186358
rect 86966 186414 87030 186418
rect 86966 186358 86970 186414
rect 86970 186358 87026 186414
rect 87026 186358 87030 186414
rect 86966 186354 87030 186358
rect 87046 186414 87110 186418
rect 87046 186358 87050 186414
rect 87050 186358 87106 186414
rect 87106 186358 87110 186414
rect 87046 186354 87110 186358
rect 87126 186414 87190 186418
rect 87126 186358 87130 186414
rect 87130 186358 87186 186414
rect 87186 186358 87190 186414
rect 87126 186354 87190 186358
rect 886 185870 950 185874
rect 886 185814 890 185870
rect 890 185814 946 185870
rect 946 185814 950 185870
rect 886 185810 950 185814
rect 966 185870 1030 185874
rect 966 185814 970 185870
rect 970 185814 1026 185870
rect 1026 185814 1030 185870
rect 966 185810 1030 185814
rect 1046 185870 1110 185874
rect 1046 185814 1050 185870
rect 1050 185814 1106 185870
rect 1106 185814 1110 185870
rect 1046 185810 1110 185814
rect 1126 185870 1190 185874
rect 1126 185814 1130 185870
rect 1130 185814 1186 185870
rect 1186 185814 1190 185870
rect 1126 185810 1190 185814
rect 84886 185870 84950 185874
rect 84886 185814 84890 185870
rect 84890 185814 84946 185870
rect 84946 185814 84950 185870
rect 84886 185810 84950 185814
rect 84966 185870 85030 185874
rect 84966 185814 84970 185870
rect 84970 185814 85026 185870
rect 85026 185814 85030 185870
rect 84966 185810 85030 185814
rect 85046 185870 85110 185874
rect 85046 185814 85050 185870
rect 85050 185814 85106 185870
rect 85106 185814 85110 185870
rect 85046 185810 85110 185814
rect 85126 185870 85190 185874
rect 85126 185814 85130 185870
rect 85130 185814 85186 185870
rect 85186 185814 85190 185870
rect 85126 185810 85190 185814
rect 2886 185326 2950 185330
rect 2886 185270 2890 185326
rect 2890 185270 2946 185326
rect 2946 185270 2950 185326
rect 2886 185266 2950 185270
rect 2966 185326 3030 185330
rect 2966 185270 2970 185326
rect 2970 185270 3026 185326
rect 3026 185270 3030 185326
rect 2966 185266 3030 185270
rect 3046 185326 3110 185330
rect 3046 185270 3050 185326
rect 3050 185270 3106 185326
rect 3106 185270 3110 185326
rect 3046 185266 3110 185270
rect 3126 185326 3190 185330
rect 3126 185270 3130 185326
rect 3130 185270 3186 185326
rect 3186 185270 3190 185326
rect 3126 185266 3190 185270
rect 86886 185326 86950 185330
rect 86886 185270 86890 185326
rect 86890 185270 86946 185326
rect 86946 185270 86950 185326
rect 86886 185266 86950 185270
rect 86966 185326 87030 185330
rect 86966 185270 86970 185326
rect 86970 185270 87026 185326
rect 87026 185270 87030 185326
rect 86966 185266 87030 185270
rect 87046 185326 87110 185330
rect 87046 185270 87050 185326
rect 87050 185270 87106 185326
rect 87106 185270 87110 185326
rect 87046 185266 87110 185270
rect 87126 185326 87190 185330
rect 87126 185270 87130 185326
rect 87130 185270 87186 185326
rect 87186 185270 87190 185326
rect 87126 185266 87190 185270
rect 886 184782 950 184786
rect 886 184726 890 184782
rect 890 184726 946 184782
rect 946 184726 950 184782
rect 886 184722 950 184726
rect 966 184782 1030 184786
rect 966 184726 970 184782
rect 970 184726 1026 184782
rect 1026 184726 1030 184782
rect 966 184722 1030 184726
rect 1046 184782 1110 184786
rect 1046 184726 1050 184782
rect 1050 184726 1106 184782
rect 1106 184726 1110 184782
rect 1046 184722 1110 184726
rect 1126 184782 1190 184786
rect 1126 184726 1130 184782
rect 1130 184726 1186 184782
rect 1186 184726 1190 184782
rect 1126 184722 1190 184726
rect 84886 184782 84950 184786
rect 84886 184726 84890 184782
rect 84890 184726 84946 184782
rect 84946 184726 84950 184782
rect 84886 184722 84950 184726
rect 84966 184782 85030 184786
rect 84966 184726 84970 184782
rect 84970 184726 85026 184782
rect 85026 184726 85030 184782
rect 84966 184722 85030 184726
rect 85046 184782 85110 184786
rect 85046 184726 85050 184782
rect 85050 184726 85106 184782
rect 85106 184726 85110 184782
rect 85046 184722 85110 184726
rect 85126 184782 85190 184786
rect 85126 184726 85130 184782
rect 85130 184726 85186 184782
rect 85186 184726 85190 184782
rect 85126 184722 85190 184726
rect 84738 184382 84802 184446
rect 2886 184238 2950 184242
rect 2886 184182 2890 184238
rect 2890 184182 2946 184238
rect 2946 184182 2950 184238
rect 2886 184178 2950 184182
rect 2966 184238 3030 184242
rect 2966 184182 2970 184238
rect 2970 184182 3026 184238
rect 3026 184182 3030 184238
rect 2966 184178 3030 184182
rect 3046 184238 3110 184242
rect 3046 184182 3050 184238
rect 3050 184182 3106 184238
rect 3106 184182 3110 184238
rect 3046 184178 3110 184182
rect 3126 184238 3190 184242
rect 3126 184182 3130 184238
rect 3130 184182 3186 184238
rect 3186 184182 3190 184238
rect 3126 184178 3190 184182
rect 86886 184238 86950 184242
rect 86886 184182 86890 184238
rect 86890 184182 86946 184238
rect 86946 184182 86950 184238
rect 86886 184178 86950 184182
rect 86966 184238 87030 184242
rect 86966 184182 86970 184238
rect 86970 184182 87026 184238
rect 87026 184182 87030 184238
rect 86966 184178 87030 184182
rect 87046 184238 87110 184242
rect 87046 184182 87050 184238
rect 87050 184182 87106 184238
rect 87106 184182 87110 184238
rect 87046 184178 87110 184182
rect 87126 184238 87190 184242
rect 87126 184182 87130 184238
rect 87130 184182 87186 184238
rect 87186 184182 87190 184238
rect 87126 184178 87190 184182
rect 886 183694 950 183698
rect 886 183638 890 183694
rect 890 183638 946 183694
rect 946 183638 950 183694
rect 886 183634 950 183638
rect 966 183694 1030 183698
rect 966 183638 970 183694
rect 970 183638 1026 183694
rect 1026 183638 1030 183694
rect 966 183634 1030 183638
rect 1046 183694 1110 183698
rect 1046 183638 1050 183694
rect 1050 183638 1106 183694
rect 1106 183638 1110 183694
rect 1046 183634 1110 183638
rect 1126 183694 1190 183698
rect 1126 183638 1130 183694
rect 1130 183638 1186 183694
rect 1186 183638 1190 183694
rect 1126 183634 1190 183638
rect 84886 183694 84950 183698
rect 84886 183638 84890 183694
rect 84890 183638 84946 183694
rect 84946 183638 84950 183694
rect 84886 183634 84950 183638
rect 84966 183694 85030 183698
rect 84966 183638 84970 183694
rect 84970 183638 85026 183694
rect 85026 183638 85030 183694
rect 84966 183634 85030 183638
rect 85046 183694 85110 183698
rect 85046 183638 85050 183694
rect 85050 183638 85106 183694
rect 85106 183638 85110 183694
rect 85046 183634 85110 183638
rect 85126 183694 85190 183698
rect 85126 183638 85130 183694
rect 85130 183638 85186 183694
rect 85186 183638 85190 183694
rect 85126 183634 85190 183638
rect 84554 183294 84618 183358
rect 2886 183150 2950 183154
rect 2886 183094 2890 183150
rect 2890 183094 2946 183150
rect 2946 183094 2950 183150
rect 2886 183090 2950 183094
rect 2966 183150 3030 183154
rect 2966 183094 2970 183150
rect 2970 183094 3026 183150
rect 3026 183094 3030 183150
rect 2966 183090 3030 183094
rect 3046 183150 3110 183154
rect 3046 183094 3050 183150
rect 3050 183094 3106 183150
rect 3106 183094 3110 183150
rect 3046 183090 3110 183094
rect 3126 183150 3190 183154
rect 3126 183094 3130 183150
rect 3130 183094 3186 183150
rect 3186 183094 3190 183150
rect 3126 183090 3190 183094
rect 86886 183150 86950 183154
rect 86886 183094 86890 183150
rect 86890 183094 86946 183150
rect 86946 183094 86950 183150
rect 86886 183090 86950 183094
rect 86966 183150 87030 183154
rect 86966 183094 86970 183150
rect 86970 183094 87026 183150
rect 87026 183094 87030 183150
rect 86966 183090 87030 183094
rect 87046 183150 87110 183154
rect 87046 183094 87050 183150
rect 87050 183094 87106 183150
rect 87106 183094 87110 183150
rect 87046 183090 87110 183094
rect 87126 183150 87190 183154
rect 87126 183094 87130 183150
rect 87130 183094 87186 183150
rect 87186 183094 87190 183150
rect 87126 183090 87190 183094
rect 886 182606 950 182610
rect 886 182550 890 182606
rect 890 182550 946 182606
rect 946 182550 950 182606
rect 886 182546 950 182550
rect 966 182606 1030 182610
rect 966 182550 970 182606
rect 970 182550 1026 182606
rect 1026 182550 1030 182606
rect 966 182546 1030 182550
rect 1046 182606 1110 182610
rect 1046 182550 1050 182606
rect 1050 182550 1106 182606
rect 1106 182550 1110 182606
rect 1046 182546 1110 182550
rect 1126 182606 1190 182610
rect 1126 182550 1130 182606
rect 1130 182550 1186 182606
rect 1186 182550 1190 182606
rect 1126 182546 1190 182550
rect 84886 182606 84950 182610
rect 84886 182550 84890 182606
rect 84890 182550 84946 182606
rect 84946 182550 84950 182606
rect 84886 182546 84950 182550
rect 84966 182606 85030 182610
rect 84966 182550 84970 182606
rect 84970 182550 85026 182606
rect 85026 182550 85030 182606
rect 84966 182546 85030 182550
rect 85046 182606 85110 182610
rect 85046 182550 85050 182606
rect 85050 182550 85106 182606
rect 85106 182550 85110 182606
rect 85046 182546 85110 182550
rect 85126 182606 85190 182610
rect 85126 182550 85130 182606
rect 85130 182550 85186 182606
rect 85186 182550 85190 182606
rect 85126 182546 85190 182550
rect 84554 182206 84618 182270
rect 2886 182062 2950 182066
rect 2886 182006 2890 182062
rect 2890 182006 2946 182062
rect 2946 182006 2950 182062
rect 2886 182002 2950 182006
rect 2966 182062 3030 182066
rect 2966 182006 2970 182062
rect 2970 182006 3026 182062
rect 3026 182006 3030 182062
rect 2966 182002 3030 182006
rect 3046 182062 3110 182066
rect 3046 182006 3050 182062
rect 3050 182006 3106 182062
rect 3106 182006 3110 182062
rect 3046 182002 3110 182006
rect 3126 182062 3190 182066
rect 3126 182006 3130 182062
rect 3130 182006 3186 182062
rect 3186 182006 3190 182062
rect 3126 182002 3190 182006
rect 86886 182062 86950 182066
rect 86886 182006 86890 182062
rect 86890 182006 86946 182062
rect 86946 182006 86950 182062
rect 86886 182002 86950 182006
rect 86966 182062 87030 182066
rect 86966 182006 86970 182062
rect 86970 182006 87026 182062
rect 87026 182006 87030 182062
rect 86966 182002 87030 182006
rect 87046 182062 87110 182066
rect 87046 182006 87050 182062
rect 87050 182006 87106 182062
rect 87106 182006 87110 182062
rect 87046 182002 87110 182006
rect 87126 182062 87190 182066
rect 87126 182006 87130 182062
rect 87130 182006 87186 182062
rect 87186 182006 87190 182062
rect 87126 182002 87190 182006
rect 886 181518 950 181522
rect 886 181462 890 181518
rect 890 181462 946 181518
rect 946 181462 950 181518
rect 886 181458 950 181462
rect 966 181518 1030 181522
rect 966 181462 970 181518
rect 970 181462 1026 181518
rect 1026 181462 1030 181518
rect 966 181458 1030 181462
rect 1046 181518 1110 181522
rect 1046 181462 1050 181518
rect 1050 181462 1106 181518
rect 1106 181462 1110 181518
rect 1046 181458 1110 181462
rect 1126 181518 1190 181522
rect 1126 181462 1130 181518
rect 1130 181462 1186 181518
rect 1186 181462 1190 181518
rect 1126 181458 1190 181462
rect 84886 181518 84950 181522
rect 84886 181462 84890 181518
rect 84890 181462 84946 181518
rect 84946 181462 84950 181518
rect 84886 181458 84950 181462
rect 84966 181518 85030 181522
rect 84966 181462 84970 181518
rect 84970 181462 85026 181518
rect 85026 181462 85030 181518
rect 84966 181458 85030 181462
rect 85046 181518 85110 181522
rect 85046 181462 85050 181518
rect 85050 181462 85106 181518
rect 85106 181462 85110 181518
rect 85046 181458 85110 181462
rect 85126 181518 85190 181522
rect 85126 181462 85130 181518
rect 85130 181462 85186 181518
rect 85186 181462 85190 181518
rect 85126 181458 85190 181462
rect 2886 180974 2950 180978
rect 2886 180918 2890 180974
rect 2890 180918 2946 180974
rect 2946 180918 2950 180974
rect 2886 180914 2950 180918
rect 2966 180974 3030 180978
rect 2966 180918 2970 180974
rect 2970 180918 3026 180974
rect 3026 180918 3030 180974
rect 2966 180914 3030 180918
rect 3046 180974 3110 180978
rect 3046 180918 3050 180974
rect 3050 180918 3106 180974
rect 3106 180918 3110 180974
rect 3046 180914 3110 180918
rect 3126 180974 3190 180978
rect 3126 180918 3130 180974
rect 3130 180918 3186 180974
rect 3186 180918 3190 180974
rect 3126 180914 3190 180918
rect 86886 180974 86950 180978
rect 86886 180918 86890 180974
rect 86890 180918 86946 180974
rect 86946 180918 86950 180974
rect 86886 180914 86950 180918
rect 86966 180974 87030 180978
rect 86966 180918 86970 180974
rect 86970 180918 87026 180974
rect 87026 180918 87030 180974
rect 86966 180914 87030 180918
rect 87046 180974 87110 180978
rect 87046 180918 87050 180974
rect 87050 180918 87106 180974
rect 87106 180918 87110 180974
rect 87046 180914 87110 180918
rect 87126 180974 87190 180978
rect 87126 180918 87130 180974
rect 87130 180918 87186 180974
rect 87186 180918 87190 180974
rect 87126 180914 87190 180918
rect 886 180430 950 180434
rect 886 180374 890 180430
rect 890 180374 946 180430
rect 946 180374 950 180430
rect 886 180370 950 180374
rect 966 180430 1030 180434
rect 966 180374 970 180430
rect 970 180374 1026 180430
rect 1026 180374 1030 180430
rect 966 180370 1030 180374
rect 1046 180430 1110 180434
rect 1046 180374 1050 180430
rect 1050 180374 1106 180430
rect 1106 180374 1110 180430
rect 1046 180370 1110 180374
rect 1126 180430 1190 180434
rect 1126 180374 1130 180430
rect 1130 180374 1186 180430
rect 1186 180374 1190 180430
rect 1126 180370 1190 180374
rect 84886 180430 84950 180434
rect 84886 180374 84890 180430
rect 84890 180374 84946 180430
rect 84946 180374 84950 180430
rect 84886 180370 84950 180374
rect 84966 180430 85030 180434
rect 84966 180374 84970 180430
rect 84970 180374 85026 180430
rect 85026 180374 85030 180430
rect 84966 180370 85030 180374
rect 85046 180430 85110 180434
rect 85046 180374 85050 180430
rect 85050 180374 85106 180430
rect 85106 180374 85110 180430
rect 85046 180370 85110 180374
rect 85126 180430 85190 180434
rect 85126 180374 85130 180430
rect 85130 180374 85186 180430
rect 85186 180374 85190 180430
rect 85126 180370 85190 180374
rect 2886 179886 2950 179890
rect 2886 179830 2890 179886
rect 2890 179830 2946 179886
rect 2946 179830 2950 179886
rect 2886 179826 2950 179830
rect 2966 179886 3030 179890
rect 2966 179830 2970 179886
rect 2970 179830 3026 179886
rect 3026 179830 3030 179886
rect 2966 179826 3030 179830
rect 3046 179886 3110 179890
rect 3046 179830 3050 179886
rect 3050 179830 3106 179886
rect 3106 179830 3110 179886
rect 3046 179826 3110 179830
rect 3126 179886 3190 179890
rect 3126 179830 3130 179886
rect 3130 179830 3186 179886
rect 3186 179830 3190 179886
rect 3126 179826 3190 179830
rect 86886 179886 86950 179890
rect 86886 179830 86890 179886
rect 86890 179830 86946 179886
rect 86946 179830 86950 179886
rect 86886 179826 86950 179830
rect 86966 179886 87030 179890
rect 86966 179830 86970 179886
rect 86970 179830 87026 179886
rect 87026 179830 87030 179886
rect 86966 179826 87030 179830
rect 87046 179886 87110 179890
rect 87046 179830 87050 179886
rect 87050 179830 87106 179886
rect 87106 179830 87110 179886
rect 87046 179826 87110 179830
rect 87126 179886 87190 179890
rect 87126 179830 87130 179886
rect 87130 179830 87186 179886
rect 87186 179830 87190 179886
rect 87126 179826 87190 179830
rect 886 179342 950 179346
rect 886 179286 890 179342
rect 890 179286 946 179342
rect 946 179286 950 179342
rect 886 179282 950 179286
rect 966 179342 1030 179346
rect 966 179286 970 179342
rect 970 179286 1026 179342
rect 1026 179286 1030 179342
rect 966 179282 1030 179286
rect 1046 179342 1110 179346
rect 1046 179286 1050 179342
rect 1050 179286 1106 179342
rect 1106 179286 1110 179342
rect 1046 179282 1110 179286
rect 1126 179342 1190 179346
rect 1126 179286 1130 179342
rect 1130 179286 1186 179342
rect 1186 179286 1190 179342
rect 1126 179282 1190 179286
rect 84886 179342 84950 179346
rect 84886 179286 84890 179342
rect 84890 179286 84946 179342
rect 84946 179286 84950 179342
rect 84886 179282 84950 179286
rect 84966 179342 85030 179346
rect 84966 179286 84970 179342
rect 84970 179286 85026 179342
rect 85026 179286 85030 179342
rect 84966 179282 85030 179286
rect 85046 179342 85110 179346
rect 85046 179286 85050 179342
rect 85050 179286 85106 179342
rect 85106 179286 85110 179342
rect 85046 179282 85110 179286
rect 85126 179342 85190 179346
rect 85126 179286 85130 179342
rect 85130 179286 85186 179342
rect 85186 179286 85190 179342
rect 85126 179282 85190 179286
rect 2886 178798 2950 178802
rect 2886 178742 2890 178798
rect 2890 178742 2946 178798
rect 2946 178742 2950 178798
rect 2886 178738 2950 178742
rect 2966 178798 3030 178802
rect 2966 178742 2970 178798
rect 2970 178742 3026 178798
rect 3026 178742 3030 178798
rect 2966 178738 3030 178742
rect 3046 178798 3110 178802
rect 3046 178742 3050 178798
rect 3050 178742 3106 178798
rect 3106 178742 3110 178798
rect 3046 178738 3110 178742
rect 3126 178798 3190 178802
rect 3126 178742 3130 178798
rect 3130 178742 3186 178798
rect 3186 178742 3190 178798
rect 3126 178738 3190 178742
rect 86886 178798 86950 178802
rect 86886 178742 86890 178798
rect 86890 178742 86946 178798
rect 86946 178742 86950 178798
rect 86886 178738 86950 178742
rect 86966 178798 87030 178802
rect 86966 178742 86970 178798
rect 86970 178742 87026 178798
rect 87026 178742 87030 178798
rect 86966 178738 87030 178742
rect 87046 178798 87110 178802
rect 87046 178742 87050 178798
rect 87050 178742 87106 178798
rect 87106 178742 87110 178798
rect 87046 178738 87110 178742
rect 87126 178798 87190 178802
rect 87126 178742 87130 178798
rect 87130 178742 87186 178798
rect 87186 178742 87190 178798
rect 87126 178738 87190 178742
rect 886 178254 950 178258
rect 886 178198 890 178254
rect 890 178198 946 178254
rect 946 178198 950 178254
rect 886 178194 950 178198
rect 966 178254 1030 178258
rect 966 178198 970 178254
rect 970 178198 1026 178254
rect 1026 178198 1030 178254
rect 966 178194 1030 178198
rect 1046 178254 1110 178258
rect 1046 178198 1050 178254
rect 1050 178198 1106 178254
rect 1106 178198 1110 178254
rect 1046 178194 1110 178198
rect 1126 178254 1190 178258
rect 1126 178198 1130 178254
rect 1130 178198 1186 178254
rect 1186 178198 1190 178254
rect 1126 178194 1190 178198
rect 84886 178254 84950 178258
rect 84886 178198 84890 178254
rect 84890 178198 84946 178254
rect 84946 178198 84950 178254
rect 84886 178194 84950 178198
rect 84966 178254 85030 178258
rect 84966 178198 84970 178254
rect 84970 178198 85026 178254
rect 85026 178198 85030 178254
rect 84966 178194 85030 178198
rect 85046 178254 85110 178258
rect 85046 178198 85050 178254
rect 85050 178198 85106 178254
rect 85106 178198 85110 178254
rect 85046 178194 85110 178198
rect 85126 178254 85190 178258
rect 85126 178198 85130 178254
rect 85130 178198 85186 178254
rect 85186 178198 85190 178254
rect 85126 178194 85190 178198
rect 2886 177710 2950 177714
rect 2886 177654 2890 177710
rect 2890 177654 2946 177710
rect 2946 177654 2950 177710
rect 2886 177650 2950 177654
rect 2966 177710 3030 177714
rect 2966 177654 2970 177710
rect 2970 177654 3026 177710
rect 3026 177654 3030 177710
rect 2966 177650 3030 177654
rect 3046 177710 3110 177714
rect 3046 177654 3050 177710
rect 3050 177654 3106 177710
rect 3106 177654 3110 177710
rect 3046 177650 3110 177654
rect 3126 177710 3190 177714
rect 3126 177654 3130 177710
rect 3130 177654 3186 177710
rect 3186 177654 3190 177710
rect 3126 177650 3190 177654
rect 86886 177710 86950 177714
rect 86886 177654 86890 177710
rect 86890 177654 86946 177710
rect 86946 177654 86950 177710
rect 86886 177650 86950 177654
rect 86966 177710 87030 177714
rect 86966 177654 86970 177710
rect 86970 177654 87026 177710
rect 87026 177654 87030 177710
rect 86966 177650 87030 177654
rect 87046 177710 87110 177714
rect 87046 177654 87050 177710
rect 87050 177654 87106 177710
rect 87106 177654 87110 177710
rect 87046 177650 87110 177654
rect 87126 177710 87190 177714
rect 87126 177654 87130 177710
rect 87130 177654 87186 177710
rect 87186 177654 87190 177710
rect 87126 177650 87190 177654
rect 886 177166 950 177170
rect 886 177110 890 177166
rect 890 177110 946 177166
rect 946 177110 950 177166
rect 886 177106 950 177110
rect 966 177166 1030 177170
rect 966 177110 970 177166
rect 970 177110 1026 177166
rect 1026 177110 1030 177166
rect 966 177106 1030 177110
rect 1046 177166 1110 177170
rect 1046 177110 1050 177166
rect 1050 177110 1106 177166
rect 1106 177110 1110 177166
rect 1046 177106 1110 177110
rect 1126 177166 1190 177170
rect 1126 177110 1130 177166
rect 1130 177110 1186 177166
rect 1186 177110 1190 177166
rect 1126 177106 1190 177110
rect 84886 177166 84950 177170
rect 84886 177110 84890 177166
rect 84890 177110 84946 177166
rect 84946 177110 84950 177166
rect 84886 177106 84950 177110
rect 84966 177166 85030 177170
rect 84966 177110 84970 177166
rect 84970 177110 85026 177166
rect 85026 177110 85030 177166
rect 84966 177106 85030 177110
rect 85046 177166 85110 177170
rect 85046 177110 85050 177166
rect 85050 177110 85106 177166
rect 85106 177110 85110 177166
rect 85046 177106 85110 177110
rect 85126 177166 85190 177170
rect 85126 177110 85130 177166
rect 85130 177110 85186 177166
rect 85186 177110 85190 177166
rect 85126 177106 85190 177110
rect 2886 176622 2950 176626
rect 2886 176566 2890 176622
rect 2890 176566 2946 176622
rect 2946 176566 2950 176622
rect 2886 176562 2950 176566
rect 2966 176622 3030 176626
rect 2966 176566 2970 176622
rect 2970 176566 3026 176622
rect 3026 176566 3030 176622
rect 2966 176562 3030 176566
rect 3046 176622 3110 176626
rect 3046 176566 3050 176622
rect 3050 176566 3106 176622
rect 3106 176566 3110 176622
rect 3046 176562 3110 176566
rect 3126 176622 3190 176626
rect 3126 176566 3130 176622
rect 3130 176566 3186 176622
rect 3186 176566 3190 176622
rect 3126 176562 3190 176566
rect 86886 176622 86950 176626
rect 86886 176566 86890 176622
rect 86890 176566 86946 176622
rect 86946 176566 86950 176622
rect 86886 176562 86950 176566
rect 86966 176622 87030 176626
rect 86966 176566 86970 176622
rect 86970 176566 87026 176622
rect 87026 176566 87030 176622
rect 86966 176562 87030 176566
rect 87046 176622 87110 176626
rect 87046 176566 87050 176622
rect 87050 176566 87106 176622
rect 87106 176566 87110 176622
rect 87046 176562 87110 176566
rect 87126 176622 87190 176626
rect 87126 176566 87130 176622
rect 87130 176566 87186 176622
rect 87186 176566 87190 176622
rect 87126 176562 87190 176566
rect 886 176078 950 176082
rect 886 176022 890 176078
rect 890 176022 946 176078
rect 946 176022 950 176078
rect 886 176018 950 176022
rect 966 176078 1030 176082
rect 966 176022 970 176078
rect 970 176022 1026 176078
rect 1026 176022 1030 176078
rect 966 176018 1030 176022
rect 1046 176078 1110 176082
rect 1046 176022 1050 176078
rect 1050 176022 1106 176078
rect 1106 176022 1110 176078
rect 1046 176018 1110 176022
rect 1126 176078 1190 176082
rect 1126 176022 1130 176078
rect 1130 176022 1186 176078
rect 1186 176022 1190 176078
rect 1126 176018 1190 176022
rect 84886 176078 84950 176082
rect 84886 176022 84890 176078
rect 84890 176022 84946 176078
rect 84946 176022 84950 176078
rect 84886 176018 84950 176022
rect 84966 176078 85030 176082
rect 84966 176022 84970 176078
rect 84970 176022 85026 176078
rect 85026 176022 85030 176078
rect 84966 176018 85030 176022
rect 85046 176078 85110 176082
rect 85046 176022 85050 176078
rect 85050 176022 85106 176078
rect 85106 176022 85110 176078
rect 85046 176018 85110 176022
rect 85126 176078 85190 176082
rect 85126 176022 85130 176078
rect 85130 176022 85186 176078
rect 85186 176022 85190 176078
rect 85126 176018 85190 176022
rect 2886 175534 2950 175538
rect 2886 175478 2890 175534
rect 2890 175478 2946 175534
rect 2946 175478 2950 175534
rect 2886 175474 2950 175478
rect 2966 175534 3030 175538
rect 2966 175478 2970 175534
rect 2970 175478 3026 175534
rect 3026 175478 3030 175534
rect 2966 175474 3030 175478
rect 3046 175534 3110 175538
rect 3046 175478 3050 175534
rect 3050 175478 3106 175534
rect 3106 175478 3110 175534
rect 3046 175474 3110 175478
rect 3126 175534 3190 175538
rect 3126 175478 3130 175534
rect 3130 175478 3186 175534
rect 3186 175478 3190 175534
rect 3126 175474 3190 175478
rect 86886 175534 86950 175538
rect 86886 175478 86890 175534
rect 86890 175478 86946 175534
rect 86946 175478 86950 175534
rect 86886 175474 86950 175478
rect 86966 175534 87030 175538
rect 86966 175478 86970 175534
rect 86970 175478 87026 175534
rect 87026 175478 87030 175534
rect 86966 175474 87030 175478
rect 87046 175534 87110 175538
rect 87046 175478 87050 175534
rect 87050 175478 87106 175534
rect 87106 175478 87110 175534
rect 87046 175474 87110 175478
rect 87126 175534 87190 175538
rect 87126 175478 87130 175534
rect 87130 175478 87186 175534
rect 87186 175478 87190 175534
rect 87126 175474 87190 175478
rect 886 174990 950 174994
rect 886 174934 890 174990
rect 890 174934 946 174990
rect 946 174934 950 174990
rect 886 174930 950 174934
rect 966 174990 1030 174994
rect 966 174934 970 174990
rect 970 174934 1026 174990
rect 1026 174934 1030 174990
rect 966 174930 1030 174934
rect 1046 174990 1110 174994
rect 1046 174934 1050 174990
rect 1050 174934 1106 174990
rect 1106 174934 1110 174990
rect 1046 174930 1110 174934
rect 1126 174990 1190 174994
rect 1126 174934 1130 174990
rect 1130 174934 1186 174990
rect 1186 174934 1190 174990
rect 1126 174930 1190 174934
rect 84886 174990 84950 174994
rect 84886 174934 84890 174990
rect 84890 174934 84946 174990
rect 84946 174934 84950 174990
rect 84886 174930 84950 174934
rect 84966 174990 85030 174994
rect 84966 174934 84970 174990
rect 84970 174934 85026 174990
rect 85026 174934 85030 174990
rect 84966 174930 85030 174934
rect 85046 174990 85110 174994
rect 85046 174934 85050 174990
rect 85050 174934 85106 174990
rect 85106 174934 85110 174990
rect 85046 174930 85110 174934
rect 85126 174990 85190 174994
rect 85126 174934 85130 174990
rect 85130 174934 85186 174990
rect 85186 174934 85190 174990
rect 85126 174930 85190 174934
rect 2886 174446 2950 174450
rect 2886 174390 2890 174446
rect 2890 174390 2946 174446
rect 2946 174390 2950 174446
rect 2886 174386 2950 174390
rect 2966 174446 3030 174450
rect 2966 174390 2970 174446
rect 2970 174390 3026 174446
rect 3026 174390 3030 174446
rect 2966 174386 3030 174390
rect 3046 174446 3110 174450
rect 3046 174390 3050 174446
rect 3050 174390 3106 174446
rect 3106 174390 3110 174446
rect 3046 174386 3110 174390
rect 3126 174446 3190 174450
rect 3126 174390 3130 174446
rect 3130 174390 3186 174446
rect 3186 174390 3190 174446
rect 3126 174386 3190 174390
rect 86886 174446 86950 174450
rect 86886 174390 86890 174446
rect 86890 174390 86946 174446
rect 86946 174390 86950 174446
rect 86886 174386 86950 174390
rect 86966 174446 87030 174450
rect 86966 174390 86970 174446
rect 86970 174390 87026 174446
rect 87026 174390 87030 174446
rect 86966 174386 87030 174390
rect 87046 174446 87110 174450
rect 87046 174390 87050 174446
rect 87050 174390 87106 174446
rect 87106 174390 87110 174446
rect 87046 174386 87110 174390
rect 87126 174446 87190 174450
rect 87126 174390 87130 174446
rect 87130 174390 87186 174446
rect 87186 174390 87190 174446
rect 87126 174386 87190 174390
rect 886 173902 950 173906
rect 886 173846 890 173902
rect 890 173846 946 173902
rect 946 173846 950 173902
rect 886 173842 950 173846
rect 966 173902 1030 173906
rect 966 173846 970 173902
rect 970 173846 1026 173902
rect 1026 173846 1030 173902
rect 966 173842 1030 173846
rect 1046 173902 1110 173906
rect 1046 173846 1050 173902
rect 1050 173846 1106 173902
rect 1106 173846 1110 173902
rect 1046 173842 1110 173846
rect 1126 173902 1190 173906
rect 1126 173846 1130 173902
rect 1130 173846 1186 173902
rect 1186 173846 1190 173902
rect 1126 173842 1190 173846
rect 84886 173902 84950 173906
rect 84886 173846 84890 173902
rect 84890 173846 84946 173902
rect 84946 173846 84950 173902
rect 84886 173842 84950 173846
rect 84966 173902 85030 173906
rect 84966 173846 84970 173902
rect 84970 173846 85026 173902
rect 85026 173846 85030 173902
rect 84966 173842 85030 173846
rect 85046 173902 85110 173906
rect 85046 173846 85050 173902
rect 85050 173846 85106 173902
rect 85106 173846 85110 173902
rect 85046 173842 85110 173846
rect 85126 173902 85190 173906
rect 85126 173846 85130 173902
rect 85130 173846 85186 173902
rect 85186 173846 85190 173902
rect 85126 173842 85190 173846
rect 2886 173358 2950 173362
rect 2886 173302 2890 173358
rect 2890 173302 2946 173358
rect 2946 173302 2950 173358
rect 2886 173298 2950 173302
rect 2966 173358 3030 173362
rect 2966 173302 2970 173358
rect 2970 173302 3026 173358
rect 3026 173302 3030 173358
rect 2966 173298 3030 173302
rect 3046 173358 3110 173362
rect 3046 173302 3050 173358
rect 3050 173302 3106 173358
rect 3106 173302 3110 173358
rect 3046 173298 3110 173302
rect 3126 173358 3190 173362
rect 3126 173302 3130 173358
rect 3130 173302 3186 173358
rect 3186 173302 3190 173358
rect 3126 173298 3190 173302
rect 86886 173358 86950 173362
rect 86886 173302 86890 173358
rect 86890 173302 86946 173358
rect 86946 173302 86950 173358
rect 86886 173298 86950 173302
rect 86966 173358 87030 173362
rect 86966 173302 86970 173358
rect 86970 173302 87026 173358
rect 87026 173302 87030 173358
rect 86966 173298 87030 173302
rect 87046 173358 87110 173362
rect 87046 173302 87050 173358
rect 87050 173302 87106 173358
rect 87106 173302 87110 173358
rect 87046 173298 87110 173302
rect 87126 173358 87190 173362
rect 87126 173302 87130 173358
rect 87130 173302 87186 173358
rect 87186 173302 87190 173358
rect 87126 173298 87190 173302
rect 886 172814 950 172818
rect 886 172758 890 172814
rect 890 172758 946 172814
rect 946 172758 950 172814
rect 886 172754 950 172758
rect 966 172814 1030 172818
rect 966 172758 970 172814
rect 970 172758 1026 172814
rect 1026 172758 1030 172814
rect 966 172754 1030 172758
rect 1046 172814 1110 172818
rect 1046 172758 1050 172814
rect 1050 172758 1106 172814
rect 1106 172758 1110 172814
rect 1046 172754 1110 172758
rect 1126 172814 1190 172818
rect 1126 172758 1130 172814
rect 1130 172758 1186 172814
rect 1186 172758 1190 172814
rect 1126 172754 1190 172758
rect 84886 172814 84950 172818
rect 84886 172758 84890 172814
rect 84890 172758 84946 172814
rect 84946 172758 84950 172814
rect 84886 172754 84950 172758
rect 84966 172814 85030 172818
rect 84966 172758 84970 172814
rect 84970 172758 85026 172814
rect 85026 172758 85030 172814
rect 84966 172754 85030 172758
rect 85046 172814 85110 172818
rect 85046 172758 85050 172814
rect 85050 172758 85106 172814
rect 85106 172758 85110 172814
rect 85046 172754 85110 172758
rect 85126 172814 85190 172818
rect 85126 172758 85130 172814
rect 85130 172758 85186 172814
rect 85186 172758 85190 172814
rect 85126 172754 85190 172758
rect 2886 172270 2950 172274
rect 2886 172214 2890 172270
rect 2890 172214 2946 172270
rect 2946 172214 2950 172270
rect 2886 172210 2950 172214
rect 2966 172270 3030 172274
rect 2966 172214 2970 172270
rect 2970 172214 3026 172270
rect 3026 172214 3030 172270
rect 2966 172210 3030 172214
rect 3046 172270 3110 172274
rect 3046 172214 3050 172270
rect 3050 172214 3106 172270
rect 3106 172214 3110 172270
rect 3046 172210 3110 172214
rect 3126 172270 3190 172274
rect 3126 172214 3130 172270
rect 3130 172214 3186 172270
rect 3186 172214 3190 172270
rect 3126 172210 3190 172214
rect 86886 172270 86950 172274
rect 86886 172214 86890 172270
rect 86890 172214 86946 172270
rect 86946 172214 86950 172270
rect 86886 172210 86950 172214
rect 86966 172270 87030 172274
rect 86966 172214 86970 172270
rect 86970 172214 87026 172270
rect 87026 172214 87030 172270
rect 86966 172210 87030 172214
rect 87046 172270 87110 172274
rect 87046 172214 87050 172270
rect 87050 172214 87106 172270
rect 87106 172214 87110 172270
rect 87046 172210 87110 172214
rect 87126 172270 87190 172274
rect 87126 172214 87130 172270
rect 87130 172214 87186 172270
rect 87186 172214 87190 172270
rect 87126 172210 87190 172214
rect 84738 172006 84802 172070
rect 886 171726 950 171730
rect 886 171670 890 171726
rect 890 171670 946 171726
rect 946 171670 950 171726
rect 886 171666 950 171670
rect 966 171726 1030 171730
rect 966 171670 970 171726
rect 970 171670 1026 171726
rect 1026 171670 1030 171726
rect 966 171666 1030 171670
rect 1046 171726 1110 171730
rect 1046 171670 1050 171726
rect 1050 171670 1106 171726
rect 1106 171670 1110 171726
rect 1046 171666 1110 171670
rect 1126 171726 1190 171730
rect 1126 171670 1130 171726
rect 1130 171670 1186 171726
rect 1186 171670 1190 171726
rect 1126 171666 1190 171670
rect 84886 171726 84950 171730
rect 84886 171670 84890 171726
rect 84890 171670 84946 171726
rect 84946 171670 84950 171726
rect 84886 171666 84950 171670
rect 84966 171726 85030 171730
rect 84966 171670 84970 171726
rect 84970 171670 85026 171726
rect 85026 171670 85030 171726
rect 84966 171666 85030 171670
rect 85046 171726 85110 171730
rect 85046 171670 85050 171726
rect 85050 171670 85106 171726
rect 85106 171670 85110 171726
rect 85046 171666 85110 171670
rect 85126 171726 85190 171730
rect 85126 171670 85130 171726
rect 85130 171670 85186 171726
rect 85186 171670 85190 171726
rect 85126 171666 85190 171670
rect 2886 171182 2950 171186
rect 2886 171126 2890 171182
rect 2890 171126 2946 171182
rect 2946 171126 2950 171182
rect 2886 171122 2950 171126
rect 2966 171182 3030 171186
rect 2966 171126 2970 171182
rect 2970 171126 3026 171182
rect 3026 171126 3030 171182
rect 2966 171122 3030 171126
rect 3046 171182 3110 171186
rect 3046 171126 3050 171182
rect 3050 171126 3106 171182
rect 3106 171126 3110 171182
rect 3046 171122 3110 171126
rect 3126 171182 3190 171186
rect 3126 171126 3130 171182
rect 3130 171126 3186 171182
rect 3186 171126 3190 171182
rect 3126 171122 3190 171126
rect 86886 171182 86950 171186
rect 86886 171126 86890 171182
rect 86890 171126 86946 171182
rect 86946 171126 86950 171182
rect 86886 171122 86950 171126
rect 86966 171182 87030 171186
rect 86966 171126 86970 171182
rect 86970 171126 87026 171182
rect 87026 171126 87030 171182
rect 86966 171122 87030 171126
rect 87046 171182 87110 171186
rect 87046 171126 87050 171182
rect 87050 171126 87106 171182
rect 87106 171126 87110 171182
rect 87046 171122 87110 171126
rect 87126 171182 87190 171186
rect 87126 171126 87130 171182
rect 87130 171126 87186 171182
rect 87186 171126 87190 171182
rect 87126 171122 87190 171126
rect 886 170638 950 170642
rect 886 170582 890 170638
rect 890 170582 946 170638
rect 946 170582 950 170638
rect 886 170578 950 170582
rect 966 170638 1030 170642
rect 966 170582 970 170638
rect 970 170582 1026 170638
rect 1026 170582 1030 170638
rect 966 170578 1030 170582
rect 1046 170638 1110 170642
rect 1046 170582 1050 170638
rect 1050 170582 1106 170638
rect 1106 170582 1110 170638
rect 1046 170578 1110 170582
rect 1126 170638 1190 170642
rect 1126 170582 1130 170638
rect 1130 170582 1186 170638
rect 1186 170582 1190 170638
rect 1126 170578 1190 170582
rect 84886 170638 84950 170642
rect 84886 170582 84890 170638
rect 84890 170582 84946 170638
rect 84946 170582 84950 170638
rect 84886 170578 84950 170582
rect 84966 170638 85030 170642
rect 84966 170582 84970 170638
rect 84970 170582 85026 170638
rect 85026 170582 85030 170638
rect 84966 170578 85030 170582
rect 85046 170638 85110 170642
rect 85046 170582 85050 170638
rect 85050 170582 85106 170638
rect 85106 170582 85110 170638
rect 85046 170578 85110 170582
rect 85126 170638 85190 170642
rect 85126 170582 85130 170638
rect 85130 170582 85186 170638
rect 85186 170582 85190 170638
rect 85126 170578 85190 170582
rect 2886 170094 2950 170098
rect 2886 170038 2890 170094
rect 2890 170038 2946 170094
rect 2946 170038 2950 170094
rect 2886 170034 2950 170038
rect 2966 170094 3030 170098
rect 2966 170038 2970 170094
rect 2970 170038 3026 170094
rect 3026 170038 3030 170094
rect 2966 170034 3030 170038
rect 3046 170094 3110 170098
rect 3046 170038 3050 170094
rect 3050 170038 3106 170094
rect 3106 170038 3110 170094
rect 3046 170034 3110 170038
rect 3126 170094 3190 170098
rect 3126 170038 3130 170094
rect 3130 170038 3186 170094
rect 3186 170038 3190 170094
rect 3126 170034 3190 170038
rect 86886 170094 86950 170098
rect 86886 170038 86890 170094
rect 86890 170038 86946 170094
rect 86946 170038 86950 170094
rect 86886 170034 86950 170038
rect 86966 170094 87030 170098
rect 86966 170038 86970 170094
rect 86970 170038 87026 170094
rect 87026 170038 87030 170094
rect 86966 170034 87030 170038
rect 87046 170094 87110 170098
rect 87046 170038 87050 170094
rect 87050 170038 87106 170094
rect 87106 170038 87110 170094
rect 87046 170034 87110 170038
rect 87126 170094 87190 170098
rect 87126 170038 87130 170094
rect 87130 170038 87186 170094
rect 87186 170038 87190 170094
rect 87126 170034 87190 170038
rect 83818 169830 83882 169894
rect 886 169550 950 169554
rect 886 169494 890 169550
rect 890 169494 946 169550
rect 946 169494 950 169550
rect 886 169490 950 169494
rect 966 169550 1030 169554
rect 966 169494 970 169550
rect 970 169494 1026 169550
rect 1026 169494 1030 169550
rect 966 169490 1030 169494
rect 1046 169550 1110 169554
rect 1046 169494 1050 169550
rect 1050 169494 1106 169550
rect 1106 169494 1110 169550
rect 1046 169490 1110 169494
rect 1126 169550 1190 169554
rect 1126 169494 1130 169550
rect 1130 169494 1186 169550
rect 1186 169494 1190 169550
rect 1126 169490 1190 169494
rect 84886 169550 84950 169554
rect 84886 169494 84890 169550
rect 84890 169494 84946 169550
rect 84946 169494 84950 169550
rect 84886 169490 84950 169494
rect 84966 169550 85030 169554
rect 84966 169494 84970 169550
rect 84970 169494 85026 169550
rect 85026 169494 85030 169550
rect 84966 169490 85030 169494
rect 85046 169550 85110 169554
rect 85046 169494 85050 169550
rect 85050 169494 85106 169550
rect 85106 169494 85110 169550
rect 85046 169490 85110 169494
rect 85126 169550 85190 169554
rect 85126 169494 85130 169550
rect 85130 169494 85186 169550
rect 85186 169494 85190 169550
rect 85126 169490 85190 169494
rect 2886 169006 2950 169010
rect 2886 168950 2890 169006
rect 2890 168950 2946 169006
rect 2946 168950 2950 169006
rect 2886 168946 2950 168950
rect 2966 169006 3030 169010
rect 2966 168950 2970 169006
rect 2970 168950 3026 169006
rect 3026 168950 3030 169006
rect 2966 168946 3030 168950
rect 3046 169006 3110 169010
rect 3046 168950 3050 169006
rect 3050 168950 3106 169006
rect 3106 168950 3110 169006
rect 3046 168946 3110 168950
rect 3126 169006 3190 169010
rect 3126 168950 3130 169006
rect 3130 168950 3186 169006
rect 3186 168950 3190 169006
rect 3126 168946 3190 168950
rect 86886 169006 86950 169010
rect 86886 168950 86890 169006
rect 86890 168950 86946 169006
rect 86946 168950 86950 169006
rect 86886 168946 86950 168950
rect 86966 169006 87030 169010
rect 86966 168950 86970 169006
rect 86970 168950 87026 169006
rect 87026 168950 87030 169006
rect 86966 168946 87030 168950
rect 87046 169006 87110 169010
rect 87046 168950 87050 169006
rect 87050 168950 87106 169006
rect 87106 168950 87110 169006
rect 87046 168946 87110 168950
rect 87126 169006 87190 169010
rect 87126 168950 87130 169006
rect 87130 168950 87186 169006
rect 87186 168950 87190 169006
rect 87126 168946 87190 168950
rect 83634 168606 83698 168670
rect 886 168462 950 168466
rect 886 168406 890 168462
rect 890 168406 946 168462
rect 946 168406 950 168462
rect 886 168402 950 168406
rect 966 168462 1030 168466
rect 966 168406 970 168462
rect 970 168406 1026 168462
rect 1026 168406 1030 168462
rect 966 168402 1030 168406
rect 1046 168462 1110 168466
rect 1046 168406 1050 168462
rect 1050 168406 1106 168462
rect 1106 168406 1110 168462
rect 1046 168402 1110 168406
rect 1126 168462 1190 168466
rect 1126 168406 1130 168462
rect 1130 168406 1186 168462
rect 1186 168406 1190 168462
rect 1126 168402 1190 168406
rect 84886 168462 84950 168466
rect 84886 168406 84890 168462
rect 84890 168406 84946 168462
rect 84946 168406 84950 168462
rect 84886 168402 84950 168406
rect 84966 168462 85030 168466
rect 84966 168406 84970 168462
rect 84970 168406 85026 168462
rect 85026 168406 85030 168462
rect 84966 168402 85030 168406
rect 85046 168462 85110 168466
rect 85046 168406 85050 168462
rect 85050 168406 85106 168462
rect 85106 168406 85110 168462
rect 85046 168402 85110 168406
rect 85126 168462 85190 168466
rect 85126 168406 85130 168462
rect 85130 168406 85186 168462
rect 85186 168406 85190 168462
rect 85126 168402 85190 168406
rect 2886 167918 2950 167922
rect 2886 167862 2890 167918
rect 2890 167862 2946 167918
rect 2946 167862 2950 167918
rect 2886 167858 2950 167862
rect 2966 167918 3030 167922
rect 2966 167862 2970 167918
rect 2970 167862 3026 167918
rect 3026 167862 3030 167918
rect 2966 167858 3030 167862
rect 3046 167918 3110 167922
rect 3046 167862 3050 167918
rect 3050 167862 3106 167918
rect 3106 167862 3110 167918
rect 3046 167858 3110 167862
rect 3126 167918 3190 167922
rect 3126 167862 3130 167918
rect 3130 167862 3186 167918
rect 3186 167862 3190 167918
rect 3126 167858 3190 167862
rect 86886 167918 86950 167922
rect 86886 167862 86890 167918
rect 86890 167862 86946 167918
rect 86946 167862 86950 167918
rect 86886 167858 86950 167862
rect 86966 167918 87030 167922
rect 86966 167862 86970 167918
rect 86970 167862 87026 167918
rect 87026 167862 87030 167918
rect 86966 167858 87030 167862
rect 87046 167918 87110 167922
rect 87046 167862 87050 167918
rect 87050 167862 87106 167918
rect 87106 167862 87110 167918
rect 87046 167858 87110 167862
rect 87126 167918 87190 167922
rect 87126 167862 87130 167918
rect 87130 167862 87186 167918
rect 87186 167862 87190 167918
rect 87126 167858 87190 167862
rect 84186 167518 84250 167582
rect 886 167374 950 167378
rect 886 167318 890 167374
rect 890 167318 946 167374
rect 946 167318 950 167374
rect 886 167314 950 167318
rect 966 167374 1030 167378
rect 966 167318 970 167374
rect 970 167318 1026 167374
rect 1026 167318 1030 167374
rect 966 167314 1030 167318
rect 1046 167374 1110 167378
rect 1046 167318 1050 167374
rect 1050 167318 1106 167374
rect 1106 167318 1110 167374
rect 1046 167314 1110 167318
rect 1126 167374 1190 167378
rect 1126 167318 1130 167374
rect 1130 167318 1186 167374
rect 1186 167318 1190 167374
rect 1126 167314 1190 167318
rect 84886 167374 84950 167378
rect 84886 167318 84890 167374
rect 84890 167318 84946 167374
rect 84946 167318 84950 167374
rect 84886 167314 84950 167318
rect 84966 167374 85030 167378
rect 84966 167318 84970 167374
rect 84970 167318 85026 167374
rect 85026 167318 85030 167374
rect 84966 167314 85030 167318
rect 85046 167374 85110 167378
rect 85046 167318 85050 167374
rect 85050 167318 85106 167374
rect 85106 167318 85110 167374
rect 85046 167314 85110 167318
rect 85126 167374 85190 167378
rect 85126 167318 85130 167374
rect 85130 167318 85186 167374
rect 85186 167318 85190 167374
rect 85126 167314 85190 167318
rect 2886 166830 2950 166834
rect 2886 166774 2890 166830
rect 2890 166774 2946 166830
rect 2946 166774 2950 166830
rect 2886 166770 2950 166774
rect 2966 166830 3030 166834
rect 2966 166774 2970 166830
rect 2970 166774 3026 166830
rect 3026 166774 3030 166830
rect 2966 166770 3030 166774
rect 3046 166830 3110 166834
rect 3046 166774 3050 166830
rect 3050 166774 3106 166830
rect 3106 166774 3110 166830
rect 3046 166770 3110 166774
rect 3126 166830 3190 166834
rect 3126 166774 3130 166830
rect 3130 166774 3186 166830
rect 3186 166774 3190 166830
rect 3126 166770 3190 166774
rect 86886 166830 86950 166834
rect 86886 166774 86890 166830
rect 86890 166774 86946 166830
rect 86946 166774 86950 166830
rect 86886 166770 86950 166774
rect 86966 166830 87030 166834
rect 86966 166774 86970 166830
rect 86970 166774 87026 166830
rect 87026 166774 87030 166830
rect 86966 166770 87030 166774
rect 87046 166830 87110 166834
rect 87046 166774 87050 166830
rect 87050 166774 87106 166830
rect 87106 166774 87110 166830
rect 87046 166770 87110 166774
rect 87126 166830 87190 166834
rect 87126 166774 87130 166830
rect 87130 166774 87186 166830
rect 87186 166774 87190 166830
rect 87126 166770 87190 166774
rect 886 166286 950 166290
rect 886 166230 890 166286
rect 890 166230 946 166286
rect 946 166230 950 166286
rect 886 166226 950 166230
rect 966 166286 1030 166290
rect 966 166230 970 166286
rect 970 166230 1026 166286
rect 1026 166230 1030 166286
rect 966 166226 1030 166230
rect 1046 166286 1110 166290
rect 1046 166230 1050 166286
rect 1050 166230 1106 166286
rect 1106 166230 1110 166286
rect 1046 166226 1110 166230
rect 1126 166286 1190 166290
rect 1126 166230 1130 166286
rect 1130 166230 1186 166286
rect 1186 166230 1190 166286
rect 1126 166226 1190 166230
rect 84886 166286 84950 166290
rect 84886 166230 84890 166286
rect 84890 166230 84946 166286
rect 84946 166230 84950 166286
rect 84886 166226 84950 166230
rect 84966 166286 85030 166290
rect 84966 166230 84970 166286
rect 84970 166230 85026 166286
rect 85026 166230 85030 166286
rect 84966 166226 85030 166230
rect 85046 166286 85110 166290
rect 85046 166230 85050 166286
rect 85050 166230 85106 166286
rect 85106 166230 85110 166286
rect 85046 166226 85110 166230
rect 85126 166286 85190 166290
rect 85126 166230 85130 166286
rect 85130 166230 85186 166286
rect 85186 166230 85190 166286
rect 85126 166226 85190 166230
rect 83450 166022 83514 166086
rect 2886 165742 2950 165746
rect 2886 165686 2890 165742
rect 2890 165686 2946 165742
rect 2946 165686 2950 165742
rect 2886 165682 2950 165686
rect 2966 165742 3030 165746
rect 2966 165686 2970 165742
rect 2970 165686 3026 165742
rect 3026 165686 3030 165742
rect 2966 165682 3030 165686
rect 3046 165742 3110 165746
rect 3046 165686 3050 165742
rect 3050 165686 3106 165742
rect 3106 165686 3110 165742
rect 3046 165682 3110 165686
rect 3126 165742 3190 165746
rect 3126 165686 3130 165742
rect 3130 165686 3186 165742
rect 3186 165686 3190 165742
rect 3126 165682 3190 165686
rect 86886 165742 86950 165746
rect 86886 165686 86890 165742
rect 86890 165686 86946 165742
rect 86946 165686 86950 165742
rect 86886 165682 86950 165686
rect 86966 165742 87030 165746
rect 86966 165686 86970 165742
rect 86970 165686 87026 165742
rect 87026 165686 87030 165742
rect 86966 165682 87030 165686
rect 87046 165742 87110 165746
rect 87046 165686 87050 165742
rect 87050 165686 87106 165742
rect 87106 165686 87110 165742
rect 87046 165682 87110 165686
rect 87126 165742 87190 165746
rect 87126 165686 87130 165742
rect 87130 165686 87186 165742
rect 87186 165686 87190 165742
rect 87126 165682 87190 165686
rect 886 165198 950 165202
rect 886 165142 890 165198
rect 890 165142 946 165198
rect 946 165142 950 165198
rect 886 165138 950 165142
rect 966 165198 1030 165202
rect 966 165142 970 165198
rect 970 165142 1026 165198
rect 1026 165142 1030 165198
rect 966 165138 1030 165142
rect 1046 165198 1110 165202
rect 1046 165142 1050 165198
rect 1050 165142 1106 165198
rect 1106 165142 1110 165198
rect 1046 165138 1110 165142
rect 1126 165198 1190 165202
rect 1126 165142 1130 165198
rect 1130 165142 1186 165198
rect 1186 165142 1190 165198
rect 1126 165138 1190 165142
rect 84886 165198 84950 165202
rect 84886 165142 84890 165198
rect 84890 165142 84946 165198
rect 84946 165142 84950 165198
rect 84886 165138 84950 165142
rect 84966 165198 85030 165202
rect 84966 165142 84970 165198
rect 84970 165142 85026 165198
rect 85026 165142 85030 165198
rect 84966 165138 85030 165142
rect 85046 165198 85110 165202
rect 85046 165142 85050 165198
rect 85050 165142 85106 165198
rect 85106 165142 85110 165198
rect 85046 165138 85110 165142
rect 85126 165198 85190 165202
rect 85126 165142 85130 165198
rect 85130 165142 85186 165198
rect 85186 165142 85190 165198
rect 85126 165138 85190 165142
rect 84370 164994 84434 164998
rect 84370 164938 84420 164994
rect 84420 164938 84434 164994
rect 84370 164934 84434 164938
rect 84554 164858 84618 164862
rect 84554 164802 84604 164858
rect 84604 164802 84618 164858
rect 84554 164798 84618 164802
rect 2886 164654 2950 164658
rect 2886 164598 2890 164654
rect 2890 164598 2946 164654
rect 2946 164598 2950 164654
rect 2886 164594 2950 164598
rect 2966 164654 3030 164658
rect 2966 164598 2970 164654
rect 2970 164598 3026 164654
rect 3026 164598 3030 164654
rect 2966 164594 3030 164598
rect 3046 164654 3110 164658
rect 3046 164598 3050 164654
rect 3050 164598 3106 164654
rect 3106 164598 3110 164654
rect 3046 164594 3110 164598
rect 3126 164654 3190 164658
rect 3126 164598 3130 164654
rect 3130 164598 3186 164654
rect 3186 164598 3190 164654
rect 3126 164594 3190 164598
rect 86886 164654 86950 164658
rect 86886 164598 86890 164654
rect 86890 164598 86946 164654
rect 86946 164598 86950 164654
rect 86886 164594 86950 164598
rect 86966 164654 87030 164658
rect 86966 164598 86970 164654
rect 86970 164598 87026 164654
rect 87026 164598 87030 164654
rect 86966 164594 87030 164598
rect 87046 164654 87110 164658
rect 87046 164598 87050 164654
rect 87050 164598 87106 164654
rect 87106 164598 87110 164654
rect 87046 164594 87110 164598
rect 87126 164654 87190 164658
rect 87126 164598 87130 164654
rect 87130 164598 87186 164654
rect 87186 164598 87190 164654
rect 87126 164594 87190 164598
rect 84370 164390 84434 164454
rect 84554 164254 84618 164318
rect 886 164110 950 164114
rect 886 164054 890 164110
rect 890 164054 946 164110
rect 946 164054 950 164110
rect 886 164050 950 164054
rect 966 164110 1030 164114
rect 966 164054 970 164110
rect 970 164054 1026 164110
rect 1026 164054 1030 164110
rect 966 164050 1030 164054
rect 1046 164110 1110 164114
rect 1046 164054 1050 164110
rect 1050 164054 1106 164110
rect 1106 164054 1110 164110
rect 1046 164050 1110 164054
rect 1126 164110 1190 164114
rect 1126 164054 1130 164110
rect 1130 164054 1186 164110
rect 1186 164054 1190 164110
rect 1126 164050 1190 164054
rect 84886 164110 84950 164114
rect 84886 164054 84890 164110
rect 84890 164054 84946 164110
rect 84946 164054 84950 164110
rect 84886 164050 84950 164054
rect 84966 164110 85030 164114
rect 84966 164054 84970 164110
rect 84970 164054 85026 164110
rect 85026 164054 85030 164110
rect 84966 164050 85030 164054
rect 85046 164110 85110 164114
rect 85046 164054 85050 164110
rect 85050 164054 85106 164110
rect 85106 164054 85110 164110
rect 85046 164050 85110 164054
rect 85126 164110 85190 164114
rect 85126 164054 85130 164110
rect 85130 164054 85186 164110
rect 85186 164054 85190 164110
rect 85126 164050 85190 164054
rect 2886 163566 2950 163570
rect 2886 163510 2890 163566
rect 2890 163510 2946 163566
rect 2946 163510 2950 163566
rect 2886 163506 2950 163510
rect 2966 163566 3030 163570
rect 2966 163510 2970 163566
rect 2970 163510 3026 163566
rect 3026 163510 3030 163566
rect 2966 163506 3030 163510
rect 3046 163566 3110 163570
rect 3046 163510 3050 163566
rect 3050 163510 3106 163566
rect 3106 163510 3110 163566
rect 3046 163506 3110 163510
rect 3126 163566 3190 163570
rect 3126 163510 3130 163566
rect 3130 163510 3186 163566
rect 3186 163510 3190 163566
rect 3126 163506 3190 163510
rect 86886 163566 86950 163570
rect 86886 163510 86890 163566
rect 86890 163510 86946 163566
rect 86946 163510 86950 163566
rect 86886 163506 86950 163510
rect 86966 163566 87030 163570
rect 86966 163510 86970 163566
rect 86970 163510 87026 163566
rect 87026 163510 87030 163566
rect 86966 163506 87030 163510
rect 87046 163566 87110 163570
rect 87046 163510 87050 163566
rect 87050 163510 87106 163566
rect 87106 163510 87110 163566
rect 87046 163506 87110 163510
rect 87126 163566 87190 163570
rect 87126 163510 87130 163566
rect 87130 163510 87186 163566
rect 87186 163510 87190 163566
rect 87126 163506 87190 163510
rect 886 163022 950 163026
rect 886 162966 890 163022
rect 890 162966 946 163022
rect 946 162966 950 163022
rect 886 162962 950 162966
rect 966 163022 1030 163026
rect 966 162966 970 163022
rect 970 162966 1026 163022
rect 1026 162966 1030 163022
rect 966 162962 1030 162966
rect 1046 163022 1110 163026
rect 1046 162966 1050 163022
rect 1050 162966 1106 163022
rect 1106 162966 1110 163022
rect 1046 162962 1110 162966
rect 1126 163022 1190 163026
rect 1126 162966 1130 163022
rect 1130 162966 1186 163022
rect 1186 162966 1190 163022
rect 1126 162962 1190 162966
rect 84886 163022 84950 163026
rect 84886 162966 84890 163022
rect 84890 162966 84946 163022
rect 84946 162966 84950 163022
rect 84886 162962 84950 162966
rect 84966 163022 85030 163026
rect 84966 162966 84970 163022
rect 84970 162966 85026 163022
rect 85026 162966 85030 163022
rect 84966 162962 85030 162966
rect 85046 163022 85110 163026
rect 85046 162966 85050 163022
rect 85050 162966 85106 163022
rect 85106 162966 85110 163022
rect 85046 162962 85110 162966
rect 85126 163022 85190 163026
rect 85126 162966 85130 163022
rect 85130 162966 85186 163022
rect 85186 162966 85190 163022
rect 85126 162962 85190 162966
rect 2886 162478 2950 162482
rect 2886 162422 2890 162478
rect 2890 162422 2946 162478
rect 2946 162422 2950 162478
rect 2886 162418 2950 162422
rect 2966 162478 3030 162482
rect 2966 162422 2970 162478
rect 2970 162422 3026 162478
rect 3026 162422 3030 162478
rect 2966 162418 3030 162422
rect 3046 162478 3110 162482
rect 3046 162422 3050 162478
rect 3050 162422 3106 162478
rect 3106 162422 3110 162478
rect 3046 162418 3110 162422
rect 3126 162478 3190 162482
rect 3126 162422 3130 162478
rect 3130 162422 3186 162478
rect 3186 162422 3190 162478
rect 3126 162418 3190 162422
rect 86886 162478 86950 162482
rect 86886 162422 86890 162478
rect 86890 162422 86946 162478
rect 86946 162422 86950 162478
rect 86886 162418 86950 162422
rect 86966 162478 87030 162482
rect 86966 162422 86970 162478
rect 86970 162422 87026 162478
rect 87026 162422 87030 162478
rect 86966 162418 87030 162422
rect 87046 162478 87110 162482
rect 87046 162422 87050 162478
rect 87050 162422 87106 162478
rect 87106 162422 87110 162478
rect 87046 162418 87110 162422
rect 87126 162478 87190 162482
rect 87126 162422 87130 162478
rect 87130 162422 87186 162478
rect 87186 162422 87190 162478
rect 87126 162418 87190 162422
rect 886 161934 950 161938
rect 886 161878 890 161934
rect 890 161878 946 161934
rect 946 161878 950 161934
rect 886 161874 950 161878
rect 966 161934 1030 161938
rect 966 161878 970 161934
rect 970 161878 1026 161934
rect 1026 161878 1030 161934
rect 966 161874 1030 161878
rect 1046 161934 1110 161938
rect 1046 161878 1050 161934
rect 1050 161878 1106 161934
rect 1106 161878 1110 161934
rect 1046 161874 1110 161878
rect 1126 161934 1190 161938
rect 1126 161878 1130 161934
rect 1130 161878 1186 161934
rect 1186 161878 1190 161934
rect 1126 161874 1190 161878
rect 84886 161934 84950 161938
rect 84886 161878 84890 161934
rect 84890 161878 84946 161934
rect 84946 161878 84950 161934
rect 84886 161874 84950 161878
rect 84966 161934 85030 161938
rect 84966 161878 84970 161934
rect 84970 161878 85026 161934
rect 85026 161878 85030 161934
rect 84966 161874 85030 161878
rect 85046 161934 85110 161938
rect 85046 161878 85050 161934
rect 85050 161878 85106 161934
rect 85106 161878 85110 161934
rect 85046 161874 85110 161878
rect 85126 161934 85190 161938
rect 85126 161878 85130 161934
rect 85130 161878 85186 161934
rect 85186 161878 85190 161934
rect 85126 161874 85190 161878
rect 2886 161390 2950 161394
rect 2886 161334 2890 161390
rect 2890 161334 2946 161390
rect 2946 161334 2950 161390
rect 2886 161330 2950 161334
rect 2966 161390 3030 161394
rect 2966 161334 2970 161390
rect 2970 161334 3026 161390
rect 3026 161334 3030 161390
rect 2966 161330 3030 161334
rect 3046 161390 3110 161394
rect 3046 161334 3050 161390
rect 3050 161334 3106 161390
rect 3106 161334 3110 161390
rect 3046 161330 3110 161334
rect 3126 161390 3190 161394
rect 3126 161334 3130 161390
rect 3130 161334 3186 161390
rect 3186 161334 3190 161390
rect 3126 161330 3190 161334
rect 86886 161390 86950 161394
rect 86886 161334 86890 161390
rect 86890 161334 86946 161390
rect 86946 161334 86950 161390
rect 86886 161330 86950 161334
rect 86966 161390 87030 161394
rect 86966 161334 86970 161390
rect 86970 161334 87026 161390
rect 87026 161334 87030 161390
rect 86966 161330 87030 161334
rect 87046 161390 87110 161394
rect 87046 161334 87050 161390
rect 87050 161334 87106 161390
rect 87106 161334 87110 161390
rect 87046 161330 87110 161334
rect 87126 161390 87190 161394
rect 87126 161334 87130 161390
rect 87130 161334 87186 161390
rect 87186 161334 87190 161390
rect 87126 161330 87190 161334
rect 886 160846 950 160850
rect 886 160790 890 160846
rect 890 160790 946 160846
rect 946 160790 950 160846
rect 886 160786 950 160790
rect 966 160846 1030 160850
rect 966 160790 970 160846
rect 970 160790 1026 160846
rect 1026 160790 1030 160846
rect 966 160786 1030 160790
rect 1046 160846 1110 160850
rect 1046 160790 1050 160846
rect 1050 160790 1106 160846
rect 1106 160790 1110 160846
rect 1046 160786 1110 160790
rect 1126 160846 1190 160850
rect 1126 160790 1130 160846
rect 1130 160790 1186 160846
rect 1186 160790 1190 160846
rect 1126 160786 1190 160790
rect 84886 160846 84950 160850
rect 84886 160790 84890 160846
rect 84890 160790 84946 160846
rect 84946 160790 84950 160846
rect 84886 160786 84950 160790
rect 84966 160846 85030 160850
rect 84966 160790 84970 160846
rect 84970 160790 85026 160846
rect 85026 160790 85030 160846
rect 84966 160786 85030 160790
rect 85046 160846 85110 160850
rect 85046 160790 85050 160846
rect 85050 160790 85106 160846
rect 85106 160790 85110 160846
rect 85046 160786 85110 160790
rect 85126 160846 85190 160850
rect 85126 160790 85130 160846
rect 85130 160790 85186 160846
rect 85186 160790 85190 160846
rect 85126 160786 85190 160790
rect 2886 160302 2950 160306
rect 2886 160246 2890 160302
rect 2890 160246 2946 160302
rect 2946 160246 2950 160302
rect 2886 160242 2950 160246
rect 2966 160302 3030 160306
rect 2966 160246 2970 160302
rect 2970 160246 3026 160302
rect 3026 160246 3030 160302
rect 2966 160242 3030 160246
rect 3046 160302 3110 160306
rect 3046 160246 3050 160302
rect 3050 160246 3106 160302
rect 3106 160246 3110 160302
rect 3046 160242 3110 160246
rect 3126 160302 3190 160306
rect 3126 160246 3130 160302
rect 3130 160246 3186 160302
rect 3186 160246 3190 160302
rect 3126 160242 3190 160246
rect 86886 160302 86950 160306
rect 86886 160246 86890 160302
rect 86890 160246 86946 160302
rect 86946 160246 86950 160302
rect 86886 160242 86950 160246
rect 86966 160302 87030 160306
rect 86966 160246 86970 160302
rect 86970 160246 87026 160302
rect 87026 160246 87030 160302
rect 86966 160242 87030 160246
rect 87046 160302 87110 160306
rect 87046 160246 87050 160302
rect 87050 160246 87106 160302
rect 87106 160246 87110 160302
rect 87046 160242 87110 160246
rect 87126 160302 87190 160306
rect 87126 160246 87130 160302
rect 87130 160246 87186 160302
rect 87186 160246 87190 160302
rect 87126 160242 87190 160246
rect 886 159758 950 159762
rect 886 159702 890 159758
rect 890 159702 946 159758
rect 946 159702 950 159758
rect 886 159698 950 159702
rect 966 159758 1030 159762
rect 966 159702 970 159758
rect 970 159702 1026 159758
rect 1026 159702 1030 159758
rect 966 159698 1030 159702
rect 1046 159758 1110 159762
rect 1046 159702 1050 159758
rect 1050 159702 1106 159758
rect 1106 159702 1110 159758
rect 1046 159698 1110 159702
rect 1126 159758 1190 159762
rect 1126 159702 1130 159758
rect 1130 159702 1186 159758
rect 1186 159702 1190 159758
rect 1126 159698 1190 159702
rect 84886 159758 84950 159762
rect 84886 159702 84890 159758
rect 84890 159702 84946 159758
rect 84946 159702 84950 159758
rect 84886 159698 84950 159702
rect 84966 159758 85030 159762
rect 84966 159702 84970 159758
rect 84970 159702 85026 159758
rect 85026 159702 85030 159758
rect 84966 159698 85030 159702
rect 85046 159758 85110 159762
rect 85046 159702 85050 159758
rect 85050 159702 85106 159758
rect 85106 159702 85110 159758
rect 85046 159698 85110 159702
rect 85126 159758 85190 159762
rect 85126 159702 85130 159758
rect 85130 159702 85186 159758
rect 85186 159702 85190 159758
rect 85126 159698 85190 159702
rect 2886 159214 2950 159218
rect 2886 159158 2890 159214
rect 2890 159158 2946 159214
rect 2946 159158 2950 159214
rect 2886 159154 2950 159158
rect 2966 159214 3030 159218
rect 2966 159158 2970 159214
rect 2970 159158 3026 159214
rect 3026 159158 3030 159214
rect 2966 159154 3030 159158
rect 3046 159214 3110 159218
rect 3046 159158 3050 159214
rect 3050 159158 3106 159214
rect 3106 159158 3110 159214
rect 3046 159154 3110 159158
rect 3126 159214 3190 159218
rect 3126 159158 3130 159214
rect 3130 159158 3186 159214
rect 3186 159158 3190 159214
rect 3126 159154 3190 159158
rect 86886 159214 86950 159218
rect 86886 159158 86890 159214
rect 86890 159158 86946 159214
rect 86946 159158 86950 159214
rect 86886 159154 86950 159158
rect 86966 159214 87030 159218
rect 86966 159158 86970 159214
rect 86970 159158 87026 159214
rect 87026 159158 87030 159214
rect 86966 159154 87030 159158
rect 87046 159214 87110 159218
rect 87046 159158 87050 159214
rect 87050 159158 87106 159214
rect 87106 159158 87110 159214
rect 87046 159154 87110 159158
rect 87126 159214 87190 159218
rect 87126 159158 87130 159214
rect 87130 159158 87186 159214
rect 87186 159158 87190 159214
rect 87126 159154 87190 159158
rect 886 158670 950 158674
rect 886 158614 890 158670
rect 890 158614 946 158670
rect 946 158614 950 158670
rect 886 158610 950 158614
rect 966 158670 1030 158674
rect 966 158614 970 158670
rect 970 158614 1026 158670
rect 1026 158614 1030 158670
rect 966 158610 1030 158614
rect 1046 158670 1110 158674
rect 1046 158614 1050 158670
rect 1050 158614 1106 158670
rect 1106 158614 1110 158670
rect 1046 158610 1110 158614
rect 1126 158670 1190 158674
rect 1126 158614 1130 158670
rect 1130 158614 1186 158670
rect 1186 158614 1190 158670
rect 1126 158610 1190 158614
rect 84886 158670 84950 158674
rect 84886 158614 84890 158670
rect 84890 158614 84946 158670
rect 84946 158614 84950 158670
rect 84886 158610 84950 158614
rect 84966 158670 85030 158674
rect 84966 158614 84970 158670
rect 84970 158614 85026 158670
rect 85026 158614 85030 158670
rect 84966 158610 85030 158614
rect 85046 158670 85110 158674
rect 85046 158614 85050 158670
rect 85050 158614 85106 158670
rect 85106 158614 85110 158670
rect 85046 158610 85110 158614
rect 85126 158670 85190 158674
rect 85126 158614 85130 158670
rect 85130 158614 85186 158670
rect 85186 158614 85190 158670
rect 85126 158610 85190 158614
rect 2886 158126 2950 158130
rect 2886 158070 2890 158126
rect 2890 158070 2946 158126
rect 2946 158070 2950 158126
rect 2886 158066 2950 158070
rect 2966 158126 3030 158130
rect 2966 158070 2970 158126
rect 2970 158070 3026 158126
rect 3026 158070 3030 158126
rect 2966 158066 3030 158070
rect 3046 158126 3110 158130
rect 3046 158070 3050 158126
rect 3050 158070 3106 158126
rect 3106 158070 3110 158126
rect 3046 158066 3110 158070
rect 3126 158126 3190 158130
rect 3126 158070 3130 158126
rect 3130 158070 3186 158126
rect 3186 158070 3190 158126
rect 3126 158066 3190 158070
rect 86886 158126 86950 158130
rect 86886 158070 86890 158126
rect 86890 158070 86946 158126
rect 86946 158070 86950 158126
rect 86886 158066 86950 158070
rect 86966 158126 87030 158130
rect 86966 158070 86970 158126
rect 86970 158070 87026 158126
rect 87026 158070 87030 158126
rect 86966 158066 87030 158070
rect 87046 158126 87110 158130
rect 87046 158070 87050 158126
rect 87050 158070 87106 158126
rect 87106 158070 87110 158126
rect 87046 158066 87110 158070
rect 87126 158126 87190 158130
rect 87126 158070 87130 158126
rect 87130 158070 87186 158126
rect 87186 158070 87190 158126
rect 87126 158066 87190 158070
rect 886 157582 950 157586
rect 886 157526 890 157582
rect 890 157526 946 157582
rect 946 157526 950 157582
rect 886 157522 950 157526
rect 966 157582 1030 157586
rect 966 157526 970 157582
rect 970 157526 1026 157582
rect 1026 157526 1030 157582
rect 966 157522 1030 157526
rect 1046 157582 1110 157586
rect 1046 157526 1050 157582
rect 1050 157526 1106 157582
rect 1106 157526 1110 157582
rect 1046 157522 1110 157526
rect 1126 157582 1190 157586
rect 1126 157526 1130 157582
rect 1130 157526 1186 157582
rect 1186 157526 1190 157582
rect 1126 157522 1190 157526
rect 84886 157582 84950 157586
rect 84886 157526 84890 157582
rect 84890 157526 84946 157582
rect 84946 157526 84950 157582
rect 84886 157522 84950 157526
rect 84966 157582 85030 157586
rect 84966 157526 84970 157582
rect 84970 157526 85026 157582
rect 85026 157526 85030 157582
rect 84966 157522 85030 157526
rect 85046 157582 85110 157586
rect 85046 157526 85050 157582
rect 85050 157526 85106 157582
rect 85106 157526 85110 157582
rect 85046 157522 85110 157526
rect 85126 157582 85190 157586
rect 85126 157526 85130 157582
rect 85130 157526 85186 157582
rect 85186 157526 85190 157582
rect 85126 157522 85190 157526
rect 2886 157038 2950 157042
rect 2886 156982 2890 157038
rect 2890 156982 2946 157038
rect 2946 156982 2950 157038
rect 2886 156978 2950 156982
rect 2966 157038 3030 157042
rect 2966 156982 2970 157038
rect 2970 156982 3026 157038
rect 3026 156982 3030 157038
rect 2966 156978 3030 156982
rect 3046 157038 3110 157042
rect 3046 156982 3050 157038
rect 3050 156982 3106 157038
rect 3106 156982 3110 157038
rect 3046 156978 3110 156982
rect 3126 157038 3190 157042
rect 3126 156982 3130 157038
rect 3130 156982 3186 157038
rect 3186 156982 3190 157038
rect 3126 156978 3190 156982
rect 86886 157038 86950 157042
rect 86886 156982 86890 157038
rect 86890 156982 86946 157038
rect 86946 156982 86950 157038
rect 86886 156978 86950 156982
rect 86966 157038 87030 157042
rect 86966 156982 86970 157038
rect 86970 156982 87026 157038
rect 87026 156982 87030 157038
rect 86966 156978 87030 156982
rect 87046 157038 87110 157042
rect 87046 156982 87050 157038
rect 87050 156982 87106 157038
rect 87106 156982 87110 157038
rect 87046 156978 87110 156982
rect 87126 157038 87190 157042
rect 87126 156982 87130 157038
rect 87130 156982 87186 157038
rect 87186 156982 87190 157038
rect 87126 156978 87190 156982
rect 886 156494 950 156498
rect 886 156438 890 156494
rect 890 156438 946 156494
rect 946 156438 950 156494
rect 886 156434 950 156438
rect 966 156494 1030 156498
rect 966 156438 970 156494
rect 970 156438 1026 156494
rect 1026 156438 1030 156494
rect 966 156434 1030 156438
rect 1046 156494 1110 156498
rect 1046 156438 1050 156494
rect 1050 156438 1106 156494
rect 1106 156438 1110 156494
rect 1046 156434 1110 156438
rect 1126 156494 1190 156498
rect 1126 156438 1130 156494
rect 1130 156438 1186 156494
rect 1186 156438 1190 156494
rect 1126 156434 1190 156438
rect 84886 156494 84950 156498
rect 84886 156438 84890 156494
rect 84890 156438 84946 156494
rect 84946 156438 84950 156494
rect 84886 156434 84950 156438
rect 84966 156494 85030 156498
rect 84966 156438 84970 156494
rect 84970 156438 85026 156494
rect 85026 156438 85030 156494
rect 84966 156434 85030 156438
rect 85046 156494 85110 156498
rect 85046 156438 85050 156494
rect 85050 156438 85106 156494
rect 85106 156438 85110 156494
rect 85046 156434 85110 156438
rect 85126 156494 85190 156498
rect 85126 156438 85130 156494
rect 85130 156438 85186 156494
rect 85186 156438 85190 156494
rect 85126 156434 85190 156438
rect 2886 155950 2950 155954
rect 2886 155894 2890 155950
rect 2890 155894 2946 155950
rect 2946 155894 2950 155950
rect 2886 155890 2950 155894
rect 2966 155950 3030 155954
rect 2966 155894 2970 155950
rect 2970 155894 3026 155950
rect 3026 155894 3030 155950
rect 2966 155890 3030 155894
rect 3046 155950 3110 155954
rect 3046 155894 3050 155950
rect 3050 155894 3106 155950
rect 3106 155894 3110 155950
rect 3046 155890 3110 155894
rect 3126 155950 3190 155954
rect 3126 155894 3130 155950
rect 3130 155894 3186 155950
rect 3186 155894 3190 155950
rect 3126 155890 3190 155894
rect 86886 155950 86950 155954
rect 86886 155894 86890 155950
rect 86890 155894 86946 155950
rect 86946 155894 86950 155950
rect 86886 155890 86950 155894
rect 86966 155950 87030 155954
rect 86966 155894 86970 155950
rect 86970 155894 87026 155950
rect 87026 155894 87030 155950
rect 86966 155890 87030 155894
rect 87046 155950 87110 155954
rect 87046 155894 87050 155950
rect 87050 155894 87106 155950
rect 87106 155894 87110 155950
rect 87046 155890 87110 155894
rect 87126 155950 87190 155954
rect 87126 155894 87130 155950
rect 87130 155894 87186 155950
rect 87186 155894 87190 155950
rect 87126 155890 87190 155894
rect 886 155406 950 155410
rect 886 155350 890 155406
rect 890 155350 946 155406
rect 946 155350 950 155406
rect 886 155346 950 155350
rect 966 155406 1030 155410
rect 966 155350 970 155406
rect 970 155350 1026 155406
rect 1026 155350 1030 155406
rect 966 155346 1030 155350
rect 1046 155406 1110 155410
rect 1046 155350 1050 155406
rect 1050 155350 1106 155406
rect 1106 155350 1110 155406
rect 1046 155346 1110 155350
rect 1126 155406 1190 155410
rect 1126 155350 1130 155406
rect 1130 155350 1186 155406
rect 1186 155350 1190 155406
rect 1126 155346 1190 155350
rect 84886 155406 84950 155410
rect 84886 155350 84890 155406
rect 84890 155350 84946 155406
rect 84946 155350 84950 155406
rect 84886 155346 84950 155350
rect 84966 155406 85030 155410
rect 84966 155350 84970 155406
rect 84970 155350 85026 155406
rect 85026 155350 85030 155406
rect 84966 155346 85030 155350
rect 85046 155406 85110 155410
rect 85046 155350 85050 155406
rect 85050 155350 85106 155406
rect 85106 155350 85110 155406
rect 85046 155346 85110 155350
rect 85126 155406 85190 155410
rect 85126 155350 85130 155406
rect 85130 155350 85186 155406
rect 85186 155350 85190 155406
rect 85126 155346 85190 155350
rect 2886 154862 2950 154866
rect 2886 154806 2890 154862
rect 2890 154806 2946 154862
rect 2946 154806 2950 154862
rect 2886 154802 2950 154806
rect 2966 154862 3030 154866
rect 2966 154806 2970 154862
rect 2970 154806 3026 154862
rect 3026 154806 3030 154862
rect 2966 154802 3030 154806
rect 3046 154862 3110 154866
rect 3046 154806 3050 154862
rect 3050 154806 3106 154862
rect 3106 154806 3110 154862
rect 3046 154802 3110 154806
rect 3126 154862 3190 154866
rect 3126 154806 3130 154862
rect 3130 154806 3186 154862
rect 3186 154806 3190 154862
rect 3126 154802 3190 154806
rect 86886 154862 86950 154866
rect 86886 154806 86890 154862
rect 86890 154806 86946 154862
rect 86946 154806 86950 154862
rect 86886 154802 86950 154806
rect 86966 154862 87030 154866
rect 86966 154806 86970 154862
rect 86970 154806 87026 154862
rect 87026 154806 87030 154862
rect 86966 154802 87030 154806
rect 87046 154862 87110 154866
rect 87046 154806 87050 154862
rect 87050 154806 87106 154862
rect 87106 154806 87110 154862
rect 87046 154802 87110 154806
rect 87126 154862 87190 154866
rect 87126 154806 87130 154862
rect 87130 154806 87186 154862
rect 87186 154806 87190 154862
rect 87126 154802 87190 154806
rect 886 154318 950 154322
rect 886 154262 890 154318
rect 890 154262 946 154318
rect 946 154262 950 154318
rect 886 154258 950 154262
rect 966 154318 1030 154322
rect 966 154262 970 154318
rect 970 154262 1026 154318
rect 1026 154262 1030 154318
rect 966 154258 1030 154262
rect 1046 154318 1110 154322
rect 1046 154262 1050 154318
rect 1050 154262 1106 154318
rect 1106 154262 1110 154318
rect 1046 154258 1110 154262
rect 1126 154318 1190 154322
rect 1126 154262 1130 154318
rect 1130 154262 1186 154318
rect 1186 154262 1190 154318
rect 1126 154258 1190 154262
rect 84886 154318 84950 154322
rect 84886 154262 84890 154318
rect 84890 154262 84946 154318
rect 84946 154262 84950 154318
rect 84886 154258 84950 154262
rect 84966 154318 85030 154322
rect 84966 154262 84970 154318
rect 84970 154262 85026 154318
rect 85026 154262 85030 154318
rect 84966 154258 85030 154262
rect 85046 154318 85110 154322
rect 85046 154262 85050 154318
rect 85050 154262 85106 154318
rect 85106 154262 85110 154318
rect 85046 154258 85110 154262
rect 85126 154318 85190 154322
rect 85126 154262 85130 154318
rect 85130 154262 85186 154318
rect 85186 154262 85190 154318
rect 85126 154258 85190 154262
rect 2886 153774 2950 153778
rect 2886 153718 2890 153774
rect 2890 153718 2946 153774
rect 2946 153718 2950 153774
rect 2886 153714 2950 153718
rect 2966 153774 3030 153778
rect 2966 153718 2970 153774
rect 2970 153718 3026 153774
rect 3026 153718 3030 153774
rect 2966 153714 3030 153718
rect 3046 153774 3110 153778
rect 3046 153718 3050 153774
rect 3050 153718 3106 153774
rect 3106 153718 3110 153774
rect 3046 153714 3110 153718
rect 3126 153774 3190 153778
rect 3126 153718 3130 153774
rect 3130 153718 3186 153774
rect 3186 153718 3190 153774
rect 3126 153714 3190 153718
rect 86886 153774 86950 153778
rect 86886 153718 86890 153774
rect 86890 153718 86946 153774
rect 86946 153718 86950 153774
rect 86886 153714 86950 153718
rect 86966 153774 87030 153778
rect 86966 153718 86970 153774
rect 86970 153718 87026 153774
rect 87026 153718 87030 153774
rect 86966 153714 87030 153718
rect 87046 153774 87110 153778
rect 87046 153718 87050 153774
rect 87050 153718 87106 153774
rect 87106 153718 87110 153774
rect 87046 153714 87110 153718
rect 87126 153774 87190 153778
rect 87126 153718 87130 153774
rect 87130 153718 87186 153774
rect 87186 153718 87190 153774
rect 87126 153714 87190 153718
rect 886 153230 950 153234
rect 886 153174 890 153230
rect 890 153174 946 153230
rect 946 153174 950 153230
rect 886 153170 950 153174
rect 966 153230 1030 153234
rect 966 153174 970 153230
rect 970 153174 1026 153230
rect 1026 153174 1030 153230
rect 966 153170 1030 153174
rect 1046 153230 1110 153234
rect 1046 153174 1050 153230
rect 1050 153174 1106 153230
rect 1106 153174 1110 153230
rect 1046 153170 1110 153174
rect 1126 153230 1190 153234
rect 1126 153174 1130 153230
rect 1130 153174 1186 153230
rect 1186 153174 1190 153230
rect 1126 153170 1190 153174
rect 84886 153230 84950 153234
rect 84886 153174 84890 153230
rect 84890 153174 84946 153230
rect 84946 153174 84950 153230
rect 84886 153170 84950 153174
rect 84966 153230 85030 153234
rect 84966 153174 84970 153230
rect 84970 153174 85026 153230
rect 85026 153174 85030 153230
rect 84966 153170 85030 153174
rect 85046 153230 85110 153234
rect 85046 153174 85050 153230
rect 85050 153174 85106 153230
rect 85106 153174 85110 153230
rect 85046 153170 85110 153174
rect 85126 153230 85190 153234
rect 85126 153174 85130 153230
rect 85130 153174 85186 153230
rect 85186 153174 85190 153230
rect 85126 153170 85190 153174
rect 2886 152686 2950 152690
rect 2886 152630 2890 152686
rect 2890 152630 2946 152686
rect 2946 152630 2950 152686
rect 2886 152626 2950 152630
rect 2966 152686 3030 152690
rect 2966 152630 2970 152686
rect 2970 152630 3026 152686
rect 3026 152630 3030 152686
rect 2966 152626 3030 152630
rect 3046 152686 3110 152690
rect 3046 152630 3050 152686
rect 3050 152630 3106 152686
rect 3106 152630 3110 152686
rect 3046 152626 3110 152630
rect 3126 152686 3190 152690
rect 3126 152630 3130 152686
rect 3130 152630 3186 152686
rect 3186 152630 3190 152686
rect 3126 152626 3190 152630
rect 86886 152686 86950 152690
rect 86886 152630 86890 152686
rect 86890 152630 86946 152686
rect 86946 152630 86950 152686
rect 86886 152626 86950 152630
rect 86966 152686 87030 152690
rect 86966 152630 86970 152686
rect 86970 152630 87026 152686
rect 87026 152630 87030 152686
rect 86966 152626 87030 152630
rect 87046 152686 87110 152690
rect 87046 152630 87050 152686
rect 87050 152630 87106 152686
rect 87106 152630 87110 152686
rect 87046 152626 87110 152630
rect 87126 152686 87190 152690
rect 87126 152630 87130 152686
rect 87130 152630 87186 152686
rect 87186 152630 87190 152686
rect 87126 152626 87190 152630
rect 886 152142 950 152146
rect 886 152086 890 152142
rect 890 152086 946 152142
rect 946 152086 950 152142
rect 886 152082 950 152086
rect 966 152142 1030 152146
rect 966 152086 970 152142
rect 970 152086 1026 152142
rect 1026 152086 1030 152142
rect 966 152082 1030 152086
rect 1046 152142 1110 152146
rect 1046 152086 1050 152142
rect 1050 152086 1106 152142
rect 1106 152086 1110 152142
rect 1046 152082 1110 152086
rect 1126 152142 1190 152146
rect 1126 152086 1130 152142
rect 1130 152086 1186 152142
rect 1186 152086 1190 152142
rect 1126 152082 1190 152086
rect 84886 152142 84950 152146
rect 84886 152086 84890 152142
rect 84890 152086 84946 152142
rect 84946 152086 84950 152142
rect 84886 152082 84950 152086
rect 84966 152142 85030 152146
rect 84966 152086 84970 152142
rect 84970 152086 85026 152142
rect 85026 152086 85030 152142
rect 84966 152082 85030 152086
rect 85046 152142 85110 152146
rect 85046 152086 85050 152142
rect 85050 152086 85106 152142
rect 85106 152086 85110 152142
rect 85046 152082 85110 152086
rect 85126 152142 85190 152146
rect 85126 152086 85130 152142
rect 85130 152086 85186 152142
rect 85186 152086 85190 152142
rect 85126 152082 85190 152086
rect 5618 151802 5682 151806
rect 5618 151746 5632 151802
rect 5632 151746 5682 151802
rect 5618 151742 5682 151746
rect 82346 151742 82410 151806
rect 2886 151598 2950 151602
rect 2886 151542 2890 151598
rect 2890 151542 2946 151598
rect 2946 151542 2950 151598
rect 2886 151538 2950 151542
rect 2966 151598 3030 151602
rect 2966 151542 2970 151598
rect 2970 151542 3026 151598
rect 3026 151542 3030 151598
rect 2966 151538 3030 151542
rect 3046 151598 3110 151602
rect 3046 151542 3050 151598
rect 3050 151542 3106 151598
rect 3106 151542 3110 151598
rect 3046 151538 3110 151542
rect 3126 151598 3190 151602
rect 3126 151542 3130 151598
rect 3130 151542 3186 151598
rect 3186 151542 3190 151598
rect 3126 151538 3190 151542
rect 86886 151598 86950 151602
rect 86886 151542 86890 151598
rect 86890 151542 86946 151598
rect 86946 151542 86950 151598
rect 86886 151538 86950 151542
rect 86966 151598 87030 151602
rect 86966 151542 86970 151598
rect 86970 151542 87026 151598
rect 87026 151542 87030 151598
rect 86966 151538 87030 151542
rect 87046 151598 87110 151602
rect 87046 151542 87050 151598
rect 87050 151542 87106 151598
rect 87106 151542 87110 151598
rect 87046 151538 87110 151542
rect 87126 151598 87190 151602
rect 87126 151542 87130 151598
rect 87130 151542 87186 151598
rect 87186 151542 87190 151598
rect 87126 151538 87190 151542
rect 886 151054 950 151058
rect 886 150998 890 151054
rect 890 150998 946 151054
rect 946 150998 950 151054
rect 886 150994 950 150998
rect 966 151054 1030 151058
rect 966 150998 970 151054
rect 970 150998 1026 151054
rect 1026 150998 1030 151054
rect 966 150994 1030 150998
rect 1046 151054 1110 151058
rect 1046 150998 1050 151054
rect 1050 150998 1106 151054
rect 1106 150998 1110 151054
rect 1046 150994 1110 150998
rect 1126 151054 1190 151058
rect 1126 150998 1130 151054
rect 1130 150998 1186 151054
rect 1186 150998 1190 151054
rect 1126 150994 1190 150998
rect 84886 151054 84950 151058
rect 84886 150998 84890 151054
rect 84890 150998 84946 151054
rect 84946 150998 84950 151054
rect 84886 150994 84950 150998
rect 84966 151054 85030 151058
rect 84966 150998 84970 151054
rect 84970 150998 85026 151054
rect 85026 150998 85030 151054
rect 84966 150994 85030 150998
rect 85046 151054 85110 151058
rect 85046 150998 85050 151054
rect 85050 150998 85106 151054
rect 85106 150998 85110 151054
rect 85046 150994 85110 150998
rect 85126 151054 85190 151058
rect 85126 150998 85130 151054
rect 85130 150998 85186 151054
rect 85186 150998 85190 151054
rect 85126 150994 85190 150998
rect 2886 150510 2950 150514
rect 2886 150454 2890 150510
rect 2890 150454 2946 150510
rect 2946 150454 2950 150510
rect 2886 150450 2950 150454
rect 2966 150510 3030 150514
rect 2966 150454 2970 150510
rect 2970 150454 3026 150510
rect 3026 150454 3030 150510
rect 2966 150450 3030 150454
rect 3046 150510 3110 150514
rect 3046 150454 3050 150510
rect 3050 150454 3106 150510
rect 3106 150454 3110 150510
rect 3046 150450 3110 150454
rect 3126 150510 3190 150514
rect 3126 150454 3130 150510
rect 3130 150454 3186 150510
rect 3186 150454 3190 150510
rect 3126 150450 3190 150454
rect 86886 150510 86950 150514
rect 86886 150454 86890 150510
rect 86890 150454 86946 150510
rect 86946 150454 86950 150510
rect 86886 150450 86950 150454
rect 86966 150510 87030 150514
rect 86966 150454 86970 150510
rect 86970 150454 87026 150510
rect 87026 150454 87030 150510
rect 86966 150450 87030 150454
rect 87046 150510 87110 150514
rect 87046 150454 87050 150510
rect 87050 150454 87106 150510
rect 87106 150454 87110 150510
rect 87046 150450 87110 150454
rect 87126 150510 87190 150514
rect 87126 150454 87130 150510
rect 87130 150454 87186 150510
rect 87186 150454 87190 150510
rect 87126 150450 87190 150454
rect 886 149966 950 149970
rect 886 149910 890 149966
rect 890 149910 946 149966
rect 946 149910 950 149966
rect 886 149906 950 149910
rect 966 149966 1030 149970
rect 966 149910 970 149966
rect 970 149910 1026 149966
rect 1026 149910 1030 149966
rect 966 149906 1030 149910
rect 1046 149966 1110 149970
rect 1046 149910 1050 149966
rect 1050 149910 1106 149966
rect 1106 149910 1110 149966
rect 1046 149906 1110 149910
rect 1126 149966 1190 149970
rect 1126 149910 1130 149966
rect 1130 149910 1186 149966
rect 1186 149910 1190 149966
rect 1126 149906 1190 149910
rect 84886 149966 84950 149970
rect 84886 149910 84890 149966
rect 84890 149910 84946 149966
rect 84946 149910 84950 149966
rect 84886 149906 84950 149910
rect 84966 149966 85030 149970
rect 84966 149910 84970 149966
rect 84970 149910 85026 149966
rect 85026 149910 85030 149966
rect 84966 149906 85030 149910
rect 85046 149966 85110 149970
rect 85046 149910 85050 149966
rect 85050 149910 85106 149966
rect 85106 149910 85110 149966
rect 85046 149906 85110 149910
rect 85126 149966 85190 149970
rect 85126 149910 85130 149966
rect 85130 149910 85186 149966
rect 85186 149910 85190 149966
rect 85126 149906 85190 149910
rect 2886 149422 2950 149426
rect 2886 149366 2890 149422
rect 2890 149366 2946 149422
rect 2946 149366 2950 149422
rect 2886 149362 2950 149366
rect 2966 149422 3030 149426
rect 2966 149366 2970 149422
rect 2970 149366 3026 149422
rect 3026 149366 3030 149422
rect 2966 149362 3030 149366
rect 3046 149422 3110 149426
rect 3046 149366 3050 149422
rect 3050 149366 3106 149422
rect 3106 149366 3110 149422
rect 3046 149362 3110 149366
rect 3126 149422 3190 149426
rect 3126 149366 3130 149422
rect 3130 149366 3186 149422
rect 3186 149366 3190 149422
rect 3126 149362 3190 149366
rect 86886 149422 86950 149426
rect 86886 149366 86890 149422
rect 86890 149366 86946 149422
rect 86946 149366 86950 149422
rect 86886 149362 86950 149366
rect 86966 149422 87030 149426
rect 86966 149366 86970 149422
rect 86970 149366 87026 149422
rect 87026 149366 87030 149422
rect 86966 149362 87030 149366
rect 87046 149422 87110 149426
rect 87046 149366 87050 149422
rect 87050 149366 87106 149422
rect 87106 149366 87110 149422
rect 87046 149362 87110 149366
rect 87126 149422 87190 149426
rect 87126 149366 87130 149422
rect 87130 149366 87186 149422
rect 87186 149366 87190 149422
rect 87126 149362 87190 149366
rect 886 148878 950 148882
rect 886 148822 890 148878
rect 890 148822 946 148878
rect 946 148822 950 148878
rect 886 148818 950 148822
rect 966 148878 1030 148882
rect 966 148822 970 148878
rect 970 148822 1026 148878
rect 1026 148822 1030 148878
rect 966 148818 1030 148822
rect 1046 148878 1110 148882
rect 1046 148822 1050 148878
rect 1050 148822 1106 148878
rect 1106 148822 1110 148878
rect 1046 148818 1110 148822
rect 1126 148878 1190 148882
rect 1126 148822 1130 148878
rect 1130 148822 1186 148878
rect 1186 148822 1190 148878
rect 1126 148818 1190 148822
rect 84886 148878 84950 148882
rect 84886 148822 84890 148878
rect 84890 148822 84946 148878
rect 84946 148822 84950 148878
rect 84886 148818 84950 148822
rect 84966 148878 85030 148882
rect 84966 148822 84970 148878
rect 84970 148822 85026 148878
rect 85026 148822 85030 148878
rect 84966 148818 85030 148822
rect 85046 148878 85110 148882
rect 85046 148822 85050 148878
rect 85050 148822 85106 148878
rect 85106 148822 85110 148878
rect 85046 148818 85110 148822
rect 85126 148878 85190 148882
rect 85126 148822 85130 148878
rect 85130 148822 85186 148878
rect 85186 148822 85190 148878
rect 85126 148818 85190 148822
rect 2886 148334 2950 148338
rect 2886 148278 2890 148334
rect 2890 148278 2946 148334
rect 2946 148278 2950 148334
rect 2886 148274 2950 148278
rect 2966 148334 3030 148338
rect 2966 148278 2970 148334
rect 2970 148278 3026 148334
rect 3026 148278 3030 148334
rect 2966 148274 3030 148278
rect 3046 148334 3110 148338
rect 3046 148278 3050 148334
rect 3050 148278 3106 148334
rect 3106 148278 3110 148334
rect 3046 148274 3110 148278
rect 3126 148334 3190 148338
rect 3126 148278 3130 148334
rect 3130 148278 3186 148334
rect 3186 148278 3190 148334
rect 3126 148274 3190 148278
rect 86886 148334 86950 148338
rect 86886 148278 86890 148334
rect 86890 148278 86946 148334
rect 86946 148278 86950 148334
rect 86886 148274 86950 148278
rect 86966 148334 87030 148338
rect 86966 148278 86970 148334
rect 86970 148278 87026 148334
rect 87026 148278 87030 148334
rect 86966 148274 87030 148278
rect 87046 148334 87110 148338
rect 87046 148278 87050 148334
rect 87050 148278 87106 148334
rect 87106 148278 87110 148334
rect 87046 148274 87110 148278
rect 87126 148334 87190 148338
rect 87126 148278 87130 148334
rect 87130 148278 87186 148334
rect 87186 148278 87190 148334
rect 87126 148274 87190 148278
rect 886 147790 950 147794
rect 886 147734 890 147790
rect 890 147734 946 147790
rect 946 147734 950 147790
rect 886 147730 950 147734
rect 966 147790 1030 147794
rect 966 147734 970 147790
rect 970 147734 1026 147790
rect 1026 147734 1030 147790
rect 966 147730 1030 147734
rect 1046 147790 1110 147794
rect 1046 147734 1050 147790
rect 1050 147734 1106 147790
rect 1106 147734 1110 147790
rect 1046 147730 1110 147734
rect 1126 147790 1190 147794
rect 1126 147734 1130 147790
rect 1130 147734 1186 147790
rect 1186 147734 1190 147790
rect 1126 147730 1190 147734
rect 84886 147790 84950 147794
rect 84886 147734 84890 147790
rect 84890 147734 84946 147790
rect 84946 147734 84950 147790
rect 84886 147730 84950 147734
rect 84966 147790 85030 147794
rect 84966 147734 84970 147790
rect 84970 147734 85026 147790
rect 85026 147734 85030 147790
rect 84966 147730 85030 147734
rect 85046 147790 85110 147794
rect 85046 147734 85050 147790
rect 85050 147734 85106 147790
rect 85106 147734 85110 147790
rect 85046 147730 85110 147734
rect 85126 147790 85190 147794
rect 85126 147734 85130 147790
rect 85130 147734 85186 147790
rect 85186 147734 85190 147790
rect 85126 147730 85190 147734
rect 2886 147246 2950 147250
rect 2886 147190 2890 147246
rect 2890 147190 2946 147246
rect 2946 147190 2950 147246
rect 2886 147186 2950 147190
rect 2966 147246 3030 147250
rect 2966 147190 2970 147246
rect 2970 147190 3026 147246
rect 3026 147190 3030 147246
rect 2966 147186 3030 147190
rect 3046 147246 3110 147250
rect 3046 147190 3050 147246
rect 3050 147190 3106 147246
rect 3106 147190 3110 147246
rect 3046 147186 3110 147190
rect 3126 147246 3190 147250
rect 3126 147190 3130 147246
rect 3130 147190 3186 147246
rect 3186 147190 3190 147246
rect 3126 147186 3190 147190
rect 86886 147246 86950 147250
rect 86886 147190 86890 147246
rect 86890 147190 86946 147246
rect 86946 147190 86950 147246
rect 86886 147186 86950 147190
rect 86966 147246 87030 147250
rect 86966 147190 86970 147246
rect 86970 147190 87026 147246
rect 87026 147190 87030 147246
rect 86966 147186 87030 147190
rect 87046 147246 87110 147250
rect 87046 147190 87050 147246
rect 87050 147190 87106 147246
rect 87106 147190 87110 147246
rect 87046 147186 87110 147190
rect 87126 147246 87190 147250
rect 87126 147190 87130 147246
rect 87130 147190 87186 147246
rect 87186 147190 87190 147246
rect 87126 147186 87190 147190
rect 886 146702 950 146706
rect 886 146646 890 146702
rect 890 146646 946 146702
rect 946 146646 950 146702
rect 886 146642 950 146646
rect 966 146702 1030 146706
rect 966 146646 970 146702
rect 970 146646 1026 146702
rect 1026 146646 1030 146702
rect 966 146642 1030 146646
rect 1046 146702 1110 146706
rect 1046 146646 1050 146702
rect 1050 146646 1106 146702
rect 1106 146646 1110 146702
rect 1046 146642 1110 146646
rect 1126 146702 1190 146706
rect 1126 146646 1130 146702
rect 1130 146646 1186 146702
rect 1186 146646 1190 146702
rect 1126 146642 1190 146646
rect 84886 146702 84950 146706
rect 84886 146646 84890 146702
rect 84890 146646 84946 146702
rect 84946 146646 84950 146702
rect 84886 146642 84950 146646
rect 84966 146702 85030 146706
rect 84966 146646 84970 146702
rect 84970 146646 85026 146702
rect 85026 146646 85030 146702
rect 84966 146642 85030 146646
rect 85046 146702 85110 146706
rect 85046 146646 85050 146702
rect 85050 146646 85106 146702
rect 85106 146646 85110 146702
rect 85046 146642 85110 146646
rect 85126 146702 85190 146706
rect 85126 146646 85130 146702
rect 85130 146646 85186 146702
rect 85186 146646 85190 146702
rect 85126 146642 85190 146646
rect 2886 146158 2950 146162
rect 2886 146102 2890 146158
rect 2890 146102 2946 146158
rect 2946 146102 2950 146158
rect 2886 146098 2950 146102
rect 2966 146158 3030 146162
rect 2966 146102 2970 146158
rect 2970 146102 3026 146158
rect 3026 146102 3030 146158
rect 2966 146098 3030 146102
rect 3046 146158 3110 146162
rect 3046 146102 3050 146158
rect 3050 146102 3106 146158
rect 3106 146102 3110 146158
rect 3046 146098 3110 146102
rect 3126 146158 3190 146162
rect 3126 146102 3130 146158
rect 3130 146102 3186 146158
rect 3186 146102 3190 146158
rect 3126 146098 3190 146102
rect 86886 146158 86950 146162
rect 86886 146102 86890 146158
rect 86890 146102 86946 146158
rect 86946 146102 86950 146158
rect 86886 146098 86950 146102
rect 86966 146158 87030 146162
rect 86966 146102 86970 146158
rect 86970 146102 87026 146158
rect 87026 146102 87030 146158
rect 86966 146098 87030 146102
rect 87046 146158 87110 146162
rect 87046 146102 87050 146158
rect 87050 146102 87106 146158
rect 87106 146102 87110 146158
rect 87046 146098 87110 146102
rect 87126 146158 87190 146162
rect 87126 146102 87130 146158
rect 87130 146102 87186 146158
rect 87186 146102 87190 146158
rect 87126 146098 87190 146102
rect 886 145614 950 145618
rect 886 145558 890 145614
rect 890 145558 946 145614
rect 946 145558 950 145614
rect 886 145554 950 145558
rect 966 145614 1030 145618
rect 966 145558 970 145614
rect 970 145558 1026 145614
rect 1026 145558 1030 145614
rect 966 145554 1030 145558
rect 1046 145614 1110 145618
rect 1046 145558 1050 145614
rect 1050 145558 1106 145614
rect 1106 145558 1110 145614
rect 1046 145554 1110 145558
rect 1126 145614 1190 145618
rect 1126 145558 1130 145614
rect 1130 145558 1186 145614
rect 1186 145558 1190 145614
rect 1126 145554 1190 145558
rect 84886 145614 84950 145618
rect 84886 145558 84890 145614
rect 84890 145558 84946 145614
rect 84946 145558 84950 145614
rect 84886 145554 84950 145558
rect 84966 145614 85030 145618
rect 84966 145558 84970 145614
rect 84970 145558 85026 145614
rect 85026 145558 85030 145614
rect 84966 145554 85030 145558
rect 85046 145614 85110 145618
rect 85046 145558 85050 145614
rect 85050 145558 85106 145614
rect 85106 145558 85110 145614
rect 85046 145554 85110 145558
rect 85126 145614 85190 145618
rect 85126 145558 85130 145614
rect 85130 145558 85186 145614
rect 85186 145558 85190 145614
rect 85126 145554 85190 145558
rect 2886 145070 2950 145074
rect 2886 145014 2890 145070
rect 2890 145014 2946 145070
rect 2946 145014 2950 145070
rect 2886 145010 2950 145014
rect 2966 145070 3030 145074
rect 2966 145014 2970 145070
rect 2970 145014 3026 145070
rect 3026 145014 3030 145070
rect 2966 145010 3030 145014
rect 3046 145070 3110 145074
rect 3046 145014 3050 145070
rect 3050 145014 3106 145070
rect 3106 145014 3110 145070
rect 3046 145010 3110 145014
rect 3126 145070 3190 145074
rect 3126 145014 3130 145070
rect 3130 145014 3186 145070
rect 3186 145014 3190 145070
rect 3126 145010 3190 145014
rect 86886 145070 86950 145074
rect 86886 145014 86890 145070
rect 86890 145014 86946 145070
rect 86946 145014 86950 145070
rect 86886 145010 86950 145014
rect 86966 145070 87030 145074
rect 86966 145014 86970 145070
rect 86970 145014 87026 145070
rect 87026 145014 87030 145070
rect 86966 145010 87030 145014
rect 87046 145070 87110 145074
rect 87046 145014 87050 145070
rect 87050 145014 87106 145070
rect 87106 145014 87110 145070
rect 87046 145010 87110 145014
rect 87126 145070 87190 145074
rect 87126 145014 87130 145070
rect 87130 145014 87186 145070
rect 87186 145014 87190 145070
rect 87126 145010 87190 145014
rect 886 144526 950 144530
rect 886 144470 890 144526
rect 890 144470 946 144526
rect 946 144470 950 144526
rect 886 144466 950 144470
rect 966 144526 1030 144530
rect 966 144470 970 144526
rect 970 144470 1026 144526
rect 1026 144470 1030 144526
rect 966 144466 1030 144470
rect 1046 144526 1110 144530
rect 1046 144470 1050 144526
rect 1050 144470 1106 144526
rect 1106 144470 1110 144526
rect 1046 144466 1110 144470
rect 1126 144526 1190 144530
rect 1126 144470 1130 144526
rect 1130 144470 1186 144526
rect 1186 144470 1190 144526
rect 1126 144466 1190 144470
rect 84886 144526 84950 144530
rect 84886 144470 84890 144526
rect 84890 144470 84946 144526
rect 84946 144470 84950 144526
rect 84886 144466 84950 144470
rect 84966 144526 85030 144530
rect 84966 144470 84970 144526
rect 84970 144470 85026 144526
rect 85026 144470 85030 144526
rect 84966 144466 85030 144470
rect 85046 144526 85110 144530
rect 85046 144470 85050 144526
rect 85050 144470 85106 144526
rect 85106 144470 85110 144526
rect 85046 144466 85110 144470
rect 85126 144526 85190 144530
rect 85126 144470 85130 144526
rect 85130 144470 85186 144526
rect 85186 144470 85190 144526
rect 85126 144466 85190 144470
rect 2886 143982 2950 143986
rect 2886 143926 2890 143982
rect 2890 143926 2946 143982
rect 2946 143926 2950 143982
rect 2886 143922 2950 143926
rect 2966 143982 3030 143986
rect 2966 143926 2970 143982
rect 2970 143926 3026 143982
rect 3026 143926 3030 143982
rect 2966 143922 3030 143926
rect 3046 143982 3110 143986
rect 3046 143926 3050 143982
rect 3050 143926 3106 143982
rect 3106 143926 3110 143982
rect 3046 143922 3110 143926
rect 3126 143982 3190 143986
rect 3126 143926 3130 143982
rect 3130 143926 3186 143982
rect 3186 143926 3190 143982
rect 3126 143922 3190 143926
rect 86886 143982 86950 143986
rect 86886 143926 86890 143982
rect 86890 143926 86946 143982
rect 86946 143926 86950 143982
rect 86886 143922 86950 143926
rect 86966 143982 87030 143986
rect 86966 143926 86970 143982
rect 86970 143926 87026 143982
rect 87026 143926 87030 143982
rect 86966 143922 87030 143926
rect 87046 143982 87110 143986
rect 87046 143926 87050 143982
rect 87050 143926 87106 143982
rect 87106 143926 87110 143982
rect 87046 143922 87110 143926
rect 87126 143982 87190 143986
rect 87126 143926 87130 143982
rect 87130 143926 87186 143982
rect 87186 143926 87190 143982
rect 87126 143922 87190 143926
rect 886 143438 950 143442
rect 886 143382 890 143438
rect 890 143382 946 143438
rect 946 143382 950 143438
rect 886 143378 950 143382
rect 966 143438 1030 143442
rect 966 143382 970 143438
rect 970 143382 1026 143438
rect 1026 143382 1030 143438
rect 966 143378 1030 143382
rect 1046 143438 1110 143442
rect 1046 143382 1050 143438
rect 1050 143382 1106 143438
rect 1106 143382 1110 143438
rect 1046 143378 1110 143382
rect 1126 143438 1190 143442
rect 1126 143382 1130 143438
rect 1130 143382 1186 143438
rect 1186 143382 1190 143438
rect 1126 143378 1190 143382
rect 84886 143438 84950 143442
rect 84886 143382 84890 143438
rect 84890 143382 84946 143438
rect 84946 143382 84950 143438
rect 84886 143378 84950 143382
rect 84966 143438 85030 143442
rect 84966 143382 84970 143438
rect 84970 143382 85026 143438
rect 85026 143382 85030 143438
rect 84966 143378 85030 143382
rect 85046 143438 85110 143442
rect 85046 143382 85050 143438
rect 85050 143382 85106 143438
rect 85106 143382 85110 143438
rect 85046 143378 85110 143382
rect 85126 143438 85190 143442
rect 85126 143382 85130 143438
rect 85130 143382 85186 143438
rect 85186 143382 85190 143438
rect 85126 143378 85190 143382
rect 2886 142894 2950 142898
rect 2886 142838 2890 142894
rect 2890 142838 2946 142894
rect 2946 142838 2950 142894
rect 2886 142834 2950 142838
rect 2966 142894 3030 142898
rect 2966 142838 2970 142894
rect 2970 142838 3026 142894
rect 3026 142838 3030 142894
rect 2966 142834 3030 142838
rect 3046 142894 3110 142898
rect 3046 142838 3050 142894
rect 3050 142838 3106 142894
rect 3106 142838 3110 142894
rect 3046 142834 3110 142838
rect 3126 142894 3190 142898
rect 3126 142838 3130 142894
rect 3130 142838 3186 142894
rect 3186 142838 3190 142894
rect 3126 142834 3190 142838
rect 86886 142894 86950 142898
rect 86886 142838 86890 142894
rect 86890 142838 86946 142894
rect 86946 142838 86950 142894
rect 86886 142834 86950 142838
rect 86966 142894 87030 142898
rect 86966 142838 86970 142894
rect 86970 142838 87026 142894
rect 87026 142838 87030 142894
rect 86966 142834 87030 142838
rect 87046 142894 87110 142898
rect 87046 142838 87050 142894
rect 87050 142838 87106 142894
rect 87106 142838 87110 142894
rect 87046 142834 87110 142838
rect 87126 142894 87190 142898
rect 87126 142838 87130 142894
rect 87130 142838 87186 142894
rect 87186 142838 87190 142894
rect 87126 142834 87190 142838
rect 886 142350 950 142354
rect 886 142294 890 142350
rect 890 142294 946 142350
rect 946 142294 950 142350
rect 886 142290 950 142294
rect 966 142350 1030 142354
rect 966 142294 970 142350
rect 970 142294 1026 142350
rect 1026 142294 1030 142350
rect 966 142290 1030 142294
rect 1046 142350 1110 142354
rect 1046 142294 1050 142350
rect 1050 142294 1106 142350
rect 1106 142294 1110 142350
rect 1046 142290 1110 142294
rect 1126 142350 1190 142354
rect 1126 142294 1130 142350
rect 1130 142294 1186 142350
rect 1186 142294 1190 142350
rect 1126 142290 1190 142294
rect 84886 142350 84950 142354
rect 84886 142294 84890 142350
rect 84890 142294 84946 142350
rect 84946 142294 84950 142350
rect 84886 142290 84950 142294
rect 84966 142350 85030 142354
rect 84966 142294 84970 142350
rect 84970 142294 85026 142350
rect 85026 142294 85030 142350
rect 84966 142290 85030 142294
rect 85046 142350 85110 142354
rect 85046 142294 85050 142350
rect 85050 142294 85106 142350
rect 85106 142294 85110 142350
rect 85046 142290 85110 142294
rect 85126 142350 85190 142354
rect 85126 142294 85130 142350
rect 85130 142294 85186 142350
rect 85186 142294 85190 142350
rect 85126 142290 85190 142294
rect 2886 141806 2950 141810
rect 2886 141750 2890 141806
rect 2890 141750 2946 141806
rect 2946 141750 2950 141806
rect 2886 141746 2950 141750
rect 2966 141806 3030 141810
rect 2966 141750 2970 141806
rect 2970 141750 3026 141806
rect 3026 141750 3030 141806
rect 2966 141746 3030 141750
rect 3046 141806 3110 141810
rect 3046 141750 3050 141806
rect 3050 141750 3106 141806
rect 3106 141750 3110 141806
rect 3046 141746 3110 141750
rect 3126 141806 3190 141810
rect 3126 141750 3130 141806
rect 3130 141750 3186 141806
rect 3186 141750 3190 141806
rect 3126 141746 3190 141750
rect 86886 141806 86950 141810
rect 86886 141750 86890 141806
rect 86890 141750 86946 141806
rect 86946 141750 86950 141806
rect 86886 141746 86950 141750
rect 86966 141806 87030 141810
rect 86966 141750 86970 141806
rect 86970 141750 87026 141806
rect 87026 141750 87030 141806
rect 86966 141746 87030 141750
rect 87046 141806 87110 141810
rect 87046 141750 87050 141806
rect 87050 141750 87106 141806
rect 87106 141750 87110 141806
rect 87046 141746 87110 141750
rect 87126 141806 87190 141810
rect 87126 141750 87130 141806
rect 87130 141750 87186 141806
rect 87186 141750 87190 141806
rect 87126 141746 87190 141750
rect 886 141262 950 141266
rect 886 141206 890 141262
rect 890 141206 946 141262
rect 946 141206 950 141262
rect 886 141202 950 141206
rect 966 141262 1030 141266
rect 966 141206 970 141262
rect 970 141206 1026 141262
rect 1026 141206 1030 141262
rect 966 141202 1030 141206
rect 1046 141262 1110 141266
rect 1046 141206 1050 141262
rect 1050 141206 1106 141262
rect 1106 141206 1110 141262
rect 1046 141202 1110 141206
rect 1126 141262 1190 141266
rect 1126 141206 1130 141262
rect 1130 141206 1186 141262
rect 1186 141206 1190 141262
rect 1126 141202 1190 141206
rect 84886 141262 84950 141266
rect 84886 141206 84890 141262
rect 84890 141206 84946 141262
rect 84946 141206 84950 141262
rect 84886 141202 84950 141206
rect 84966 141262 85030 141266
rect 84966 141206 84970 141262
rect 84970 141206 85026 141262
rect 85026 141206 85030 141262
rect 84966 141202 85030 141206
rect 85046 141262 85110 141266
rect 85046 141206 85050 141262
rect 85050 141206 85106 141262
rect 85106 141206 85110 141262
rect 85046 141202 85110 141206
rect 85126 141262 85190 141266
rect 85126 141206 85130 141262
rect 85130 141206 85186 141262
rect 85186 141206 85190 141262
rect 85126 141202 85190 141206
rect 82346 140998 82410 141062
rect 2886 140718 2950 140722
rect 2886 140662 2890 140718
rect 2890 140662 2946 140718
rect 2946 140662 2950 140718
rect 2886 140658 2950 140662
rect 2966 140718 3030 140722
rect 2966 140662 2970 140718
rect 2970 140662 3026 140718
rect 3026 140662 3030 140718
rect 2966 140658 3030 140662
rect 3046 140718 3110 140722
rect 3046 140662 3050 140718
rect 3050 140662 3106 140718
rect 3106 140662 3110 140718
rect 3046 140658 3110 140662
rect 3126 140718 3190 140722
rect 3126 140662 3130 140718
rect 3130 140662 3186 140718
rect 3186 140662 3190 140718
rect 3126 140658 3190 140662
rect 86886 140718 86950 140722
rect 86886 140662 86890 140718
rect 86890 140662 86946 140718
rect 86946 140662 86950 140718
rect 86886 140658 86950 140662
rect 86966 140718 87030 140722
rect 86966 140662 86970 140718
rect 86970 140662 87026 140718
rect 87026 140662 87030 140718
rect 86966 140658 87030 140662
rect 87046 140718 87110 140722
rect 87046 140662 87050 140718
rect 87050 140662 87106 140718
rect 87106 140662 87110 140718
rect 87046 140658 87110 140662
rect 87126 140718 87190 140722
rect 87126 140662 87130 140718
rect 87130 140662 87186 140718
rect 87186 140662 87190 140718
rect 87126 140658 87190 140662
rect 886 140174 950 140178
rect 886 140118 890 140174
rect 890 140118 946 140174
rect 946 140118 950 140174
rect 886 140114 950 140118
rect 966 140174 1030 140178
rect 966 140118 970 140174
rect 970 140118 1026 140174
rect 1026 140118 1030 140174
rect 966 140114 1030 140118
rect 1046 140174 1110 140178
rect 1046 140118 1050 140174
rect 1050 140118 1106 140174
rect 1106 140118 1110 140174
rect 1046 140114 1110 140118
rect 1126 140174 1190 140178
rect 1126 140118 1130 140174
rect 1130 140118 1186 140174
rect 1186 140118 1190 140174
rect 1126 140114 1190 140118
rect 84886 140174 84950 140178
rect 84886 140118 84890 140174
rect 84890 140118 84946 140174
rect 84946 140118 84950 140174
rect 84886 140114 84950 140118
rect 84966 140174 85030 140178
rect 84966 140118 84970 140174
rect 84970 140118 85026 140174
rect 85026 140118 85030 140174
rect 84966 140114 85030 140118
rect 85046 140174 85110 140178
rect 85046 140118 85050 140174
rect 85050 140118 85106 140174
rect 85106 140118 85110 140174
rect 85046 140114 85110 140118
rect 85126 140174 85190 140178
rect 85126 140118 85130 140174
rect 85130 140118 85186 140174
rect 85186 140118 85190 140174
rect 85126 140114 85190 140118
rect 2886 139630 2950 139634
rect 2886 139574 2890 139630
rect 2890 139574 2946 139630
rect 2946 139574 2950 139630
rect 2886 139570 2950 139574
rect 2966 139630 3030 139634
rect 2966 139574 2970 139630
rect 2970 139574 3026 139630
rect 3026 139574 3030 139630
rect 2966 139570 3030 139574
rect 3046 139630 3110 139634
rect 3046 139574 3050 139630
rect 3050 139574 3106 139630
rect 3106 139574 3110 139630
rect 3046 139570 3110 139574
rect 3126 139630 3190 139634
rect 3126 139574 3130 139630
rect 3130 139574 3186 139630
rect 3186 139574 3190 139630
rect 3126 139570 3190 139574
rect 86886 139630 86950 139634
rect 86886 139574 86890 139630
rect 86890 139574 86946 139630
rect 86946 139574 86950 139630
rect 86886 139570 86950 139574
rect 86966 139630 87030 139634
rect 86966 139574 86970 139630
rect 86970 139574 87026 139630
rect 87026 139574 87030 139630
rect 86966 139570 87030 139574
rect 87046 139630 87110 139634
rect 87046 139574 87050 139630
rect 87050 139574 87106 139630
rect 87106 139574 87110 139630
rect 87046 139570 87110 139574
rect 87126 139630 87190 139634
rect 87126 139574 87130 139630
rect 87130 139574 87186 139630
rect 87186 139574 87190 139630
rect 87126 139570 87190 139574
rect 886 139086 950 139090
rect 886 139030 890 139086
rect 890 139030 946 139086
rect 946 139030 950 139086
rect 886 139026 950 139030
rect 966 139086 1030 139090
rect 966 139030 970 139086
rect 970 139030 1026 139086
rect 1026 139030 1030 139086
rect 966 139026 1030 139030
rect 1046 139086 1110 139090
rect 1046 139030 1050 139086
rect 1050 139030 1106 139086
rect 1106 139030 1110 139086
rect 1046 139026 1110 139030
rect 1126 139086 1190 139090
rect 1126 139030 1130 139086
rect 1130 139030 1186 139086
rect 1186 139030 1190 139086
rect 1126 139026 1190 139030
rect 84886 139086 84950 139090
rect 84886 139030 84890 139086
rect 84890 139030 84946 139086
rect 84946 139030 84950 139086
rect 84886 139026 84950 139030
rect 84966 139086 85030 139090
rect 84966 139030 84970 139086
rect 84970 139030 85026 139086
rect 85026 139030 85030 139086
rect 84966 139026 85030 139030
rect 85046 139086 85110 139090
rect 85046 139030 85050 139086
rect 85050 139030 85106 139086
rect 85106 139030 85110 139086
rect 85046 139026 85110 139030
rect 85126 139086 85190 139090
rect 85126 139030 85130 139086
rect 85130 139030 85186 139086
rect 85186 139030 85190 139086
rect 85126 139026 85190 139030
rect 2886 138542 2950 138546
rect 2886 138486 2890 138542
rect 2890 138486 2946 138542
rect 2946 138486 2950 138542
rect 2886 138482 2950 138486
rect 2966 138542 3030 138546
rect 2966 138486 2970 138542
rect 2970 138486 3026 138542
rect 3026 138486 3030 138542
rect 2966 138482 3030 138486
rect 3046 138542 3110 138546
rect 3046 138486 3050 138542
rect 3050 138486 3106 138542
rect 3106 138486 3110 138542
rect 3046 138482 3110 138486
rect 3126 138542 3190 138546
rect 3126 138486 3130 138542
rect 3130 138486 3186 138542
rect 3186 138486 3190 138542
rect 3126 138482 3190 138486
rect 86886 138542 86950 138546
rect 86886 138486 86890 138542
rect 86890 138486 86946 138542
rect 86946 138486 86950 138542
rect 86886 138482 86950 138486
rect 86966 138542 87030 138546
rect 86966 138486 86970 138542
rect 86970 138486 87026 138542
rect 87026 138486 87030 138542
rect 86966 138482 87030 138486
rect 87046 138542 87110 138546
rect 87046 138486 87050 138542
rect 87050 138486 87106 138542
rect 87106 138486 87110 138542
rect 87046 138482 87110 138486
rect 87126 138542 87190 138546
rect 87126 138486 87130 138542
rect 87130 138486 87186 138542
rect 87186 138486 87190 138542
rect 87126 138482 87190 138486
rect 886 137998 950 138002
rect 886 137942 890 137998
rect 890 137942 946 137998
rect 946 137942 950 137998
rect 886 137938 950 137942
rect 966 137998 1030 138002
rect 966 137942 970 137998
rect 970 137942 1026 137998
rect 1026 137942 1030 137998
rect 966 137938 1030 137942
rect 1046 137998 1110 138002
rect 1046 137942 1050 137998
rect 1050 137942 1106 137998
rect 1106 137942 1110 137998
rect 1046 137938 1110 137942
rect 1126 137998 1190 138002
rect 1126 137942 1130 137998
rect 1130 137942 1186 137998
rect 1186 137942 1190 137998
rect 1126 137938 1190 137942
rect 84886 137998 84950 138002
rect 84886 137942 84890 137998
rect 84890 137942 84946 137998
rect 84946 137942 84950 137998
rect 84886 137938 84950 137942
rect 84966 137998 85030 138002
rect 84966 137942 84970 137998
rect 84970 137942 85026 137998
rect 85026 137942 85030 137998
rect 84966 137938 85030 137942
rect 85046 137998 85110 138002
rect 85046 137942 85050 137998
rect 85050 137942 85106 137998
rect 85106 137942 85110 137998
rect 85046 137938 85110 137942
rect 85126 137998 85190 138002
rect 85126 137942 85130 137998
rect 85130 137942 85186 137998
rect 85186 137942 85190 137998
rect 85126 137938 85190 137942
rect 2886 137454 2950 137458
rect 2886 137398 2890 137454
rect 2890 137398 2946 137454
rect 2946 137398 2950 137454
rect 2886 137394 2950 137398
rect 2966 137454 3030 137458
rect 2966 137398 2970 137454
rect 2970 137398 3026 137454
rect 3026 137398 3030 137454
rect 2966 137394 3030 137398
rect 3046 137454 3110 137458
rect 3046 137398 3050 137454
rect 3050 137398 3106 137454
rect 3106 137398 3110 137454
rect 3046 137394 3110 137398
rect 3126 137454 3190 137458
rect 3126 137398 3130 137454
rect 3130 137398 3186 137454
rect 3186 137398 3190 137454
rect 3126 137394 3190 137398
rect 86886 137454 86950 137458
rect 86886 137398 86890 137454
rect 86890 137398 86946 137454
rect 86946 137398 86950 137454
rect 86886 137394 86950 137398
rect 86966 137454 87030 137458
rect 86966 137398 86970 137454
rect 86970 137398 87026 137454
rect 87026 137398 87030 137454
rect 86966 137394 87030 137398
rect 87046 137454 87110 137458
rect 87046 137398 87050 137454
rect 87050 137398 87106 137454
rect 87106 137398 87110 137454
rect 87046 137394 87110 137398
rect 87126 137454 87190 137458
rect 87126 137398 87130 137454
rect 87130 137398 87186 137454
rect 87186 137398 87190 137454
rect 87126 137394 87190 137398
rect 886 136910 950 136914
rect 886 136854 890 136910
rect 890 136854 946 136910
rect 946 136854 950 136910
rect 886 136850 950 136854
rect 966 136910 1030 136914
rect 966 136854 970 136910
rect 970 136854 1026 136910
rect 1026 136854 1030 136910
rect 966 136850 1030 136854
rect 1046 136910 1110 136914
rect 1046 136854 1050 136910
rect 1050 136854 1106 136910
rect 1106 136854 1110 136910
rect 1046 136850 1110 136854
rect 1126 136910 1190 136914
rect 1126 136854 1130 136910
rect 1130 136854 1186 136910
rect 1186 136854 1190 136910
rect 1126 136850 1190 136854
rect 84886 136910 84950 136914
rect 84886 136854 84890 136910
rect 84890 136854 84946 136910
rect 84946 136854 84950 136910
rect 84886 136850 84950 136854
rect 84966 136910 85030 136914
rect 84966 136854 84970 136910
rect 84970 136854 85026 136910
rect 85026 136854 85030 136910
rect 84966 136850 85030 136854
rect 85046 136910 85110 136914
rect 85046 136854 85050 136910
rect 85050 136854 85106 136910
rect 85106 136854 85110 136910
rect 85046 136850 85110 136854
rect 85126 136910 85190 136914
rect 85126 136854 85130 136910
rect 85130 136854 85186 136910
rect 85186 136854 85190 136910
rect 85126 136850 85190 136854
rect 2886 136366 2950 136370
rect 2886 136310 2890 136366
rect 2890 136310 2946 136366
rect 2946 136310 2950 136366
rect 2886 136306 2950 136310
rect 2966 136366 3030 136370
rect 2966 136310 2970 136366
rect 2970 136310 3026 136366
rect 3026 136310 3030 136366
rect 2966 136306 3030 136310
rect 3046 136366 3110 136370
rect 3046 136310 3050 136366
rect 3050 136310 3106 136366
rect 3106 136310 3110 136366
rect 3046 136306 3110 136310
rect 3126 136366 3190 136370
rect 3126 136310 3130 136366
rect 3130 136310 3186 136366
rect 3186 136310 3190 136366
rect 3126 136306 3190 136310
rect 86886 136366 86950 136370
rect 86886 136310 86890 136366
rect 86890 136310 86946 136366
rect 86946 136310 86950 136366
rect 86886 136306 86950 136310
rect 86966 136366 87030 136370
rect 86966 136310 86970 136366
rect 86970 136310 87026 136366
rect 87026 136310 87030 136366
rect 86966 136306 87030 136310
rect 87046 136366 87110 136370
rect 87046 136310 87050 136366
rect 87050 136310 87106 136366
rect 87106 136310 87110 136366
rect 87046 136306 87110 136310
rect 87126 136366 87190 136370
rect 87126 136310 87130 136366
rect 87130 136310 87186 136366
rect 87186 136310 87190 136366
rect 87126 136306 87190 136310
rect 886 135822 950 135826
rect 886 135766 890 135822
rect 890 135766 946 135822
rect 946 135766 950 135822
rect 886 135762 950 135766
rect 966 135822 1030 135826
rect 966 135766 970 135822
rect 970 135766 1026 135822
rect 1026 135766 1030 135822
rect 966 135762 1030 135766
rect 1046 135822 1110 135826
rect 1046 135766 1050 135822
rect 1050 135766 1106 135822
rect 1106 135766 1110 135822
rect 1046 135762 1110 135766
rect 1126 135822 1190 135826
rect 1126 135766 1130 135822
rect 1130 135766 1186 135822
rect 1186 135766 1190 135822
rect 1126 135762 1190 135766
rect 84886 135822 84950 135826
rect 84886 135766 84890 135822
rect 84890 135766 84946 135822
rect 84946 135766 84950 135822
rect 84886 135762 84950 135766
rect 84966 135822 85030 135826
rect 84966 135766 84970 135822
rect 84970 135766 85026 135822
rect 85026 135766 85030 135822
rect 84966 135762 85030 135766
rect 85046 135822 85110 135826
rect 85046 135766 85050 135822
rect 85050 135766 85106 135822
rect 85106 135766 85110 135822
rect 85046 135762 85110 135766
rect 85126 135822 85190 135826
rect 85126 135766 85130 135822
rect 85130 135766 85186 135822
rect 85186 135766 85190 135822
rect 85126 135762 85190 135766
rect 2886 135278 2950 135282
rect 2886 135222 2890 135278
rect 2890 135222 2946 135278
rect 2946 135222 2950 135278
rect 2886 135218 2950 135222
rect 2966 135278 3030 135282
rect 2966 135222 2970 135278
rect 2970 135222 3026 135278
rect 3026 135222 3030 135278
rect 2966 135218 3030 135222
rect 3046 135278 3110 135282
rect 3046 135222 3050 135278
rect 3050 135222 3106 135278
rect 3106 135222 3110 135278
rect 3046 135218 3110 135222
rect 3126 135278 3190 135282
rect 3126 135222 3130 135278
rect 3130 135222 3186 135278
rect 3186 135222 3190 135278
rect 3126 135218 3190 135222
rect 86886 135278 86950 135282
rect 86886 135222 86890 135278
rect 86890 135222 86946 135278
rect 86946 135222 86950 135278
rect 86886 135218 86950 135222
rect 86966 135278 87030 135282
rect 86966 135222 86970 135278
rect 86970 135222 87026 135278
rect 87026 135222 87030 135278
rect 86966 135218 87030 135222
rect 87046 135278 87110 135282
rect 87046 135222 87050 135278
rect 87050 135222 87106 135278
rect 87106 135222 87110 135278
rect 87046 135218 87110 135222
rect 87126 135278 87190 135282
rect 87126 135222 87130 135278
rect 87130 135222 87186 135278
rect 87186 135222 87190 135278
rect 87126 135218 87190 135222
rect 886 134734 950 134738
rect 886 134678 890 134734
rect 890 134678 946 134734
rect 946 134678 950 134734
rect 886 134674 950 134678
rect 966 134734 1030 134738
rect 966 134678 970 134734
rect 970 134678 1026 134734
rect 1026 134678 1030 134734
rect 966 134674 1030 134678
rect 1046 134734 1110 134738
rect 1046 134678 1050 134734
rect 1050 134678 1106 134734
rect 1106 134678 1110 134734
rect 1046 134674 1110 134678
rect 1126 134734 1190 134738
rect 1126 134678 1130 134734
rect 1130 134678 1186 134734
rect 1186 134678 1190 134734
rect 1126 134674 1190 134678
rect 84886 134734 84950 134738
rect 84886 134678 84890 134734
rect 84890 134678 84946 134734
rect 84946 134678 84950 134734
rect 84886 134674 84950 134678
rect 84966 134734 85030 134738
rect 84966 134678 84970 134734
rect 84970 134678 85026 134734
rect 85026 134678 85030 134734
rect 84966 134674 85030 134678
rect 85046 134734 85110 134738
rect 85046 134678 85050 134734
rect 85050 134678 85106 134734
rect 85106 134678 85110 134734
rect 85046 134674 85110 134678
rect 85126 134734 85190 134738
rect 85126 134678 85130 134734
rect 85130 134678 85186 134734
rect 85186 134678 85190 134734
rect 85126 134674 85190 134678
rect 2886 134190 2950 134194
rect 2886 134134 2890 134190
rect 2890 134134 2946 134190
rect 2946 134134 2950 134190
rect 2886 134130 2950 134134
rect 2966 134190 3030 134194
rect 2966 134134 2970 134190
rect 2970 134134 3026 134190
rect 3026 134134 3030 134190
rect 2966 134130 3030 134134
rect 3046 134190 3110 134194
rect 3046 134134 3050 134190
rect 3050 134134 3106 134190
rect 3106 134134 3110 134190
rect 3046 134130 3110 134134
rect 3126 134190 3190 134194
rect 3126 134134 3130 134190
rect 3130 134134 3186 134190
rect 3186 134134 3190 134190
rect 3126 134130 3190 134134
rect 86886 134190 86950 134194
rect 86886 134134 86890 134190
rect 86890 134134 86946 134190
rect 86946 134134 86950 134190
rect 86886 134130 86950 134134
rect 86966 134190 87030 134194
rect 86966 134134 86970 134190
rect 86970 134134 87026 134190
rect 87026 134134 87030 134190
rect 86966 134130 87030 134134
rect 87046 134190 87110 134194
rect 87046 134134 87050 134190
rect 87050 134134 87106 134190
rect 87106 134134 87110 134190
rect 87046 134130 87110 134134
rect 87126 134190 87190 134194
rect 87126 134134 87130 134190
rect 87130 134134 87186 134190
rect 87186 134134 87190 134190
rect 87126 134130 87190 134134
rect 886 133646 950 133650
rect 886 133590 890 133646
rect 890 133590 946 133646
rect 946 133590 950 133646
rect 886 133586 950 133590
rect 966 133646 1030 133650
rect 966 133590 970 133646
rect 970 133590 1026 133646
rect 1026 133590 1030 133646
rect 966 133586 1030 133590
rect 1046 133646 1110 133650
rect 1046 133590 1050 133646
rect 1050 133590 1106 133646
rect 1106 133590 1110 133646
rect 1046 133586 1110 133590
rect 1126 133646 1190 133650
rect 1126 133590 1130 133646
rect 1130 133590 1186 133646
rect 1186 133590 1190 133646
rect 1126 133586 1190 133590
rect 84886 133646 84950 133650
rect 84886 133590 84890 133646
rect 84890 133590 84946 133646
rect 84946 133590 84950 133646
rect 84886 133586 84950 133590
rect 84966 133646 85030 133650
rect 84966 133590 84970 133646
rect 84970 133590 85026 133646
rect 85026 133590 85030 133646
rect 84966 133586 85030 133590
rect 85046 133646 85110 133650
rect 85046 133590 85050 133646
rect 85050 133590 85106 133646
rect 85106 133590 85110 133646
rect 85046 133586 85110 133590
rect 85126 133646 85190 133650
rect 85126 133590 85130 133646
rect 85130 133590 85186 133646
rect 85186 133590 85190 133646
rect 85126 133586 85190 133590
rect 2886 133102 2950 133106
rect 2886 133046 2890 133102
rect 2890 133046 2946 133102
rect 2946 133046 2950 133102
rect 2886 133042 2950 133046
rect 2966 133102 3030 133106
rect 2966 133046 2970 133102
rect 2970 133046 3026 133102
rect 3026 133046 3030 133102
rect 2966 133042 3030 133046
rect 3046 133102 3110 133106
rect 3046 133046 3050 133102
rect 3050 133046 3106 133102
rect 3106 133046 3110 133102
rect 3046 133042 3110 133046
rect 3126 133102 3190 133106
rect 3126 133046 3130 133102
rect 3130 133046 3186 133102
rect 3186 133046 3190 133102
rect 3126 133042 3190 133046
rect 86886 133102 86950 133106
rect 86886 133046 86890 133102
rect 86890 133046 86946 133102
rect 86946 133046 86950 133102
rect 86886 133042 86950 133046
rect 86966 133102 87030 133106
rect 86966 133046 86970 133102
rect 86970 133046 87026 133102
rect 87026 133046 87030 133102
rect 86966 133042 87030 133046
rect 87046 133102 87110 133106
rect 87046 133046 87050 133102
rect 87050 133046 87106 133102
rect 87106 133046 87110 133102
rect 87046 133042 87110 133046
rect 87126 133102 87190 133106
rect 87126 133046 87130 133102
rect 87130 133046 87186 133102
rect 87186 133046 87190 133102
rect 87126 133042 87190 133046
rect 886 132558 950 132562
rect 886 132502 890 132558
rect 890 132502 946 132558
rect 946 132502 950 132558
rect 886 132498 950 132502
rect 966 132558 1030 132562
rect 966 132502 970 132558
rect 970 132502 1026 132558
rect 1026 132502 1030 132558
rect 966 132498 1030 132502
rect 1046 132558 1110 132562
rect 1046 132502 1050 132558
rect 1050 132502 1106 132558
rect 1106 132502 1110 132558
rect 1046 132498 1110 132502
rect 1126 132558 1190 132562
rect 1126 132502 1130 132558
rect 1130 132502 1186 132558
rect 1186 132502 1190 132558
rect 1126 132498 1190 132502
rect 84886 132558 84950 132562
rect 84886 132502 84890 132558
rect 84890 132502 84946 132558
rect 84946 132502 84950 132558
rect 84886 132498 84950 132502
rect 84966 132558 85030 132562
rect 84966 132502 84970 132558
rect 84970 132502 85026 132558
rect 85026 132502 85030 132558
rect 84966 132498 85030 132502
rect 85046 132558 85110 132562
rect 85046 132502 85050 132558
rect 85050 132502 85106 132558
rect 85106 132502 85110 132558
rect 85046 132498 85110 132502
rect 85126 132558 85190 132562
rect 85126 132502 85130 132558
rect 85130 132502 85186 132558
rect 85186 132502 85190 132558
rect 85126 132498 85190 132502
rect 2886 132014 2950 132018
rect 2886 131958 2890 132014
rect 2890 131958 2946 132014
rect 2946 131958 2950 132014
rect 2886 131954 2950 131958
rect 2966 132014 3030 132018
rect 2966 131958 2970 132014
rect 2970 131958 3026 132014
rect 3026 131958 3030 132014
rect 2966 131954 3030 131958
rect 3046 132014 3110 132018
rect 3046 131958 3050 132014
rect 3050 131958 3106 132014
rect 3106 131958 3110 132014
rect 3046 131954 3110 131958
rect 3126 132014 3190 132018
rect 3126 131958 3130 132014
rect 3130 131958 3186 132014
rect 3186 131958 3190 132014
rect 3126 131954 3190 131958
rect 86886 132014 86950 132018
rect 86886 131958 86890 132014
rect 86890 131958 86946 132014
rect 86946 131958 86950 132014
rect 86886 131954 86950 131958
rect 86966 132014 87030 132018
rect 86966 131958 86970 132014
rect 86970 131958 87026 132014
rect 87026 131958 87030 132014
rect 86966 131954 87030 131958
rect 87046 132014 87110 132018
rect 87046 131958 87050 132014
rect 87050 131958 87106 132014
rect 87106 131958 87110 132014
rect 87046 131954 87110 131958
rect 87126 132014 87190 132018
rect 87126 131958 87130 132014
rect 87130 131958 87186 132014
rect 87186 131958 87190 132014
rect 87126 131954 87190 131958
rect 886 131470 950 131474
rect 886 131414 890 131470
rect 890 131414 946 131470
rect 946 131414 950 131470
rect 886 131410 950 131414
rect 966 131470 1030 131474
rect 966 131414 970 131470
rect 970 131414 1026 131470
rect 1026 131414 1030 131470
rect 966 131410 1030 131414
rect 1046 131470 1110 131474
rect 1046 131414 1050 131470
rect 1050 131414 1106 131470
rect 1106 131414 1110 131470
rect 1046 131410 1110 131414
rect 1126 131470 1190 131474
rect 1126 131414 1130 131470
rect 1130 131414 1186 131470
rect 1186 131414 1190 131470
rect 1126 131410 1190 131414
rect 84886 131470 84950 131474
rect 84886 131414 84890 131470
rect 84890 131414 84946 131470
rect 84946 131414 84950 131470
rect 84886 131410 84950 131414
rect 84966 131470 85030 131474
rect 84966 131414 84970 131470
rect 84970 131414 85026 131470
rect 85026 131414 85030 131470
rect 84966 131410 85030 131414
rect 85046 131470 85110 131474
rect 85046 131414 85050 131470
rect 85050 131414 85106 131470
rect 85106 131414 85110 131470
rect 85046 131410 85110 131414
rect 85126 131470 85190 131474
rect 85126 131414 85130 131470
rect 85130 131414 85186 131470
rect 85186 131414 85190 131470
rect 85126 131410 85190 131414
rect 2886 130926 2950 130930
rect 2886 130870 2890 130926
rect 2890 130870 2946 130926
rect 2946 130870 2950 130926
rect 2886 130866 2950 130870
rect 2966 130926 3030 130930
rect 2966 130870 2970 130926
rect 2970 130870 3026 130926
rect 3026 130870 3030 130926
rect 2966 130866 3030 130870
rect 3046 130926 3110 130930
rect 3046 130870 3050 130926
rect 3050 130870 3106 130926
rect 3106 130870 3110 130926
rect 3046 130866 3110 130870
rect 3126 130926 3190 130930
rect 3126 130870 3130 130926
rect 3130 130870 3186 130926
rect 3186 130870 3190 130926
rect 3126 130866 3190 130870
rect 86886 130926 86950 130930
rect 86886 130870 86890 130926
rect 86890 130870 86946 130926
rect 86946 130870 86950 130926
rect 86886 130866 86950 130870
rect 86966 130926 87030 130930
rect 86966 130870 86970 130926
rect 86970 130870 87026 130926
rect 87026 130870 87030 130926
rect 86966 130866 87030 130870
rect 87046 130926 87110 130930
rect 87046 130870 87050 130926
rect 87050 130870 87106 130926
rect 87106 130870 87110 130926
rect 87046 130866 87110 130870
rect 87126 130926 87190 130930
rect 87126 130870 87130 130926
rect 87130 130870 87186 130926
rect 87186 130870 87190 130926
rect 87126 130866 87190 130870
rect 886 130382 950 130386
rect 886 130326 890 130382
rect 890 130326 946 130382
rect 946 130326 950 130382
rect 886 130322 950 130326
rect 966 130382 1030 130386
rect 966 130326 970 130382
rect 970 130326 1026 130382
rect 1026 130326 1030 130382
rect 966 130322 1030 130326
rect 1046 130382 1110 130386
rect 1046 130326 1050 130382
rect 1050 130326 1106 130382
rect 1106 130326 1110 130382
rect 1046 130322 1110 130326
rect 1126 130382 1190 130386
rect 1126 130326 1130 130382
rect 1130 130326 1186 130382
rect 1186 130326 1190 130382
rect 1126 130322 1190 130326
rect 84886 130382 84950 130386
rect 84886 130326 84890 130382
rect 84890 130326 84946 130382
rect 84946 130326 84950 130382
rect 84886 130322 84950 130326
rect 84966 130382 85030 130386
rect 84966 130326 84970 130382
rect 84970 130326 85026 130382
rect 85026 130326 85030 130382
rect 84966 130322 85030 130326
rect 85046 130382 85110 130386
rect 85046 130326 85050 130382
rect 85050 130326 85106 130382
rect 85106 130326 85110 130382
rect 85046 130322 85110 130326
rect 85126 130382 85190 130386
rect 85126 130326 85130 130382
rect 85130 130326 85186 130382
rect 85186 130326 85190 130382
rect 85126 130322 85190 130326
rect 2886 129838 2950 129842
rect 2886 129782 2890 129838
rect 2890 129782 2946 129838
rect 2946 129782 2950 129838
rect 2886 129778 2950 129782
rect 2966 129838 3030 129842
rect 2966 129782 2970 129838
rect 2970 129782 3026 129838
rect 3026 129782 3030 129838
rect 2966 129778 3030 129782
rect 3046 129838 3110 129842
rect 3046 129782 3050 129838
rect 3050 129782 3106 129838
rect 3106 129782 3110 129838
rect 3046 129778 3110 129782
rect 3126 129838 3190 129842
rect 3126 129782 3130 129838
rect 3130 129782 3186 129838
rect 3186 129782 3190 129838
rect 3126 129778 3190 129782
rect 86886 129838 86950 129842
rect 86886 129782 86890 129838
rect 86890 129782 86946 129838
rect 86946 129782 86950 129838
rect 86886 129778 86950 129782
rect 86966 129838 87030 129842
rect 86966 129782 86970 129838
rect 86970 129782 87026 129838
rect 87026 129782 87030 129838
rect 86966 129778 87030 129782
rect 87046 129838 87110 129842
rect 87046 129782 87050 129838
rect 87050 129782 87106 129838
rect 87106 129782 87110 129838
rect 87046 129778 87110 129782
rect 87126 129838 87190 129842
rect 87126 129782 87130 129838
rect 87130 129782 87186 129838
rect 87186 129782 87190 129838
rect 87126 129778 87190 129782
rect 886 129294 950 129298
rect 886 129238 890 129294
rect 890 129238 946 129294
rect 946 129238 950 129294
rect 886 129234 950 129238
rect 966 129294 1030 129298
rect 966 129238 970 129294
rect 970 129238 1026 129294
rect 1026 129238 1030 129294
rect 966 129234 1030 129238
rect 1046 129294 1110 129298
rect 1046 129238 1050 129294
rect 1050 129238 1106 129294
rect 1106 129238 1110 129294
rect 1046 129234 1110 129238
rect 1126 129294 1190 129298
rect 1126 129238 1130 129294
rect 1130 129238 1186 129294
rect 1186 129238 1190 129294
rect 1126 129234 1190 129238
rect 84886 129294 84950 129298
rect 84886 129238 84890 129294
rect 84890 129238 84946 129294
rect 84946 129238 84950 129294
rect 84886 129234 84950 129238
rect 84966 129294 85030 129298
rect 84966 129238 84970 129294
rect 84970 129238 85026 129294
rect 85026 129238 85030 129294
rect 84966 129234 85030 129238
rect 85046 129294 85110 129298
rect 85046 129238 85050 129294
rect 85050 129238 85106 129294
rect 85106 129238 85110 129294
rect 85046 129234 85110 129238
rect 85126 129294 85190 129298
rect 85126 129238 85130 129294
rect 85130 129238 85186 129294
rect 85186 129238 85190 129294
rect 85126 129234 85190 129238
rect 2886 128750 2950 128754
rect 2886 128694 2890 128750
rect 2890 128694 2946 128750
rect 2946 128694 2950 128750
rect 2886 128690 2950 128694
rect 2966 128750 3030 128754
rect 2966 128694 2970 128750
rect 2970 128694 3026 128750
rect 3026 128694 3030 128750
rect 2966 128690 3030 128694
rect 3046 128750 3110 128754
rect 3046 128694 3050 128750
rect 3050 128694 3106 128750
rect 3106 128694 3110 128750
rect 3046 128690 3110 128694
rect 3126 128750 3190 128754
rect 3126 128694 3130 128750
rect 3130 128694 3186 128750
rect 3186 128694 3190 128750
rect 3126 128690 3190 128694
rect 86886 128750 86950 128754
rect 86886 128694 86890 128750
rect 86890 128694 86946 128750
rect 86946 128694 86950 128750
rect 86886 128690 86950 128694
rect 86966 128750 87030 128754
rect 86966 128694 86970 128750
rect 86970 128694 87026 128750
rect 87026 128694 87030 128750
rect 86966 128690 87030 128694
rect 87046 128750 87110 128754
rect 87046 128694 87050 128750
rect 87050 128694 87106 128750
rect 87106 128694 87110 128750
rect 87046 128690 87110 128694
rect 87126 128750 87190 128754
rect 87126 128694 87130 128750
rect 87130 128694 87186 128750
rect 87186 128694 87190 128750
rect 87126 128690 87190 128694
rect 886 128206 950 128210
rect 886 128150 890 128206
rect 890 128150 946 128206
rect 946 128150 950 128206
rect 886 128146 950 128150
rect 966 128206 1030 128210
rect 966 128150 970 128206
rect 970 128150 1026 128206
rect 1026 128150 1030 128206
rect 966 128146 1030 128150
rect 1046 128206 1110 128210
rect 1046 128150 1050 128206
rect 1050 128150 1106 128206
rect 1106 128150 1110 128206
rect 1046 128146 1110 128150
rect 1126 128206 1190 128210
rect 1126 128150 1130 128206
rect 1130 128150 1186 128206
rect 1186 128150 1190 128206
rect 1126 128146 1190 128150
rect 84886 128206 84950 128210
rect 84886 128150 84890 128206
rect 84890 128150 84946 128206
rect 84946 128150 84950 128206
rect 84886 128146 84950 128150
rect 84966 128206 85030 128210
rect 84966 128150 84970 128206
rect 84970 128150 85026 128206
rect 85026 128150 85030 128206
rect 84966 128146 85030 128150
rect 85046 128206 85110 128210
rect 85046 128150 85050 128206
rect 85050 128150 85106 128206
rect 85106 128150 85110 128206
rect 85046 128146 85110 128150
rect 85126 128206 85190 128210
rect 85126 128150 85130 128206
rect 85130 128150 85186 128206
rect 85186 128150 85190 128206
rect 85126 128146 85190 128150
rect 2886 127662 2950 127666
rect 2886 127606 2890 127662
rect 2890 127606 2946 127662
rect 2946 127606 2950 127662
rect 2886 127602 2950 127606
rect 2966 127662 3030 127666
rect 2966 127606 2970 127662
rect 2970 127606 3026 127662
rect 3026 127606 3030 127662
rect 2966 127602 3030 127606
rect 3046 127662 3110 127666
rect 3046 127606 3050 127662
rect 3050 127606 3106 127662
rect 3106 127606 3110 127662
rect 3046 127602 3110 127606
rect 3126 127662 3190 127666
rect 3126 127606 3130 127662
rect 3130 127606 3186 127662
rect 3186 127606 3190 127662
rect 3126 127602 3190 127606
rect 86886 127662 86950 127666
rect 86886 127606 86890 127662
rect 86890 127606 86946 127662
rect 86946 127606 86950 127662
rect 86886 127602 86950 127606
rect 86966 127662 87030 127666
rect 86966 127606 86970 127662
rect 86970 127606 87026 127662
rect 87026 127606 87030 127662
rect 86966 127602 87030 127606
rect 87046 127662 87110 127666
rect 87046 127606 87050 127662
rect 87050 127606 87106 127662
rect 87106 127606 87110 127662
rect 87046 127602 87110 127606
rect 87126 127662 87190 127666
rect 87126 127606 87130 127662
rect 87130 127606 87186 127662
rect 87186 127606 87190 127662
rect 87126 127602 87190 127606
rect 886 127118 950 127122
rect 886 127062 890 127118
rect 890 127062 946 127118
rect 946 127062 950 127118
rect 886 127058 950 127062
rect 966 127118 1030 127122
rect 966 127062 970 127118
rect 970 127062 1026 127118
rect 1026 127062 1030 127118
rect 966 127058 1030 127062
rect 1046 127118 1110 127122
rect 1046 127062 1050 127118
rect 1050 127062 1106 127118
rect 1106 127062 1110 127118
rect 1046 127058 1110 127062
rect 1126 127118 1190 127122
rect 1126 127062 1130 127118
rect 1130 127062 1186 127118
rect 1186 127062 1190 127118
rect 1126 127058 1190 127062
rect 84886 127118 84950 127122
rect 84886 127062 84890 127118
rect 84890 127062 84946 127118
rect 84946 127062 84950 127118
rect 84886 127058 84950 127062
rect 84966 127118 85030 127122
rect 84966 127062 84970 127118
rect 84970 127062 85026 127118
rect 85026 127062 85030 127118
rect 84966 127058 85030 127062
rect 85046 127118 85110 127122
rect 85046 127062 85050 127118
rect 85050 127062 85106 127118
rect 85106 127062 85110 127118
rect 85046 127058 85110 127062
rect 85126 127118 85190 127122
rect 85126 127062 85130 127118
rect 85130 127062 85186 127118
rect 85186 127062 85190 127118
rect 85126 127058 85190 127062
rect 2886 126574 2950 126578
rect 2886 126518 2890 126574
rect 2890 126518 2946 126574
rect 2946 126518 2950 126574
rect 2886 126514 2950 126518
rect 2966 126574 3030 126578
rect 2966 126518 2970 126574
rect 2970 126518 3026 126574
rect 3026 126518 3030 126574
rect 2966 126514 3030 126518
rect 3046 126574 3110 126578
rect 3046 126518 3050 126574
rect 3050 126518 3106 126574
rect 3106 126518 3110 126574
rect 3046 126514 3110 126518
rect 3126 126574 3190 126578
rect 3126 126518 3130 126574
rect 3130 126518 3186 126574
rect 3186 126518 3190 126574
rect 3126 126514 3190 126518
rect 86886 126574 86950 126578
rect 86886 126518 86890 126574
rect 86890 126518 86946 126574
rect 86946 126518 86950 126574
rect 86886 126514 86950 126518
rect 86966 126574 87030 126578
rect 86966 126518 86970 126574
rect 86970 126518 87026 126574
rect 87026 126518 87030 126574
rect 86966 126514 87030 126518
rect 87046 126574 87110 126578
rect 87046 126518 87050 126574
rect 87050 126518 87106 126574
rect 87106 126518 87110 126574
rect 87046 126514 87110 126518
rect 87126 126574 87190 126578
rect 87126 126518 87130 126574
rect 87130 126518 87186 126574
rect 87186 126518 87190 126574
rect 87126 126514 87190 126518
rect 886 126030 950 126034
rect 886 125974 890 126030
rect 890 125974 946 126030
rect 946 125974 950 126030
rect 886 125970 950 125974
rect 966 126030 1030 126034
rect 966 125974 970 126030
rect 970 125974 1026 126030
rect 1026 125974 1030 126030
rect 966 125970 1030 125974
rect 1046 126030 1110 126034
rect 1046 125974 1050 126030
rect 1050 125974 1106 126030
rect 1106 125974 1110 126030
rect 1046 125970 1110 125974
rect 1126 126030 1190 126034
rect 1126 125974 1130 126030
rect 1130 125974 1186 126030
rect 1186 125974 1190 126030
rect 1126 125970 1190 125974
rect 84886 126030 84950 126034
rect 84886 125974 84890 126030
rect 84890 125974 84946 126030
rect 84946 125974 84950 126030
rect 84886 125970 84950 125974
rect 84966 126030 85030 126034
rect 84966 125974 84970 126030
rect 84970 125974 85026 126030
rect 85026 125974 85030 126030
rect 84966 125970 85030 125974
rect 85046 126030 85110 126034
rect 85046 125974 85050 126030
rect 85050 125974 85106 126030
rect 85106 125974 85110 126030
rect 85046 125970 85110 125974
rect 85126 126030 85190 126034
rect 85126 125974 85130 126030
rect 85130 125974 85186 126030
rect 85186 125974 85190 126030
rect 85126 125970 85190 125974
rect 2886 125486 2950 125490
rect 2886 125430 2890 125486
rect 2890 125430 2946 125486
rect 2946 125430 2950 125486
rect 2886 125426 2950 125430
rect 2966 125486 3030 125490
rect 2966 125430 2970 125486
rect 2970 125430 3026 125486
rect 3026 125430 3030 125486
rect 2966 125426 3030 125430
rect 3046 125486 3110 125490
rect 3046 125430 3050 125486
rect 3050 125430 3106 125486
rect 3106 125430 3110 125486
rect 3046 125426 3110 125430
rect 3126 125486 3190 125490
rect 3126 125430 3130 125486
rect 3130 125430 3186 125486
rect 3186 125430 3190 125486
rect 3126 125426 3190 125430
rect 86886 125486 86950 125490
rect 86886 125430 86890 125486
rect 86890 125430 86946 125486
rect 86946 125430 86950 125486
rect 86886 125426 86950 125430
rect 86966 125486 87030 125490
rect 86966 125430 86970 125486
rect 86970 125430 87026 125486
rect 87026 125430 87030 125486
rect 86966 125426 87030 125430
rect 87046 125486 87110 125490
rect 87046 125430 87050 125486
rect 87050 125430 87106 125486
rect 87106 125430 87110 125486
rect 87046 125426 87110 125430
rect 87126 125486 87190 125490
rect 87126 125430 87130 125486
rect 87130 125430 87186 125486
rect 87186 125430 87190 125486
rect 87126 125426 87190 125430
rect 886 124942 950 124946
rect 886 124886 890 124942
rect 890 124886 946 124942
rect 946 124886 950 124942
rect 886 124882 950 124886
rect 966 124942 1030 124946
rect 966 124886 970 124942
rect 970 124886 1026 124942
rect 1026 124886 1030 124942
rect 966 124882 1030 124886
rect 1046 124942 1110 124946
rect 1046 124886 1050 124942
rect 1050 124886 1106 124942
rect 1106 124886 1110 124942
rect 1046 124882 1110 124886
rect 1126 124942 1190 124946
rect 1126 124886 1130 124942
rect 1130 124886 1186 124942
rect 1186 124886 1190 124942
rect 1126 124882 1190 124886
rect 84886 124942 84950 124946
rect 84886 124886 84890 124942
rect 84890 124886 84946 124942
rect 84946 124886 84950 124942
rect 84886 124882 84950 124886
rect 84966 124942 85030 124946
rect 84966 124886 84970 124942
rect 84970 124886 85026 124942
rect 85026 124886 85030 124942
rect 84966 124882 85030 124886
rect 85046 124942 85110 124946
rect 85046 124886 85050 124942
rect 85050 124886 85106 124942
rect 85106 124886 85110 124942
rect 85046 124882 85110 124886
rect 85126 124942 85190 124946
rect 85126 124886 85130 124942
rect 85130 124886 85186 124942
rect 85186 124886 85190 124942
rect 85126 124882 85190 124886
rect 2306 124678 2370 124742
rect 2886 124398 2950 124402
rect 2886 124342 2890 124398
rect 2890 124342 2946 124398
rect 2946 124342 2950 124398
rect 2886 124338 2950 124342
rect 2966 124398 3030 124402
rect 2966 124342 2970 124398
rect 2970 124342 3026 124398
rect 3026 124342 3030 124398
rect 2966 124338 3030 124342
rect 3046 124398 3110 124402
rect 3046 124342 3050 124398
rect 3050 124342 3106 124398
rect 3106 124342 3110 124398
rect 3046 124338 3110 124342
rect 3126 124398 3190 124402
rect 3126 124342 3130 124398
rect 3130 124342 3186 124398
rect 3186 124342 3190 124398
rect 3126 124338 3190 124342
rect 86886 124398 86950 124402
rect 86886 124342 86890 124398
rect 86890 124342 86946 124398
rect 86946 124342 86950 124398
rect 86886 124338 86950 124342
rect 86966 124398 87030 124402
rect 86966 124342 86970 124398
rect 86970 124342 87026 124398
rect 87026 124342 87030 124398
rect 86966 124338 87030 124342
rect 87046 124398 87110 124402
rect 87046 124342 87050 124398
rect 87050 124342 87106 124398
rect 87106 124342 87110 124398
rect 87046 124338 87110 124342
rect 87126 124398 87190 124402
rect 87126 124342 87130 124398
rect 87130 124342 87186 124398
rect 87186 124342 87190 124398
rect 87126 124338 87190 124342
rect 886 123854 950 123858
rect 886 123798 890 123854
rect 890 123798 946 123854
rect 946 123798 950 123854
rect 886 123794 950 123798
rect 966 123854 1030 123858
rect 966 123798 970 123854
rect 970 123798 1026 123854
rect 1026 123798 1030 123854
rect 966 123794 1030 123798
rect 1046 123854 1110 123858
rect 1046 123798 1050 123854
rect 1050 123798 1106 123854
rect 1106 123798 1110 123854
rect 1046 123794 1110 123798
rect 1126 123854 1190 123858
rect 1126 123798 1130 123854
rect 1130 123798 1186 123854
rect 1186 123798 1190 123854
rect 1126 123794 1190 123798
rect 84886 123854 84950 123858
rect 84886 123798 84890 123854
rect 84890 123798 84946 123854
rect 84946 123798 84950 123854
rect 84886 123794 84950 123798
rect 84966 123854 85030 123858
rect 84966 123798 84970 123854
rect 84970 123798 85026 123854
rect 85026 123798 85030 123854
rect 84966 123794 85030 123798
rect 85046 123854 85110 123858
rect 85046 123798 85050 123854
rect 85050 123798 85106 123854
rect 85106 123798 85110 123854
rect 85046 123794 85110 123798
rect 85126 123854 85190 123858
rect 85126 123798 85130 123854
rect 85130 123798 85186 123854
rect 85186 123798 85190 123854
rect 85126 123794 85190 123798
rect 2886 123310 2950 123314
rect 2886 123254 2890 123310
rect 2890 123254 2946 123310
rect 2946 123254 2950 123310
rect 2886 123250 2950 123254
rect 2966 123310 3030 123314
rect 2966 123254 2970 123310
rect 2970 123254 3026 123310
rect 3026 123254 3030 123310
rect 2966 123250 3030 123254
rect 3046 123310 3110 123314
rect 3046 123254 3050 123310
rect 3050 123254 3106 123310
rect 3106 123254 3110 123310
rect 3046 123250 3110 123254
rect 3126 123310 3190 123314
rect 3126 123254 3130 123310
rect 3130 123254 3186 123310
rect 3186 123254 3190 123310
rect 3126 123250 3190 123254
rect 86886 123310 86950 123314
rect 86886 123254 86890 123310
rect 86890 123254 86946 123310
rect 86946 123254 86950 123310
rect 86886 123250 86950 123254
rect 86966 123310 87030 123314
rect 86966 123254 86970 123310
rect 86970 123254 87026 123310
rect 87026 123254 87030 123310
rect 86966 123250 87030 123254
rect 87046 123310 87110 123314
rect 87046 123254 87050 123310
rect 87050 123254 87106 123310
rect 87106 123254 87110 123310
rect 87046 123250 87110 123254
rect 87126 123310 87190 123314
rect 87126 123254 87130 123310
rect 87130 123254 87186 123310
rect 87186 123254 87190 123310
rect 87126 123250 87190 123254
rect 886 122766 950 122770
rect 886 122710 890 122766
rect 890 122710 946 122766
rect 946 122710 950 122766
rect 886 122706 950 122710
rect 966 122766 1030 122770
rect 966 122710 970 122766
rect 970 122710 1026 122766
rect 1026 122710 1030 122766
rect 966 122706 1030 122710
rect 1046 122766 1110 122770
rect 1046 122710 1050 122766
rect 1050 122710 1106 122766
rect 1106 122710 1110 122766
rect 1046 122706 1110 122710
rect 1126 122766 1190 122770
rect 1126 122710 1130 122766
rect 1130 122710 1186 122766
rect 1186 122710 1190 122766
rect 1126 122706 1190 122710
rect 84886 122766 84950 122770
rect 84886 122710 84890 122766
rect 84890 122710 84946 122766
rect 84946 122710 84950 122766
rect 84886 122706 84950 122710
rect 84966 122766 85030 122770
rect 84966 122710 84970 122766
rect 84970 122710 85026 122766
rect 85026 122710 85030 122766
rect 84966 122706 85030 122710
rect 85046 122766 85110 122770
rect 85046 122710 85050 122766
rect 85050 122710 85106 122766
rect 85106 122710 85110 122766
rect 85046 122706 85110 122710
rect 85126 122766 85190 122770
rect 85126 122710 85130 122766
rect 85130 122710 85186 122766
rect 85186 122710 85190 122766
rect 85126 122706 85190 122710
rect 2886 122222 2950 122226
rect 2886 122166 2890 122222
rect 2890 122166 2946 122222
rect 2946 122166 2950 122222
rect 2886 122162 2950 122166
rect 2966 122222 3030 122226
rect 2966 122166 2970 122222
rect 2970 122166 3026 122222
rect 3026 122166 3030 122222
rect 2966 122162 3030 122166
rect 3046 122222 3110 122226
rect 3046 122166 3050 122222
rect 3050 122166 3106 122222
rect 3106 122166 3110 122222
rect 3046 122162 3110 122166
rect 3126 122222 3190 122226
rect 3126 122166 3130 122222
rect 3130 122166 3186 122222
rect 3186 122166 3190 122222
rect 3126 122162 3190 122166
rect 86886 122222 86950 122226
rect 86886 122166 86890 122222
rect 86890 122166 86946 122222
rect 86946 122166 86950 122222
rect 86886 122162 86950 122166
rect 86966 122222 87030 122226
rect 86966 122166 86970 122222
rect 86970 122166 87026 122222
rect 87026 122166 87030 122222
rect 86966 122162 87030 122166
rect 87046 122222 87110 122226
rect 87046 122166 87050 122222
rect 87050 122166 87106 122222
rect 87106 122166 87110 122222
rect 87046 122162 87110 122166
rect 87126 122222 87190 122226
rect 87126 122166 87130 122222
rect 87130 122166 87186 122222
rect 87186 122166 87190 122222
rect 87126 122162 87190 122166
rect 886 121678 950 121682
rect 886 121622 890 121678
rect 890 121622 946 121678
rect 946 121622 950 121678
rect 886 121618 950 121622
rect 966 121678 1030 121682
rect 966 121622 970 121678
rect 970 121622 1026 121678
rect 1026 121622 1030 121678
rect 966 121618 1030 121622
rect 1046 121678 1110 121682
rect 1046 121622 1050 121678
rect 1050 121622 1106 121678
rect 1106 121622 1110 121678
rect 1046 121618 1110 121622
rect 1126 121678 1190 121682
rect 1126 121622 1130 121678
rect 1130 121622 1186 121678
rect 1186 121622 1190 121678
rect 1126 121618 1190 121622
rect 84886 121678 84950 121682
rect 84886 121622 84890 121678
rect 84890 121622 84946 121678
rect 84946 121622 84950 121678
rect 84886 121618 84950 121622
rect 84966 121678 85030 121682
rect 84966 121622 84970 121678
rect 84970 121622 85026 121678
rect 85026 121622 85030 121678
rect 84966 121618 85030 121622
rect 85046 121678 85110 121682
rect 85046 121622 85050 121678
rect 85050 121622 85106 121678
rect 85106 121622 85110 121678
rect 85046 121618 85110 121622
rect 85126 121678 85190 121682
rect 85126 121622 85130 121678
rect 85130 121622 85186 121678
rect 85186 121622 85190 121678
rect 85126 121618 85190 121622
rect 2886 121134 2950 121138
rect 2886 121078 2890 121134
rect 2890 121078 2946 121134
rect 2946 121078 2950 121134
rect 2886 121074 2950 121078
rect 2966 121134 3030 121138
rect 2966 121078 2970 121134
rect 2970 121078 3026 121134
rect 3026 121078 3030 121134
rect 2966 121074 3030 121078
rect 3046 121134 3110 121138
rect 3046 121078 3050 121134
rect 3050 121078 3106 121134
rect 3106 121078 3110 121134
rect 3046 121074 3110 121078
rect 3126 121134 3190 121138
rect 3126 121078 3130 121134
rect 3130 121078 3186 121134
rect 3186 121078 3190 121134
rect 3126 121074 3190 121078
rect 86886 121134 86950 121138
rect 86886 121078 86890 121134
rect 86890 121078 86946 121134
rect 86946 121078 86950 121134
rect 86886 121074 86950 121078
rect 86966 121134 87030 121138
rect 86966 121078 86970 121134
rect 86970 121078 87026 121134
rect 87026 121078 87030 121134
rect 86966 121074 87030 121078
rect 87046 121134 87110 121138
rect 87046 121078 87050 121134
rect 87050 121078 87106 121134
rect 87106 121078 87110 121134
rect 87046 121074 87110 121078
rect 87126 121134 87190 121138
rect 87126 121078 87130 121134
rect 87130 121078 87186 121134
rect 87186 121078 87190 121134
rect 87126 121074 87190 121078
rect 886 120590 950 120594
rect 886 120534 890 120590
rect 890 120534 946 120590
rect 946 120534 950 120590
rect 886 120530 950 120534
rect 966 120590 1030 120594
rect 966 120534 970 120590
rect 970 120534 1026 120590
rect 1026 120534 1030 120590
rect 966 120530 1030 120534
rect 1046 120590 1110 120594
rect 1046 120534 1050 120590
rect 1050 120534 1106 120590
rect 1106 120534 1110 120590
rect 1046 120530 1110 120534
rect 1126 120590 1190 120594
rect 1126 120534 1130 120590
rect 1130 120534 1186 120590
rect 1186 120534 1190 120590
rect 1126 120530 1190 120534
rect 84886 120590 84950 120594
rect 84886 120534 84890 120590
rect 84890 120534 84946 120590
rect 84946 120534 84950 120590
rect 84886 120530 84950 120534
rect 84966 120590 85030 120594
rect 84966 120534 84970 120590
rect 84970 120534 85026 120590
rect 85026 120534 85030 120590
rect 84966 120530 85030 120534
rect 85046 120590 85110 120594
rect 85046 120534 85050 120590
rect 85050 120534 85106 120590
rect 85106 120534 85110 120590
rect 85046 120530 85110 120534
rect 85126 120590 85190 120594
rect 85126 120534 85130 120590
rect 85130 120534 85186 120590
rect 85186 120534 85190 120590
rect 85126 120530 85190 120534
rect 2886 120046 2950 120050
rect 2886 119990 2890 120046
rect 2890 119990 2946 120046
rect 2946 119990 2950 120046
rect 2886 119986 2950 119990
rect 2966 120046 3030 120050
rect 2966 119990 2970 120046
rect 2970 119990 3026 120046
rect 3026 119990 3030 120046
rect 2966 119986 3030 119990
rect 3046 120046 3110 120050
rect 3046 119990 3050 120046
rect 3050 119990 3106 120046
rect 3106 119990 3110 120046
rect 3046 119986 3110 119990
rect 3126 120046 3190 120050
rect 3126 119990 3130 120046
rect 3130 119990 3186 120046
rect 3186 119990 3190 120046
rect 3126 119986 3190 119990
rect 86886 120046 86950 120050
rect 86886 119990 86890 120046
rect 86890 119990 86946 120046
rect 86946 119990 86950 120046
rect 86886 119986 86950 119990
rect 86966 120046 87030 120050
rect 86966 119990 86970 120046
rect 86970 119990 87026 120046
rect 87026 119990 87030 120046
rect 86966 119986 87030 119990
rect 87046 120046 87110 120050
rect 87046 119990 87050 120046
rect 87050 119990 87106 120046
rect 87106 119990 87110 120046
rect 87046 119986 87110 119990
rect 87126 120046 87190 120050
rect 87126 119990 87130 120046
rect 87130 119990 87186 120046
rect 87186 119990 87190 120046
rect 87126 119986 87190 119990
rect 886 119502 950 119506
rect 886 119446 890 119502
rect 890 119446 946 119502
rect 946 119446 950 119502
rect 886 119442 950 119446
rect 966 119502 1030 119506
rect 966 119446 970 119502
rect 970 119446 1026 119502
rect 1026 119446 1030 119502
rect 966 119442 1030 119446
rect 1046 119502 1110 119506
rect 1046 119446 1050 119502
rect 1050 119446 1106 119502
rect 1106 119446 1110 119502
rect 1046 119442 1110 119446
rect 1126 119502 1190 119506
rect 1126 119446 1130 119502
rect 1130 119446 1186 119502
rect 1186 119446 1190 119502
rect 1126 119442 1190 119446
rect 84886 119502 84950 119506
rect 84886 119446 84890 119502
rect 84890 119446 84946 119502
rect 84946 119446 84950 119502
rect 84886 119442 84950 119446
rect 84966 119502 85030 119506
rect 84966 119446 84970 119502
rect 84970 119446 85026 119502
rect 85026 119446 85030 119502
rect 84966 119442 85030 119446
rect 85046 119502 85110 119506
rect 85046 119446 85050 119502
rect 85050 119446 85106 119502
rect 85106 119446 85110 119502
rect 85046 119442 85110 119446
rect 85126 119502 85190 119506
rect 85126 119446 85130 119502
rect 85130 119446 85186 119502
rect 85186 119446 85190 119502
rect 85126 119442 85190 119446
rect 2886 118958 2950 118962
rect 2886 118902 2890 118958
rect 2890 118902 2946 118958
rect 2946 118902 2950 118958
rect 2886 118898 2950 118902
rect 2966 118958 3030 118962
rect 2966 118902 2970 118958
rect 2970 118902 3026 118958
rect 3026 118902 3030 118958
rect 2966 118898 3030 118902
rect 3046 118958 3110 118962
rect 3046 118902 3050 118958
rect 3050 118902 3106 118958
rect 3106 118902 3110 118958
rect 3046 118898 3110 118902
rect 3126 118958 3190 118962
rect 3126 118902 3130 118958
rect 3130 118902 3186 118958
rect 3186 118902 3190 118958
rect 3126 118898 3190 118902
rect 86886 118958 86950 118962
rect 86886 118902 86890 118958
rect 86890 118902 86946 118958
rect 86946 118902 86950 118958
rect 86886 118898 86950 118902
rect 86966 118958 87030 118962
rect 86966 118902 86970 118958
rect 86970 118902 87026 118958
rect 87026 118902 87030 118958
rect 86966 118898 87030 118902
rect 87046 118958 87110 118962
rect 87046 118902 87050 118958
rect 87050 118902 87106 118958
rect 87106 118902 87110 118958
rect 87046 118898 87110 118902
rect 87126 118958 87190 118962
rect 87126 118902 87130 118958
rect 87130 118902 87186 118958
rect 87186 118902 87190 118958
rect 87126 118898 87190 118902
rect 886 118414 950 118418
rect 886 118358 890 118414
rect 890 118358 946 118414
rect 946 118358 950 118414
rect 886 118354 950 118358
rect 966 118414 1030 118418
rect 966 118358 970 118414
rect 970 118358 1026 118414
rect 1026 118358 1030 118414
rect 966 118354 1030 118358
rect 1046 118414 1110 118418
rect 1046 118358 1050 118414
rect 1050 118358 1106 118414
rect 1106 118358 1110 118414
rect 1046 118354 1110 118358
rect 1126 118414 1190 118418
rect 1126 118358 1130 118414
rect 1130 118358 1186 118414
rect 1186 118358 1190 118414
rect 1126 118354 1190 118358
rect 84886 118414 84950 118418
rect 84886 118358 84890 118414
rect 84890 118358 84946 118414
rect 84946 118358 84950 118414
rect 84886 118354 84950 118358
rect 84966 118414 85030 118418
rect 84966 118358 84970 118414
rect 84970 118358 85026 118414
rect 85026 118358 85030 118414
rect 84966 118354 85030 118358
rect 85046 118414 85110 118418
rect 85046 118358 85050 118414
rect 85050 118358 85106 118414
rect 85106 118358 85110 118414
rect 85046 118354 85110 118358
rect 85126 118414 85190 118418
rect 85126 118358 85130 118414
rect 85130 118358 85186 118414
rect 85186 118358 85190 118414
rect 85126 118354 85190 118358
rect 2886 117870 2950 117874
rect 2886 117814 2890 117870
rect 2890 117814 2946 117870
rect 2946 117814 2950 117870
rect 2886 117810 2950 117814
rect 2966 117870 3030 117874
rect 2966 117814 2970 117870
rect 2970 117814 3026 117870
rect 3026 117814 3030 117870
rect 2966 117810 3030 117814
rect 3046 117870 3110 117874
rect 3046 117814 3050 117870
rect 3050 117814 3106 117870
rect 3106 117814 3110 117870
rect 3046 117810 3110 117814
rect 3126 117870 3190 117874
rect 3126 117814 3130 117870
rect 3130 117814 3186 117870
rect 3186 117814 3190 117870
rect 3126 117810 3190 117814
rect 86886 117870 86950 117874
rect 86886 117814 86890 117870
rect 86890 117814 86946 117870
rect 86946 117814 86950 117870
rect 86886 117810 86950 117814
rect 86966 117870 87030 117874
rect 86966 117814 86970 117870
rect 86970 117814 87026 117870
rect 87026 117814 87030 117870
rect 86966 117810 87030 117814
rect 87046 117870 87110 117874
rect 87046 117814 87050 117870
rect 87050 117814 87106 117870
rect 87106 117814 87110 117870
rect 87046 117810 87110 117814
rect 87126 117870 87190 117874
rect 87126 117814 87130 117870
rect 87130 117814 87186 117870
rect 87186 117814 87190 117870
rect 87126 117810 87190 117814
rect 886 117326 950 117330
rect 886 117270 890 117326
rect 890 117270 946 117326
rect 946 117270 950 117326
rect 886 117266 950 117270
rect 966 117326 1030 117330
rect 966 117270 970 117326
rect 970 117270 1026 117326
rect 1026 117270 1030 117326
rect 966 117266 1030 117270
rect 1046 117326 1110 117330
rect 1046 117270 1050 117326
rect 1050 117270 1106 117326
rect 1106 117270 1110 117326
rect 1046 117266 1110 117270
rect 1126 117326 1190 117330
rect 1126 117270 1130 117326
rect 1130 117270 1186 117326
rect 1186 117270 1190 117326
rect 1126 117266 1190 117270
rect 84886 117326 84950 117330
rect 84886 117270 84890 117326
rect 84890 117270 84946 117326
rect 84946 117270 84950 117326
rect 84886 117266 84950 117270
rect 84966 117326 85030 117330
rect 84966 117270 84970 117326
rect 84970 117270 85026 117326
rect 85026 117270 85030 117326
rect 84966 117266 85030 117270
rect 85046 117326 85110 117330
rect 85046 117270 85050 117326
rect 85050 117270 85106 117326
rect 85106 117270 85110 117326
rect 85046 117266 85110 117270
rect 85126 117326 85190 117330
rect 85126 117270 85130 117326
rect 85130 117270 85186 117326
rect 85186 117270 85190 117326
rect 85126 117266 85190 117270
rect 2886 116782 2950 116786
rect 2886 116726 2890 116782
rect 2890 116726 2946 116782
rect 2946 116726 2950 116782
rect 2886 116722 2950 116726
rect 2966 116782 3030 116786
rect 2966 116726 2970 116782
rect 2970 116726 3026 116782
rect 3026 116726 3030 116782
rect 2966 116722 3030 116726
rect 3046 116782 3110 116786
rect 3046 116726 3050 116782
rect 3050 116726 3106 116782
rect 3106 116726 3110 116782
rect 3046 116722 3110 116726
rect 3126 116782 3190 116786
rect 3126 116726 3130 116782
rect 3130 116726 3186 116782
rect 3186 116726 3190 116782
rect 3126 116722 3190 116726
rect 86886 116782 86950 116786
rect 86886 116726 86890 116782
rect 86890 116726 86946 116782
rect 86946 116726 86950 116782
rect 86886 116722 86950 116726
rect 86966 116782 87030 116786
rect 86966 116726 86970 116782
rect 86970 116726 87026 116782
rect 87026 116726 87030 116782
rect 86966 116722 87030 116726
rect 87046 116782 87110 116786
rect 87046 116726 87050 116782
rect 87050 116726 87106 116782
rect 87106 116726 87110 116782
rect 87046 116722 87110 116726
rect 87126 116782 87190 116786
rect 87126 116726 87130 116782
rect 87130 116726 87186 116782
rect 87186 116726 87190 116782
rect 87126 116722 87190 116726
rect 886 116238 950 116242
rect 886 116182 890 116238
rect 890 116182 946 116238
rect 946 116182 950 116238
rect 886 116178 950 116182
rect 966 116238 1030 116242
rect 966 116182 970 116238
rect 970 116182 1026 116238
rect 1026 116182 1030 116238
rect 966 116178 1030 116182
rect 1046 116238 1110 116242
rect 1046 116182 1050 116238
rect 1050 116182 1106 116238
rect 1106 116182 1110 116238
rect 1046 116178 1110 116182
rect 1126 116238 1190 116242
rect 1126 116182 1130 116238
rect 1130 116182 1186 116238
rect 1186 116182 1190 116238
rect 1126 116178 1190 116182
rect 84886 116238 84950 116242
rect 84886 116182 84890 116238
rect 84890 116182 84946 116238
rect 84946 116182 84950 116238
rect 84886 116178 84950 116182
rect 84966 116238 85030 116242
rect 84966 116182 84970 116238
rect 84970 116182 85026 116238
rect 85026 116182 85030 116238
rect 84966 116178 85030 116182
rect 85046 116238 85110 116242
rect 85046 116182 85050 116238
rect 85050 116182 85106 116238
rect 85106 116182 85110 116238
rect 85046 116178 85110 116182
rect 85126 116238 85190 116242
rect 85126 116182 85130 116238
rect 85130 116182 85186 116238
rect 85186 116182 85190 116238
rect 85126 116178 85190 116182
rect 2886 115694 2950 115698
rect 2886 115638 2890 115694
rect 2890 115638 2946 115694
rect 2946 115638 2950 115694
rect 2886 115634 2950 115638
rect 2966 115694 3030 115698
rect 2966 115638 2970 115694
rect 2970 115638 3026 115694
rect 3026 115638 3030 115694
rect 2966 115634 3030 115638
rect 3046 115694 3110 115698
rect 3046 115638 3050 115694
rect 3050 115638 3106 115694
rect 3106 115638 3110 115694
rect 3046 115634 3110 115638
rect 3126 115694 3190 115698
rect 3126 115638 3130 115694
rect 3130 115638 3186 115694
rect 3186 115638 3190 115694
rect 3126 115634 3190 115638
rect 86886 115694 86950 115698
rect 86886 115638 86890 115694
rect 86890 115638 86946 115694
rect 86946 115638 86950 115694
rect 86886 115634 86950 115638
rect 86966 115694 87030 115698
rect 86966 115638 86970 115694
rect 86970 115638 87026 115694
rect 87026 115638 87030 115694
rect 86966 115634 87030 115638
rect 87046 115694 87110 115698
rect 87046 115638 87050 115694
rect 87050 115638 87106 115694
rect 87106 115638 87110 115694
rect 87046 115634 87110 115638
rect 87126 115694 87190 115698
rect 87126 115638 87130 115694
rect 87130 115638 87186 115694
rect 87186 115638 87190 115694
rect 87126 115634 87190 115638
rect 886 115150 950 115154
rect 886 115094 890 115150
rect 890 115094 946 115150
rect 946 115094 950 115150
rect 886 115090 950 115094
rect 966 115150 1030 115154
rect 966 115094 970 115150
rect 970 115094 1026 115150
rect 1026 115094 1030 115150
rect 966 115090 1030 115094
rect 1046 115150 1110 115154
rect 1046 115094 1050 115150
rect 1050 115094 1106 115150
rect 1106 115094 1110 115150
rect 1046 115090 1110 115094
rect 1126 115150 1190 115154
rect 1126 115094 1130 115150
rect 1130 115094 1186 115150
rect 1186 115094 1190 115150
rect 1126 115090 1190 115094
rect 84886 115150 84950 115154
rect 84886 115094 84890 115150
rect 84890 115094 84946 115150
rect 84946 115094 84950 115150
rect 84886 115090 84950 115094
rect 84966 115150 85030 115154
rect 84966 115094 84970 115150
rect 84970 115094 85026 115150
rect 85026 115094 85030 115150
rect 84966 115090 85030 115094
rect 85046 115150 85110 115154
rect 85046 115094 85050 115150
rect 85050 115094 85106 115150
rect 85106 115094 85110 115150
rect 85046 115090 85110 115094
rect 85126 115150 85190 115154
rect 85126 115094 85130 115150
rect 85130 115094 85186 115150
rect 85186 115094 85190 115150
rect 85126 115090 85190 115094
rect 2886 114606 2950 114610
rect 2886 114550 2890 114606
rect 2890 114550 2946 114606
rect 2946 114550 2950 114606
rect 2886 114546 2950 114550
rect 2966 114606 3030 114610
rect 2966 114550 2970 114606
rect 2970 114550 3026 114606
rect 3026 114550 3030 114606
rect 2966 114546 3030 114550
rect 3046 114606 3110 114610
rect 3046 114550 3050 114606
rect 3050 114550 3106 114606
rect 3106 114550 3110 114606
rect 3046 114546 3110 114550
rect 3126 114606 3190 114610
rect 3126 114550 3130 114606
rect 3130 114550 3186 114606
rect 3186 114550 3190 114606
rect 3126 114546 3190 114550
rect 86886 114606 86950 114610
rect 86886 114550 86890 114606
rect 86890 114550 86946 114606
rect 86946 114550 86950 114606
rect 86886 114546 86950 114550
rect 86966 114606 87030 114610
rect 86966 114550 86970 114606
rect 86970 114550 87026 114606
rect 87026 114550 87030 114606
rect 86966 114546 87030 114550
rect 87046 114606 87110 114610
rect 87046 114550 87050 114606
rect 87050 114550 87106 114606
rect 87106 114550 87110 114606
rect 87046 114546 87110 114550
rect 87126 114606 87190 114610
rect 87126 114550 87130 114606
rect 87130 114550 87186 114606
rect 87186 114550 87190 114606
rect 87126 114546 87190 114550
rect 886 114062 950 114066
rect 886 114006 890 114062
rect 890 114006 946 114062
rect 946 114006 950 114062
rect 886 114002 950 114006
rect 966 114062 1030 114066
rect 966 114006 970 114062
rect 970 114006 1026 114062
rect 1026 114006 1030 114062
rect 966 114002 1030 114006
rect 1046 114062 1110 114066
rect 1046 114006 1050 114062
rect 1050 114006 1106 114062
rect 1106 114006 1110 114062
rect 1046 114002 1110 114006
rect 1126 114062 1190 114066
rect 1126 114006 1130 114062
rect 1130 114006 1186 114062
rect 1186 114006 1190 114062
rect 1126 114002 1190 114006
rect 84886 114062 84950 114066
rect 84886 114006 84890 114062
rect 84890 114006 84946 114062
rect 84946 114006 84950 114062
rect 84886 114002 84950 114006
rect 84966 114062 85030 114066
rect 84966 114006 84970 114062
rect 84970 114006 85026 114062
rect 85026 114006 85030 114062
rect 84966 114002 85030 114006
rect 85046 114062 85110 114066
rect 85046 114006 85050 114062
rect 85050 114006 85106 114062
rect 85106 114006 85110 114062
rect 85046 114002 85110 114006
rect 85126 114062 85190 114066
rect 85126 114006 85130 114062
rect 85130 114006 85186 114062
rect 85186 114006 85190 114062
rect 85126 114002 85190 114006
rect 2886 113518 2950 113522
rect 2886 113462 2890 113518
rect 2890 113462 2946 113518
rect 2946 113462 2950 113518
rect 2886 113458 2950 113462
rect 2966 113518 3030 113522
rect 2966 113462 2970 113518
rect 2970 113462 3026 113518
rect 3026 113462 3030 113518
rect 2966 113458 3030 113462
rect 3046 113518 3110 113522
rect 3046 113462 3050 113518
rect 3050 113462 3106 113518
rect 3106 113462 3110 113518
rect 3046 113458 3110 113462
rect 3126 113518 3190 113522
rect 3126 113462 3130 113518
rect 3130 113462 3186 113518
rect 3186 113462 3190 113518
rect 3126 113458 3190 113462
rect 86886 113518 86950 113522
rect 86886 113462 86890 113518
rect 86890 113462 86946 113518
rect 86946 113462 86950 113518
rect 86886 113458 86950 113462
rect 86966 113518 87030 113522
rect 86966 113462 86970 113518
rect 86970 113462 87026 113518
rect 87026 113462 87030 113518
rect 86966 113458 87030 113462
rect 87046 113518 87110 113522
rect 87046 113462 87050 113518
rect 87050 113462 87106 113518
rect 87106 113462 87110 113518
rect 87046 113458 87110 113462
rect 87126 113518 87190 113522
rect 87126 113462 87130 113518
rect 87130 113462 87186 113518
rect 87186 113462 87190 113518
rect 87126 113458 87190 113462
rect 886 112974 950 112978
rect 886 112918 890 112974
rect 890 112918 946 112974
rect 946 112918 950 112974
rect 886 112914 950 112918
rect 966 112974 1030 112978
rect 966 112918 970 112974
rect 970 112918 1026 112974
rect 1026 112918 1030 112974
rect 966 112914 1030 112918
rect 1046 112974 1110 112978
rect 1046 112918 1050 112974
rect 1050 112918 1106 112974
rect 1106 112918 1110 112974
rect 1046 112914 1110 112918
rect 1126 112974 1190 112978
rect 1126 112918 1130 112974
rect 1130 112918 1186 112974
rect 1186 112918 1190 112974
rect 1126 112914 1190 112918
rect 84886 112974 84950 112978
rect 84886 112918 84890 112974
rect 84890 112918 84946 112974
rect 84946 112918 84950 112974
rect 84886 112914 84950 112918
rect 84966 112974 85030 112978
rect 84966 112918 84970 112974
rect 84970 112918 85026 112974
rect 85026 112918 85030 112974
rect 84966 112914 85030 112918
rect 85046 112974 85110 112978
rect 85046 112918 85050 112974
rect 85050 112918 85106 112974
rect 85106 112918 85110 112974
rect 85046 112914 85110 112918
rect 85126 112974 85190 112978
rect 85126 112918 85130 112974
rect 85130 112918 85186 112974
rect 85186 112918 85190 112974
rect 85126 112914 85190 112918
rect 2886 112430 2950 112434
rect 2886 112374 2890 112430
rect 2890 112374 2946 112430
rect 2946 112374 2950 112430
rect 2886 112370 2950 112374
rect 2966 112430 3030 112434
rect 2966 112374 2970 112430
rect 2970 112374 3026 112430
rect 3026 112374 3030 112430
rect 2966 112370 3030 112374
rect 3046 112430 3110 112434
rect 3046 112374 3050 112430
rect 3050 112374 3106 112430
rect 3106 112374 3110 112430
rect 3046 112370 3110 112374
rect 3126 112430 3190 112434
rect 3126 112374 3130 112430
rect 3130 112374 3186 112430
rect 3186 112374 3190 112430
rect 3126 112370 3190 112374
rect 86886 112430 86950 112434
rect 86886 112374 86890 112430
rect 86890 112374 86946 112430
rect 86946 112374 86950 112430
rect 86886 112370 86950 112374
rect 86966 112430 87030 112434
rect 86966 112374 86970 112430
rect 86970 112374 87026 112430
rect 87026 112374 87030 112430
rect 86966 112370 87030 112374
rect 87046 112430 87110 112434
rect 87046 112374 87050 112430
rect 87050 112374 87106 112430
rect 87106 112374 87110 112430
rect 87046 112370 87110 112374
rect 87126 112430 87190 112434
rect 87126 112374 87130 112430
rect 87130 112374 87186 112430
rect 87186 112374 87190 112430
rect 87126 112370 87190 112374
rect 886 111886 950 111890
rect 886 111830 890 111886
rect 890 111830 946 111886
rect 946 111830 950 111886
rect 886 111826 950 111830
rect 966 111886 1030 111890
rect 966 111830 970 111886
rect 970 111830 1026 111886
rect 1026 111830 1030 111886
rect 966 111826 1030 111830
rect 1046 111886 1110 111890
rect 1046 111830 1050 111886
rect 1050 111830 1106 111886
rect 1106 111830 1110 111886
rect 1046 111826 1110 111830
rect 1126 111886 1190 111890
rect 1126 111830 1130 111886
rect 1130 111830 1186 111886
rect 1186 111830 1190 111886
rect 1126 111826 1190 111830
rect 84886 111886 84950 111890
rect 84886 111830 84890 111886
rect 84890 111830 84946 111886
rect 84946 111830 84950 111886
rect 84886 111826 84950 111830
rect 84966 111886 85030 111890
rect 84966 111830 84970 111886
rect 84970 111830 85026 111886
rect 85026 111830 85030 111886
rect 84966 111826 85030 111830
rect 85046 111886 85110 111890
rect 85046 111830 85050 111886
rect 85050 111830 85106 111886
rect 85106 111830 85110 111886
rect 85046 111826 85110 111830
rect 85126 111886 85190 111890
rect 85126 111830 85130 111886
rect 85130 111830 85186 111886
rect 85186 111830 85190 111886
rect 85126 111826 85190 111830
rect 2886 111342 2950 111346
rect 2886 111286 2890 111342
rect 2890 111286 2946 111342
rect 2946 111286 2950 111342
rect 2886 111282 2950 111286
rect 2966 111342 3030 111346
rect 2966 111286 2970 111342
rect 2970 111286 3026 111342
rect 3026 111286 3030 111342
rect 2966 111282 3030 111286
rect 3046 111342 3110 111346
rect 3046 111286 3050 111342
rect 3050 111286 3106 111342
rect 3106 111286 3110 111342
rect 3046 111282 3110 111286
rect 3126 111342 3190 111346
rect 3126 111286 3130 111342
rect 3130 111286 3186 111342
rect 3186 111286 3190 111342
rect 3126 111282 3190 111286
rect 86886 111342 86950 111346
rect 86886 111286 86890 111342
rect 86890 111286 86946 111342
rect 86946 111286 86950 111342
rect 86886 111282 86950 111286
rect 86966 111342 87030 111346
rect 86966 111286 86970 111342
rect 86970 111286 87026 111342
rect 87026 111286 87030 111342
rect 86966 111282 87030 111286
rect 87046 111342 87110 111346
rect 87046 111286 87050 111342
rect 87050 111286 87106 111342
rect 87106 111286 87110 111342
rect 87046 111282 87110 111286
rect 87126 111342 87190 111346
rect 87126 111286 87130 111342
rect 87130 111286 87186 111342
rect 87186 111286 87190 111342
rect 87126 111282 87190 111286
rect 886 110798 950 110802
rect 886 110742 890 110798
rect 890 110742 946 110798
rect 946 110742 950 110798
rect 886 110738 950 110742
rect 966 110798 1030 110802
rect 966 110742 970 110798
rect 970 110742 1026 110798
rect 1026 110742 1030 110798
rect 966 110738 1030 110742
rect 1046 110798 1110 110802
rect 1046 110742 1050 110798
rect 1050 110742 1106 110798
rect 1106 110742 1110 110798
rect 1046 110738 1110 110742
rect 1126 110798 1190 110802
rect 1126 110742 1130 110798
rect 1130 110742 1186 110798
rect 1186 110742 1190 110798
rect 1126 110738 1190 110742
rect 84886 110798 84950 110802
rect 84886 110742 84890 110798
rect 84890 110742 84946 110798
rect 84946 110742 84950 110798
rect 84886 110738 84950 110742
rect 84966 110798 85030 110802
rect 84966 110742 84970 110798
rect 84970 110742 85026 110798
rect 85026 110742 85030 110798
rect 84966 110738 85030 110742
rect 85046 110798 85110 110802
rect 85046 110742 85050 110798
rect 85050 110742 85106 110798
rect 85106 110742 85110 110798
rect 85046 110738 85110 110742
rect 85126 110798 85190 110802
rect 85126 110742 85130 110798
rect 85130 110742 85186 110798
rect 85186 110742 85190 110798
rect 85126 110738 85190 110742
rect 2886 110254 2950 110258
rect 2886 110198 2890 110254
rect 2890 110198 2946 110254
rect 2946 110198 2950 110254
rect 2886 110194 2950 110198
rect 2966 110254 3030 110258
rect 2966 110198 2970 110254
rect 2970 110198 3026 110254
rect 3026 110198 3030 110254
rect 2966 110194 3030 110198
rect 3046 110254 3110 110258
rect 3046 110198 3050 110254
rect 3050 110198 3106 110254
rect 3106 110198 3110 110254
rect 3046 110194 3110 110198
rect 3126 110254 3190 110258
rect 3126 110198 3130 110254
rect 3130 110198 3186 110254
rect 3186 110198 3190 110254
rect 3126 110194 3190 110198
rect 86886 110254 86950 110258
rect 86886 110198 86890 110254
rect 86890 110198 86946 110254
rect 86946 110198 86950 110254
rect 86886 110194 86950 110198
rect 86966 110254 87030 110258
rect 86966 110198 86970 110254
rect 86970 110198 87026 110254
rect 87026 110198 87030 110254
rect 86966 110194 87030 110198
rect 87046 110254 87110 110258
rect 87046 110198 87050 110254
rect 87050 110198 87106 110254
rect 87106 110198 87110 110254
rect 87046 110194 87110 110198
rect 87126 110254 87190 110258
rect 87126 110198 87130 110254
rect 87130 110198 87186 110254
rect 87186 110198 87190 110254
rect 87126 110194 87190 110198
rect 886 109710 950 109714
rect 886 109654 890 109710
rect 890 109654 946 109710
rect 946 109654 950 109710
rect 886 109650 950 109654
rect 966 109710 1030 109714
rect 966 109654 970 109710
rect 970 109654 1026 109710
rect 1026 109654 1030 109710
rect 966 109650 1030 109654
rect 1046 109710 1110 109714
rect 1046 109654 1050 109710
rect 1050 109654 1106 109710
rect 1106 109654 1110 109710
rect 1046 109650 1110 109654
rect 1126 109710 1190 109714
rect 1126 109654 1130 109710
rect 1130 109654 1186 109710
rect 1186 109654 1190 109710
rect 1126 109650 1190 109654
rect 84886 109710 84950 109714
rect 84886 109654 84890 109710
rect 84890 109654 84946 109710
rect 84946 109654 84950 109710
rect 84886 109650 84950 109654
rect 84966 109710 85030 109714
rect 84966 109654 84970 109710
rect 84970 109654 85026 109710
rect 85026 109654 85030 109710
rect 84966 109650 85030 109654
rect 85046 109710 85110 109714
rect 85046 109654 85050 109710
rect 85050 109654 85106 109710
rect 85106 109654 85110 109710
rect 85046 109650 85110 109654
rect 85126 109710 85190 109714
rect 85126 109654 85130 109710
rect 85130 109654 85186 109710
rect 85186 109654 85190 109710
rect 85126 109650 85190 109654
rect 2886 109166 2950 109170
rect 2886 109110 2890 109166
rect 2890 109110 2946 109166
rect 2946 109110 2950 109166
rect 2886 109106 2950 109110
rect 2966 109166 3030 109170
rect 2966 109110 2970 109166
rect 2970 109110 3026 109166
rect 3026 109110 3030 109166
rect 2966 109106 3030 109110
rect 3046 109166 3110 109170
rect 3046 109110 3050 109166
rect 3050 109110 3106 109166
rect 3106 109110 3110 109166
rect 3046 109106 3110 109110
rect 3126 109166 3190 109170
rect 3126 109110 3130 109166
rect 3130 109110 3186 109166
rect 3186 109110 3190 109166
rect 3126 109106 3190 109110
rect 86886 109166 86950 109170
rect 86886 109110 86890 109166
rect 86890 109110 86946 109166
rect 86946 109110 86950 109166
rect 86886 109106 86950 109110
rect 86966 109166 87030 109170
rect 86966 109110 86970 109166
rect 86970 109110 87026 109166
rect 87026 109110 87030 109166
rect 86966 109106 87030 109110
rect 87046 109166 87110 109170
rect 87046 109110 87050 109166
rect 87050 109110 87106 109166
rect 87106 109110 87110 109166
rect 87046 109106 87110 109110
rect 87126 109166 87190 109170
rect 87126 109110 87130 109166
rect 87130 109110 87186 109166
rect 87186 109110 87190 109166
rect 87126 109106 87190 109110
rect 886 108622 950 108626
rect 886 108566 890 108622
rect 890 108566 946 108622
rect 946 108566 950 108622
rect 886 108562 950 108566
rect 966 108622 1030 108626
rect 966 108566 970 108622
rect 970 108566 1026 108622
rect 1026 108566 1030 108622
rect 966 108562 1030 108566
rect 1046 108622 1110 108626
rect 1046 108566 1050 108622
rect 1050 108566 1106 108622
rect 1106 108566 1110 108622
rect 1046 108562 1110 108566
rect 1126 108622 1190 108626
rect 1126 108566 1130 108622
rect 1130 108566 1186 108622
rect 1186 108566 1190 108622
rect 1126 108562 1190 108566
rect 84886 108622 84950 108626
rect 84886 108566 84890 108622
rect 84890 108566 84946 108622
rect 84946 108566 84950 108622
rect 84886 108562 84950 108566
rect 84966 108622 85030 108626
rect 84966 108566 84970 108622
rect 84970 108566 85026 108622
rect 85026 108566 85030 108622
rect 84966 108562 85030 108566
rect 85046 108622 85110 108626
rect 85046 108566 85050 108622
rect 85050 108566 85106 108622
rect 85106 108566 85110 108622
rect 85046 108562 85110 108566
rect 85126 108622 85190 108626
rect 85126 108566 85130 108622
rect 85130 108566 85186 108622
rect 85186 108566 85190 108622
rect 85126 108562 85190 108566
rect 2306 108086 2370 108150
rect 2886 108078 2950 108082
rect 2886 108022 2890 108078
rect 2890 108022 2946 108078
rect 2946 108022 2950 108078
rect 2886 108018 2950 108022
rect 2966 108078 3030 108082
rect 2966 108022 2970 108078
rect 2970 108022 3026 108078
rect 3026 108022 3030 108078
rect 2966 108018 3030 108022
rect 3046 108078 3110 108082
rect 3046 108022 3050 108078
rect 3050 108022 3106 108078
rect 3106 108022 3110 108078
rect 3046 108018 3110 108022
rect 3126 108078 3190 108082
rect 3126 108022 3130 108078
rect 3130 108022 3186 108078
rect 3186 108022 3190 108078
rect 3126 108018 3190 108022
rect 86886 108078 86950 108082
rect 86886 108022 86890 108078
rect 86890 108022 86946 108078
rect 86946 108022 86950 108078
rect 86886 108018 86950 108022
rect 86966 108078 87030 108082
rect 86966 108022 86970 108078
rect 86970 108022 87026 108078
rect 87026 108022 87030 108078
rect 86966 108018 87030 108022
rect 87046 108078 87110 108082
rect 87046 108022 87050 108078
rect 87050 108022 87106 108078
rect 87106 108022 87110 108078
rect 87046 108018 87110 108022
rect 87126 108078 87190 108082
rect 87126 108022 87130 108078
rect 87130 108022 87186 108078
rect 87186 108022 87190 108078
rect 87126 108018 87190 108022
rect 886 107534 950 107538
rect 886 107478 890 107534
rect 890 107478 946 107534
rect 946 107478 950 107534
rect 886 107474 950 107478
rect 966 107534 1030 107538
rect 966 107478 970 107534
rect 970 107478 1026 107534
rect 1026 107478 1030 107534
rect 966 107474 1030 107478
rect 1046 107534 1110 107538
rect 1046 107478 1050 107534
rect 1050 107478 1106 107534
rect 1106 107478 1110 107534
rect 1046 107474 1110 107478
rect 1126 107534 1190 107538
rect 1126 107478 1130 107534
rect 1130 107478 1186 107534
rect 1186 107478 1190 107534
rect 1126 107474 1190 107478
rect 84886 107534 84950 107538
rect 84886 107478 84890 107534
rect 84890 107478 84946 107534
rect 84946 107478 84950 107534
rect 84886 107474 84950 107478
rect 84966 107534 85030 107538
rect 84966 107478 84970 107534
rect 84970 107478 85026 107534
rect 85026 107478 85030 107534
rect 84966 107474 85030 107478
rect 85046 107534 85110 107538
rect 85046 107478 85050 107534
rect 85050 107478 85106 107534
rect 85106 107478 85110 107534
rect 85046 107474 85110 107478
rect 85126 107534 85190 107538
rect 85126 107478 85130 107534
rect 85130 107478 85186 107534
rect 85186 107478 85190 107534
rect 85126 107474 85190 107478
rect 2886 106990 2950 106994
rect 2886 106934 2890 106990
rect 2890 106934 2946 106990
rect 2946 106934 2950 106990
rect 2886 106930 2950 106934
rect 2966 106990 3030 106994
rect 2966 106934 2970 106990
rect 2970 106934 3026 106990
rect 3026 106934 3030 106990
rect 2966 106930 3030 106934
rect 3046 106990 3110 106994
rect 3046 106934 3050 106990
rect 3050 106934 3106 106990
rect 3106 106934 3110 106990
rect 3046 106930 3110 106934
rect 3126 106990 3190 106994
rect 3126 106934 3130 106990
rect 3130 106934 3186 106990
rect 3186 106934 3190 106990
rect 3126 106930 3190 106934
rect 86886 106990 86950 106994
rect 86886 106934 86890 106990
rect 86890 106934 86946 106990
rect 86946 106934 86950 106990
rect 86886 106930 86950 106934
rect 86966 106990 87030 106994
rect 86966 106934 86970 106990
rect 86970 106934 87026 106990
rect 87026 106934 87030 106990
rect 86966 106930 87030 106934
rect 87046 106990 87110 106994
rect 87046 106934 87050 106990
rect 87050 106934 87106 106990
rect 87106 106934 87110 106990
rect 87046 106930 87110 106934
rect 87126 106990 87190 106994
rect 87126 106934 87130 106990
rect 87130 106934 87186 106990
rect 87186 106934 87190 106990
rect 87126 106930 87190 106934
rect 886 106446 950 106450
rect 886 106390 890 106446
rect 890 106390 946 106446
rect 946 106390 950 106446
rect 886 106386 950 106390
rect 966 106446 1030 106450
rect 966 106390 970 106446
rect 970 106390 1026 106446
rect 1026 106390 1030 106446
rect 966 106386 1030 106390
rect 1046 106446 1110 106450
rect 1046 106390 1050 106446
rect 1050 106390 1106 106446
rect 1106 106390 1110 106446
rect 1046 106386 1110 106390
rect 1126 106446 1190 106450
rect 1126 106390 1130 106446
rect 1130 106390 1186 106446
rect 1186 106390 1190 106446
rect 1126 106386 1190 106390
rect 84886 106446 84950 106450
rect 84886 106390 84890 106446
rect 84890 106390 84946 106446
rect 84946 106390 84950 106446
rect 84886 106386 84950 106390
rect 84966 106446 85030 106450
rect 84966 106390 84970 106446
rect 84970 106390 85026 106446
rect 85026 106390 85030 106446
rect 84966 106386 85030 106390
rect 85046 106446 85110 106450
rect 85046 106390 85050 106446
rect 85050 106390 85106 106446
rect 85106 106390 85110 106446
rect 85046 106386 85110 106390
rect 85126 106446 85190 106450
rect 85126 106390 85130 106446
rect 85130 106390 85186 106446
rect 85186 106390 85190 106446
rect 85126 106386 85190 106390
rect 2886 105902 2950 105906
rect 2886 105846 2890 105902
rect 2890 105846 2946 105902
rect 2946 105846 2950 105902
rect 2886 105842 2950 105846
rect 2966 105902 3030 105906
rect 2966 105846 2970 105902
rect 2970 105846 3026 105902
rect 3026 105846 3030 105902
rect 2966 105842 3030 105846
rect 3046 105902 3110 105906
rect 3046 105846 3050 105902
rect 3050 105846 3106 105902
rect 3106 105846 3110 105902
rect 3046 105842 3110 105846
rect 3126 105902 3190 105906
rect 3126 105846 3130 105902
rect 3130 105846 3186 105902
rect 3186 105846 3190 105902
rect 3126 105842 3190 105846
rect 86886 105902 86950 105906
rect 86886 105846 86890 105902
rect 86890 105846 86946 105902
rect 86946 105846 86950 105902
rect 86886 105842 86950 105846
rect 86966 105902 87030 105906
rect 86966 105846 86970 105902
rect 86970 105846 87026 105902
rect 87026 105846 87030 105902
rect 86966 105842 87030 105846
rect 87046 105902 87110 105906
rect 87046 105846 87050 105902
rect 87050 105846 87106 105902
rect 87106 105846 87110 105902
rect 87046 105842 87110 105846
rect 87126 105902 87190 105906
rect 87126 105846 87130 105902
rect 87130 105846 87186 105902
rect 87186 105846 87190 105902
rect 87126 105842 87190 105846
rect 886 105358 950 105362
rect 886 105302 890 105358
rect 890 105302 946 105358
rect 946 105302 950 105358
rect 886 105298 950 105302
rect 966 105358 1030 105362
rect 966 105302 970 105358
rect 970 105302 1026 105358
rect 1026 105302 1030 105358
rect 966 105298 1030 105302
rect 1046 105358 1110 105362
rect 1046 105302 1050 105358
rect 1050 105302 1106 105358
rect 1106 105302 1110 105358
rect 1046 105298 1110 105302
rect 1126 105358 1190 105362
rect 1126 105302 1130 105358
rect 1130 105302 1186 105358
rect 1186 105302 1190 105358
rect 1126 105298 1190 105302
rect 84886 105358 84950 105362
rect 84886 105302 84890 105358
rect 84890 105302 84946 105358
rect 84946 105302 84950 105358
rect 84886 105298 84950 105302
rect 84966 105358 85030 105362
rect 84966 105302 84970 105358
rect 84970 105302 85026 105358
rect 85026 105302 85030 105358
rect 84966 105298 85030 105302
rect 85046 105358 85110 105362
rect 85046 105302 85050 105358
rect 85050 105302 85106 105358
rect 85106 105302 85110 105358
rect 85046 105298 85110 105302
rect 85126 105358 85190 105362
rect 85126 105302 85130 105358
rect 85130 105302 85186 105358
rect 85186 105302 85190 105358
rect 85126 105298 85190 105302
rect 2886 104814 2950 104818
rect 2886 104758 2890 104814
rect 2890 104758 2946 104814
rect 2946 104758 2950 104814
rect 2886 104754 2950 104758
rect 2966 104814 3030 104818
rect 2966 104758 2970 104814
rect 2970 104758 3026 104814
rect 3026 104758 3030 104814
rect 2966 104754 3030 104758
rect 3046 104814 3110 104818
rect 3046 104758 3050 104814
rect 3050 104758 3106 104814
rect 3106 104758 3110 104814
rect 3046 104754 3110 104758
rect 3126 104814 3190 104818
rect 3126 104758 3130 104814
rect 3130 104758 3186 104814
rect 3186 104758 3190 104814
rect 3126 104754 3190 104758
rect 86886 104814 86950 104818
rect 86886 104758 86890 104814
rect 86890 104758 86946 104814
rect 86946 104758 86950 104814
rect 86886 104754 86950 104758
rect 86966 104814 87030 104818
rect 86966 104758 86970 104814
rect 86970 104758 87026 104814
rect 87026 104758 87030 104814
rect 86966 104754 87030 104758
rect 87046 104814 87110 104818
rect 87046 104758 87050 104814
rect 87050 104758 87106 104814
rect 87106 104758 87110 104814
rect 87046 104754 87110 104758
rect 87126 104814 87190 104818
rect 87126 104758 87130 104814
rect 87130 104758 87186 104814
rect 87186 104758 87190 104814
rect 87126 104754 87190 104758
rect 886 104270 950 104274
rect 886 104214 890 104270
rect 890 104214 946 104270
rect 946 104214 950 104270
rect 886 104210 950 104214
rect 966 104270 1030 104274
rect 966 104214 970 104270
rect 970 104214 1026 104270
rect 1026 104214 1030 104270
rect 966 104210 1030 104214
rect 1046 104270 1110 104274
rect 1046 104214 1050 104270
rect 1050 104214 1106 104270
rect 1106 104214 1110 104270
rect 1046 104210 1110 104214
rect 1126 104270 1190 104274
rect 1126 104214 1130 104270
rect 1130 104214 1186 104270
rect 1186 104214 1190 104270
rect 1126 104210 1190 104214
rect 84886 104270 84950 104274
rect 84886 104214 84890 104270
rect 84890 104214 84946 104270
rect 84946 104214 84950 104270
rect 84886 104210 84950 104214
rect 84966 104270 85030 104274
rect 84966 104214 84970 104270
rect 84970 104214 85026 104270
rect 85026 104214 85030 104270
rect 84966 104210 85030 104214
rect 85046 104270 85110 104274
rect 85046 104214 85050 104270
rect 85050 104214 85106 104270
rect 85106 104214 85110 104270
rect 85046 104210 85110 104214
rect 85126 104270 85190 104274
rect 85126 104214 85130 104270
rect 85130 104214 85186 104270
rect 85186 104214 85190 104270
rect 85126 104210 85190 104214
rect 2886 103726 2950 103730
rect 2886 103670 2890 103726
rect 2890 103670 2946 103726
rect 2946 103670 2950 103726
rect 2886 103666 2950 103670
rect 2966 103726 3030 103730
rect 2966 103670 2970 103726
rect 2970 103670 3026 103726
rect 3026 103670 3030 103726
rect 2966 103666 3030 103670
rect 3046 103726 3110 103730
rect 3046 103670 3050 103726
rect 3050 103670 3106 103726
rect 3106 103670 3110 103726
rect 3046 103666 3110 103670
rect 3126 103726 3190 103730
rect 3126 103670 3130 103726
rect 3130 103670 3186 103726
rect 3186 103670 3190 103726
rect 3126 103666 3190 103670
rect 86886 103726 86950 103730
rect 86886 103670 86890 103726
rect 86890 103670 86946 103726
rect 86946 103670 86950 103726
rect 86886 103666 86950 103670
rect 86966 103726 87030 103730
rect 86966 103670 86970 103726
rect 86970 103670 87026 103726
rect 87026 103670 87030 103726
rect 86966 103666 87030 103670
rect 87046 103726 87110 103730
rect 87046 103670 87050 103726
rect 87050 103670 87106 103726
rect 87106 103670 87110 103726
rect 87046 103666 87110 103670
rect 87126 103726 87190 103730
rect 87126 103670 87130 103726
rect 87130 103670 87186 103726
rect 87186 103670 87190 103726
rect 87126 103666 87190 103670
rect 886 103182 950 103186
rect 886 103126 890 103182
rect 890 103126 946 103182
rect 946 103126 950 103182
rect 886 103122 950 103126
rect 966 103182 1030 103186
rect 966 103126 970 103182
rect 970 103126 1026 103182
rect 1026 103126 1030 103182
rect 966 103122 1030 103126
rect 1046 103182 1110 103186
rect 1046 103126 1050 103182
rect 1050 103126 1106 103182
rect 1106 103126 1110 103182
rect 1046 103122 1110 103126
rect 1126 103182 1190 103186
rect 1126 103126 1130 103182
rect 1130 103126 1186 103182
rect 1186 103126 1190 103182
rect 1126 103122 1190 103126
rect 84886 103182 84950 103186
rect 84886 103126 84890 103182
rect 84890 103126 84946 103182
rect 84946 103126 84950 103182
rect 84886 103122 84950 103126
rect 84966 103182 85030 103186
rect 84966 103126 84970 103182
rect 84970 103126 85026 103182
rect 85026 103126 85030 103182
rect 84966 103122 85030 103126
rect 85046 103182 85110 103186
rect 85046 103126 85050 103182
rect 85050 103126 85106 103182
rect 85106 103126 85110 103182
rect 85046 103122 85110 103126
rect 85126 103182 85190 103186
rect 85126 103126 85130 103182
rect 85130 103126 85186 103182
rect 85186 103126 85190 103182
rect 85126 103122 85190 103126
rect 2886 102638 2950 102642
rect 2886 102582 2890 102638
rect 2890 102582 2946 102638
rect 2946 102582 2950 102638
rect 2886 102578 2950 102582
rect 2966 102638 3030 102642
rect 2966 102582 2970 102638
rect 2970 102582 3026 102638
rect 3026 102582 3030 102638
rect 2966 102578 3030 102582
rect 3046 102638 3110 102642
rect 3046 102582 3050 102638
rect 3050 102582 3106 102638
rect 3106 102582 3110 102638
rect 3046 102578 3110 102582
rect 3126 102638 3190 102642
rect 3126 102582 3130 102638
rect 3130 102582 3186 102638
rect 3186 102582 3190 102638
rect 3126 102578 3190 102582
rect 86886 102638 86950 102642
rect 86886 102582 86890 102638
rect 86890 102582 86946 102638
rect 86946 102582 86950 102638
rect 86886 102578 86950 102582
rect 86966 102638 87030 102642
rect 86966 102582 86970 102638
rect 86970 102582 87026 102638
rect 87026 102582 87030 102638
rect 86966 102578 87030 102582
rect 87046 102638 87110 102642
rect 87046 102582 87050 102638
rect 87050 102582 87106 102638
rect 87106 102582 87110 102638
rect 87046 102578 87110 102582
rect 87126 102638 87190 102642
rect 87126 102582 87130 102638
rect 87130 102582 87186 102638
rect 87186 102582 87190 102638
rect 87126 102578 87190 102582
rect 886 102094 950 102098
rect 886 102038 890 102094
rect 890 102038 946 102094
rect 946 102038 950 102094
rect 886 102034 950 102038
rect 966 102094 1030 102098
rect 966 102038 970 102094
rect 970 102038 1026 102094
rect 1026 102038 1030 102094
rect 966 102034 1030 102038
rect 1046 102094 1110 102098
rect 1046 102038 1050 102094
rect 1050 102038 1106 102094
rect 1106 102038 1110 102094
rect 1046 102034 1110 102038
rect 1126 102094 1190 102098
rect 1126 102038 1130 102094
rect 1130 102038 1186 102094
rect 1186 102038 1190 102094
rect 1126 102034 1190 102038
rect 84886 102094 84950 102098
rect 84886 102038 84890 102094
rect 84890 102038 84946 102094
rect 84946 102038 84950 102094
rect 84886 102034 84950 102038
rect 84966 102094 85030 102098
rect 84966 102038 84970 102094
rect 84970 102038 85026 102094
rect 85026 102038 85030 102094
rect 84966 102034 85030 102038
rect 85046 102094 85110 102098
rect 85046 102038 85050 102094
rect 85050 102038 85106 102094
rect 85106 102038 85110 102094
rect 85046 102034 85110 102038
rect 85126 102094 85190 102098
rect 85126 102038 85130 102094
rect 85130 102038 85186 102094
rect 85186 102038 85190 102094
rect 85126 102034 85190 102038
rect 2886 101550 2950 101554
rect 2886 101494 2890 101550
rect 2890 101494 2946 101550
rect 2946 101494 2950 101550
rect 2886 101490 2950 101494
rect 2966 101550 3030 101554
rect 2966 101494 2970 101550
rect 2970 101494 3026 101550
rect 3026 101494 3030 101550
rect 2966 101490 3030 101494
rect 3046 101550 3110 101554
rect 3046 101494 3050 101550
rect 3050 101494 3106 101550
rect 3106 101494 3110 101550
rect 3046 101490 3110 101494
rect 3126 101550 3190 101554
rect 3126 101494 3130 101550
rect 3130 101494 3186 101550
rect 3186 101494 3190 101550
rect 3126 101490 3190 101494
rect 86886 101550 86950 101554
rect 86886 101494 86890 101550
rect 86890 101494 86946 101550
rect 86946 101494 86950 101550
rect 86886 101490 86950 101494
rect 86966 101550 87030 101554
rect 86966 101494 86970 101550
rect 86970 101494 87026 101550
rect 87026 101494 87030 101550
rect 86966 101490 87030 101494
rect 87046 101550 87110 101554
rect 87046 101494 87050 101550
rect 87050 101494 87106 101550
rect 87106 101494 87110 101550
rect 87046 101490 87110 101494
rect 87126 101550 87190 101554
rect 87126 101494 87130 101550
rect 87130 101494 87186 101550
rect 87186 101494 87190 101550
rect 87126 101490 87190 101494
rect 886 101006 950 101010
rect 886 100950 890 101006
rect 890 100950 946 101006
rect 946 100950 950 101006
rect 886 100946 950 100950
rect 966 101006 1030 101010
rect 966 100950 970 101006
rect 970 100950 1026 101006
rect 1026 100950 1030 101006
rect 966 100946 1030 100950
rect 1046 101006 1110 101010
rect 1046 100950 1050 101006
rect 1050 100950 1106 101006
rect 1106 100950 1110 101006
rect 1046 100946 1110 100950
rect 1126 101006 1190 101010
rect 1126 100950 1130 101006
rect 1130 100950 1186 101006
rect 1186 100950 1190 101006
rect 1126 100946 1190 100950
rect 84886 101006 84950 101010
rect 84886 100950 84890 101006
rect 84890 100950 84946 101006
rect 84946 100950 84950 101006
rect 84886 100946 84950 100950
rect 84966 101006 85030 101010
rect 84966 100950 84970 101006
rect 84970 100950 85026 101006
rect 85026 100950 85030 101006
rect 84966 100946 85030 100950
rect 85046 101006 85110 101010
rect 85046 100950 85050 101006
rect 85050 100950 85106 101006
rect 85106 100950 85110 101006
rect 85046 100946 85110 100950
rect 85126 101006 85190 101010
rect 85126 100950 85130 101006
rect 85130 100950 85186 101006
rect 85186 100950 85190 101006
rect 85126 100946 85190 100950
rect 2886 100462 2950 100466
rect 2886 100406 2890 100462
rect 2890 100406 2946 100462
rect 2946 100406 2950 100462
rect 2886 100402 2950 100406
rect 2966 100462 3030 100466
rect 2966 100406 2970 100462
rect 2970 100406 3026 100462
rect 3026 100406 3030 100462
rect 2966 100402 3030 100406
rect 3046 100462 3110 100466
rect 3046 100406 3050 100462
rect 3050 100406 3106 100462
rect 3106 100406 3110 100462
rect 3046 100402 3110 100406
rect 3126 100462 3190 100466
rect 3126 100406 3130 100462
rect 3130 100406 3186 100462
rect 3186 100406 3190 100462
rect 3126 100402 3190 100406
rect 86886 100462 86950 100466
rect 86886 100406 86890 100462
rect 86890 100406 86946 100462
rect 86946 100406 86950 100462
rect 86886 100402 86950 100406
rect 86966 100462 87030 100466
rect 86966 100406 86970 100462
rect 86970 100406 87026 100462
rect 87026 100406 87030 100462
rect 86966 100402 87030 100406
rect 87046 100462 87110 100466
rect 87046 100406 87050 100462
rect 87050 100406 87106 100462
rect 87106 100406 87110 100462
rect 87046 100402 87110 100406
rect 87126 100462 87190 100466
rect 87126 100406 87130 100462
rect 87130 100406 87186 100462
rect 87186 100406 87190 100462
rect 87126 100402 87190 100406
rect 886 99918 950 99922
rect 886 99862 890 99918
rect 890 99862 946 99918
rect 946 99862 950 99918
rect 886 99858 950 99862
rect 966 99918 1030 99922
rect 966 99862 970 99918
rect 970 99862 1026 99918
rect 1026 99862 1030 99918
rect 966 99858 1030 99862
rect 1046 99918 1110 99922
rect 1046 99862 1050 99918
rect 1050 99862 1106 99918
rect 1106 99862 1110 99918
rect 1046 99858 1110 99862
rect 1126 99918 1190 99922
rect 1126 99862 1130 99918
rect 1130 99862 1186 99918
rect 1186 99862 1190 99918
rect 1126 99858 1190 99862
rect 84886 99918 84950 99922
rect 84886 99862 84890 99918
rect 84890 99862 84946 99918
rect 84946 99862 84950 99918
rect 84886 99858 84950 99862
rect 84966 99918 85030 99922
rect 84966 99862 84970 99918
rect 84970 99862 85026 99918
rect 85026 99862 85030 99918
rect 84966 99858 85030 99862
rect 85046 99918 85110 99922
rect 85046 99862 85050 99918
rect 85050 99862 85106 99918
rect 85106 99862 85110 99918
rect 85046 99858 85110 99862
rect 85126 99918 85190 99922
rect 85126 99862 85130 99918
rect 85130 99862 85186 99918
rect 85186 99862 85190 99918
rect 85126 99858 85190 99862
rect 2886 99374 2950 99378
rect 2886 99318 2890 99374
rect 2890 99318 2946 99374
rect 2946 99318 2950 99374
rect 2886 99314 2950 99318
rect 2966 99374 3030 99378
rect 2966 99318 2970 99374
rect 2970 99318 3026 99374
rect 3026 99318 3030 99374
rect 2966 99314 3030 99318
rect 3046 99374 3110 99378
rect 3046 99318 3050 99374
rect 3050 99318 3106 99374
rect 3106 99318 3110 99374
rect 3046 99314 3110 99318
rect 3126 99374 3190 99378
rect 3126 99318 3130 99374
rect 3130 99318 3186 99374
rect 3186 99318 3190 99374
rect 3126 99314 3190 99318
rect 86886 99374 86950 99378
rect 86886 99318 86890 99374
rect 86890 99318 86946 99374
rect 86946 99318 86950 99374
rect 86886 99314 86950 99318
rect 86966 99374 87030 99378
rect 86966 99318 86970 99374
rect 86970 99318 87026 99374
rect 87026 99318 87030 99374
rect 86966 99314 87030 99318
rect 87046 99374 87110 99378
rect 87046 99318 87050 99374
rect 87050 99318 87106 99374
rect 87106 99318 87110 99374
rect 87046 99314 87110 99318
rect 87126 99374 87190 99378
rect 87126 99318 87130 99374
rect 87130 99318 87186 99374
rect 87186 99318 87190 99374
rect 87126 99314 87190 99318
rect 886 98830 950 98834
rect 886 98774 890 98830
rect 890 98774 946 98830
rect 946 98774 950 98830
rect 886 98770 950 98774
rect 966 98830 1030 98834
rect 966 98774 970 98830
rect 970 98774 1026 98830
rect 1026 98774 1030 98830
rect 966 98770 1030 98774
rect 1046 98830 1110 98834
rect 1046 98774 1050 98830
rect 1050 98774 1106 98830
rect 1106 98774 1110 98830
rect 1046 98770 1110 98774
rect 1126 98830 1190 98834
rect 1126 98774 1130 98830
rect 1130 98774 1186 98830
rect 1186 98774 1190 98830
rect 1126 98770 1190 98774
rect 84886 98830 84950 98834
rect 84886 98774 84890 98830
rect 84890 98774 84946 98830
rect 84946 98774 84950 98830
rect 84886 98770 84950 98774
rect 84966 98830 85030 98834
rect 84966 98774 84970 98830
rect 84970 98774 85026 98830
rect 85026 98774 85030 98830
rect 84966 98770 85030 98774
rect 85046 98830 85110 98834
rect 85046 98774 85050 98830
rect 85050 98774 85106 98830
rect 85106 98774 85110 98830
rect 85046 98770 85110 98774
rect 85126 98830 85190 98834
rect 85126 98774 85130 98830
rect 85130 98774 85186 98830
rect 85186 98774 85190 98830
rect 85126 98770 85190 98774
rect 4330 98294 4394 98358
rect 2886 98286 2950 98290
rect 2886 98230 2890 98286
rect 2890 98230 2946 98286
rect 2946 98230 2950 98286
rect 2886 98226 2950 98230
rect 2966 98286 3030 98290
rect 2966 98230 2970 98286
rect 2970 98230 3026 98286
rect 3026 98230 3030 98286
rect 2966 98226 3030 98230
rect 3046 98286 3110 98290
rect 3046 98230 3050 98286
rect 3050 98230 3106 98286
rect 3106 98230 3110 98286
rect 3046 98226 3110 98230
rect 3126 98286 3190 98290
rect 3126 98230 3130 98286
rect 3130 98230 3186 98286
rect 3186 98230 3190 98286
rect 3126 98226 3190 98230
rect 86886 98286 86950 98290
rect 86886 98230 86890 98286
rect 86890 98230 86946 98286
rect 86946 98230 86950 98286
rect 86886 98226 86950 98230
rect 86966 98286 87030 98290
rect 86966 98230 86970 98286
rect 86970 98230 87026 98286
rect 87026 98230 87030 98286
rect 86966 98226 87030 98230
rect 87046 98286 87110 98290
rect 87046 98230 87050 98286
rect 87050 98230 87106 98286
rect 87106 98230 87110 98286
rect 87046 98226 87110 98230
rect 87126 98286 87190 98290
rect 87126 98230 87130 98286
rect 87130 98230 87186 98286
rect 87186 98230 87190 98286
rect 87126 98226 87190 98230
rect 3778 98158 3842 98222
rect 886 97742 950 97746
rect 886 97686 890 97742
rect 890 97686 946 97742
rect 946 97686 950 97742
rect 886 97682 950 97686
rect 966 97742 1030 97746
rect 966 97686 970 97742
rect 970 97686 1026 97742
rect 1026 97686 1030 97742
rect 966 97682 1030 97686
rect 1046 97742 1110 97746
rect 1046 97686 1050 97742
rect 1050 97686 1106 97742
rect 1106 97686 1110 97742
rect 1046 97682 1110 97686
rect 1126 97742 1190 97746
rect 1126 97686 1130 97742
rect 1130 97686 1186 97742
rect 1186 97686 1190 97742
rect 1126 97682 1190 97686
rect 84886 97742 84950 97746
rect 84886 97686 84890 97742
rect 84890 97686 84946 97742
rect 84946 97686 84950 97742
rect 84886 97682 84950 97686
rect 84966 97742 85030 97746
rect 84966 97686 84970 97742
rect 84970 97686 85026 97742
rect 85026 97686 85030 97742
rect 84966 97682 85030 97686
rect 85046 97742 85110 97746
rect 85046 97686 85050 97742
rect 85050 97686 85106 97742
rect 85106 97686 85110 97742
rect 85046 97682 85110 97686
rect 85126 97742 85190 97746
rect 85126 97686 85130 97742
rect 85130 97686 85186 97742
rect 85186 97686 85190 97742
rect 85126 97682 85190 97686
rect 83634 97614 83698 97678
rect 2886 97198 2950 97202
rect 2886 97142 2890 97198
rect 2890 97142 2946 97198
rect 2946 97142 2950 97198
rect 2886 97138 2950 97142
rect 2966 97198 3030 97202
rect 2966 97142 2970 97198
rect 2970 97142 3026 97198
rect 3026 97142 3030 97198
rect 2966 97138 3030 97142
rect 3046 97198 3110 97202
rect 3046 97142 3050 97198
rect 3050 97142 3106 97198
rect 3106 97142 3110 97198
rect 3046 97138 3110 97142
rect 3126 97198 3190 97202
rect 3126 97142 3130 97198
rect 3130 97142 3186 97198
rect 3186 97142 3190 97198
rect 3126 97138 3190 97142
rect 86886 97198 86950 97202
rect 86886 97142 86890 97198
rect 86890 97142 86946 97198
rect 86946 97142 86950 97198
rect 86886 97138 86950 97142
rect 86966 97198 87030 97202
rect 86966 97142 86970 97198
rect 86970 97142 87026 97198
rect 87026 97142 87030 97198
rect 86966 97138 87030 97142
rect 87046 97198 87110 97202
rect 87046 97142 87050 97198
rect 87050 97142 87106 97198
rect 87106 97142 87110 97198
rect 87046 97138 87110 97142
rect 87126 97198 87190 97202
rect 87126 97142 87130 97198
rect 87130 97142 87186 97198
rect 87186 97142 87190 97198
rect 87126 97138 87190 97142
rect 84186 97130 84250 97134
rect 84186 97074 84200 97130
rect 84200 97074 84250 97130
rect 39106 96934 39170 96998
rect 14634 96858 14698 96862
rect 14634 96802 14648 96858
rect 14648 96802 14698 96858
rect 14634 96798 14698 96802
rect 84186 97070 84250 97074
rect 82346 96934 82410 96998
rect 33402 96798 33466 96862
rect 45362 96798 45426 96862
rect 3410 96662 3474 96726
rect 15738 96662 15802 96726
rect 21994 96662 22058 96726
rect 25306 96722 25370 96726
rect 25306 96666 25320 96722
rect 25320 96666 25370 96722
rect 25306 96662 25370 96666
rect 28986 96722 29050 96726
rect 28986 96666 29000 96722
rect 29000 96666 29050 96722
rect 28986 96662 29050 96666
rect 29977 96722 30041 96726
rect 29977 96666 30012 96722
rect 30012 96666 30041 96722
rect 29977 96662 30041 96666
rect 34969 96722 35033 96726
rect 34969 96666 35016 96722
rect 35016 96666 35033 96722
rect 34969 96662 35033 96666
rect 36898 96722 36962 96726
rect 36898 96666 36912 96722
rect 36912 96666 36962 96722
rect 36898 96662 36962 96666
rect 886 96654 950 96658
rect 886 96598 890 96654
rect 890 96598 946 96654
rect 946 96598 950 96654
rect 886 96594 950 96598
rect 966 96654 1030 96658
rect 966 96598 970 96654
rect 970 96598 1026 96654
rect 1026 96598 1030 96654
rect 966 96594 1030 96598
rect 1046 96654 1110 96658
rect 1046 96598 1050 96654
rect 1050 96598 1106 96654
rect 1106 96598 1110 96654
rect 1046 96594 1110 96598
rect 1126 96654 1190 96658
rect 1126 96598 1130 96654
rect 1130 96598 1186 96654
rect 1186 96598 1190 96654
rect 1126 96594 1190 96598
rect 5250 96526 5314 96590
rect 44258 96662 44322 96726
rect 48858 96722 48922 96726
rect 48858 96666 48908 96722
rect 48908 96666 48922 96722
rect 48858 96662 48922 96666
rect 50146 96722 50210 96726
rect 83450 96858 83514 96862
rect 83450 96802 83500 96858
rect 83500 96802 83514 96858
rect 83450 96798 83514 96802
rect 84738 96798 84802 96862
rect 50146 96666 50196 96722
rect 50196 96666 50210 96722
rect 50146 96662 50210 96666
rect 82162 96662 82226 96726
rect 84886 96654 84950 96658
rect 84886 96598 84890 96654
rect 84890 96598 84946 96654
rect 84946 96598 84950 96654
rect 84886 96594 84950 96598
rect 84966 96654 85030 96658
rect 84966 96598 84970 96654
rect 84970 96598 85026 96654
rect 85026 96598 85030 96654
rect 84966 96594 85030 96598
rect 85046 96654 85110 96658
rect 85046 96598 85050 96654
rect 85050 96598 85106 96654
rect 85106 96598 85110 96654
rect 85046 96594 85110 96598
rect 85126 96654 85190 96658
rect 85126 96598 85130 96654
rect 85130 96598 85186 96654
rect 85186 96598 85190 96654
rect 85126 96594 85190 96598
rect 4514 96390 4578 96454
rect 3778 96254 3842 96318
rect 40394 96390 40458 96454
rect 82530 96526 82594 96590
rect 83818 96314 83882 96318
rect 83818 96258 83832 96314
rect 83832 96258 83882 96314
rect 83818 96254 83882 96258
rect 38186 96178 38250 96182
rect 38186 96122 38200 96178
rect 38200 96122 38250 96178
rect 38186 96118 38250 96122
rect 47018 96118 47082 96182
rect 47570 96178 47634 96182
rect 47570 96122 47620 96178
rect 47620 96122 47634 96178
rect 47570 96118 47634 96122
rect 2886 96110 2950 96114
rect 2886 96054 2890 96110
rect 2890 96054 2946 96110
rect 2946 96054 2950 96110
rect 2886 96050 2950 96054
rect 2966 96110 3030 96114
rect 2966 96054 2970 96110
rect 2970 96054 3026 96110
rect 3026 96054 3030 96110
rect 2966 96050 3030 96054
rect 3046 96110 3110 96114
rect 3046 96054 3050 96110
rect 3050 96054 3106 96110
rect 3106 96054 3110 96110
rect 3046 96050 3110 96054
rect 3126 96110 3190 96114
rect 3126 96054 3130 96110
rect 3130 96054 3186 96110
rect 3186 96054 3190 96110
rect 3126 96050 3190 96054
rect 86886 96110 86950 96114
rect 86886 96054 86890 96110
rect 86890 96054 86946 96110
rect 86946 96054 86950 96110
rect 86886 96050 86950 96054
rect 86966 96110 87030 96114
rect 86966 96054 86970 96110
rect 86970 96054 87026 96110
rect 87026 96054 87030 96110
rect 86966 96050 87030 96054
rect 87046 96110 87110 96114
rect 87046 96054 87050 96110
rect 87050 96054 87106 96110
rect 87106 96054 87110 96110
rect 87046 96050 87110 96054
rect 87126 96110 87190 96114
rect 87126 96054 87130 96110
rect 87130 96054 87186 96110
rect 87186 96054 87190 96110
rect 87126 96050 87190 96054
rect 18498 95982 18562 96046
rect 23414 96042 23478 96046
rect 23414 95986 23424 96042
rect 23424 95986 23478 96042
rect 23414 95982 23478 95986
rect 32666 95982 32730 96046
rect 14070 95906 14134 95910
rect 14070 95850 14096 95906
rect 14096 95850 14134 95906
rect 14070 95846 14134 95850
rect 17574 95846 17638 95910
rect 24018 95906 24082 95910
rect 24018 95850 24032 95906
rect 24032 95850 24082 95906
rect 24018 95846 24082 95850
rect 31746 95846 31810 95910
rect 19786 95770 19850 95774
rect 19786 95714 19836 95770
rect 19836 95714 19850 95770
rect 19786 95710 19850 95714
rect 29354 95710 29418 95774
rect 27146 95634 27210 95638
rect 27146 95578 27196 95634
rect 27196 95578 27210 95634
rect 27146 95574 27210 95578
rect 51434 95634 51498 95638
rect 51434 95578 51484 95634
rect 51484 95578 51498 95634
rect 51434 95574 51498 95578
rect 886 95566 950 95570
rect 886 95510 890 95566
rect 890 95510 946 95566
rect 946 95510 950 95566
rect 886 95506 950 95510
rect 966 95566 1030 95570
rect 966 95510 970 95566
rect 970 95510 1026 95566
rect 1026 95510 1030 95566
rect 966 95506 1030 95510
rect 1046 95566 1110 95570
rect 1046 95510 1050 95566
rect 1050 95510 1106 95566
rect 1106 95510 1110 95566
rect 1046 95506 1110 95510
rect 1126 95566 1190 95570
rect 1126 95510 1130 95566
rect 1130 95510 1186 95566
rect 1186 95510 1190 95566
rect 1126 95506 1190 95510
rect 84886 95566 84950 95570
rect 84886 95510 84890 95566
rect 84890 95510 84946 95566
rect 84946 95510 84950 95566
rect 84886 95506 84950 95510
rect 84966 95566 85030 95570
rect 84966 95510 84970 95566
rect 84970 95510 85026 95566
rect 85026 95510 85030 95566
rect 84966 95506 85030 95510
rect 85046 95566 85110 95570
rect 85046 95510 85050 95566
rect 85050 95510 85106 95566
rect 85106 95510 85110 95566
rect 85046 95506 85110 95510
rect 85126 95566 85190 95570
rect 85126 95510 85130 95566
rect 85130 95510 85186 95566
rect 85186 95510 85190 95566
rect 85126 95506 85190 95510
rect 24386 95226 24450 95230
rect 24386 95170 24436 95226
rect 24436 95170 24450 95226
rect 24386 95166 24450 95170
rect 25674 95226 25738 95230
rect 25674 95170 25724 95226
rect 25724 95170 25738 95226
rect 25674 95166 25738 95170
rect 26594 95226 26658 95230
rect 26594 95170 26644 95226
rect 26644 95170 26658 95226
rect 26594 95166 26658 95170
rect 34322 95166 34386 95230
rect 35610 95226 35674 95230
rect 35610 95170 35660 95226
rect 35660 95170 35674 95226
rect 35610 95166 35674 95170
rect 36162 95226 36226 95230
rect 36162 95170 36212 95226
rect 36212 95170 36226 95226
rect 36162 95166 36226 95170
rect 37450 95226 37514 95230
rect 37450 95170 37500 95226
rect 37500 95170 37514 95226
rect 37450 95166 37514 95170
rect 38554 95226 38618 95230
rect 38554 95170 38604 95226
rect 38604 95170 38618 95226
rect 38554 95166 38618 95170
rect 41866 95226 41930 95230
rect 41866 95170 41880 95226
rect 41880 95170 41930 95226
rect 41866 95166 41930 95170
rect 43706 95226 43770 95230
rect 43706 95170 43756 95226
rect 43756 95170 43770 95226
rect 43706 95166 43770 95170
rect 44442 95226 44506 95230
rect 44442 95170 44492 95226
rect 44492 95170 44506 95226
rect 44442 95166 44506 95170
rect 46466 95226 46530 95230
rect 46466 95170 46516 95226
rect 46516 95170 46530 95226
rect 46466 95166 46530 95170
rect 47754 95226 47818 95230
rect 47754 95170 47804 95226
rect 47804 95170 47818 95226
rect 47754 95166 47818 95170
rect 48674 95226 48738 95230
rect 48674 95170 48724 95226
rect 48724 95170 48738 95226
rect 48674 95166 48738 95170
rect 50146 95226 50210 95230
rect 50146 95170 50196 95226
rect 50196 95170 50210 95226
rect 50146 95166 50210 95170
rect 51434 95166 51498 95230
rect 56586 95226 56650 95230
rect 56586 95170 56636 95226
rect 56636 95170 56650 95226
rect 56586 95166 56650 95170
rect 57874 95226 57938 95230
rect 57874 95170 57924 95226
rect 57924 95170 57938 95226
rect 57874 95166 57938 95170
rect 59346 95226 59410 95230
rect 59346 95170 59396 95226
rect 59396 95170 59410 95226
rect 59346 95166 59410 95170
rect 61738 95226 61802 95230
rect 61738 95170 61788 95226
rect 61788 95170 61802 95226
rect 61738 95166 61802 95170
rect 62658 95166 62722 95230
rect 4330 95090 4394 95094
rect 4330 95034 4344 95090
rect 4344 95034 4394 95090
rect 4330 95030 4394 95034
rect 8194 95090 8258 95094
rect 8194 95034 8208 95090
rect 8208 95034 8258 95090
rect 8194 95030 8258 95034
rect 12242 95030 12306 95094
rect 31378 95030 31442 95094
rect 36346 95090 36410 95094
rect 36346 95034 36360 95090
rect 36360 95034 36410 95090
rect 36346 95030 36410 95034
rect 36714 95030 36778 95094
rect 38738 95090 38802 95094
rect 38738 95034 38788 95090
rect 38788 95034 38802 95090
rect 38738 95030 38802 95034
rect 43338 95030 43402 95094
rect 47938 95030 48002 95094
rect 50330 95090 50394 95094
rect 50330 95034 50380 95090
rect 50380 95034 50394 95090
rect 50330 95030 50394 95034
rect 54194 95090 54258 95094
rect 54194 95034 54244 95090
rect 54244 95034 54258 95090
rect 54194 95030 54258 95034
rect 2886 95022 2950 95026
rect 2886 94966 2890 95022
rect 2890 94966 2946 95022
rect 2946 94966 2950 95022
rect 2886 94962 2950 94966
rect 2966 95022 3030 95026
rect 2966 94966 2970 95022
rect 2970 94966 3026 95022
rect 3026 94966 3030 95022
rect 2966 94962 3030 94966
rect 3046 95022 3110 95026
rect 3046 94966 3050 95022
rect 3050 94966 3106 95022
rect 3106 94966 3110 95022
rect 3046 94962 3110 94966
rect 3126 95022 3190 95026
rect 3126 94966 3130 95022
rect 3130 94966 3186 95022
rect 3186 94966 3190 95022
rect 3126 94962 3190 94966
rect 86886 95022 86950 95026
rect 86886 94966 86890 95022
rect 86890 94966 86946 95022
rect 86946 94966 86950 95022
rect 86886 94962 86950 94966
rect 86966 95022 87030 95026
rect 86966 94966 86970 95022
rect 86970 94966 87026 95022
rect 87026 94966 87030 95022
rect 86966 94962 87030 94966
rect 87046 95022 87110 95026
rect 87046 94966 87050 95022
rect 87050 94966 87106 95022
rect 87106 94966 87110 95022
rect 87046 94962 87110 94966
rect 87126 95022 87190 95026
rect 87126 94966 87130 95022
rect 87130 94966 87186 95022
rect 87186 94966 87190 95022
rect 87126 94962 87190 94966
rect 11322 94894 11386 94958
rect 22730 94894 22794 94958
rect 25306 94894 25370 94958
rect 18130 94818 18194 94822
rect 18130 94762 18180 94818
rect 18180 94762 18194 94818
rect 18130 94758 18194 94762
rect 19970 94758 20034 94822
rect 21442 94758 21506 94822
rect 26410 94758 26474 94822
rect 49778 94758 49842 94822
rect 52354 94758 52418 94822
rect 27514 94622 27578 94686
rect 32482 94682 32546 94686
rect 32482 94626 32496 94682
rect 32496 94626 32546 94682
rect 32482 94622 32546 94626
rect 48490 94622 48554 94686
rect 52722 94622 52786 94686
rect 83818 94622 83882 94686
rect 40026 94546 40090 94550
rect 40026 94490 40076 94546
rect 40076 94490 40090 94546
rect 40026 94486 40090 94490
rect 41498 94546 41562 94550
rect 41498 94490 41512 94546
rect 41512 94490 41562 94546
rect 41498 94486 41562 94490
rect 42602 94546 42666 94550
rect 42602 94490 42652 94546
rect 42652 94490 42666 94546
rect 42602 94486 42666 94490
rect 53826 94486 53890 94550
rect 886 94478 950 94482
rect 886 94422 890 94478
rect 890 94422 946 94478
rect 946 94422 950 94478
rect 886 94418 950 94422
rect 966 94478 1030 94482
rect 966 94422 970 94478
rect 970 94422 1026 94478
rect 1026 94422 1030 94478
rect 966 94418 1030 94422
rect 1046 94478 1110 94482
rect 1046 94422 1050 94478
rect 1050 94422 1106 94478
rect 1106 94422 1110 94478
rect 1046 94418 1110 94422
rect 1126 94478 1190 94482
rect 1126 94422 1130 94478
rect 1130 94422 1186 94478
rect 1186 94422 1190 94478
rect 1126 94418 1190 94422
rect 84886 94478 84950 94482
rect 84886 94422 84890 94478
rect 84890 94422 84946 94478
rect 84946 94422 84950 94478
rect 84886 94418 84950 94422
rect 84966 94478 85030 94482
rect 84966 94422 84970 94478
rect 84970 94422 85026 94478
rect 85026 94422 85030 94478
rect 84966 94418 85030 94422
rect 85046 94478 85110 94482
rect 85046 94422 85050 94478
rect 85050 94422 85106 94478
rect 85106 94422 85110 94478
rect 85046 94418 85110 94422
rect 85126 94478 85190 94482
rect 85126 94422 85130 94478
rect 85130 94422 85186 94478
rect 85186 94422 85190 94478
rect 85126 94418 85190 94422
rect 18682 94350 18746 94414
rect 29722 94410 29786 94414
rect 29722 94354 29772 94410
rect 29772 94354 29786 94410
rect 29722 94350 29786 94354
rect 41314 94410 41378 94414
rect 41314 94354 41328 94410
rect 41328 94354 41378 94410
rect 41314 94350 41378 94354
rect 41682 94410 41746 94414
rect 41682 94354 41732 94410
rect 41732 94354 41746 94410
rect 41682 94350 41746 94354
rect 43890 94410 43954 94414
rect 43890 94354 43940 94410
rect 43940 94354 43954 94410
rect 43890 94350 43954 94354
rect 44626 94350 44690 94414
rect 51618 94410 51682 94414
rect 51618 94354 51668 94410
rect 51668 94354 51682 94410
rect 51618 94350 51682 94354
rect 69834 94350 69898 94414
rect 21810 94214 21874 94278
rect 23834 94078 23898 94142
rect 28250 94078 28314 94142
rect 30642 93942 30706 94006
rect 45730 93942 45794 94006
rect 52906 93942 52970 94006
rect 2886 93934 2950 93938
rect 2886 93878 2890 93934
rect 2890 93878 2946 93934
rect 2946 93878 2950 93934
rect 2886 93874 2950 93878
rect 2966 93934 3030 93938
rect 2966 93878 2970 93934
rect 2970 93878 3026 93934
rect 3026 93878 3030 93934
rect 2966 93874 3030 93878
rect 3046 93934 3110 93938
rect 3046 93878 3050 93934
rect 3050 93878 3106 93934
rect 3106 93878 3110 93934
rect 3046 93874 3110 93878
rect 3126 93934 3190 93938
rect 3126 93878 3130 93934
rect 3130 93878 3186 93934
rect 3186 93878 3190 93934
rect 3126 93874 3190 93878
rect 30642 93866 30706 93870
rect 30642 93810 30692 93866
rect 30692 93810 30706 93866
rect 30642 93806 30706 93810
rect 32298 93866 32362 93870
rect 32298 93810 32348 93866
rect 32348 93810 32362 93866
rect 32298 93806 32362 93810
rect 33402 93806 33466 93870
rect 34690 93806 34754 93870
rect 35794 93806 35858 93870
rect 38002 93806 38066 93870
rect 39961 93806 40025 93870
rect 53689 93866 53753 93870
rect 53689 93810 53692 93866
rect 53692 93810 53748 93866
rect 53748 93810 53753 93866
rect 53689 93806 53753 93810
rect 69834 93806 69898 93870
rect 82714 93942 82778 94006
rect 86886 93934 86950 93938
rect 86886 93878 86890 93934
rect 86890 93878 86946 93934
rect 86946 93878 86950 93934
rect 86886 93874 86950 93878
rect 86966 93934 87030 93938
rect 86966 93878 86970 93934
rect 86970 93878 87026 93934
rect 87026 93878 87030 93934
rect 86966 93874 87030 93878
rect 87046 93934 87110 93938
rect 87046 93878 87050 93934
rect 87050 93878 87106 93934
rect 87106 93878 87110 93934
rect 87046 93874 87110 93878
rect 87126 93934 87190 93938
rect 87126 93878 87130 93934
rect 87130 93878 87186 93934
rect 87186 93878 87190 93934
rect 87126 93874 87190 93878
rect 78482 93866 78546 93870
rect 78482 93810 78496 93866
rect 78496 93810 78546 93866
rect 78482 93806 78546 93810
rect 27481 93534 27545 93598
rect 886 93390 950 93394
rect 886 93334 890 93390
rect 890 93334 946 93390
rect 946 93334 950 93390
rect 886 93330 950 93334
rect 966 93390 1030 93394
rect 966 93334 970 93390
rect 970 93334 1026 93390
rect 1026 93334 1030 93390
rect 966 93330 1030 93334
rect 1046 93390 1110 93394
rect 1046 93334 1050 93390
rect 1050 93334 1106 93390
rect 1106 93334 1110 93390
rect 1046 93330 1110 93334
rect 1126 93390 1190 93394
rect 1126 93334 1130 93390
rect 1130 93334 1186 93390
rect 1186 93334 1190 93390
rect 1126 93330 1190 93334
rect 84886 93390 84950 93394
rect 84886 93334 84890 93390
rect 84890 93334 84946 93390
rect 84946 93334 84950 93390
rect 84886 93330 84950 93334
rect 84966 93390 85030 93394
rect 84966 93334 84970 93390
rect 84970 93334 85026 93390
rect 85026 93334 85030 93390
rect 84966 93330 85030 93334
rect 85046 93390 85110 93394
rect 85046 93334 85050 93390
rect 85050 93334 85106 93390
rect 85106 93334 85110 93390
rect 85046 93330 85110 93334
rect 85126 93390 85190 93394
rect 85126 93334 85130 93390
rect 85130 93334 85186 93390
rect 85186 93334 85190 93390
rect 85126 93330 85190 93334
rect 25858 93126 25922 93190
rect 2886 92846 2950 92850
rect 2886 92790 2890 92846
rect 2890 92790 2946 92846
rect 2946 92790 2950 92846
rect 2886 92786 2950 92790
rect 2966 92846 3030 92850
rect 2966 92790 2970 92846
rect 2970 92790 3026 92846
rect 3026 92790 3030 92846
rect 2966 92786 3030 92790
rect 3046 92846 3110 92850
rect 3046 92790 3050 92846
rect 3050 92790 3106 92846
rect 3106 92790 3110 92846
rect 3046 92786 3110 92790
rect 3126 92846 3190 92850
rect 3126 92790 3130 92846
rect 3130 92790 3186 92846
rect 3186 92790 3190 92846
rect 3126 92786 3190 92790
rect 86886 92846 86950 92850
rect 86886 92790 86890 92846
rect 86890 92790 86946 92846
rect 86946 92790 86950 92846
rect 86886 92786 86950 92790
rect 86966 92846 87030 92850
rect 86966 92790 86970 92846
rect 86970 92790 87026 92846
rect 87026 92790 87030 92846
rect 86966 92786 87030 92790
rect 87046 92846 87110 92850
rect 87046 92790 87050 92846
rect 87050 92790 87106 92846
rect 87106 92790 87110 92846
rect 87046 92786 87110 92790
rect 87126 92846 87190 92850
rect 87126 92790 87130 92846
rect 87130 92790 87186 92846
rect 87186 92790 87190 92846
rect 87126 92786 87190 92790
rect 55298 92642 55362 92646
rect 55298 92586 55348 92642
rect 55348 92586 55362 92642
rect 55298 92582 55362 92586
rect 60450 92642 60514 92646
rect 60450 92586 60500 92642
rect 60500 92586 60514 92642
rect 60450 92582 60514 92586
rect 73698 92642 73762 92646
rect 73698 92586 73748 92642
rect 73748 92586 73762 92642
rect 73698 92582 73762 92586
rect 886 92302 950 92306
rect 886 92246 890 92302
rect 890 92246 946 92302
rect 946 92246 950 92302
rect 886 92242 950 92246
rect 966 92302 1030 92306
rect 966 92246 970 92302
rect 970 92246 1026 92302
rect 1026 92246 1030 92302
rect 966 92242 1030 92246
rect 1046 92302 1110 92306
rect 1046 92246 1050 92302
rect 1050 92246 1106 92302
rect 1106 92246 1110 92302
rect 1046 92242 1110 92246
rect 1126 92302 1190 92306
rect 1126 92246 1130 92302
rect 1130 92246 1186 92302
rect 1186 92246 1190 92302
rect 1126 92242 1190 92246
rect 84886 92302 84950 92306
rect 84886 92246 84890 92302
rect 84890 92246 84946 92302
rect 84946 92246 84950 92302
rect 84886 92242 84950 92246
rect 84966 92302 85030 92306
rect 84966 92246 84970 92302
rect 84970 92246 85026 92302
rect 85026 92246 85030 92302
rect 84966 92242 85030 92246
rect 85046 92302 85110 92306
rect 85046 92246 85050 92302
rect 85050 92246 85106 92302
rect 85106 92246 85110 92302
rect 85046 92242 85110 92246
rect 85126 92302 85190 92306
rect 85126 92246 85130 92302
rect 85130 92246 85186 92302
rect 85186 92246 85190 92302
rect 85126 92242 85190 92246
rect 2886 91758 2950 91762
rect 2886 91702 2890 91758
rect 2890 91702 2946 91758
rect 2946 91702 2950 91758
rect 2886 91698 2950 91702
rect 2966 91758 3030 91762
rect 2966 91702 2970 91758
rect 2970 91702 3026 91758
rect 3026 91702 3030 91758
rect 2966 91698 3030 91702
rect 3046 91758 3110 91762
rect 3046 91702 3050 91758
rect 3050 91702 3106 91758
rect 3106 91702 3110 91758
rect 3046 91698 3110 91702
rect 3126 91758 3190 91762
rect 3126 91702 3130 91758
rect 3130 91702 3186 91758
rect 3186 91702 3190 91758
rect 3126 91698 3190 91702
rect 86886 91758 86950 91762
rect 86886 91702 86890 91758
rect 86890 91702 86946 91758
rect 86946 91702 86950 91758
rect 86886 91698 86950 91702
rect 86966 91758 87030 91762
rect 86966 91702 86970 91758
rect 86970 91702 87026 91758
rect 87026 91702 87030 91758
rect 86966 91698 87030 91702
rect 87046 91758 87110 91762
rect 87046 91702 87050 91758
rect 87050 91702 87106 91758
rect 87106 91702 87110 91758
rect 87046 91698 87110 91702
rect 87126 91758 87190 91762
rect 87126 91702 87130 91758
rect 87130 91702 87186 91758
rect 87186 91702 87190 91758
rect 87126 91698 87190 91702
rect 886 91214 950 91218
rect 886 91158 890 91214
rect 890 91158 946 91214
rect 946 91158 950 91214
rect 886 91154 950 91158
rect 966 91214 1030 91218
rect 966 91158 970 91214
rect 970 91158 1026 91214
rect 1026 91158 1030 91214
rect 966 91154 1030 91158
rect 1046 91214 1110 91218
rect 1046 91158 1050 91214
rect 1050 91158 1106 91214
rect 1106 91158 1110 91214
rect 1046 91154 1110 91158
rect 1126 91214 1190 91218
rect 1126 91158 1130 91214
rect 1130 91158 1186 91214
rect 1186 91158 1190 91214
rect 1126 91154 1190 91158
rect 84886 91214 84950 91218
rect 84886 91158 84890 91214
rect 84890 91158 84946 91214
rect 84946 91158 84950 91214
rect 84886 91154 84950 91158
rect 84966 91214 85030 91218
rect 84966 91158 84970 91214
rect 84970 91158 85026 91214
rect 85026 91158 85030 91214
rect 84966 91154 85030 91158
rect 85046 91214 85110 91218
rect 85046 91158 85050 91214
rect 85050 91158 85106 91214
rect 85106 91158 85110 91214
rect 85046 91154 85110 91158
rect 85126 91214 85190 91218
rect 85126 91158 85130 91214
rect 85130 91158 85186 91214
rect 85186 91158 85190 91214
rect 85126 91154 85190 91158
rect 2886 90670 2950 90674
rect 2886 90614 2890 90670
rect 2890 90614 2946 90670
rect 2946 90614 2950 90670
rect 2886 90610 2950 90614
rect 2966 90670 3030 90674
rect 2966 90614 2970 90670
rect 2970 90614 3026 90670
rect 3026 90614 3030 90670
rect 2966 90610 3030 90614
rect 3046 90670 3110 90674
rect 3046 90614 3050 90670
rect 3050 90614 3106 90670
rect 3106 90614 3110 90670
rect 3046 90610 3110 90614
rect 3126 90670 3190 90674
rect 3126 90614 3130 90670
rect 3130 90614 3186 90670
rect 3186 90614 3190 90670
rect 3126 90610 3190 90614
rect 86886 90670 86950 90674
rect 86886 90614 86890 90670
rect 86890 90614 86946 90670
rect 86946 90614 86950 90670
rect 86886 90610 86950 90614
rect 86966 90670 87030 90674
rect 86966 90614 86970 90670
rect 86970 90614 87026 90670
rect 87026 90614 87030 90670
rect 86966 90610 87030 90614
rect 87046 90670 87110 90674
rect 87046 90614 87050 90670
rect 87050 90614 87106 90670
rect 87106 90614 87110 90670
rect 87046 90610 87110 90614
rect 87126 90670 87190 90674
rect 87126 90614 87130 90670
rect 87130 90614 87186 90670
rect 87186 90614 87190 90670
rect 87126 90610 87190 90614
rect 886 90126 950 90130
rect 886 90070 890 90126
rect 890 90070 946 90126
rect 946 90070 950 90126
rect 886 90066 950 90070
rect 966 90126 1030 90130
rect 966 90070 970 90126
rect 970 90070 1026 90126
rect 1026 90070 1030 90126
rect 966 90066 1030 90070
rect 1046 90126 1110 90130
rect 1046 90070 1050 90126
rect 1050 90070 1106 90126
rect 1106 90070 1110 90126
rect 1046 90066 1110 90070
rect 1126 90126 1190 90130
rect 1126 90070 1130 90126
rect 1130 90070 1186 90126
rect 1186 90070 1190 90126
rect 1126 90066 1190 90070
rect 84886 90126 84950 90130
rect 84886 90070 84890 90126
rect 84890 90070 84946 90126
rect 84946 90070 84950 90126
rect 84886 90066 84950 90070
rect 84966 90126 85030 90130
rect 84966 90070 84970 90126
rect 84970 90070 85026 90126
rect 85026 90070 85030 90126
rect 84966 90066 85030 90070
rect 85046 90126 85110 90130
rect 85046 90070 85050 90126
rect 85050 90070 85106 90126
rect 85106 90070 85110 90126
rect 85046 90066 85110 90070
rect 85126 90126 85190 90130
rect 85126 90070 85130 90126
rect 85130 90070 85186 90126
rect 85186 90070 85190 90126
rect 85126 90066 85190 90070
rect 2886 89582 2950 89586
rect 2886 89526 2890 89582
rect 2890 89526 2946 89582
rect 2946 89526 2950 89582
rect 2886 89522 2950 89526
rect 2966 89582 3030 89586
rect 2966 89526 2970 89582
rect 2970 89526 3026 89582
rect 3026 89526 3030 89582
rect 2966 89522 3030 89526
rect 3046 89582 3110 89586
rect 3046 89526 3050 89582
rect 3050 89526 3106 89582
rect 3106 89526 3110 89582
rect 3046 89522 3110 89526
rect 3126 89582 3190 89586
rect 3126 89526 3130 89582
rect 3130 89526 3186 89582
rect 3186 89526 3190 89582
rect 3126 89522 3190 89526
rect 86886 89582 86950 89586
rect 86886 89526 86890 89582
rect 86890 89526 86946 89582
rect 86946 89526 86950 89582
rect 86886 89522 86950 89526
rect 86966 89582 87030 89586
rect 86966 89526 86970 89582
rect 86970 89526 87026 89582
rect 87026 89526 87030 89582
rect 86966 89522 87030 89526
rect 87046 89582 87110 89586
rect 87046 89526 87050 89582
rect 87050 89526 87106 89582
rect 87106 89526 87110 89582
rect 87046 89522 87110 89526
rect 87126 89582 87190 89586
rect 87126 89526 87130 89582
rect 87130 89526 87186 89582
rect 87186 89526 87190 89582
rect 87126 89522 87190 89526
rect 886 89038 950 89042
rect 886 88982 890 89038
rect 890 88982 946 89038
rect 946 88982 950 89038
rect 886 88978 950 88982
rect 966 89038 1030 89042
rect 966 88982 970 89038
rect 970 88982 1026 89038
rect 1026 88982 1030 89038
rect 966 88978 1030 88982
rect 1046 89038 1110 89042
rect 1046 88982 1050 89038
rect 1050 88982 1106 89038
rect 1106 88982 1110 89038
rect 1046 88978 1110 88982
rect 1126 89038 1190 89042
rect 1126 88982 1130 89038
rect 1130 88982 1186 89038
rect 1186 88982 1190 89038
rect 1126 88978 1190 88982
rect 84886 89038 84950 89042
rect 84886 88982 84890 89038
rect 84890 88982 84946 89038
rect 84946 88982 84950 89038
rect 84886 88978 84950 88982
rect 84966 89038 85030 89042
rect 84966 88982 84970 89038
rect 84970 88982 85026 89038
rect 85026 88982 85030 89038
rect 84966 88978 85030 88982
rect 85046 89038 85110 89042
rect 85046 88982 85050 89038
rect 85050 88982 85106 89038
rect 85106 88982 85110 89038
rect 85046 88978 85110 88982
rect 85126 89038 85190 89042
rect 85126 88982 85130 89038
rect 85130 88982 85186 89038
rect 85186 88982 85190 89038
rect 85126 88978 85190 88982
rect 2886 88494 2950 88498
rect 2886 88438 2890 88494
rect 2890 88438 2946 88494
rect 2946 88438 2950 88494
rect 2886 88434 2950 88438
rect 2966 88494 3030 88498
rect 2966 88438 2970 88494
rect 2970 88438 3026 88494
rect 3026 88438 3030 88494
rect 2966 88434 3030 88438
rect 3046 88494 3110 88498
rect 3046 88438 3050 88494
rect 3050 88438 3106 88494
rect 3106 88438 3110 88494
rect 3046 88434 3110 88438
rect 3126 88494 3190 88498
rect 3126 88438 3130 88494
rect 3130 88438 3186 88494
rect 3186 88438 3190 88494
rect 3126 88434 3190 88438
rect 86886 88494 86950 88498
rect 86886 88438 86890 88494
rect 86890 88438 86946 88494
rect 86946 88438 86950 88494
rect 86886 88434 86950 88438
rect 86966 88494 87030 88498
rect 86966 88438 86970 88494
rect 86970 88438 87026 88494
rect 87026 88438 87030 88494
rect 86966 88434 87030 88438
rect 87046 88494 87110 88498
rect 87046 88438 87050 88494
rect 87050 88438 87106 88494
rect 87106 88438 87110 88494
rect 87046 88434 87110 88438
rect 87126 88494 87190 88498
rect 87126 88438 87130 88494
rect 87130 88438 87186 88494
rect 87186 88438 87190 88494
rect 87126 88434 87190 88438
rect 886 87950 950 87954
rect 886 87894 890 87950
rect 890 87894 946 87950
rect 946 87894 950 87950
rect 886 87890 950 87894
rect 966 87950 1030 87954
rect 966 87894 970 87950
rect 970 87894 1026 87950
rect 1026 87894 1030 87950
rect 966 87890 1030 87894
rect 1046 87950 1110 87954
rect 1046 87894 1050 87950
rect 1050 87894 1106 87950
rect 1106 87894 1110 87950
rect 1046 87890 1110 87894
rect 1126 87950 1190 87954
rect 1126 87894 1130 87950
rect 1130 87894 1186 87950
rect 1186 87894 1190 87950
rect 1126 87890 1190 87894
rect 84886 87950 84950 87954
rect 84886 87894 84890 87950
rect 84890 87894 84946 87950
rect 84946 87894 84950 87950
rect 84886 87890 84950 87894
rect 84966 87950 85030 87954
rect 84966 87894 84970 87950
rect 84970 87894 85026 87950
rect 85026 87894 85030 87950
rect 84966 87890 85030 87894
rect 85046 87950 85110 87954
rect 85046 87894 85050 87950
rect 85050 87894 85106 87950
rect 85106 87894 85110 87950
rect 85046 87890 85110 87894
rect 85126 87950 85190 87954
rect 85126 87894 85130 87950
rect 85130 87894 85186 87950
rect 85186 87894 85190 87950
rect 85126 87890 85190 87894
rect 2886 87406 2950 87410
rect 2886 87350 2890 87406
rect 2890 87350 2946 87406
rect 2946 87350 2950 87406
rect 2886 87346 2950 87350
rect 2966 87406 3030 87410
rect 2966 87350 2970 87406
rect 2970 87350 3026 87406
rect 3026 87350 3030 87406
rect 2966 87346 3030 87350
rect 3046 87406 3110 87410
rect 3046 87350 3050 87406
rect 3050 87350 3106 87406
rect 3106 87350 3110 87406
rect 3046 87346 3110 87350
rect 3126 87406 3190 87410
rect 3126 87350 3130 87406
rect 3130 87350 3186 87406
rect 3186 87350 3190 87406
rect 3126 87346 3190 87350
rect 86886 87406 86950 87410
rect 86886 87350 86890 87406
rect 86890 87350 86946 87406
rect 86946 87350 86950 87406
rect 86886 87346 86950 87350
rect 86966 87406 87030 87410
rect 86966 87350 86970 87406
rect 86970 87350 87026 87406
rect 87026 87350 87030 87406
rect 86966 87346 87030 87350
rect 87046 87406 87110 87410
rect 87046 87350 87050 87406
rect 87050 87350 87106 87406
rect 87106 87350 87110 87406
rect 87046 87346 87110 87350
rect 87126 87406 87190 87410
rect 87126 87350 87130 87406
rect 87130 87350 87186 87406
rect 87186 87350 87190 87406
rect 87126 87346 87190 87350
rect 886 86862 950 86866
rect 886 86806 890 86862
rect 890 86806 946 86862
rect 946 86806 950 86862
rect 886 86802 950 86806
rect 966 86862 1030 86866
rect 966 86806 970 86862
rect 970 86806 1026 86862
rect 1026 86806 1030 86862
rect 966 86802 1030 86806
rect 1046 86862 1110 86866
rect 1046 86806 1050 86862
rect 1050 86806 1106 86862
rect 1106 86806 1110 86862
rect 1046 86802 1110 86806
rect 1126 86862 1190 86866
rect 1126 86806 1130 86862
rect 1130 86806 1186 86862
rect 1186 86806 1190 86862
rect 1126 86802 1190 86806
rect 84886 86862 84950 86866
rect 84886 86806 84890 86862
rect 84890 86806 84946 86862
rect 84946 86806 84950 86862
rect 84886 86802 84950 86806
rect 84966 86862 85030 86866
rect 84966 86806 84970 86862
rect 84970 86806 85026 86862
rect 85026 86806 85030 86862
rect 84966 86802 85030 86806
rect 85046 86862 85110 86866
rect 85046 86806 85050 86862
rect 85050 86806 85106 86862
rect 85106 86806 85110 86862
rect 85046 86802 85110 86806
rect 85126 86862 85190 86866
rect 85126 86806 85130 86862
rect 85130 86806 85186 86862
rect 85186 86806 85190 86862
rect 85126 86802 85190 86806
rect 2886 86318 2950 86322
rect 2886 86262 2890 86318
rect 2890 86262 2946 86318
rect 2946 86262 2950 86318
rect 2886 86258 2950 86262
rect 2966 86318 3030 86322
rect 2966 86262 2970 86318
rect 2970 86262 3026 86318
rect 3026 86262 3030 86318
rect 2966 86258 3030 86262
rect 3046 86318 3110 86322
rect 3046 86262 3050 86318
rect 3050 86262 3106 86318
rect 3106 86262 3110 86318
rect 3046 86258 3110 86262
rect 3126 86318 3190 86322
rect 3126 86262 3130 86318
rect 3130 86262 3186 86318
rect 3186 86262 3190 86318
rect 3126 86258 3190 86262
rect 86886 86318 86950 86322
rect 86886 86262 86890 86318
rect 86890 86262 86946 86318
rect 86946 86262 86950 86318
rect 86886 86258 86950 86262
rect 86966 86318 87030 86322
rect 86966 86262 86970 86318
rect 86970 86262 87026 86318
rect 87026 86262 87030 86318
rect 86966 86258 87030 86262
rect 87046 86318 87110 86322
rect 87046 86262 87050 86318
rect 87050 86262 87106 86318
rect 87106 86262 87110 86318
rect 87046 86258 87110 86262
rect 87126 86318 87190 86322
rect 87126 86262 87130 86318
rect 87130 86262 87186 86318
rect 87186 86262 87190 86318
rect 87126 86258 87190 86262
rect 886 85774 950 85778
rect 886 85718 890 85774
rect 890 85718 946 85774
rect 946 85718 950 85774
rect 886 85714 950 85718
rect 966 85774 1030 85778
rect 966 85718 970 85774
rect 970 85718 1026 85774
rect 1026 85718 1030 85774
rect 966 85714 1030 85718
rect 1046 85774 1110 85778
rect 1046 85718 1050 85774
rect 1050 85718 1106 85774
rect 1106 85718 1110 85774
rect 1046 85714 1110 85718
rect 1126 85774 1190 85778
rect 1126 85718 1130 85774
rect 1130 85718 1186 85774
rect 1186 85718 1190 85774
rect 1126 85714 1190 85718
rect 84886 85774 84950 85778
rect 84886 85718 84890 85774
rect 84890 85718 84946 85774
rect 84946 85718 84950 85774
rect 84886 85714 84950 85718
rect 84966 85774 85030 85778
rect 84966 85718 84970 85774
rect 84970 85718 85026 85774
rect 85026 85718 85030 85774
rect 84966 85714 85030 85718
rect 85046 85774 85110 85778
rect 85046 85718 85050 85774
rect 85050 85718 85106 85774
rect 85106 85718 85110 85774
rect 85046 85714 85110 85718
rect 85126 85774 85190 85778
rect 85126 85718 85130 85774
rect 85130 85718 85186 85774
rect 85186 85718 85190 85774
rect 85126 85714 85190 85718
rect 2886 85230 2950 85234
rect 2886 85174 2890 85230
rect 2890 85174 2946 85230
rect 2946 85174 2950 85230
rect 2886 85170 2950 85174
rect 2966 85230 3030 85234
rect 2966 85174 2970 85230
rect 2970 85174 3026 85230
rect 3026 85174 3030 85230
rect 2966 85170 3030 85174
rect 3046 85230 3110 85234
rect 3046 85174 3050 85230
rect 3050 85174 3106 85230
rect 3106 85174 3110 85230
rect 3046 85170 3110 85174
rect 3126 85230 3190 85234
rect 3126 85174 3130 85230
rect 3130 85174 3186 85230
rect 3186 85174 3190 85230
rect 3126 85170 3190 85174
rect 86886 85230 86950 85234
rect 86886 85174 86890 85230
rect 86890 85174 86946 85230
rect 86946 85174 86950 85230
rect 86886 85170 86950 85174
rect 86966 85230 87030 85234
rect 86966 85174 86970 85230
rect 86970 85174 87026 85230
rect 87026 85174 87030 85230
rect 86966 85170 87030 85174
rect 87046 85230 87110 85234
rect 87046 85174 87050 85230
rect 87050 85174 87106 85230
rect 87106 85174 87110 85230
rect 87046 85170 87110 85174
rect 87126 85230 87190 85234
rect 87126 85174 87130 85230
rect 87130 85174 87186 85230
rect 87186 85174 87190 85230
rect 87126 85170 87190 85174
rect 886 84686 950 84690
rect 886 84630 890 84686
rect 890 84630 946 84686
rect 946 84630 950 84686
rect 886 84626 950 84630
rect 966 84686 1030 84690
rect 966 84630 970 84686
rect 970 84630 1026 84686
rect 1026 84630 1030 84686
rect 966 84626 1030 84630
rect 1046 84686 1110 84690
rect 1046 84630 1050 84686
rect 1050 84630 1106 84686
rect 1106 84630 1110 84686
rect 1046 84626 1110 84630
rect 1126 84686 1190 84690
rect 1126 84630 1130 84686
rect 1130 84630 1186 84686
rect 1186 84630 1190 84686
rect 1126 84626 1190 84630
rect 84886 84686 84950 84690
rect 84886 84630 84890 84686
rect 84890 84630 84946 84686
rect 84946 84630 84950 84686
rect 84886 84626 84950 84630
rect 84966 84686 85030 84690
rect 84966 84630 84970 84686
rect 84970 84630 85026 84686
rect 85026 84630 85030 84686
rect 84966 84626 85030 84630
rect 85046 84686 85110 84690
rect 85046 84630 85050 84686
rect 85050 84630 85106 84686
rect 85106 84630 85110 84686
rect 85046 84626 85110 84630
rect 85126 84686 85190 84690
rect 85126 84630 85130 84686
rect 85130 84630 85186 84686
rect 85186 84630 85190 84686
rect 85126 84626 85190 84630
rect 2886 84142 2950 84146
rect 2886 84086 2890 84142
rect 2890 84086 2946 84142
rect 2946 84086 2950 84142
rect 2886 84082 2950 84086
rect 2966 84142 3030 84146
rect 2966 84086 2970 84142
rect 2970 84086 3026 84142
rect 3026 84086 3030 84142
rect 2966 84082 3030 84086
rect 3046 84142 3110 84146
rect 3046 84086 3050 84142
rect 3050 84086 3106 84142
rect 3106 84086 3110 84142
rect 3046 84082 3110 84086
rect 3126 84142 3190 84146
rect 3126 84086 3130 84142
rect 3130 84086 3186 84142
rect 3186 84086 3190 84142
rect 3126 84082 3190 84086
rect 86886 84142 86950 84146
rect 86886 84086 86890 84142
rect 86890 84086 86946 84142
rect 86946 84086 86950 84142
rect 86886 84082 86950 84086
rect 86966 84142 87030 84146
rect 86966 84086 86970 84142
rect 86970 84086 87026 84142
rect 87026 84086 87030 84142
rect 86966 84082 87030 84086
rect 87046 84142 87110 84146
rect 87046 84086 87050 84142
rect 87050 84086 87106 84142
rect 87106 84086 87110 84142
rect 87046 84082 87110 84086
rect 87126 84142 87190 84146
rect 87126 84086 87130 84142
rect 87130 84086 87186 84142
rect 87186 84086 87190 84142
rect 87126 84082 87190 84086
rect 4698 83606 4762 83670
rect 886 83598 950 83602
rect 886 83542 890 83598
rect 890 83542 946 83598
rect 946 83542 950 83598
rect 886 83538 950 83542
rect 966 83598 1030 83602
rect 966 83542 970 83598
rect 970 83542 1026 83598
rect 1026 83542 1030 83598
rect 966 83538 1030 83542
rect 1046 83598 1110 83602
rect 1046 83542 1050 83598
rect 1050 83542 1106 83598
rect 1106 83542 1110 83598
rect 1046 83538 1110 83542
rect 1126 83598 1190 83602
rect 1126 83542 1130 83598
rect 1130 83542 1186 83598
rect 1186 83542 1190 83598
rect 1126 83538 1190 83542
rect 84886 83598 84950 83602
rect 84886 83542 84890 83598
rect 84890 83542 84946 83598
rect 84946 83542 84950 83598
rect 84886 83538 84950 83542
rect 84966 83598 85030 83602
rect 84966 83542 84970 83598
rect 84970 83542 85026 83598
rect 85026 83542 85030 83598
rect 84966 83538 85030 83542
rect 85046 83598 85110 83602
rect 85046 83542 85050 83598
rect 85050 83542 85106 83598
rect 85106 83542 85110 83598
rect 85046 83538 85110 83542
rect 85126 83598 85190 83602
rect 85126 83542 85130 83598
rect 85130 83542 85186 83598
rect 85186 83542 85190 83598
rect 85126 83538 85190 83542
rect 4698 83334 4762 83398
rect 2886 83054 2950 83058
rect 2886 82998 2890 83054
rect 2890 82998 2946 83054
rect 2946 82998 2950 83054
rect 2886 82994 2950 82998
rect 2966 83054 3030 83058
rect 2966 82998 2970 83054
rect 2970 82998 3026 83054
rect 3026 82998 3030 83054
rect 2966 82994 3030 82998
rect 3046 83054 3110 83058
rect 3046 82998 3050 83054
rect 3050 82998 3106 83054
rect 3106 82998 3110 83054
rect 3046 82994 3110 82998
rect 3126 83054 3190 83058
rect 3126 82998 3130 83054
rect 3130 82998 3186 83054
rect 3186 82998 3190 83054
rect 3126 82994 3190 82998
rect 86886 83054 86950 83058
rect 86886 82998 86890 83054
rect 86890 82998 86946 83054
rect 86946 82998 86950 83054
rect 86886 82994 86950 82998
rect 86966 83054 87030 83058
rect 86966 82998 86970 83054
rect 86970 82998 87026 83054
rect 87026 82998 87030 83054
rect 86966 82994 87030 82998
rect 87046 83054 87110 83058
rect 87046 82998 87050 83054
rect 87050 82998 87106 83054
rect 87106 82998 87110 83054
rect 87046 82994 87110 82998
rect 87126 83054 87190 83058
rect 87126 82998 87130 83054
rect 87130 82998 87186 83054
rect 87186 82998 87190 83054
rect 87126 82994 87190 82998
rect 886 82510 950 82514
rect 886 82454 890 82510
rect 890 82454 946 82510
rect 946 82454 950 82510
rect 886 82450 950 82454
rect 966 82510 1030 82514
rect 966 82454 970 82510
rect 970 82454 1026 82510
rect 1026 82454 1030 82510
rect 966 82450 1030 82454
rect 1046 82510 1110 82514
rect 1046 82454 1050 82510
rect 1050 82454 1106 82510
rect 1106 82454 1110 82510
rect 1046 82450 1110 82454
rect 1126 82510 1190 82514
rect 1126 82454 1130 82510
rect 1130 82454 1186 82510
rect 1186 82454 1190 82510
rect 1126 82450 1190 82454
rect 84886 82510 84950 82514
rect 84886 82454 84890 82510
rect 84890 82454 84946 82510
rect 84946 82454 84950 82510
rect 84886 82450 84950 82454
rect 84966 82510 85030 82514
rect 84966 82454 84970 82510
rect 84970 82454 85026 82510
rect 85026 82454 85030 82510
rect 84966 82450 85030 82454
rect 85046 82510 85110 82514
rect 85046 82454 85050 82510
rect 85050 82454 85106 82510
rect 85106 82454 85110 82510
rect 85046 82450 85110 82454
rect 85126 82510 85190 82514
rect 85126 82454 85130 82510
rect 85130 82454 85186 82510
rect 85186 82454 85190 82510
rect 85126 82450 85190 82454
rect 2886 81966 2950 81970
rect 2886 81910 2890 81966
rect 2890 81910 2946 81966
rect 2946 81910 2950 81966
rect 2886 81906 2950 81910
rect 2966 81966 3030 81970
rect 2966 81910 2970 81966
rect 2970 81910 3026 81966
rect 3026 81910 3030 81966
rect 2966 81906 3030 81910
rect 3046 81966 3110 81970
rect 3046 81910 3050 81966
rect 3050 81910 3106 81966
rect 3106 81910 3110 81966
rect 3046 81906 3110 81910
rect 3126 81966 3190 81970
rect 3126 81910 3130 81966
rect 3130 81910 3186 81966
rect 3186 81910 3190 81966
rect 3126 81906 3190 81910
rect 86886 81966 86950 81970
rect 86886 81910 86890 81966
rect 86890 81910 86946 81966
rect 86946 81910 86950 81966
rect 86886 81906 86950 81910
rect 86966 81966 87030 81970
rect 86966 81910 86970 81966
rect 86970 81910 87026 81966
rect 87026 81910 87030 81966
rect 86966 81906 87030 81910
rect 87046 81966 87110 81970
rect 87046 81910 87050 81966
rect 87050 81910 87106 81966
rect 87106 81910 87110 81966
rect 87046 81906 87110 81910
rect 87126 81966 87190 81970
rect 87126 81910 87130 81966
rect 87130 81910 87186 81966
rect 87186 81910 87190 81966
rect 87126 81906 87190 81910
rect 886 81422 950 81426
rect 886 81366 890 81422
rect 890 81366 946 81422
rect 946 81366 950 81422
rect 886 81362 950 81366
rect 966 81422 1030 81426
rect 966 81366 970 81422
rect 970 81366 1026 81422
rect 1026 81366 1030 81422
rect 966 81362 1030 81366
rect 1046 81422 1110 81426
rect 1046 81366 1050 81422
rect 1050 81366 1106 81422
rect 1106 81366 1110 81422
rect 1046 81362 1110 81366
rect 1126 81422 1190 81426
rect 1126 81366 1130 81422
rect 1130 81366 1186 81422
rect 1186 81366 1190 81422
rect 1126 81362 1190 81366
rect 84886 81422 84950 81426
rect 84886 81366 84890 81422
rect 84890 81366 84946 81422
rect 84946 81366 84950 81422
rect 84886 81362 84950 81366
rect 84966 81422 85030 81426
rect 84966 81366 84970 81422
rect 84970 81366 85026 81422
rect 85026 81366 85030 81422
rect 84966 81362 85030 81366
rect 85046 81422 85110 81426
rect 85046 81366 85050 81422
rect 85050 81366 85106 81422
rect 85106 81366 85110 81422
rect 85046 81362 85110 81366
rect 85126 81422 85190 81426
rect 85126 81366 85130 81422
rect 85130 81366 85186 81422
rect 85186 81366 85190 81422
rect 85126 81362 85190 81366
rect 2886 80878 2950 80882
rect 2886 80822 2890 80878
rect 2890 80822 2946 80878
rect 2946 80822 2950 80878
rect 2886 80818 2950 80822
rect 2966 80878 3030 80882
rect 2966 80822 2970 80878
rect 2970 80822 3026 80878
rect 3026 80822 3030 80878
rect 2966 80818 3030 80822
rect 3046 80878 3110 80882
rect 3046 80822 3050 80878
rect 3050 80822 3106 80878
rect 3106 80822 3110 80878
rect 3046 80818 3110 80822
rect 3126 80878 3190 80882
rect 3126 80822 3130 80878
rect 3130 80822 3186 80878
rect 3186 80822 3190 80878
rect 3126 80818 3190 80822
rect 86886 80878 86950 80882
rect 86886 80822 86890 80878
rect 86890 80822 86946 80878
rect 86946 80822 86950 80878
rect 86886 80818 86950 80822
rect 86966 80878 87030 80882
rect 86966 80822 86970 80878
rect 86970 80822 87026 80878
rect 87026 80822 87030 80878
rect 86966 80818 87030 80822
rect 87046 80878 87110 80882
rect 87046 80822 87050 80878
rect 87050 80822 87106 80878
rect 87106 80822 87110 80878
rect 87046 80818 87110 80822
rect 87126 80878 87190 80882
rect 87126 80822 87130 80878
rect 87130 80822 87186 80878
rect 87186 80822 87190 80878
rect 87126 80818 87190 80822
rect 886 80334 950 80338
rect 886 80278 890 80334
rect 890 80278 946 80334
rect 946 80278 950 80334
rect 886 80274 950 80278
rect 966 80334 1030 80338
rect 966 80278 970 80334
rect 970 80278 1026 80334
rect 1026 80278 1030 80334
rect 966 80274 1030 80278
rect 1046 80334 1110 80338
rect 1046 80278 1050 80334
rect 1050 80278 1106 80334
rect 1106 80278 1110 80334
rect 1046 80274 1110 80278
rect 1126 80334 1190 80338
rect 1126 80278 1130 80334
rect 1130 80278 1186 80334
rect 1186 80278 1190 80334
rect 1126 80274 1190 80278
rect 84886 80334 84950 80338
rect 84886 80278 84890 80334
rect 84890 80278 84946 80334
rect 84946 80278 84950 80334
rect 84886 80274 84950 80278
rect 84966 80334 85030 80338
rect 84966 80278 84970 80334
rect 84970 80278 85026 80334
rect 85026 80278 85030 80334
rect 84966 80274 85030 80278
rect 85046 80334 85110 80338
rect 85046 80278 85050 80334
rect 85050 80278 85106 80334
rect 85106 80278 85110 80334
rect 85046 80274 85110 80278
rect 85126 80334 85190 80338
rect 85126 80278 85130 80334
rect 85130 80278 85186 80334
rect 85186 80278 85190 80334
rect 85126 80274 85190 80278
rect 2886 79790 2950 79794
rect 2886 79734 2890 79790
rect 2890 79734 2946 79790
rect 2946 79734 2950 79790
rect 2886 79730 2950 79734
rect 2966 79790 3030 79794
rect 2966 79734 2970 79790
rect 2970 79734 3026 79790
rect 3026 79734 3030 79790
rect 2966 79730 3030 79734
rect 3046 79790 3110 79794
rect 3046 79734 3050 79790
rect 3050 79734 3106 79790
rect 3106 79734 3110 79790
rect 3046 79730 3110 79734
rect 3126 79790 3190 79794
rect 3126 79734 3130 79790
rect 3130 79734 3186 79790
rect 3186 79734 3190 79790
rect 3126 79730 3190 79734
rect 86886 79790 86950 79794
rect 86886 79734 86890 79790
rect 86890 79734 86946 79790
rect 86946 79734 86950 79790
rect 86886 79730 86950 79734
rect 86966 79790 87030 79794
rect 86966 79734 86970 79790
rect 86970 79734 87026 79790
rect 87026 79734 87030 79790
rect 86966 79730 87030 79734
rect 87046 79790 87110 79794
rect 87046 79734 87050 79790
rect 87050 79734 87106 79790
rect 87106 79734 87110 79790
rect 87046 79730 87110 79734
rect 87126 79790 87190 79794
rect 87126 79734 87130 79790
rect 87130 79734 87186 79790
rect 87186 79734 87190 79790
rect 87126 79730 87190 79734
rect 886 79246 950 79250
rect 886 79190 890 79246
rect 890 79190 946 79246
rect 946 79190 950 79246
rect 886 79186 950 79190
rect 966 79246 1030 79250
rect 966 79190 970 79246
rect 970 79190 1026 79246
rect 1026 79190 1030 79246
rect 966 79186 1030 79190
rect 1046 79246 1110 79250
rect 1046 79190 1050 79246
rect 1050 79190 1106 79246
rect 1106 79190 1110 79246
rect 1046 79186 1110 79190
rect 1126 79246 1190 79250
rect 1126 79190 1130 79246
rect 1130 79190 1186 79246
rect 1186 79190 1190 79246
rect 1126 79186 1190 79190
rect 84886 79246 84950 79250
rect 84886 79190 84890 79246
rect 84890 79190 84946 79246
rect 84946 79190 84950 79246
rect 84886 79186 84950 79190
rect 84966 79246 85030 79250
rect 84966 79190 84970 79246
rect 84970 79190 85026 79246
rect 85026 79190 85030 79246
rect 84966 79186 85030 79190
rect 85046 79246 85110 79250
rect 85046 79190 85050 79246
rect 85050 79190 85106 79246
rect 85106 79190 85110 79246
rect 85046 79186 85110 79190
rect 85126 79246 85190 79250
rect 85126 79190 85130 79246
rect 85130 79190 85186 79246
rect 85186 79190 85190 79246
rect 85126 79186 85190 79190
rect 2886 78702 2950 78706
rect 2886 78646 2890 78702
rect 2890 78646 2946 78702
rect 2946 78646 2950 78702
rect 2886 78642 2950 78646
rect 2966 78702 3030 78706
rect 2966 78646 2970 78702
rect 2970 78646 3026 78702
rect 3026 78646 3030 78702
rect 2966 78642 3030 78646
rect 3046 78702 3110 78706
rect 3046 78646 3050 78702
rect 3050 78646 3106 78702
rect 3106 78646 3110 78702
rect 3046 78642 3110 78646
rect 3126 78702 3190 78706
rect 3126 78646 3130 78702
rect 3130 78646 3186 78702
rect 3186 78646 3190 78702
rect 3126 78642 3190 78646
rect 86886 78702 86950 78706
rect 86886 78646 86890 78702
rect 86890 78646 86946 78702
rect 86946 78646 86950 78702
rect 86886 78642 86950 78646
rect 86966 78702 87030 78706
rect 86966 78646 86970 78702
rect 86970 78646 87026 78702
rect 87026 78646 87030 78702
rect 86966 78642 87030 78646
rect 87046 78702 87110 78706
rect 87046 78646 87050 78702
rect 87050 78646 87106 78702
rect 87106 78646 87110 78702
rect 87046 78642 87110 78646
rect 87126 78702 87190 78706
rect 87126 78646 87130 78702
rect 87130 78646 87186 78702
rect 87186 78646 87190 78702
rect 87126 78642 87190 78646
rect 886 78158 950 78162
rect 886 78102 890 78158
rect 890 78102 946 78158
rect 946 78102 950 78158
rect 886 78098 950 78102
rect 966 78158 1030 78162
rect 966 78102 970 78158
rect 970 78102 1026 78158
rect 1026 78102 1030 78158
rect 966 78098 1030 78102
rect 1046 78158 1110 78162
rect 1046 78102 1050 78158
rect 1050 78102 1106 78158
rect 1106 78102 1110 78158
rect 1046 78098 1110 78102
rect 1126 78158 1190 78162
rect 1126 78102 1130 78158
rect 1130 78102 1186 78158
rect 1186 78102 1190 78158
rect 1126 78098 1190 78102
rect 84886 78158 84950 78162
rect 84886 78102 84890 78158
rect 84890 78102 84946 78158
rect 84946 78102 84950 78158
rect 84886 78098 84950 78102
rect 84966 78158 85030 78162
rect 84966 78102 84970 78158
rect 84970 78102 85026 78158
rect 85026 78102 85030 78158
rect 84966 78098 85030 78102
rect 85046 78158 85110 78162
rect 85046 78102 85050 78158
rect 85050 78102 85106 78158
rect 85106 78102 85110 78158
rect 85046 78098 85110 78102
rect 85126 78158 85190 78162
rect 85126 78102 85130 78158
rect 85130 78102 85186 78158
rect 85186 78102 85190 78158
rect 85126 78098 85190 78102
rect 2886 77614 2950 77618
rect 2886 77558 2890 77614
rect 2890 77558 2946 77614
rect 2946 77558 2950 77614
rect 2886 77554 2950 77558
rect 2966 77614 3030 77618
rect 2966 77558 2970 77614
rect 2970 77558 3026 77614
rect 3026 77558 3030 77614
rect 2966 77554 3030 77558
rect 3046 77614 3110 77618
rect 3046 77558 3050 77614
rect 3050 77558 3106 77614
rect 3106 77558 3110 77614
rect 3046 77554 3110 77558
rect 3126 77614 3190 77618
rect 3126 77558 3130 77614
rect 3130 77558 3186 77614
rect 3186 77558 3190 77614
rect 3126 77554 3190 77558
rect 86886 77614 86950 77618
rect 86886 77558 86890 77614
rect 86890 77558 86946 77614
rect 86946 77558 86950 77614
rect 86886 77554 86950 77558
rect 86966 77614 87030 77618
rect 86966 77558 86970 77614
rect 86970 77558 87026 77614
rect 87026 77558 87030 77614
rect 86966 77554 87030 77558
rect 87046 77614 87110 77618
rect 87046 77558 87050 77614
rect 87050 77558 87106 77614
rect 87106 77558 87110 77614
rect 87046 77554 87110 77558
rect 87126 77614 87190 77618
rect 87126 77558 87130 77614
rect 87130 77558 87186 77614
rect 87186 77558 87190 77614
rect 87126 77554 87190 77558
rect 886 77070 950 77074
rect 886 77014 890 77070
rect 890 77014 946 77070
rect 946 77014 950 77070
rect 886 77010 950 77014
rect 966 77070 1030 77074
rect 966 77014 970 77070
rect 970 77014 1026 77070
rect 1026 77014 1030 77070
rect 966 77010 1030 77014
rect 1046 77070 1110 77074
rect 1046 77014 1050 77070
rect 1050 77014 1106 77070
rect 1106 77014 1110 77070
rect 1046 77010 1110 77014
rect 1126 77070 1190 77074
rect 1126 77014 1130 77070
rect 1130 77014 1186 77070
rect 1186 77014 1190 77070
rect 1126 77010 1190 77014
rect 84886 77070 84950 77074
rect 84886 77014 84890 77070
rect 84890 77014 84946 77070
rect 84946 77014 84950 77070
rect 84886 77010 84950 77014
rect 84966 77070 85030 77074
rect 84966 77014 84970 77070
rect 84970 77014 85026 77070
rect 85026 77014 85030 77070
rect 84966 77010 85030 77014
rect 85046 77070 85110 77074
rect 85046 77014 85050 77070
rect 85050 77014 85106 77070
rect 85106 77014 85110 77070
rect 85046 77010 85110 77014
rect 85126 77070 85190 77074
rect 85126 77014 85130 77070
rect 85130 77014 85186 77070
rect 85186 77014 85190 77070
rect 85126 77010 85190 77014
rect 2886 76526 2950 76530
rect 2886 76470 2890 76526
rect 2890 76470 2946 76526
rect 2946 76470 2950 76526
rect 2886 76466 2950 76470
rect 2966 76526 3030 76530
rect 2966 76470 2970 76526
rect 2970 76470 3026 76526
rect 3026 76470 3030 76526
rect 2966 76466 3030 76470
rect 3046 76526 3110 76530
rect 3046 76470 3050 76526
rect 3050 76470 3106 76526
rect 3106 76470 3110 76526
rect 3046 76466 3110 76470
rect 3126 76526 3190 76530
rect 3126 76470 3130 76526
rect 3130 76470 3186 76526
rect 3186 76470 3190 76526
rect 3126 76466 3190 76470
rect 86886 76526 86950 76530
rect 86886 76470 86890 76526
rect 86890 76470 86946 76526
rect 86946 76470 86950 76526
rect 86886 76466 86950 76470
rect 86966 76526 87030 76530
rect 86966 76470 86970 76526
rect 86970 76470 87026 76526
rect 87026 76470 87030 76526
rect 86966 76466 87030 76470
rect 87046 76526 87110 76530
rect 87046 76470 87050 76526
rect 87050 76470 87106 76526
rect 87106 76470 87110 76526
rect 87046 76466 87110 76470
rect 87126 76526 87190 76530
rect 87126 76470 87130 76526
rect 87130 76470 87186 76526
rect 87186 76470 87190 76526
rect 87126 76466 87190 76470
rect 886 75982 950 75986
rect 886 75926 890 75982
rect 890 75926 946 75982
rect 946 75926 950 75982
rect 886 75922 950 75926
rect 966 75982 1030 75986
rect 966 75926 970 75982
rect 970 75926 1026 75982
rect 1026 75926 1030 75982
rect 966 75922 1030 75926
rect 1046 75982 1110 75986
rect 1046 75926 1050 75982
rect 1050 75926 1106 75982
rect 1106 75926 1110 75982
rect 1046 75922 1110 75926
rect 1126 75982 1190 75986
rect 1126 75926 1130 75982
rect 1130 75926 1186 75982
rect 1186 75926 1190 75982
rect 1126 75922 1190 75926
rect 84886 75982 84950 75986
rect 84886 75926 84890 75982
rect 84890 75926 84946 75982
rect 84946 75926 84950 75982
rect 84886 75922 84950 75926
rect 84966 75982 85030 75986
rect 84966 75926 84970 75982
rect 84970 75926 85026 75982
rect 85026 75926 85030 75982
rect 84966 75922 85030 75926
rect 85046 75982 85110 75986
rect 85046 75926 85050 75982
rect 85050 75926 85106 75982
rect 85106 75926 85110 75982
rect 85046 75922 85110 75926
rect 85126 75982 85190 75986
rect 85126 75926 85130 75982
rect 85130 75926 85186 75982
rect 85186 75926 85190 75982
rect 85126 75922 85190 75926
rect 2886 75438 2950 75442
rect 2886 75382 2890 75438
rect 2890 75382 2946 75438
rect 2946 75382 2950 75438
rect 2886 75378 2950 75382
rect 2966 75438 3030 75442
rect 2966 75382 2970 75438
rect 2970 75382 3026 75438
rect 3026 75382 3030 75438
rect 2966 75378 3030 75382
rect 3046 75438 3110 75442
rect 3046 75382 3050 75438
rect 3050 75382 3106 75438
rect 3106 75382 3110 75438
rect 3046 75378 3110 75382
rect 3126 75438 3190 75442
rect 3126 75382 3130 75438
rect 3130 75382 3186 75438
rect 3186 75382 3190 75438
rect 3126 75378 3190 75382
rect 86886 75438 86950 75442
rect 86886 75382 86890 75438
rect 86890 75382 86946 75438
rect 86946 75382 86950 75438
rect 86886 75378 86950 75382
rect 86966 75438 87030 75442
rect 86966 75382 86970 75438
rect 86970 75382 87026 75438
rect 87026 75382 87030 75438
rect 86966 75378 87030 75382
rect 87046 75438 87110 75442
rect 87046 75382 87050 75438
rect 87050 75382 87106 75438
rect 87106 75382 87110 75438
rect 87046 75378 87110 75382
rect 87126 75438 87190 75442
rect 87126 75382 87130 75438
rect 87130 75382 87186 75438
rect 87186 75382 87190 75438
rect 87126 75378 87190 75382
rect 886 74894 950 74898
rect 886 74838 890 74894
rect 890 74838 946 74894
rect 946 74838 950 74894
rect 886 74834 950 74838
rect 966 74894 1030 74898
rect 966 74838 970 74894
rect 970 74838 1026 74894
rect 1026 74838 1030 74894
rect 966 74834 1030 74838
rect 1046 74894 1110 74898
rect 1046 74838 1050 74894
rect 1050 74838 1106 74894
rect 1106 74838 1110 74894
rect 1046 74834 1110 74838
rect 1126 74894 1190 74898
rect 1126 74838 1130 74894
rect 1130 74838 1186 74894
rect 1186 74838 1190 74894
rect 1126 74834 1190 74838
rect 84886 74894 84950 74898
rect 84886 74838 84890 74894
rect 84890 74838 84946 74894
rect 84946 74838 84950 74894
rect 84886 74834 84950 74838
rect 84966 74894 85030 74898
rect 84966 74838 84970 74894
rect 84970 74838 85026 74894
rect 85026 74838 85030 74894
rect 84966 74834 85030 74838
rect 85046 74894 85110 74898
rect 85046 74838 85050 74894
rect 85050 74838 85106 74894
rect 85106 74838 85110 74894
rect 85046 74834 85110 74838
rect 85126 74894 85190 74898
rect 85126 74838 85130 74894
rect 85130 74838 85186 74894
rect 85186 74838 85190 74894
rect 85126 74834 85190 74838
rect 4698 74630 4762 74694
rect 4514 74358 4578 74422
rect 2886 74350 2950 74354
rect 2886 74294 2890 74350
rect 2890 74294 2946 74350
rect 2946 74294 2950 74350
rect 2886 74290 2950 74294
rect 2966 74350 3030 74354
rect 2966 74294 2970 74350
rect 2970 74294 3026 74350
rect 3026 74294 3030 74350
rect 2966 74290 3030 74294
rect 3046 74350 3110 74354
rect 3046 74294 3050 74350
rect 3050 74294 3106 74350
rect 3106 74294 3110 74350
rect 3046 74290 3110 74294
rect 3126 74350 3190 74354
rect 3126 74294 3130 74350
rect 3130 74294 3186 74350
rect 3186 74294 3190 74350
rect 3126 74290 3190 74294
rect 86886 74350 86950 74354
rect 86886 74294 86890 74350
rect 86890 74294 86946 74350
rect 86946 74294 86950 74350
rect 86886 74290 86950 74294
rect 86966 74350 87030 74354
rect 86966 74294 86970 74350
rect 86970 74294 87026 74350
rect 87026 74294 87030 74350
rect 86966 74290 87030 74294
rect 87046 74350 87110 74354
rect 87046 74294 87050 74350
rect 87050 74294 87106 74350
rect 87106 74294 87110 74350
rect 87046 74290 87110 74294
rect 87126 74350 87190 74354
rect 87126 74294 87130 74350
rect 87130 74294 87186 74350
rect 87186 74294 87190 74350
rect 87126 74290 87190 74294
rect 886 73806 950 73810
rect 886 73750 890 73806
rect 890 73750 946 73806
rect 946 73750 950 73806
rect 886 73746 950 73750
rect 966 73806 1030 73810
rect 966 73750 970 73806
rect 970 73750 1026 73806
rect 1026 73750 1030 73806
rect 966 73746 1030 73750
rect 1046 73806 1110 73810
rect 1046 73750 1050 73806
rect 1050 73750 1106 73806
rect 1106 73750 1110 73806
rect 1046 73746 1110 73750
rect 1126 73806 1190 73810
rect 1126 73750 1130 73806
rect 1130 73750 1186 73806
rect 1186 73750 1190 73806
rect 1126 73746 1190 73750
rect 84886 73806 84950 73810
rect 84886 73750 84890 73806
rect 84890 73750 84946 73806
rect 84946 73750 84950 73806
rect 84886 73746 84950 73750
rect 84966 73806 85030 73810
rect 84966 73750 84970 73806
rect 84970 73750 85026 73806
rect 85026 73750 85030 73806
rect 84966 73746 85030 73750
rect 85046 73806 85110 73810
rect 85046 73750 85050 73806
rect 85050 73750 85106 73806
rect 85106 73750 85110 73806
rect 85046 73746 85110 73750
rect 85126 73806 85190 73810
rect 85126 73750 85130 73806
rect 85130 73750 85186 73806
rect 85186 73750 85190 73806
rect 85126 73746 85190 73750
rect 2886 73262 2950 73266
rect 2886 73206 2890 73262
rect 2890 73206 2946 73262
rect 2946 73206 2950 73262
rect 2886 73202 2950 73206
rect 2966 73262 3030 73266
rect 2966 73206 2970 73262
rect 2970 73206 3026 73262
rect 3026 73206 3030 73262
rect 2966 73202 3030 73206
rect 3046 73262 3110 73266
rect 3046 73206 3050 73262
rect 3050 73206 3106 73262
rect 3106 73206 3110 73262
rect 3046 73202 3110 73206
rect 3126 73262 3190 73266
rect 3126 73206 3130 73262
rect 3130 73206 3186 73262
rect 3186 73206 3190 73262
rect 3126 73202 3190 73206
rect 86886 73262 86950 73266
rect 86886 73206 86890 73262
rect 86890 73206 86946 73262
rect 86946 73206 86950 73262
rect 86886 73202 86950 73206
rect 86966 73262 87030 73266
rect 86966 73206 86970 73262
rect 86970 73206 87026 73262
rect 87026 73206 87030 73262
rect 86966 73202 87030 73206
rect 87046 73262 87110 73266
rect 87046 73206 87050 73262
rect 87050 73206 87106 73262
rect 87106 73206 87110 73262
rect 87046 73202 87110 73206
rect 87126 73262 87190 73266
rect 87126 73206 87130 73262
rect 87130 73206 87186 73262
rect 87186 73206 87190 73262
rect 87126 73202 87190 73206
rect 886 72718 950 72722
rect 886 72662 890 72718
rect 890 72662 946 72718
rect 946 72662 950 72718
rect 886 72658 950 72662
rect 966 72718 1030 72722
rect 966 72662 970 72718
rect 970 72662 1026 72718
rect 1026 72662 1030 72718
rect 966 72658 1030 72662
rect 1046 72718 1110 72722
rect 1046 72662 1050 72718
rect 1050 72662 1106 72718
rect 1106 72662 1110 72718
rect 1046 72658 1110 72662
rect 1126 72718 1190 72722
rect 1126 72662 1130 72718
rect 1130 72662 1186 72718
rect 1186 72662 1190 72718
rect 1126 72658 1190 72662
rect 84886 72718 84950 72722
rect 84886 72662 84890 72718
rect 84890 72662 84946 72718
rect 84946 72662 84950 72718
rect 84886 72658 84950 72662
rect 84966 72718 85030 72722
rect 84966 72662 84970 72718
rect 84970 72662 85026 72718
rect 85026 72662 85030 72718
rect 84966 72658 85030 72662
rect 85046 72718 85110 72722
rect 85046 72662 85050 72718
rect 85050 72662 85106 72718
rect 85106 72662 85110 72718
rect 85046 72658 85110 72662
rect 85126 72718 85190 72722
rect 85126 72662 85130 72718
rect 85130 72662 85186 72718
rect 85186 72662 85190 72718
rect 85126 72658 85190 72662
rect 2886 72174 2950 72178
rect 2886 72118 2890 72174
rect 2890 72118 2946 72174
rect 2946 72118 2950 72174
rect 2886 72114 2950 72118
rect 2966 72174 3030 72178
rect 2966 72118 2970 72174
rect 2970 72118 3026 72174
rect 3026 72118 3030 72174
rect 2966 72114 3030 72118
rect 3046 72174 3110 72178
rect 3046 72118 3050 72174
rect 3050 72118 3106 72174
rect 3106 72118 3110 72174
rect 3046 72114 3110 72118
rect 3126 72174 3190 72178
rect 3126 72118 3130 72174
rect 3130 72118 3186 72174
rect 3186 72118 3190 72174
rect 3126 72114 3190 72118
rect 86886 72174 86950 72178
rect 86886 72118 86890 72174
rect 86890 72118 86946 72174
rect 86946 72118 86950 72174
rect 86886 72114 86950 72118
rect 86966 72174 87030 72178
rect 86966 72118 86970 72174
rect 86970 72118 87026 72174
rect 87026 72118 87030 72174
rect 86966 72114 87030 72118
rect 87046 72174 87110 72178
rect 87046 72118 87050 72174
rect 87050 72118 87106 72174
rect 87106 72118 87110 72174
rect 87046 72114 87110 72118
rect 87126 72174 87190 72178
rect 87126 72118 87130 72174
rect 87130 72118 87186 72174
rect 87186 72118 87190 72174
rect 87126 72114 87190 72118
rect 886 71630 950 71634
rect 886 71574 890 71630
rect 890 71574 946 71630
rect 946 71574 950 71630
rect 886 71570 950 71574
rect 966 71630 1030 71634
rect 966 71574 970 71630
rect 970 71574 1026 71630
rect 1026 71574 1030 71630
rect 966 71570 1030 71574
rect 1046 71630 1110 71634
rect 1046 71574 1050 71630
rect 1050 71574 1106 71630
rect 1106 71574 1110 71630
rect 1046 71570 1110 71574
rect 1126 71630 1190 71634
rect 1126 71574 1130 71630
rect 1130 71574 1186 71630
rect 1186 71574 1190 71630
rect 1126 71570 1190 71574
rect 84886 71630 84950 71634
rect 84886 71574 84890 71630
rect 84890 71574 84946 71630
rect 84946 71574 84950 71630
rect 84886 71570 84950 71574
rect 84966 71630 85030 71634
rect 84966 71574 84970 71630
rect 84970 71574 85026 71630
rect 85026 71574 85030 71630
rect 84966 71570 85030 71574
rect 85046 71630 85110 71634
rect 85046 71574 85050 71630
rect 85050 71574 85106 71630
rect 85106 71574 85110 71630
rect 85046 71570 85110 71574
rect 85126 71630 85190 71634
rect 85126 71574 85130 71630
rect 85130 71574 85186 71630
rect 85186 71574 85190 71630
rect 85126 71570 85190 71574
rect 2886 71086 2950 71090
rect 2886 71030 2890 71086
rect 2890 71030 2946 71086
rect 2946 71030 2950 71086
rect 2886 71026 2950 71030
rect 2966 71086 3030 71090
rect 2966 71030 2970 71086
rect 2970 71030 3026 71086
rect 3026 71030 3030 71086
rect 2966 71026 3030 71030
rect 3046 71086 3110 71090
rect 3046 71030 3050 71086
rect 3050 71030 3106 71086
rect 3106 71030 3110 71086
rect 3046 71026 3110 71030
rect 3126 71086 3190 71090
rect 3126 71030 3130 71086
rect 3130 71030 3186 71086
rect 3186 71030 3190 71086
rect 3126 71026 3190 71030
rect 86886 71086 86950 71090
rect 86886 71030 86890 71086
rect 86890 71030 86946 71086
rect 86946 71030 86950 71086
rect 86886 71026 86950 71030
rect 86966 71086 87030 71090
rect 86966 71030 86970 71086
rect 86970 71030 87026 71086
rect 87026 71030 87030 71086
rect 86966 71026 87030 71030
rect 87046 71086 87110 71090
rect 87046 71030 87050 71086
rect 87050 71030 87106 71086
rect 87106 71030 87110 71086
rect 87046 71026 87110 71030
rect 87126 71086 87190 71090
rect 87126 71030 87130 71086
rect 87130 71030 87186 71086
rect 87186 71030 87190 71086
rect 87126 71026 87190 71030
rect 886 70542 950 70546
rect 886 70486 890 70542
rect 890 70486 946 70542
rect 946 70486 950 70542
rect 886 70482 950 70486
rect 966 70542 1030 70546
rect 966 70486 970 70542
rect 970 70486 1026 70542
rect 1026 70486 1030 70542
rect 966 70482 1030 70486
rect 1046 70542 1110 70546
rect 1046 70486 1050 70542
rect 1050 70486 1106 70542
rect 1106 70486 1110 70542
rect 1046 70482 1110 70486
rect 1126 70542 1190 70546
rect 1126 70486 1130 70542
rect 1130 70486 1186 70542
rect 1186 70486 1190 70542
rect 1126 70482 1190 70486
rect 84886 70542 84950 70546
rect 84886 70486 84890 70542
rect 84890 70486 84946 70542
rect 84946 70486 84950 70542
rect 84886 70482 84950 70486
rect 84966 70542 85030 70546
rect 84966 70486 84970 70542
rect 84970 70486 85026 70542
rect 85026 70486 85030 70542
rect 84966 70482 85030 70486
rect 85046 70542 85110 70546
rect 85046 70486 85050 70542
rect 85050 70486 85106 70542
rect 85106 70486 85110 70542
rect 85046 70482 85110 70486
rect 85126 70542 85190 70546
rect 85126 70486 85130 70542
rect 85130 70486 85186 70542
rect 85186 70486 85190 70542
rect 85126 70482 85190 70486
rect 2886 69998 2950 70002
rect 2886 69942 2890 69998
rect 2890 69942 2946 69998
rect 2946 69942 2950 69998
rect 2886 69938 2950 69942
rect 2966 69998 3030 70002
rect 2966 69942 2970 69998
rect 2970 69942 3026 69998
rect 3026 69942 3030 69998
rect 2966 69938 3030 69942
rect 3046 69998 3110 70002
rect 3046 69942 3050 69998
rect 3050 69942 3106 69998
rect 3106 69942 3110 69998
rect 3046 69938 3110 69942
rect 3126 69998 3190 70002
rect 3126 69942 3130 69998
rect 3130 69942 3186 69998
rect 3186 69942 3190 69998
rect 3126 69938 3190 69942
rect 86886 69998 86950 70002
rect 86886 69942 86890 69998
rect 86890 69942 86946 69998
rect 86946 69942 86950 69998
rect 86886 69938 86950 69942
rect 86966 69998 87030 70002
rect 86966 69942 86970 69998
rect 86970 69942 87026 69998
rect 87026 69942 87030 69998
rect 86966 69938 87030 69942
rect 87046 69998 87110 70002
rect 87046 69942 87050 69998
rect 87050 69942 87106 69998
rect 87106 69942 87110 69998
rect 87046 69938 87110 69942
rect 87126 69998 87190 70002
rect 87126 69942 87130 69998
rect 87130 69942 87186 69998
rect 87186 69942 87190 69998
rect 87126 69938 87190 69942
rect 886 69454 950 69458
rect 886 69398 890 69454
rect 890 69398 946 69454
rect 946 69398 950 69454
rect 886 69394 950 69398
rect 966 69454 1030 69458
rect 966 69398 970 69454
rect 970 69398 1026 69454
rect 1026 69398 1030 69454
rect 966 69394 1030 69398
rect 1046 69454 1110 69458
rect 1046 69398 1050 69454
rect 1050 69398 1106 69454
rect 1106 69398 1110 69454
rect 1046 69394 1110 69398
rect 1126 69454 1190 69458
rect 1126 69398 1130 69454
rect 1130 69398 1186 69454
rect 1186 69398 1190 69454
rect 1126 69394 1190 69398
rect 84886 69454 84950 69458
rect 84886 69398 84890 69454
rect 84890 69398 84946 69454
rect 84946 69398 84950 69454
rect 84886 69394 84950 69398
rect 84966 69454 85030 69458
rect 84966 69398 84970 69454
rect 84970 69398 85026 69454
rect 85026 69398 85030 69454
rect 84966 69394 85030 69398
rect 85046 69454 85110 69458
rect 85046 69398 85050 69454
rect 85050 69398 85106 69454
rect 85106 69398 85110 69454
rect 85046 69394 85110 69398
rect 85126 69454 85190 69458
rect 85126 69398 85130 69454
rect 85130 69398 85186 69454
rect 85186 69398 85190 69454
rect 85126 69394 85190 69398
rect 2886 68910 2950 68914
rect 2886 68854 2890 68910
rect 2890 68854 2946 68910
rect 2946 68854 2950 68910
rect 2886 68850 2950 68854
rect 2966 68910 3030 68914
rect 2966 68854 2970 68910
rect 2970 68854 3026 68910
rect 3026 68854 3030 68910
rect 2966 68850 3030 68854
rect 3046 68910 3110 68914
rect 3046 68854 3050 68910
rect 3050 68854 3106 68910
rect 3106 68854 3110 68910
rect 3046 68850 3110 68854
rect 3126 68910 3190 68914
rect 3126 68854 3130 68910
rect 3130 68854 3186 68910
rect 3186 68854 3190 68910
rect 3126 68850 3190 68854
rect 86886 68910 86950 68914
rect 86886 68854 86890 68910
rect 86890 68854 86946 68910
rect 86946 68854 86950 68910
rect 86886 68850 86950 68854
rect 86966 68910 87030 68914
rect 86966 68854 86970 68910
rect 86970 68854 87026 68910
rect 87026 68854 87030 68910
rect 86966 68850 87030 68854
rect 87046 68910 87110 68914
rect 87046 68854 87050 68910
rect 87050 68854 87106 68910
rect 87106 68854 87110 68910
rect 87046 68850 87110 68854
rect 87126 68910 87190 68914
rect 87126 68854 87130 68910
rect 87130 68854 87186 68910
rect 87186 68854 87190 68910
rect 87126 68850 87190 68854
rect 886 68366 950 68370
rect 886 68310 890 68366
rect 890 68310 946 68366
rect 946 68310 950 68366
rect 886 68306 950 68310
rect 966 68366 1030 68370
rect 966 68310 970 68366
rect 970 68310 1026 68366
rect 1026 68310 1030 68366
rect 966 68306 1030 68310
rect 1046 68366 1110 68370
rect 1046 68310 1050 68366
rect 1050 68310 1106 68366
rect 1106 68310 1110 68366
rect 1046 68306 1110 68310
rect 1126 68366 1190 68370
rect 1126 68310 1130 68366
rect 1130 68310 1186 68366
rect 1186 68310 1190 68366
rect 1126 68306 1190 68310
rect 84886 68366 84950 68370
rect 84886 68310 84890 68366
rect 84890 68310 84946 68366
rect 84946 68310 84950 68366
rect 84886 68306 84950 68310
rect 84966 68366 85030 68370
rect 84966 68310 84970 68366
rect 84970 68310 85026 68366
rect 85026 68310 85030 68366
rect 84966 68306 85030 68310
rect 85046 68366 85110 68370
rect 85046 68310 85050 68366
rect 85050 68310 85106 68366
rect 85106 68310 85110 68366
rect 85046 68306 85110 68310
rect 85126 68366 85190 68370
rect 85126 68310 85130 68366
rect 85130 68310 85186 68366
rect 85186 68310 85190 68366
rect 85126 68306 85190 68310
rect 2886 67822 2950 67826
rect 2886 67766 2890 67822
rect 2890 67766 2946 67822
rect 2946 67766 2950 67822
rect 2886 67762 2950 67766
rect 2966 67822 3030 67826
rect 2966 67766 2970 67822
rect 2970 67766 3026 67822
rect 3026 67766 3030 67822
rect 2966 67762 3030 67766
rect 3046 67822 3110 67826
rect 3046 67766 3050 67822
rect 3050 67766 3106 67822
rect 3106 67766 3110 67822
rect 3046 67762 3110 67766
rect 3126 67822 3190 67826
rect 3126 67766 3130 67822
rect 3130 67766 3186 67822
rect 3186 67766 3190 67822
rect 3126 67762 3190 67766
rect 86886 67822 86950 67826
rect 86886 67766 86890 67822
rect 86890 67766 86946 67822
rect 86946 67766 86950 67822
rect 86886 67762 86950 67766
rect 86966 67822 87030 67826
rect 86966 67766 86970 67822
rect 86970 67766 87026 67822
rect 87026 67766 87030 67822
rect 86966 67762 87030 67766
rect 87046 67822 87110 67826
rect 87046 67766 87050 67822
rect 87050 67766 87106 67822
rect 87106 67766 87110 67822
rect 87046 67762 87110 67766
rect 87126 67822 87190 67826
rect 87126 67766 87130 67822
rect 87130 67766 87186 67822
rect 87186 67766 87190 67822
rect 87126 67762 87190 67766
rect 886 67278 950 67282
rect 886 67222 890 67278
rect 890 67222 946 67278
rect 946 67222 950 67278
rect 886 67218 950 67222
rect 966 67278 1030 67282
rect 966 67222 970 67278
rect 970 67222 1026 67278
rect 1026 67222 1030 67278
rect 966 67218 1030 67222
rect 1046 67278 1110 67282
rect 1046 67222 1050 67278
rect 1050 67222 1106 67278
rect 1106 67222 1110 67278
rect 1046 67218 1110 67222
rect 1126 67278 1190 67282
rect 1126 67222 1130 67278
rect 1130 67222 1186 67278
rect 1186 67222 1190 67278
rect 1126 67218 1190 67222
rect 84886 67278 84950 67282
rect 84886 67222 84890 67278
rect 84890 67222 84946 67278
rect 84946 67222 84950 67278
rect 84886 67218 84950 67222
rect 84966 67278 85030 67282
rect 84966 67222 84970 67278
rect 84970 67222 85026 67278
rect 85026 67222 85030 67278
rect 84966 67218 85030 67222
rect 85046 67278 85110 67282
rect 85046 67222 85050 67278
rect 85050 67222 85106 67278
rect 85106 67222 85110 67278
rect 85046 67218 85110 67222
rect 85126 67278 85190 67282
rect 85126 67222 85130 67278
rect 85130 67222 85186 67278
rect 85186 67222 85190 67278
rect 85126 67218 85190 67222
rect 2886 66734 2950 66738
rect 2886 66678 2890 66734
rect 2890 66678 2946 66734
rect 2946 66678 2950 66734
rect 2886 66674 2950 66678
rect 2966 66734 3030 66738
rect 2966 66678 2970 66734
rect 2970 66678 3026 66734
rect 3026 66678 3030 66734
rect 2966 66674 3030 66678
rect 3046 66734 3110 66738
rect 3046 66678 3050 66734
rect 3050 66678 3106 66734
rect 3106 66678 3110 66734
rect 3046 66674 3110 66678
rect 3126 66734 3190 66738
rect 3126 66678 3130 66734
rect 3130 66678 3186 66734
rect 3186 66678 3190 66734
rect 3126 66674 3190 66678
rect 86886 66734 86950 66738
rect 86886 66678 86890 66734
rect 86890 66678 86946 66734
rect 86946 66678 86950 66734
rect 86886 66674 86950 66678
rect 86966 66734 87030 66738
rect 86966 66678 86970 66734
rect 86970 66678 87026 66734
rect 87026 66678 87030 66734
rect 86966 66674 87030 66678
rect 87046 66734 87110 66738
rect 87046 66678 87050 66734
rect 87050 66678 87106 66734
rect 87106 66678 87110 66734
rect 87046 66674 87110 66678
rect 87126 66734 87190 66738
rect 87126 66678 87130 66734
rect 87130 66678 87186 66734
rect 87186 66678 87190 66734
rect 87126 66674 87190 66678
rect 886 66190 950 66194
rect 886 66134 890 66190
rect 890 66134 946 66190
rect 946 66134 950 66190
rect 886 66130 950 66134
rect 966 66190 1030 66194
rect 966 66134 970 66190
rect 970 66134 1026 66190
rect 1026 66134 1030 66190
rect 966 66130 1030 66134
rect 1046 66190 1110 66194
rect 1046 66134 1050 66190
rect 1050 66134 1106 66190
rect 1106 66134 1110 66190
rect 1046 66130 1110 66134
rect 1126 66190 1190 66194
rect 1126 66134 1130 66190
rect 1130 66134 1186 66190
rect 1186 66134 1190 66190
rect 1126 66130 1190 66134
rect 84886 66190 84950 66194
rect 84886 66134 84890 66190
rect 84890 66134 84946 66190
rect 84946 66134 84950 66190
rect 84886 66130 84950 66134
rect 84966 66190 85030 66194
rect 84966 66134 84970 66190
rect 84970 66134 85026 66190
rect 85026 66134 85030 66190
rect 84966 66130 85030 66134
rect 85046 66190 85110 66194
rect 85046 66134 85050 66190
rect 85050 66134 85106 66190
rect 85106 66134 85110 66190
rect 85046 66130 85110 66134
rect 85126 66190 85190 66194
rect 85126 66134 85130 66190
rect 85130 66134 85186 66190
rect 85186 66134 85190 66190
rect 85126 66130 85190 66134
rect 2886 65646 2950 65650
rect 2886 65590 2890 65646
rect 2890 65590 2946 65646
rect 2946 65590 2950 65646
rect 2886 65586 2950 65590
rect 2966 65646 3030 65650
rect 2966 65590 2970 65646
rect 2970 65590 3026 65646
rect 3026 65590 3030 65646
rect 2966 65586 3030 65590
rect 3046 65646 3110 65650
rect 3046 65590 3050 65646
rect 3050 65590 3106 65646
rect 3106 65590 3110 65646
rect 3046 65586 3110 65590
rect 3126 65646 3190 65650
rect 3126 65590 3130 65646
rect 3130 65590 3186 65646
rect 3186 65590 3190 65646
rect 3126 65586 3190 65590
rect 86886 65646 86950 65650
rect 86886 65590 86890 65646
rect 86890 65590 86946 65646
rect 86946 65590 86950 65646
rect 86886 65586 86950 65590
rect 86966 65646 87030 65650
rect 86966 65590 86970 65646
rect 86970 65590 87026 65646
rect 87026 65590 87030 65646
rect 86966 65586 87030 65590
rect 87046 65646 87110 65650
rect 87046 65590 87050 65646
rect 87050 65590 87106 65646
rect 87106 65590 87110 65646
rect 87046 65586 87110 65590
rect 87126 65646 87190 65650
rect 87126 65590 87130 65646
rect 87130 65590 87186 65646
rect 87186 65590 87190 65646
rect 87126 65586 87190 65590
rect 4514 65518 4578 65582
rect 4698 65246 4762 65310
rect 886 65102 950 65106
rect 886 65046 890 65102
rect 890 65046 946 65102
rect 946 65046 950 65102
rect 886 65042 950 65046
rect 966 65102 1030 65106
rect 966 65046 970 65102
rect 970 65046 1026 65102
rect 1026 65046 1030 65102
rect 966 65042 1030 65046
rect 1046 65102 1110 65106
rect 1046 65046 1050 65102
rect 1050 65046 1106 65102
rect 1106 65046 1110 65102
rect 1046 65042 1110 65046
rect 1126 65102 1190 65106
rect 1126 65046 1130 65102
rect 1130 65046 1186 65102
rect 1186 65046 1190 65102
rect 1126 65042 1190 65046
rect 84886 65102 84950 65106
rect 84886 65046 84890 65102
rect 84890 65046 84946 65102
rect 84946 65046 84950 65102
rect 84886 65042 84950 65046
rect 84966 65102 85030 65106
rect 84966 65046 84970 65102
rect 84970 65046 85026 65102
rect 85026 65046 85030 65102
rect 84966 65042 85030 65046
rect 85046 65102 85110 65106
rect 85046 65046 85050 65102
rect 85050 65046 85106 65102
rect 85106 65046 85110 65102
rect 85046 65042 85110 65046
rect 85126 65102 85190 65106
rect 85126 65046 85130 65102
rect 85130 65046 85186 65102
rect 85186 65046 85190 65102
rect 85126 65042 85190 65046
rect 2886 64558 2950 64562
rect 2886 64502 2890 64558
rect 2890 64502 2946 64558
rect 2946 64502 2950 64558
rect 2886 64498 2950 64502
rect 2966 64558 3030 64562
rect 2966 64502 2970 64558
rect 2970 64502 3026 64558
rect 3026 64502 3030 64558
rect 2966 64498 3030 64502
rect 3046 64558 3110 64562
rect 3046 64502 3050 64558
rect 3050 64502 3106 64558
rect 3106 64502 3110 64558
rect 3046 64498 3110 64502
rect 3126 64558 3190 64562
rect 3126 64502 3130 64558
rect 3130 64502 3186 64558
rect 3186 64502 3190 64558
rect 3126 64498 3190 64502
rect 86886 64558 86950 64562
rect 86886 64502 86890 64558
rect 86890 64502 86946 64558
rect 86946 64502 86950 64558
rect 86886 64498 86950 64502
rect 86966 64558 87030 64562
rect 86966 64502 86970 64558
rect 86970 64502 87026 64558
rect 87026 64502 87030 64558
rect 86966 64498 87030 64502
rect 87046 64558 87110 64562
rect 87046 64502 87050 64558
rect 87050 64502 87106 64558
rect 87106 64502 87110 64558
rect 87046 64498 87110 64502
rect 87126 64558 87190 64562
rect 87126 64502 87130 64558
rect 87130 64502 87186 64558
rect 87186 64502 87190 64558
rect 87126 64498 87190 64502
rect 886 64014 950 64018
rect 886 63958 890 64014
rect 890 63958 946 64014
rect 946 63958 950 64014
rect 886 63954 950 63958
rect 966 64014 1030 64018
rect 966 63958 970 64014
rect 970 63958 1026 64014
rect 1026 63958 1030 64014
rect 966 63954 1030 63958
rect 1046 64014 1110 64018
rect 1046 63958 1050 64014
rect 1050 63958 1106 64014
rect 1106 63958 1110 64014
rect 1046 63954 1110 63958
rect 1126 64014 1190 64018
rect 1126 63958 1130 64014
rect 1130 63958 1186 64014
rect 1186 63958 1190 64014
rect 1126 63954 1190 63958
rect 84886 64014 84950 64018
rect 84886 63958 84890 64014
rect 84890 63958 84946 64014
rect 84946 63958 84950 64014
rect 84886 63954 84950 63958
rect 84966 64014 85030 64018
rect 84966 63958 84970 64014
rect 84970 63958 85026 64014
rect 85026 63958 85030 64014
rect 84966 63954 85030 63958
rect 85046 64014 85110 64018
rect 85046 63958 85050 64014
rect 85050 63958 85106 64014
rect 85106 63958 85110 64014
rect 85046 63954 85110 63958
rect 85126 64014 85190 64018
rect 85126 63958 85130 64014
rect 85130 63958 85186 64014
rect 85186 63958 85190 64014
rect 85126 63954 85190 63958
rect 2886 63470 2950 63474
rect 2886 63414 2890 63470
rect 2890 63414 2946 63470
rect 2946 63414 2950 63470
rect 2886 63410 2950 63414
rect 2966 63470 3030 63474
rect 2966 63414 2970 63470
rect 2970 63414 3026 63470
rect 3026 63414 3030 63470
rect 2966 63410 3030 63414
rect 3046 63470 3110 63474
rect 3046 63414 3050 63470
rect 3050 63414 3106 63470
rect 3106 63414 3110 63470
rect 3046 63410 3110 63414
rect 3126 63470 3190 63474
rect 3126 63414 3130 63470
rect 3130 63414 3186 63470
rect 3186 63414 3190 63470
rect 3126 63410 3190 63414
rect 86886 63470 86950 63474
rect 86886 63414 86890 63470
rect 86890 63414 86946 63470
rect 86946 63414 86950 63470
rect 86886 63410 86950 63414
rect 86966 63470 87030 63474
rect 86966 63414 86970 63470
rect 86970 63414 87026 63470
rect 87026 63414 87030 63470
rect 86966 63410 87030 63414
rect 87046 63470 87110 63474
rect 87046 63414 87050 63470
rect 87050 63414 87106 63470
rect 87106 63414 87110 63470
rect 87046 63410 87110 63414
rect 87126 63470 87190 63474
rect 87126 63414 87130 63470
rect 87130 63414 87186 63470
rect 87186 63414 87190 63470
rect 87126 63410 87190 63414
rect 886 62926 950 62930
rect 886 62870 890 62926
rect 890 62870 946 62926
rect 946 62870 950 62926
rect 886 62866 950 62870
rect 966 62926 1030 62930
rect 966 62870 970 62926
rect 970 62870 1026 62926
rect 1026 62870 1030 62926
rect 966 62866 1030 62870
rect 1046 62926 1110 62930
rect 1046 62870 1050 62926
rect 1050 62870 1106 62926
rect 1106 62870 1110 62926
rect 1046 62866 1110 62870
rect 1126 62926 1190 62930
rect 1126 62870 1130 62926
rect 1130 62870 1186 62926
rect 1186 62870 1190 62926
rect 1126 62866 1190 62870
rect 84886 62926 84950 62930
rect 84886 62870 84890 62926
rect 84890 62870 84946 62926
rect 84946 62870 84950 62926
rect 84886 62866 84950 62870
rect 84966 62926 85030 62930
rect 84966 62870 84970 62926
rect 84970 62870 85026 62926
rect 85026 62870 85030 62926
rect 84966 62866 85030 62870
rect 85046 62926 85110 62930
rect 85046 62870 85050 62926
rect 85050 62870 85106 62926
rect 85106 62870 85110 62926
rect 85046 62866 85110 62870
rect 85126 62926 85190 62930
rect 85126 62870 85130 62926
rect 85130 62870 85186 62926
rect 85186 62870 85190 62926
rect 85126 62866 85190 62870
rect 2886 62382 2950 62386
rect 2886 62326 2890 62382
rect 2890 62326 2946 62382
rect 2946 62326 2950 62382
rect 2886 62322 2950 62326
rect 2966 62382 3030 62386
rect 2966 62326 2970 62382
rect 2970 62326 3026 62382
rect 3026 62326 3030 62382
rect 2966 62322 3030 62326
rect 3046 62382 3110 62386
rect 3046 62326 3050 62382
rect 3050 62326 3106 62382
rect 3106 62326 3110 62382
rect 3046 62322 3110 62326
rect 3126 62382 3190 62386
rect 3126 62326 3130 62382
rect 3130 62326 3186 62382
rect 3186 62326 3190 62382
rect 3126 62322 3190 62326
rect 86886 62382 86950 62386
rect 86886 62326 86890 62382
rect 86890 62326 86946 62382
rect 86946 62326 86950 62382
rect 86886 62322 86950 62326
rect 86966 62382 87030 62386
rect 86966 62326 86970 62382
rect 86970 62326 87026 62382
rect 87026 62326 87030 62382
rect 86966 62322 87030 62326
rect 87046 62382 87110 62386
rect 87046 62326 87050 62382
rect 87050 62326 87106 62382
rect 87106 62326 87110 62382
rect 87046 62322 87110 62326
rect 87126 62382 87190 62386
rect 87126 62326 87130 62382
rect 87130 62326 87186 62382
rect 87186 62326 87190 62382
rect 87126 62322 87190 62326
rect 886 61838 950 61842
rect 886 61782 890 61838
rect 890 61782 946 61838
rect 946 61782 950 61838
rect 886 61778 950 61782
rect 966 61838 1030 61842
rect 966 61782 970 61838
rect 970 61782 1026 61838
rect 1026 61782 1030 61838
rect 966 61778 1030 61782
rect 1046 61838 1110 61842
rect 1046 61782 1050 61838
rect 1050 61782 1106 61838
rect 1106 61782 1110 61838
rect 1046 61778 1110 61782
rect 1126 61838 1190 61842
rect 1126 61782 1130 61838
rect 1130 61782 1186 61838
rect 1186 61782 1190 61838
rect 1126 61778 1190 61782
rect 84886 61838 84950 61842
rect 84886 61782 84890 61838
rect 84890 61782 84946 61838
rect 84946 61782 84950 61838
rect 84886 61778 84950 61782
rect 84966 61838 85030 61842
rect 84966 61782 84970 61838
rect 84970 61782 85026 61838
rect 85026 61782 85030 61838
rect 84966 61778 85030 61782
rect 85046 61838 85110 61842
rect 85046 61782 85050 61838
rect 85050 61782 85106 61838
rect 85106 61782 85110 61838
rect 85046 61778 85110 61782
rect 85126 61838 85190 61842
rect 85126 61782 85130 61838
rect 85130 61782 85186 61838
rect 85186 61782 85190 61838
rect 85126 61778 85190 61782
rect 2886 61294 2950 61298
rect 2886 61238 2890 61294
rect 2890 61238 2946 61294
rect 2946 61238 2950 61294
rect 2886 61234 2950 61238
rect 2966 61294 3030 61298
rect 2966 61238 2970 61294
rect 2970 61238 3026 61294
rect 3026 61238 3030 61294
rect 2966 61234 3030 61238
rect 3046 61294 3110 61298
rect 3046 61238 3050 61294
rect 3050 61238 3106 61294
rect 3106 61238 3110 61294
rect 3046 61234 3110 61238
rect 3126 61294 3190 61298
rect 3126 61238 3130 61294
rect 3130 61238 3186 61294
rect 3186 61238 3190 61294
rect 3126 61234 3190 61238
rect 86886 61294 86950 61298
rect 86886 61238 86890 61294
rect 86890 61238 86946 61294
rect 86946 61238 86950 61294
rect 86886 61234 86950 61238
rect 86966 61294 87030 61298
rect 86966 61238 86970 61294
rect 86970 61238 87026 61294
rect 87026 61238 87030 61294
rect 86966 61234 87030 61238
rect 87046 61294 87110 61298
rect 87046 61238 87050 61294
rect 87050 61238 87106 61294
rect 87106 61238 87110 61294
rect 87046 61234 87110 61238
rect 87126 61294 87190 61298
rect 87126 61238 87130 61294
rect 87130 61238 87186 61294
rect 87186 61238 87190 61294
rect 87126 61234 87190 61238
rect 886 60750 950 60754
rect 886 60694 890 60750
rect 890 60694 946 60750
rect 946 60694 950 60750
rect 886 60690 950 60694
rect 966 60750 1030 60754
rect 966 60694 970 60750
rect 970 60694 1026 60750
rect 1026 60694 1030 60750
rect 966 60690 1030 60694
rect 1046 60750 1110 60754
rect 1046 60694 1050 60750
rect 1050 60694 1106 60750
rect 1106 60694 1110 60750
rect 1046 60690 1110 60694
rect 1126 60750 1190 60754
rect 1126 60694 1130 60750
rect 1130 60694 1186 60750
rect 1186 60694 1190 60750
rect 1126 60690 1190 60694
rect 84886 60750 84950 60754
rect 84886 60694 84890 60750
rect 84890 60694 84946 60750
rect 84946 60694 84950 60750
rect 84886 60690 84950 60694
rect 84966 60750 85030 60754
rect 84966 60694 84970 60750
rect 84970 60694 85026 60750
rect 85026 60694 85030 60750
rect 84966 60690 85030 60694
rect 85046 60750 85110 60754
rect 85046 60694 85050 60750
rect 85050 60694 85106 60750
rect 85106 60694 85110 60750
rect 85046 60690 85110 60694
rect 85126 60750 85190 60754
rect 85126 60694 85130 60750
rect 85130 60694 85186 60750
rect 85186 60694 85190 60750
rect 85126 60690 85190 60694
rect 2886 60206 2950 60210
rect 2886 60150 2890 60206
rect 2890 60150 2946 60206
rect 2946 60150 2950 60206
rect 2886 60146 2950 60150
rect 2966 60206 3030 60210
rect 2966 60150 2970 60206
rect 2970 60150 3026 60206
rect 3026 60150 3030 60206
rect 2966 60146 3030 60150
rect 3046 60206 3110 60210
rect 3046 60150 3050 60206
rect 3050 60150 3106 60206
rect 3106 60150 3110 60206
rect 3046 60146 3110 60150
rect 3126 60206 3190 60210
rect 3126 60150 3130 60206
rect 3130 60150 3186 60206
rect 3186 60150 3190 60206
rect 3126 60146 3190 60150
rect 86886 60206 86950 60210
rect 86886 60150 86890 60206
rect 86890 60150 86946 60206
rect 86946 60150 86950 60206
rect 86886 60146 86950 60150
rect 86966 60206 87030 60210
rect 86966 60150 86970 60206
rect 86970 60150 87026 60206
rect 87026 60150 87030 60206
rect 86966 60146 87030 60150
rect 87046 60206 87110 60210
rect 87046 60150 87050 60206
rect 87050 60150 87106 60206
rect 87106 60150 87110 60206
rect 87046 60146 87110 60150
rect 87126 60206 87190 60210
rect 87126 60150 87130 60206
rect 87130 60150 87186 60206
rect 87186 60150 87190 60206
rect 87126 60146 87190 60150
rect 886 59662 950 59666
rect 886 59606 890 59662
rect 890 59606 946 59662
rect 946 59606 950 59662
rect 886 59602 950 59606
rect 966 59662 1030 59666
rect 966 59606 970 59662
rect 970 59606 1026 59662
rect 1026 59606 1030 59662
rect 966 59602 1030 59606
rect 1046 59662 1110 59666
rect 1046 59606 1050 59662
rect 1050 59606 1106 59662
rect 1106 59606 1110 59662
rect 1046 59602 1110 59606
rect 1126 59662 1190 59666
rect 1126 59606 1130 59662
rect 1130 59606 1186 59662
rect 1186 59606 1190 59662
rect 1126 59602 1190 59606
rect 84886 59662 84950 59666
rect 84886 59606 84890 59662
rect 84890 59606 84946 59662
rect 84946 59606 84950 59662
rect 84886 59602 84950 59606
rect 84966 59662 85030 59666
rect 84966 59606 84970 59662
rect 84970 59606 85026 59662
rect 85026 59606 85030 59662
rect 84966 59602 85030 59606
rect 85046 59662 85110 59666
rect 85046 59606 85050 59662
rect 85050 59606 85106 59662
rect 85106 59606 85110 59662
rect 85046 59602 85110 59606
rect 85126 59662 85190 59666
rect 85126 59606 85130 59662
rect 85130 59606 85186 59662
rect 85186 59606 85190 59662
rect 85126 59602 85190 59606
rect 83266 59262 83330 59326
rect 2886 59118 2950 59122
rect 2886 59062 2890 59118
rect 2890 59062 2946 59118
rect 2946 59062 2950 59118
rect 2886 59058 2950 59062
rect 2966 59118 3030 59122
rect 2966 59062 2970 59118
rect 2970 59062 3026 59118
rect 3026 59062 3030 59118
rect 2966 59058 3030 59062
rect 3046 59118 3110 59122
rect 3046 59062 3050 59118
rect 3050 59062 3106 59118
rect 3106 59062 3110 59118
rect 3046 59058 3110 59062
rect 3126 59118 3190 59122
rect 3126 59062 3130 59118
rect 3130 59062 3186 59118
rect 3186 59062 3190 59118
rect 3126 59058 3190 59062
rect 86886 59118 86950 59122
rect 86886 59062 86890 59118
rect 86890 59062 86946 59118
rect 86946 59062 86950 59118
rect 86886 59058 86950 59062
rect 86966 59118 87030 59122
rect 86966 59062 86970 59118
rect 86970 59062 87026 59118
rect 87026 59062 87030 59118
rect 86966 59058 87030 59062
rect 87046 59118 87110 59122
rect 87046 59062 87050 59118
rect 87050 59062 87106 59118
rect 87106 59062 87110 59118
rect 87046 59058 87110 59062
rect 87126 59118 87190 59122
rect 87126 59062 87130 59118
rect 87130 59062 87186 59118
rect 87186 59062 87190 59118
rect 87126 59058 87190 59062
rect 886 58574 950 58578
rect 886 58518 890 58574
rect 890 58518 946 58574
rect 946 58518 950 58574
rect 886 58514 950 58518
rect 966 58574 1030 58578
rect 966 58518 970 58574
rect 970 58518 1026 58574
rect 1026 58518 1030 58574
rect 966 58514 1030 58518
rect 1046 58574 1110 58578
rect 1046 58518 1050 58574
rect 1050 58518 1106 58574
rect 1106 58518 1110 58574
rect 1046 58514 1110 58518
rect 1126 58574 1190 58578
rect 1126 58518 1130 58574
rect 1130 58518 1186 58574
rect 1186 58518 1190 58574
rect 1126 58514 1190 58518
rect 84886 58574 84950 58578
rect 84886 58518 84890 58574
rect 84890 58518 84946 58574
rect 84946 58518 84950 58574
rect 84886 58514 84950 58518
rect 84966 58574 85030 58578
rect 84966 58518 84970 58574
rect 84970 58518 85026 58574
rect 85026 58518 85030 58574
rect 84966 58514 85030 58518
rect 85046 58574 85110 58578
rect 85046 58518 85050 58574
rect 85050 58518 85106 58574
rect 85106 58518 85110 58574
rect 85046 58514 85110 58518
rect 85126 58574 85190 58578
rect 85126 58518 85130 58574
rect 85130 58518 85186 58574
rect 85186 58518 85190 58574
rect 85126 58514 85190 58518
rect 2886 58030 2950 58034
rect 2886 57974 2890 58030
rect 2890 57974 2946 58030
rect 2946 57974 2950 58030
rect 2886 57970 2950 57974
rect 2966 58030 3030 58034
rect 2966 57974 2970 58030
rect 2970 57974 3026 58030
rect 3026 57974 3030 58030
rect 2966 57970 3030 57974
rect 3046 58030 3110 58034
rect 3046 57974 3050 58030
rect 3050 57974 3106 58030
rect 3106 57974 3110 58030
rect 3046 57970 3110 57974
rect 3126 58030 3190 58034
rect 3126 57974 3130 58030
rect 3130 57974 3186 58030
rect 3186 57974 3190 58030
rect 3126 57970 3190 57974
rect 86886 58030 86950 58034
rect 86886 57974 86890 58030
rect 86890 57974 86946 58030
rect 86946 57974 86950 58030
rect 86886 57970 86950 57974
rect 86966 58030 87030 58034
rect 86966 57974 86970 58030
rect 86970 57974 87026 58030
rect 87026 57974 87030 58030
rect 86966 57970 87030 57974
rect 87046 58030 87110 58034
rect 87046 57974 87050 58030
rect 87050 57974 87106 58030
rect 87106 57974 87110 58030
rect 87046 57970 87110 57974
rect 87126 58030 87190 58034
rect 87126 57974 87130 58030
rect 87130 57974 87186 58030
rect 87186 57974 87190 58030
rect 87126 57970 87190 57974
rect 84554 57766 84618 57830
rect 886 57486 950 57490
rect 886 57430 890 57486
rect 890 57430 946 57486
rect 946 57430 950 57486
rect 886 57426 950 57430
rect 966 57486 1030 57490
rect 966 57430 970 57486
rect 970 57430 1026 57486
rect 1026 57430 1030 57486
rect 966 57426 1030 57430
rect 1046 57486 1110 57490
rect 1046 57430 1050 57486
rect 1050 57430 1106 57486
rect 1106 57430 1110 57486
rect 1046 57426 1110 57430
rect 1126 57486 1190 57490
rect 1126 57430 1130 57486
rect 1130 57430 1186 57486
rect 1186 57430 1190 57486
rect 1126 57426 1190 57430
rect 84886 57486 84950 57490
rect 84886 57430 84890 57486
rect 84890 57430 84946 57486
rect 84946 57430 84950 57486
rect 84886 57426 84950 57430
rect 84966 57486 85030 57490
rect 84966 57430 84970 57486
rect 84970 57430 85026 57486
rect 85026 57430 85030 57486
rect 84966 57426 85030 57430
rect 85046 57486 85110 57490
rect 85046 57430 85050 57486
rect 85050 57430 85106 57486
rect 85106 57430 85110 57486
rect 85046 57426 85110 57430
rect 85126 57486 85190 57490
rect 85126 57430 85130 57486
rect 85130 57430 85186 57486
rect 85186 57430 85190 57486
rect 85126 57426 85190 57430
rect 2886 56942 2950 56946
rect 2886 56886 2890 56942
rect 2890 56886 2946 56942
rect 2946 56886 2950 56942
rect 2886 56882 2950 56886
rect 2966 56942 3030 56946
rect 2966 56886 2970 56942
rect 2970 56886 3026 56942
rect 3026 56886 3030 56942
rect 2966 56882 3030 56886
rect 3046 56942 3110 56946
rect 3046 56886 3050 56942
rect 3050 56886 3106 56942
rect 3106 56886 3110 56942
rect 3046 56882 3110 56886
rect 3126 56942 3190 56946
rect 3126 56886 3130 56942
rect 3130 56886 3186 56942
rect 3186 56886 3190 56942
rect 3126 56882 3190 56886
rect 86886 56942 86950 56946
rect 86886 56886 86890 56942
rect 86890 56886 86946 56942
rect 86946 56886 86950 56942
rect 86886 56882 86950 56886
rect 86966 56942 87030 56946
rect 86966 56886 86970 56942
rect 86970 56886 87026 56942
rect 87026 56886 87030 56942
rect 86966 56882 87030 56886
rect 87046 56942 87110 56946
rect 87046 56886 87050 56942
rect 87050 56886 87106 56942
rect 87106 56886 87110 56942
rect 87046 56882 87110 56886
rect 87126 56942 87190 56946
rect 87126 56886 87130 56942
rect 87130 56886 87186 56942
rect 87186 56886 87190 56942
rect 87126 56882 87190 56886
rect 886 56398 950 56402
rect 886 56342 890 56398
rect 890 56342 946 56398
rect 946 56342 950 56398
rect 886 56338 950 56342
rect 966 56398 1030 56402
rect 966 56342 970 56398
rect 970 56342 1026 56398
rect 1026 56342 1030 56398
rect 966 56338 1030 56342
rect 1046 56398 1110 56402
rect 1046 56342 1050 56398
rect 1050 56342 1106 56398
rect 1106 56342 1110 56398
rect 1046 56338 1110 56342
rect 1126 56398 1190 56402
rect 1126 56342 1130 56398
rect 1130 56342 1186 56398
rect 1186 56342 1190 56398
rect 1126 56338 1190 56342
rect 84886 56398 84950 56402
rect 84886 56342 84890 56398
rect 84890 56342 84946 56398
rect 84946 56342 84950 56398
rect 84886 56338 84950 56342
rect 84966 56398 85030 56402
rect 84966 56342 84970 56398
rect 84970 56342 85026 56398
rect 85026 56342 85030 56398
rect 84966 56338 85030 56342
rect 85046 56398 85110 56402
rect 85046 56342 85050 56398
rect 85050 56342 85106 56398
rect 85106 56342 85110 56398
rect 85046 56338 85110 56342
rect 85126 56398 85190 56402
rect 85126 56342 85130 56398
rect 85130 56342 85186 56398
rect 85186 56342 85190 56398
rect 85126 56338 85190 56342
rect 2886 55854 2950 55858
rect 2886 55798 2890 55854
rect 2890 55798 2946 55854
rect 2946 55798 2950 55854
rect 2886 55794 2950 55798
rect 2966 55854 3030 55858
rect 2966 55798 2970 55854
rect 2970 55798 3026 55854
rect 3026 55798 3030 55854
rect 2966 55794 3030 55798
rect 3046 55854 3110 55858
rect 3046 55798 3050 55854
rect 3050 55798 3106 55854
rect 3106 55798 3110 55854
rect 3046 55794 3110 55798
rect 3126 55854 3190 55858
rect 3126 55798 3130 55854
rect 3130 55798 3186 55854
rect 3186 55798 3190 55854
rect 3126 55794 3190 55798
rect 86886 55854 86950 55858
rect 86886 55798 86890 55854
rect 86890 55798 86946 55854
rect 86946 55798 86950 55854
rect 86886 55794 86950 55798
rect 86966 55854 87030 55858
rect 86966 55798 86970 55854
rect 86970 55798 87026 55854
rect 87026 55798 87030 55854
rect 86966 55794 87030 55798
rect 87046 55854 87110 55858
rect 87046 55798 87050 55854
rect 87050 55798 87106 55854
rect 87106 55798 87110 55854
rect 87046 55794 87110 55798
rect 87126 55854 87190 55858
rect 87126 55798 87130 55854
rect 87130 55798 87186 55854
rect 87186 55798 87190 55854
rect 87126 55794 87190 55798
rect 886 55310 950 55314
rect 886 55254 890 55310
rect 890 55254 946 55310
rect 946 55254 950 55310
rect 886 55250 950 55254
rect 966 55310 1030 55314
rect 966 55254 970 55310
rect 970 55254 1026 55310
rect 1026 55254 1030 55310
rect 966 55250 1030 55254
rect 1046 55310 1110 55314
rect 1046 55254 1050 55310
rect 1050 55254 1106 55310
rect 1106 55254 1110 55310
rect 1046 55250 1110 55254
rect 1126 55310 1190 55314
rect 1126 55254 1130 55310
rect 1130 55254 1186 55310
rect 1186 55254 1190 55310
rect 1126 55250 1190 55254
rect 84886 55310 84950 55314
rect 84886 55254 84890 55310
rect 84890 55254 84946 55310
rect 84946 55254 84950 55310
rect 84886 55250 84950 55254
rect 84966 55310 85030 55314
rect 84966 55254 84970 55310
rect 84970 55254 85026 55310
rect 85026 55254 85030 55310
rect 84966 55250 85030 55254
rect 85046 55310 85110 55314
rect 85046 55254 85050 55310
rect 85050 55254 85106 55310
rect 85106 55254 85110 55310
rect 85046 55250 85110 55254
rect 85126 55310 85190 55314
rect 85126 55254 85130 55310
rect 85130 55254 85186 55310
rect 85186 55254 85190 55310
rect 85126 55250 85190 55254
rect 83450 55182 83514 55246
rect 2886 54766 2950 54770
rect 2886 54710 2890 54766
rect 2890 54710 2946 54766
rect 2946 54710 2950 54766
rect 2886 54706 2950 54710
rect 2966 54766 3030 54770
rect 2966 54710 2970 54766
rect 2970 54710 3026 54766
rect 3026 54710 3030 54766
rect 2966 54706 3030 54710
rect 3046 54766 3110 54770
rect 3046 54710 3050 54766
rect 3050 54710 3106 54766
rect 3106 54710 3110 54766
rect 3046 54706 3110 54710
rect 3126 54766 3190 54770
rect 3126 54710 3130 54766
rect 3130 54710 3186 54766
rect 3186 54710 3190 54766
rect 3126 54706 3190 54710
rect 86886 54766 86950 54770
rect 86886 54710 86890 54766
rect 86890 54710 86946 54766
rect 86946 54710 86950 54766
rect 86886 54706 86950 54710
rect 86966 54766 87030 54770
rect 86966 54710 86970 54766
rect 86970 54710 87026 54766
rect 87026 54710 87030 54766
rect 86966 54706 87030 54710
rect 87046 54766 87110 54770
rect 87046 54710 87050 54766
rect 87050 54710 87106 54766
rect 87106 54710 87110 54766
rect 87046 54706 87110 54710
rect 87126 54766 87190 54770
rect 87126 54710 87130 54766
rect 87130 54710 87186 54766
rect 87186 54710 87190 54766
rect 87126 54706 87190 54710
rect 886 54222 950 54226
rect 886 54166 890 54222
rect 890 54166 946 54222
rect 946 54166 950 54222
rect 886 54162 950 54166
rect 966 54222 1030 54226
rect 966 54166 970 54222
rect 970 54166 1026 54222
rect 1026 54166 1030 54222
rect 966 54162 1030 54166
rect 1046 54222 1110 54226
rect 1046 54166 1050 54222
rect 1050 54166 1106 54222
rect 1106 54166 1110 54222
rect 1046 54162 1110 54166
rect 1126 54222 1190 54226
rect 1126 54166 1130 54222
rect 1130 54166 1186 54222
rect 1186 54166 1190 54222
rect 1126 54162 1190 54166
rect 84886 54222 84950 54226
rect 84886 54166 84890 54222
rect 84890 54166 84946 54222
rect 84946 54166 84950 54222
rect 84886 54162 84950 54166
rect 84966 54222 85030 54226
rect 84966 54166 84970 54222
rect 84970 54166 85026 54222
rect 85026 54166 85030 54222
rect 84966 54162 85030 54166
rect 85046 54222 85110 54226
rect 85046 54166 85050 54222
rect 85050 54166 85106 54222
rect 85106 54166 85110 54222
rect 85046 54162 85110 54166
rect 85126 54222 85190 54226
rect 85126 54166 85130 54222
rect 85130 54166 85186 54222
rect 85186 54166 85190 54222
rect 85126 54162 85190 54166
rect 2886 53678 2950 53682
rect 2886 53622 2890 53678
rect 2890 53622 2946 53678
rect 2946 53622 2950 53678
rect 2886 53618 2950 53622
rect 2966 53678 3030 53682
rect 2966 53622 2970 53678
rect 2970 53622 3026 53678
rect 3026 53622 3030 53678
rect 2966 53618 3030 53622
rect 3046 53678 3110 53682
rect 3046 53622 3050 53678
rect 3050 53622 3106 53678
rect 3106 53622 3110 53678
rect 3046 53618 3110 53622
rect 3126 53678 3190 53682
rect 3126 53622 3130 53678
rect 3130 53622 3186 53678
rect 3186 53622 3190 53678
rect 3126 53618 3190 53622
rect 86886 53678 86950 53682
rect 86886 53622 86890 53678
rect 86890 53622 86946 53678
rect 86946 53622 86950 53678
rect 86886 53618 86950 53622
rect 86966 53678 87030 53682
rect 86966 53622 86970 53678
rect 86970 53622 87026 53678
rect 87026 53622 87030 53678
rect 86966 53618 87030 53622
rect 87046 53678 87110 53682
rect 87046 53622 87050 53678
rect 87050 53622 87106 53678
rect 87106 53622 87110 53678
rect 87046 53618 87110 53622
rect 87126 53678 87190 53682
rect 87126 53622 87130 53678
rect 87130 53622 87186 53678
rect 87186 53622 87190 53678
rect 87126 53618 87190 53622
rect 886 53134 950 53138
rect 886 53078 890 53134
rect 890 53078 946 53134
rect 946 53078 950 53134
rect 886 53074 950 53078
rect 966 53134 1030 53138
rect 966 53078 970 53134
rect 970 53078 1026 53134
rect 1026 53078 1030 53134
rect 966 53074 1030 53078
rect 1046 53134 1110 53138
rect 1046 53078 1050 53134
rect 1050 53078 1106 53134
rect 1106 53078 1110 53134
rect 1046 53074 1110 53078
rect 1126 53134 1190 53138
rect 1126 53078 1130 53134
rect 1130 53078 1186 53134
rect 1186 53078 1190 53134
rect 1126 53074 1190 53078
rect 84886 53134 84950 53138
rect 84886 53078 84890 53134
rect 84890 53078 84946 53134
rect 84946 53078 84950 53134
rect 84886 53074 84950 53078
rect 84966 53134 85030 53138
rect 84966 53078 84970 53134
rect 84970 53078 85026 53134
rect 85026 53078 85030 53134
rect 84966 53074 85030 53078
rect 85046 53134 85110 53138
rect 85046 53078 85050 53134
rect 85050 53078 85106 53134
rect 85106 53078 85110 53134
rect 85046 53074 85110 53078
rect 85126 53134 85190 53138
rect 85126 53078 85130 53134
rect 85130 53078 85186 53134
rect 85186 53078 85190 53134
rect 85126 53074 85190 53078
rect 2886 52590 2950 52594
rect 2886 52534 2890 52590
rect 2890 52534 2946 52590
rect 2946 52534 2950 52590
rect 2886 52530 2950 52534
rect 2966 52590 3030 52594
rect 2966 52534 2970 52590
rect 2970 52534 3026 52590
rect 3026 52534 3030 52590
rect 2966 52530 3030 52534
rect 3046 52590 3110 52594
rect 3046 52534 3050 52590
rect 3050 52534 3106 52590
rect 3106 52534 3110 52590
rect 3046 52530 3110 52534
rect 3126 52590 3190 52594
rect 3126 52534 3130 52590
rect 3130 52534 3186 52590
rect 3186 52534 3190 52590
rect 3126 52530 3190 52534
rect 86886 52590 86950 52594
rect 86886 52534 86890 52590
rect 86890 52534 86946 52590
rect 86946 52534 86950 52590
rect 86886 52530 86950 52534
rect 86966 52590 87030 52594
rect 86966 52534 86970 52590
rect 86970 52534 87026 52590
rect 87026 52534 87030 52590
rect 86966 52530 87030 52534
rect 87046 52590 87110 52594
rect 87046 52534 87050 52590
rect 87050 52534 87106 52590
rect 87106 52534 87110 52590
rect 87046 52530 87110 52534
rect 87126 52590 87190 52594
rect 87126 52534 87130 52590
rect 87130 52534 87186 52590
rect 87186 52534 87190 52590
rect 87126 52530 87190 52534
rect 886 52046 950 52050
rect 886 51990 890 52046
rect 890 51990 946 52046
rect 946 51990 950 52046
rect 886 51986 950 51990
rect 966 52046 1030 52050
rect 966 51990 970 52046
rect 970 51990 1026 52046
rect 1026 51990 1030 52046
rect 966 51986 1030 51990
rect 1046 52046 1110 52050
rect 1046 51990 1050 52046
rect 1050 51990 1106 52046
rect 1106 51990 1110 52046
rect 1046 51986 1110 51990
rect 1126 52046 1190 52050
rect 1126 51990 1130 52046
rect 1130 51990 1186 52046
rect 1186 51990 1190 52046
rect 1126 51986 1190 51990
rect 84886 52046 84950 52050
rect 84886 51990 84890 52046
rect 84890 51990 84946 52046
rect 84946 51990 84950 52046
rect 84886 51986 84950 51990
rect 84966 52046 85030 52050
rect 84966 51990 84970 52046
rect 84970 51990 85026 52046
rect 85026 51990 85030 52046
rect 84966 51986 85030 51990
rect 85046 52046 85110 52050
rect 85046 51990 85050 52046
rect 85050 51990 85106 52046
rect 85106 51990 85110 52046
rect 85046 51986 85110 51990
rect 85126 52046 85190 52050
rect 85126 51990 85130 52046
rect 85130 51990 85186 52046
rect 85186 51990 85190 52046
rect 85126 51986 85190 51990
rect 2886 51502 2950 51506
rect 2886 51446 2890 51502
rect 2890 51446 2946 51502
rect 2946 51446 2950 51502
rect 2886 51442 2950 51446
rect 2966 51502 3030 51506
rect 2966 51446 2970 51502
rect 2970 51446 3026 51502
rect 3026 51446 3030 51502
rect 2966 51442 3030 51446
rect 3046 51502 3110 51506
rect 3046 51446 3050 51502
rect 3050 51446 3106 51502
rect 3106 51446 3110 51502
rect 3046 51442 3110 51446
rect 3126 51502 3190 51506
rect 3126 51446 3130 51502
rect 3130 51446 3186 51502
rect 3186 51446 3190 51502
rect 3126 51442 3190 51446
rect 86886 51502 86950 51506
rect 86886 51446 86890 51502
rect 86890 51446 86946 51502
rect 86946 51446 86950 51502
rect 86886 51442 86950 51446
rect 86966 51502 87030 51506
rect 86966 51446 86970 51502
rect 86970 51446 87026 51502
rect 87026 51446 87030 51502
rect 86966 51442 87030 51446
rect 87046 51502 87110 51506
rect 87046 51446 87050 51502
rect 87050 51446 87106 51502
rect 87106 51446 87110 51502
rect 87046 51442 87110 51446
rect 87126 51502 87190 51506
rect 87126 51446 87130 51502
rect 87130 51446 87186 51502
rect 87186 51446 87190 51502
rect 87126 51442 87190 51446
rect 886 50958 950 50962
rect 886 50902 890 50958
rect 890 50902 946 50958
rect 946 50902 950 50958
rect 886 50898 950 50902
rect 966 50958 1030 50962
rect 966 50902 970 50958
rect 970 50902 1026 50958
rect 1026 50902 1030 50958
rect 966 50898 1030 50902
rect 1046 50958 1110 50962
rect 1046 50902 1050 50958
rect 1050 50902 1106 50958
rect 1106 50902 1110 50958
rect 1046 50898 1110 50902
rect 1126 50958 1190 50962
rect 1126 50902 1130 50958
rect 1130 50902 1186 50958
rect 1186 50902 1190 50958
rect 1126 50898 1190 50902
rect 84886 50958 84950 50962
rect 84886 50902 84890 50958
rect 84890 50902 84946 50958
rect 84946 50902 84950 50958
rect 84886 50898 84950 50902
rect 84966 50958 85030 50962
rect 84966 50902 84970 50958
rect 84970 50902 85026 50958
rect 85026 50902 85030 50958
rect 84966 50898 85030 50902
rect 85046 50958 85110 50962
rect 85046 50902 85050 50958
rect 85050 50902 85106 50958
rect 85106 50902 85110 50958
rect 85046 50898 85110 50902
rect 85126 50958 85190 50962
rect 85126 50902 85130 50958
rect 85130 50902 85186 50958
rect 85186 50902 85190 50958
rect 85126 50898 85190 50902
rect 2886 50414 2950 50418
rect 2886 50358 2890 50414
rect 2890 50358 2946 50414
rect 2946 50358 2950 50414
rect 2886 50354 2950 50358
rect 2966 50414 3030 50418
rect 2966 50358 2970 50414
rect 2970 50358 3026 50414
rect 3026 50358 3030 50414
rect 2966 50354 3030 50358
rect 3046 50414 3110 50418
rect 3046 50358 3050 50414
rect 3050 50358 3106 50414
rect 3106 50358 3110 50414
rect 3046 50354 3110 50358
rect 3126 50414 3190 50418
rect 3126 50358 3130 50414
rect 3130 50358 3186 50414
rect 3186 50358 3190 50414
rect 3126 50354 3190 50358
rect 86886 50414 86950 50418
rect 86886 50358 86890 50414
rect 86890 50358 86946 50414
rect 86946 50358 86950 50414
rect 86886 50354 86950 50358
rect 86966 50414 87030 50418
rect 86966 50358 86970 50414
rect 86970 50358 87026 50414
rect 87026 50358 87030 50414
rect 86966 50354 87030 50358
rect 87046 50414 87110 50418
rect 87046 50358 87050 50414
rect 87050 50358 87106 50414
rect 87106 50358 87110 50414
rect 87046 50354 87110 50358
rect 87126 50414 87190 50418
rect 87126 50358 87130 50414
rect 87130 50358 87186 50414
rect 87186 50358 87190 50414
rect 87126 50354 87190 50358
rect 886 49870 950 49874
rect 886 49814 890 49870
rect 890 49814 946 49870
rect 946 49814 950 49870
rect 886 49810 950 49814
rect 966 49870 1030 49874
rect 966 49814 970 49870
rect 970 49814 1026 49870
rect 1026 49814 1030 49870
rect 966 49810 1030 49814
rect 1046 49870 1110 49874
rect 1046 49814 1050 49870
rect 1050 49814 1106 49870
rect 1106 49814 1110 49870
rect 1046 49810 1110 49814
rect 1126 49870 1190 49874
rect 1126 49814 1130 49870
rect 1130 49814 1186 49870
rect 1186 49814 1190 49870
rect 1126 49810 1190 49814
rect 84886 49870 84950 49874
rect 84886 49814 84890 49870
rect 84890 49814 84946 49870
rect 84946 49814 84950 49870
rect 84886 49810 84950 49814
rect 84966 49870 85030 49874
rect 84966 49814 84970 49870
rect 84970 49814 85026 49870
rect 85026 49814 85030 49870
rect 84966 49810 85030 49814
rect 85046 49870 85110 49874
rect 85046 49814 85050 49870
rect 85050 49814 85106 49870
rect 85106 49814 85110 49870
rect 85046 49810 85110 49814
rect 85126 49870 85190 49874
rect 85126 49814 85130 49870
rect 85130 49814 85186 49870
rect 85186 49814 85190 49870
rect 85126 49810 85190 49814
rect 2886 49326 2950 49330
rect 2886 49270 2890 49326
rect 2890 49270 2946 49326
rect 2946 49270 2950 49326
rect 2886 49266 2950 49270
rect 2966 49326 3030 49330
rect 2966 49270 2970 49326
rect 2970 49270 3026 49326
rect 3026 49270 3030 49326
rect 2966 49266 3030 49270
rect 3046 49326 3110 49330
rect 3046 49270 3050 49326
rect 3050 49270 3106 49326
rect 3106 49270 3110 49326
rect 3046 49266 3110 49270
rect 3126 49326 3190 49330
rect 3126 49270 3130 49326
rect 3130 49270 3186 49326
rect 3186 49270 3190 49326
rect 3126 49266 3190 49270
rect 86886 49326 86950 49330
rect 86886 49270 86890 49326
rect 86890 49270 86946 49326
rect 86946 49270 86950 49326
rect 86886 49266 86950 49270
rect 86966 49326 87030 49330
rect 86966 49270 86970 49326
rect 86970 49270 87026 49326
rect 87026 49270 87030 49326
rect 86966 49266 87030 49270
rect 87046 49326 87110 49330
rect 87046 49270 87050 49326
rect 87050 49270 87106 49326
rect 87106 49270 87110 49326
rect 87046 49266 87110 49270
rect 87126 49326 87190 49330
rect 87126 49270 87130 49326
rect 87130 49270 87186 49326
rect 87186 49270 87190 49326
rect 87126 49266 87190 49270
rect 886 48782 950 48786
rect 886 48726 890 48782
rect 890 48726 946 48782
rect 946 48726 950 48782
rect 886 48722 950 48726
rect 966 48782 1030 48786
rect 966 48726 970 48782
rect 970 48726 1026 48782
rect 1026 48726 1030 48782
rect 966 48722 1030 48726
rect 1046 48782 1110 48786
rect 1046 48726 1050 48782
rect 1050 48726 1106 48782
rect 1106 48726 1110 48782
rect 1046 48722 1110 48726
rect 1126 48782 1190 48786
rect 1126 48726 1130 48782
rect 1130 48726 1186 48782
rect 1186 48726 1190 48782
rect 1126 48722 1190 48726
rect 84886 48782 84950 48786
rect 84886 48726 84890 48782
rect 84890 48726 84946 48782
rect 84946 48726 84950 48782
rect 84886 48722 84950 48726
rect 84966 48782 85030 48786
rect 84966 48726 84970 48782
rect 84970 48726 85026 48782
rect 85026 48726 85030 48782
rect 84966 48722 85030 48726
rect 85046 48782 85110 48786
rect 85046 48726 85050 48782
rect 85050 48726 85106 48782
rect 85106 48726 85110 48782
rect 85046 48722 85110 48726
rect 85126 48782 85190 48786
rect 85126 48726 85130 48782
rect 85130 48726 85186 48782
rect 85186 48726 85190 48782
rect 85126 48722 85190 48726
rect 2886 48238 2950 48242
rect 2886 48182 2890 48238
rect 2890 48182 2946 48238
rect 2946 48182 2950 48238
rect 2886 48178 2950 48182
rect 2966 48238 3030 48242
rect 2966 48182 2970 48238
rect 2970 48182 3026 48238
rect 3026 48182 3030 48238
rect 2966 48178 3030 48182
rect 3046 48238 3110 48242
rect 3046 48182 3050 48238
rect 3050 48182 3106 48238
rect 3106 48182 3110 48238
rect 3046 48178 3110 48182
rect 3126 48238 3190 48242
rect 3126 48182 3130 48238
rect 3130 48182 3186 48238
rect 3186 48182 3190 48238
rect 3126 48178 3190 48182
rect 86886 48238 86950 48242
rect 86886 48182 86890 48238
rect 86890 48182 86946 48238
rect 86946 48182 86950 48238
rect 86886 48178 86950 48182
rect 86966 48238 87030 48242
rect 86966 48182 86970 48238
rect 86970 48182 87026 48238
rect 87026 48182 87030 48238
rect 86966 48178 87030 48182
rect 87046 48238 87110 48242
rect 87046 48182 87050 48238
rect 87050 48182 87106 48238
rect 87106 48182 87110 48238
rect 87046 48178 87110 48182
rect 87126 48238 87190 48242
rect 87126 48182 87130 48238
rect 87130 48182 87186 48238
rect 87186 48182 87190 48238
rect 87126 48178 87190 48182
rect 886 47694 950 47698
rect 886 47638 890 47694
rect 890 47638 946 47694
rect 946 47638 950 47694
rect 886 47634 950 47638
rect 966 47694 1030 47698
rect 966 47638 970 47694
rect 970 47638 1026 47694
rect 1026 47638 1030 47694
rect 966 47634 1030 47638
rect 1046 47694 1110 47698
rect 1046 47638 1050 47694
rect 1050 47638 1106 47694
rect 1106 47638 1110 47694
rect 1046 47634 1110 47638
rect 1126 47694 1190 47698
rect 1126 47638 1130 47694
rect 1130 47638 1186 47694
rect 1186 47638 1190 47694
rect 1126 47634 1190 47638
rect 84886 47694 84950 47698
rect 84886 47638 84890 47694
rect 84890 47638 84946 47694
rect 84946 47638 84950 47694
rect 84886 47634 84950 47638
rect 84966 47694 85030 47698
rect 84966 47638 84970 47694
rect 84970 47638 85026 47694
rect 85026 47638 85030 47694
rect 84966 47634 85030 47638
rect 85046 47694 85110 47698
rect 85046 47638 85050 47694
rect 85050 47638 85106 47694
rect 85106 47638 85110 47694
rect 85046 47634 85110 47638
rect 85126 47694 85190 47698
rect 85126 47638 85130 47694
rect 85130 47638 85186 47694
rect 85186 47638 85190 47694
rect 85126 47634 85190 47638
rect 2886 47150 2950 47154
rect 2886 47094 2890 47150
rect 2890 47094 2946 47150
rect 2946 47094 2950 47150
rect 2886 47090 2950 47094
rect 2966 47150 3030 47154
rect 2966 47094 2970 47150
rect 2970 47094 3026 47150
rect 3026 47094 3030 47150
rect 2966 47090 3030 47094
rect 3046 47150 3110 47154
rect 3046 47094 3050 47150
rect 3050 47094 3106 47150
rect 3106 47094 3110 47150
rect 3046 47090 3110 47094
rect 3126 47150 3190 47154
rect 3126 47094 3130 47150
rect 3130 47094 3186 47150
rect 3186 47094 3190 47150
rect 3126 47090 3190 47094
rect 86886 47150 86950 47154
rect 86886 47094 86890 47150
rect 86890 47094 86946 47150
rect 86946 47094 86950 47150
rect 86886 47090 86950 47094
rect 86966 47150 87030 47154
rect 86966 47094 86970 47150
rect 86970 47094 87026 47150
rect 87026 47094 87030 47150
rect 86966 47090 87030 47094
rect 87046 47150 87110 47154
rect 87046 47094 87050 47150
rect 87050 47094 87106 47150
rect 87106 47094 87110 47150
rect 87046 47090 87110 47094
rect 87126 47150 87190 47154
rect 87126 47094 87130 47150
rect 87130 47094 87186 47150
rect 87186 47094 87190 47150
rect 87126 47090 87190 47094
rect 886 46606 950 46610
rect 886 46550 890 46606
rect 890 46550 946 46606
rect 946 46550 950 46606
rect 886 46546 950 46550
rect 966 46606 1030 46610
rect 966 46550 970 46606
rect 970 46550 1026 46606
rect 1026 46550 1030 46606
rect 966 46546 1030 46550
rect 1046 46606 1110 46610
rect 1046 46550 1050 46606
rect 1050 46550 1106 46606
rect 1106 46550 1110 46606
rect 1046 46546 1110 46550
rect 1126 46606 1190 46610
rect 1126 46550 1130 46606
rect 1130 46550 1186 46606
rect 1186 46550 1190 46606
rect 1126 46546 1190 46550
rect 84886 46606 84950 46610
rect 84886 46550 84890 46606
rect 84890 46550 84946 46606
rect 84946 46550 84950 46606
rect 84886 46546 84950 46550
rect 84966 46606 85030 46610
rect 84966 46550 84970 46606
rect 84970 46550 85026 46606
rect 85026 46550 85030 46606
rect 84966 46546 85030 46550
rect 85046 46606 85110 46610
rect 85046 46550 85050 46606
rect 85050 46550 85106 46606
rect 85106 46550 85110 46606
rect 85046 46546 85110 46550
rect 85126 46606 85190 46610
rect 85126 46550 85130 46606
rect 85130 46550 85186 46606
rect 85186 46550 85190 46606
rect 85126 46546 85190 46550
rect 2886 46062 2950 46066
rect 2886 46006 2890 46062
rect 2890 46006 2946 46062
rect 2946 46006 2950 46062
rect 2886 46002 2950 46006
rect 2966 46062 3030 46066
rect 2966 46006 2970 46062
rect 2970 46006 3026 46062
rect 3026 46006 3030 46062
rect 2966 46002 3030 46006
rect 3046 46062 3110 46066
rect 3046 46006 3050 46062
rect 3050 46006 3106 46062
rect 3106 46006 3110 46062
rect 3046 46002 3110 46006
rect 3126 46062 3190 46066
rect 3126 46006 3130 46062
rect 3130 46006 3186 46062
rect 3186 46006 3190 46062
rect 3126 46002 3190 46006
rect 86886 46062 86950 46066
rect 86886 46006 86890 46062
rect 86890 46006 86946 46062
rect 86946 46006 86950 46062
rect 86886 46002 86950 46006
rect 86966 46062 87030 46066
rect 86966 46006 86970 46062
rect 86970 46006 87026 46062
rect 87026 46006 87030 46062
rect 86966 46002 87030 46006
rect 87046 46062 87110 46066
rect 87046 46006 87050 46062
rect 87050 46006 87106 46062
rect 87106 46006 87110 46062
rect 87046 46002 87110 46006
rect 87126 46062 87190 46066
rect 87126 46006 87130 46062
rect 87130 46006 87186 46062
rect 87186 46006 87190 46062
rect 87126 46002 87190 46006
rect 886 45518 950 45522
rect 886 45462 890 45518
rect 890 45462 946 45518
rect 946 45462 950 45518
rect 886 45458 950 45462
rect 966 45518 1030 45522
rect 966 45462 970 45518
rect 970 45462 1026 45518
rect 1026 45462 1030 45518
rect 966 45458 1030 45462
rect 1046 45518 1110 45522
rect 1046 45462 1050 45518
rect 1050 45462 1106 45518
rect 1106 45462 1110 45518
rect 1046 45458 1110 45462
rect 1126 45518 1190 45522
rect 1126 45462 1130 45518
rect 1130 45462 1186 45518
rect 1186 45462 1190 45518
rect 1126 45458 1190 45462
rect 84886 45518 84950 45522
rect 84886 45462 84890 45518
rect 84890 45462 84946 45518
rect 84946 45462 84950 45518
rect 84886 45458 84950 45462
rect 84966 45518 85030 45522
rect 84966 45462 84970 45518
rect 84970 45462 85026 45518
rect 85026 45462 85030 45518
rect 84966 45458 85030 45462
rect 85046 45518 85110 45522
rect 85046 45462 85050 45518
rect 85050 45462 85106 45518
rect 85106 45462 85110 45518
rect 85046 45458 85110 45462
rect 85126 45518 85190 45522
rect 85126 45462 85130 45518
rect 85130 45462 85186 45518
rect 85186 45462 85190 45518
rect 85126 45458 85190 45462
rect 2886 44974 2950 44978
rect 2886 44918 2890 44974
rect 2890 44918 2946 44974
rect 2946 44918 2950 44974
rect 2886 44914 2950 44918
rect 2966 44974 3030 44978
rect 2966 44918 2970 44974
rect 2970 44918 3026 44974
rect 3026 44918 3030 44974
rect 2966 44914 3030 44918
rect 3046 44974 3110 44978
rect 3046 44918 3050 44974
rect 3050 44918 3106 44974
rect 3106 44918 3110 44974
rect 3046 44914 3110 44918
rect 3126 44974 3190 44978
rect 3126 44918 3130 44974
rect 3130 44918 3186 44974
rect 3186 44918 3190 44974
rect 3126 44914 3190 44918
rect 86886 44974 86950 44978
rect 86886 44918 86890 44974
rect 86890 44918 86946 44974
rect 86946 44918 86950 44974
rect 86886 44914 86950 44918
rect 86966 44974 87030 44978
rect 86966 44918 86970 44974
rect 86970 44918 87026 44974
rect 87026 44918 87030 44974
rect 86966 44914 87030 44918
rect 87046 44974 87110 44978
rect 87046 44918 87050 44974
rect 87050 44918 87106 44974
rect 87106 44918 87110 44974
rect 87046 44914 87110 44918
rect 87126 44974 87190 44978
rect 87126 44918 87130 44974
rect 87130 44918 87186 44974
rect 87186 44918 87190 44974
rect 87126 44914 87190 44918
rect 886 44430 950 44434
rect 886 44374 890 44430
rect 890 44374 946 44430
rect 946 44374 950 44430
rect 886 44370 950 44374
rect 966 44430 1030 44434
rect 966 44374 970 44430
rect 970 44374 1026 44430
rect 1026 44374 1030 44430
rect 966 44370 1030 44374
rect 1046 44430 1110 44434
rect 1046 44374 1050 44430
rect 1050 44374 1106 44430
rect 1106 44374 1110 44430
rect 1046 44370 1110 44374
rect 1126 44430 1190 44434
rect 1126 44374 1130 44430
rect 1130 44374 1186 44430
rect 1186 44374 1190 44430
rect 1126 44370 1190 44374
rect 84886 44430 84950 44434
rect 84886 44374 84890 44430
rect 84890 44374 84946 44430
rect 84946 44374 84950 44430
rect 84886 44370 84950 44374
rect 84966 44430 85030 44434
rect 84966 44374 84970 44430
rect 84970 44374 85026 44430
rect 85026 44374 85030 44430
rect 84966 44370 85030 44374
rect 85046 44430 85110 44434
rect 85046 44374 85050 44430
rect 85050 44374 85106 44430
rect 85106 44374 85110 44430
rect 85046 44370 85110 44374
rect 85126 44430 85190 44434
rect 85126 44374 85130 44430
rect 85130 44374 85186 44430
rect 85186 44374 85190 44430
rect 85126 44370 85190 44374
rect 2886 43886 2950 43890
rect 2886 43830 2890 43886
rect 2890 43830 2946 43886
rect 2946 43830 2950 43886
rect 2886 43826 2950 43830
rect 2966 43886 3030 43890
rect 2966 43830 2970 43886
rect 2970 43830 3026 43886
rect 3026 43830 3030 43886
rect 2966 43826 3030 43830
rect 3046 43886 3110 43890
rect 3046 43830 3050 43886
rect 3050 43830 3106 43886
rect 3106 43830 3110 43886
rect 3046 43826 3110 43830
rect 3126 43886 3190 43890
rect 3126 43830 3130 43886
rect 3130 43830 3186 43886
rect 3186 43830 3190 43886
rect 3126 43826 3190 43830
rect 86886 43886 86950 43890
rect 86886 43830 86890 43886
rect 86890 43830 86946 43886
rect 86946 43830 86950 43886
rect 86886 43826 86950 43830
rect 86966 43886 87030 43890
rect 86966 43830 86970 43886
rect 86970 43830 87026 43886
rect 87026 43830 87030 43886
rect 86966 43826 87030 43830
rect 87046 43886 87110 43890
rect 87046 43830 87050 43886
rect 87050 43830 87106 43886
rect 87106 43830 87110 43886
rect 87046 43826 87110 43830
rect 87126 43886 87190 43890
rect 87126 43830 87130 43886
rect 87130 43830 87186 43886
rect 87186 43830 87190 43886
rect 87126 43826 87190 43830
rect 886 43342 950 43346
rect 886 43286 890 43342
rect 890 43286 946 43342
rect 946 43286 950 43342
rect 886 43282 950 43286
rect 966 43342 1030 43346
rect 966 43286 970 43342
rect 970 43286 1026 43342
rect 1026 43286 1030 43342
rect 966 43282 1030 43286
rect 1046 43342 1110 43346
rect 1046 43286 1050 43342
rect 1050 43286 1106 43342
rect 1106 43286 1110 43342
rect 1046 43282 1110 43286
rect 1126 43342 1190 43346
rect 1126 43286 1130 43342
rect 1130 43286 1186 43342
rect 1186 43286 1190 43342
rect 1126 43282 1190 43286
rect 84886 43342 84950 43346
rect 84886 43286 84890 43342
rect 84890 43286 84946 43342
rect 84946 43286 84950 43342
rect 84886 43282 84950 43286
rect 84966 43342 85030 43346
rect 84966 43286 84970 43342
rect 84970 43286 85026 43342
rect 85026 43286 85030 43342
rect 84966 43282 85030 43286
rect 85046 43342 85110 43346
rect 85046 43286 85050 43342
rect 85050 43286 85106 43342
rect 85106 43286 85110 43342
rect 85046 43282 85110 43286
rect 85126 43342 85190 43346
rect 85126 43286 85130 43342
rect 85130 43286 85186 43342
rect 85186 43286 85190 43342
rect 85126 43282 85190 43286
rect 2886 42798 2950 42802
rect 2886 42742 2890 42798
rect 2890 42742 2946 42798
rect 2946 42742 2950 42798
rect 2886 42738 2950 42742
rect 2966 42798 3030 42802
rect 2966 42742 2970 42798
rect 2970 42742 3026 42798
rect 3026 42742 3030 42798
rect 2966 42738 3030 42742
rect 3046 42798 3110 42802
rect 3046 42742 3050 42798
rect 3050 42742 3106 42798
rect 3106 42742 3110 42798
rect 3046 42738 3110 42742
rect 3126 42798 3190 42802
rect 3126 42742 3130 42798
rect 3130 42742 3186 42798
rect 3186 42742 3190 42798
rect 3126 42738 3190 42742
rect 86886 42798 86950 42802
rect 86886 42742 86890 42798
rect 86890 42742 86946 42798
rect 86946 42742 86950 42798
rect 86886 42738 86950 42742
rect 86966 42798 87030 42802
rect 86966 42742 86970 42798
rect 86970 42742 87026 42798
rect 87026 42742 87030 42798
rect 86966 42738 87030 42742
rect 87046 42798 87110 42802
rect 87046 42742 87050 42798
rect 87050 42742 87106 42798
rect 87106 42742 87110 42798
rect 87046 42738 87110 42742
rect 87126 42798 87190 42802
rect 87126 42742 87130 42798
rect 87130 42742 87186 42798
rect 87186 42742 87190 42798
rect 87126 42738 87190 42742
rect 886 42254 950 42258
rect 886 42198 890 42254
rect 890 42198 946 42254
rect 946 42198 950 42254
rect 886 42194 950 42198
rect 966 42254 1030 42258
rect 966 42198 970 42254
rect 970 42198 1026 42254
rect 1026 42198 1030 42254
rect 966 42194 1030 42198
rect 1046 42254 1110 42258
rect 1046 42198 1050 42254
rect 1050 42198 1106 42254
rect 1106 42198 1110 42254
rect 1046 42194 1110 42198
rect 1126 42254 1190 42258
rect 1126 42198 1130 42254
rect 1130 42198 1186 42254
rect 1186 42198 1190 42254
rect 1126 42194 1190 42198
rect 84886 42254 84950 42258
rect 84886 42198 84890 42254
rect 84890 42198 84946 42254
rect 84946 42198 84950 42254
rect 84886 42194 84950 42198
rect 84966 42254 85030 42258
rect 84966 42198 84970 42254
rect 84970 42198 85026 42254
rect 85026 42198 85030 42254
rect 84966 42194 85030 42198
rect 85046 42254 85110 42258
rect 85046 42198 85050 42254
rect 85050 42198 85106 42254
rect 85106 42198 85110 42254
rect 85046 42194 85110 42198
rect 85126 42254 85190 42258
rect 85126 42198 85130 42254
rect 85130 42198 85186 42254
rect 85186 42198 85190 42254
rect 85126 42194 85190 42198
rect 2886 41710 2950 41714
rect 2886 41654 2890 41710
rect 2890 41654 2946 41710
rect 2946 41654 2950 41710
rect 2886 41650 2950 41654
rect 2966 41710 3030 41714
rect 2966 41654 2970 41710
rect 2970 41654 3026 41710
rect 3026 41654 3030 41710
rect 2966 41650 3030 41654
rect 3046 41710 3110 41714
rect 3046 41654 3050 41710
rect 3050 41654 3106 41710
rect 3106 41654 3110 41710
rect 3046 41650 3110 41654
rect 3126 41710 3190 41714
rect 3126 41654 3130 41710
rect 3130 41654 3186 41710
rect 3186 41654 3190 41710
rect 3126 41650 3190 41654
rect 86886 41710 86950 41714
rect 86886 41654 86890 41710
rect 86890 41654 86946 41710
rect 86946 41654 86950 41710
rect 86886 41650 86950 41654
rect 86966 41710 87030 41714
rect 86966 41654 86970 41710
rect 86970 41654 87026 41710
rect 87026 41654 87030 41710
rect 86966 41650 87030 41654
rect 87046 41710 87110 41714
rect 87046 41654 87050 41710
rect 87050 41654 87106 41710
rect 87106 41654 87110 41710
rect 87046 41650 87110 41654
rect 87126 41710 87190 41714
rect 87126 41654 87130 41710
rect 87130 41654 87186 41710
rect 87186 41654 87190 41710
rect 87126 41650 87190 41654
rect 886 41166 950 41170
rect 886 41110 890 41166
rect 890 41110 946 41166
rect 946 41110 950 41166
rect 886 41106 950 41110
rect 966 41166 1030 41170
rect 966 41110 970 41166
rect 970 41110 1026 41166
rect 1026 41110 1030 41166
rect 966 41106 1030 41110
rect 1046 41166 1110 41170
rect 1046 41110 1050 41166
rect 1050 41110 1106 41166
rect 1106 41110 1110 41166
rect 1046 41106 1110 41110
rect 1126 41166 1190 41170
rect 1126 41110 1130 41166
rect 1130 41110 1186 41166
rect 1186 41110 1190 41166
rect 1126 41106 1190 41110
rect 84886 41166 84950 41170
rect 84886 41110 84890 41166
rect 84890 41110 84946 41166
rect 84946 41110 84950 41166
rect 84886 41106 84950 41110
rect 84966 41166 85030 41170
rect 84966 41110 84970 41166
rect 84970 41110 85026 41166
rect 85026 41110 85030 41166
rect 84966 41106 85030 41110
rect 85046 41166 85110 41170
rect 85046 41110 85050 41166
rect 85050 41110 85106 41166
rect 85106 41110 85110 41166
rect 85046 41106 85110 41110
rect 85126 41166 85190 41170
rect 85126 41110 85130 41166
rect 85130 41110 85186 41166
rect 85186 41110 85190 41166
rect 85126 41106 85190 41110
rect 2886 40622 2950 40626
rect 2886 40566 2890 40622
rect 2890 40566 2946 40622
rect 2946 40566 2950 40622
rect 2886 40562 2950 40566
rect 2966 40622 3030 40626
rect 2966 40566 2970 40622
rect 2970 40566 3026 40622
rect 3026 40566 3030 40622
rect 2966 40562 3030 40566
rect 3046 40622 3110 40626
rect 3046 40566 3050 40622
rect 3050 40566 3106 40622
rect 3106 40566 3110 40622
rect 3046 40562 3110 40566
rect 3126 40622 3190 40626
rect 3126 40566 3130 40622
rect 3130 40566 3186 40622
rect 3186 40566 3190 40622
rect 3126 40562 3190 40566
rect 86886 40622 86950 40626
rect 86886 40566 86890 40622
rect 86890 40566 86946 40622
rect 86946 40566 86950 40622
rect 86886 40562 86950 40566
rect 86966 40622 87030 40626
rect 86966 40566 86970 40622
rect 86970 40566 87026 40622
rect 87026 40566 87030 40622
rect 86966 40562 87030 40566
rect 87046 40622 87110 40626
rect 87046 40566 87050 40622
rect 87050 40566 87106 40622
rect 87106 40566 87110 40622
rect 87046 40562 87110 40566
rect 87126 40622 87190 40626
rect 87126 40566 87130 40622
rect 87130 40566 87186 40622
rect 87186 40566 87190 40622
rect 87126 40562 87190 40566
rect 886 40078 950 40082
rect 886 40022 890 40078
rect 890 40022 946 40078
rect 946 40022 950 40078
rect 886 40018 950 40022
rect 966 40078 1030 40082
rect 966 40022 970 40078
rect 970 40022 1026 40078
rect 1026 40022 1030 40078
rect 966 40018 1030 40022
rect 1046 40078 1110 40082
rect 1046 40022 1050 40078
rect 1050 40022 1106 40078
rect 1106 40022 1110 40078
rect 1046 40018 1110 40022
rect 1126 40078 1190 40082
rect 1126 40022 1130 40078
rect 1130 40022 1186 40078
rect 1186 40022 1190 40078
rect 1126 40018 1190 40022
rect 84886 40078 84950 40082
rect 84886 40022 84890 40078
rect 84890 40022 84946 40078
rect 84946 40022 84950 40078
rect 84886 40018 84950 40022
rect 84966 40078 85030 40082
rect 84966 40022 84970 40078
rect 84970 40022 85026 40078
rect 85026 40022 85030 40078
rect 84966 40018 85030 40022
rect 85046 40078 85110 40082
rect 85046 40022 85050 40078
rect 85050 40022 85106 40078
rect 85106 40022 85110 40078
rect 85046 40018 85110 40022
rect 85126 40078 85190 40082
rect 85126 40022 85130 40078
rect 85130 40022 85186 40078
rect 85186 40022 85190 40078
rect 85126 40018 85190 40022
rect 2886 39534 2950 39538
rect 2886 39478 2890 39534
rect 2890 39478 2946 39534
rect 2946 39478 2950 39534
rect 2886 39474 2950 39478
rect 2966 39534 3030 39538
rect 2966 39478 2970 39534
rect 2970 39478 3026 39534
rect 3026 39478 3030 39534
rect 2966 39474 3030 39478
rect 3046 39534 3110 39538
rect 3046 39478 3050 39534
rect 3050 39478 3106 39534
rect 3106 39478 3110 39534
rect 3046 39474 3110 39478
rect 3126 39534 3190 39538
rect 3126 39478 3130 39534
rect 3130 39478 3186 39534
rect 3186 39478 3190 39534
rect 3126 39474 3190 39478
rect 86886 39534 86950 39538
rect 86886 39478 86890 39534
rect 86890 39478 86946 39534
rect 86946 39478 86950 39534
rect 86886 39474 86950 39478
rect 86966 39534 87030 39538
rect 86966 39478 86970 39534
rect 86970 39478 87026 39534
rect 87026 39478 87030 39534
rect 86966 39474 87030 39478
rect 87046 39534 87110 39538
rect 87046 39478 87050 39534
rect 87050 39478 87106 39534
rect 87106 39478 87110 39534
rect 87046 39474 87110 39478
rect 87126 39534 87190 39538
rect 87126 39478 87130 39534
rect 87130 39478 87186 39534
rect 87186 39478 87190 39534
rect 87126 39474 87190 39478
rect 886 38990 950 38994
rect 886 38934 890 38990
rect 890 38934 946 38990
rect 946 38934 950 38990
rect 886 38930 950 38934
rect 966 38990 1030 38994
rect 966 38934 970 38990
rect 970 38934 1026 38990
rect 1026 38934 1030 38990
rect 966 38930 1030 38934
rect 1046 38990 1110 38994
rect 1046 38934 1050 38990
rect 1050 38934 1106 38990
rect 1106 38934 1110 38990
rect 1046 38930 1110 38934
rect 1126 38990 1190 38994
rect 1126 38934 1130 38990
rect 1130 38934 1186 38990
rect 1186 38934 1190 38990
rect 1126 38930 1190 38934
rect 84886 38990 84950 38994
rect 84886 38934 84890 38990
rect 84890 38934 84946 38990
rect 84946 38934 84950 38990
rect 84886 38930 84950 38934
rect 84966 38990 85030 38994
rect 84966 38934 84970 38990
rect 84970 38934 85026 38990
rect 85026 38934 85030 38990
rect 84966 38930 85030 38934
rect 85046 38990 85110 38994
rect 85046 38934 85050 38990
rect 85050 38934 85106 38990
rect 85106 38934 85110 38990
rect 85046 38930 85110 38934
rect 85126 38990 85190 38994
rect 85126 38934 85130 38990
rect 85130 38934 85186 38990
rect 85186 38934 85190 38990
rect 85126 38930 85190 38934
rect 2886 38446 2950 38450
rect 2886 38390 2890 38446
rect 2890 38390 2946 38446
rect 2946 38390 2950 38446
rect 2886 38386 2950 38390
rect 2966 38446 3030 38450
rect 2966 38390 2970 38446
rect 2970 38390 3026 38446
rect 3026 38390 3030 38446
rect 2966 38386 3030 38390
rect 3046 38446 3110 38450
rect 3046 38390 3050 38446
rect 3050 38390 3106 38446
rect 3106 38390 3110 38446
rect 3046 38386 3110 38390
rect 3126 38446 3190 38450
rect 3126 38390 3130 38446
rect 3130 38390 3186 38446
rect 3186 38390 3190 38446
rect 3126 38386 3190 38390
rect 86886 38446 86950 38450
rect 86886 38390 86890 38446
rect 86890 38390 86946 38446
rect 86946 38390 86950 38446
rect 86886 38386 86950 38390
rect 86966 38446 87030 38450
rect 86966 38390 86970 38446
rect 86970 38390 87026 38446
rect 87026 38390 87030 38446
rect 86966 38386 87030 38390
rect 87046 38446 87110 38450
rect 87046 38390 87050 38446
rect 87050 38390 87106 38446
rect 87106 38390 87110 38446
rect 87046 38386 87110 38390
rect 87126 38446 87190 38450
rect 87126 38390 87130 38446
rect 87130 38390 87186 38446
rect 87186 38390 87190 38446
rect 87126 38386 87190 38390
rect 886 37902 950 37906
rect 886 37846 890 37902
rect 890 37846 946 37902
rect 946 37846 950 37902
rect 886 37842 950 37846
rect 966 37902 1030 37906
rect 966 37846 970 37902
rect 970 37846 1026 37902
rect 1026 37846 1030 37902
rect 966 37842 1030 37846
rect 1046 37902 1110 37906
rect 1046 37846 1050 37902
rect 1050 37846 1106 37902
rect 1106 37846 1110 37902
rect 1046 37842 1110 37846
rect 1126 37902 1190 37906
rect 1126 37846 1130 37902
rect 1130 37846 1186 37902
rect 1186 37846 1190 37902
rect 1126 37842 1190 37846
rect 84886 37902 84950 37906
rect 84886 37846 84890 37902
rect 84890 37846 84946 37902
rect 84946 37846 84950 37902
rect 84886 37842 84950 37846
rect 84966 37902 85030 37906
rect 84966 37846 84970 37902
rect 84970 37846 85026 37902
rect 85026 37846 85030 37902
rect 84966 37842 85030 37846
rect 85046 37902 85110 37906
rect 85046 37846 85050 37902
rect 85050 37846 85106 37902
rect 85106 37846 85110 37902
rect 85046 37842 85110 37846
rect 85126 37902 85190 37906
rect 85126 37846 85130 37902
rect 85130 37846 85186 37902
rect 85186 37846 85190 37902
rect 85126 37842 85190 37846
rect 2886 37358 2950 37362
rect 2886 37302 2890 37358
rect 2890 37302 2946 37358
rect 2946 37302 2950 37358
rect 2886 37298 2950 37302
rect 2966 37358 3030 37362
rect 2966 37302 2970 37358
rect 2970 37302 3026 37358
rect 3026 37302 3030 37358
rect 2966 37298 3030 37302
rect 3046 37358 3110 37362
rect 3046 37302 3050 37358
rect 3050 37302 3106 37358
rect 3106 37302 3110 37358
rect 3046 37298 3110 37302
rect 3126 37358 3190 37362
rect 3126 37302 3130 37358
rect 3130 37302 3186 37358
rect 3186 37302 3190 37358
rect 3126 37298 3190 37302
rect 86886 37358 86950 37362
rect 86886 37302 86890 37358
rect 86890 37302 86946 37358
rect 86946 37302 86950 37358
rect 86886 37298 86950 37302
rect 86966 37358 87030 37362
rect 86966 37302 86970 37358
rect 86970 37302 87026 37358
rect 87026 37302 87030 37358
rect 86966 37298 87030 37302
rect 87046 37358 87110 37362
rect 87046 37302 87050 37358
rect 87050 37302 87106 37358
rect 87106 37302 87110 37358
rect 87046 37298 87110 37302
rect 87126 37358 87190 37362
rect 87126 37302 87130 37358
rect 87130 37302 87186 37358
rect 87186 37302 87190 37358
rect 87126 37298 87190 37302
rect 886 36814 950 36818
rect 886 36758 890 36814
rect 890 36758 946 36814
rect 946 36758 950 36814
rect 886 36754 950 36758
rect 966 36814 1030 36818
rect 966 36758 970 36814
rect 970 36758 1026 36814
rect 1026 36758 1030 36814
rect 966 36754 1030 36758
rect 1046 36814 1110 36818
rect 1046 36758 1050 36814
rect 1050 36758 1106 36814
rect 1106 36758 1110 36814
rect 1046 36754 1110 36758
rect 1126 36814 1190 36818
rect 1126 36758 1130 36814
rect 1130 36758 1186 36814
rect 1186 36758 1190 36814
rect 1126 36754 1190 36758
rect 84886 36814 84950 36818
rect 84886 36758 84890 36814
rect 84890 36758 84946 36814
rect 84946 36758 84950 36814
rect 84886 36754 84950 36758
rect 84966 36814 85030 36818
rect 84966 36758 84970 36814
rect 84970 36758 85026 36814
rect 85026 36758 85030 36814
rect 84966 36754 85030 36758
rect 85046 36814 85110 36818
rect 85046 36758 85050 36814
rect 85050 36758 85106 36814
rect 85106 36758 85110 36814
rect 85046 36754 85110 36758
rect 85126 36814 85190 36818
rect 85126 36758 85130 36814
rect 85130 36758 85186 36814
rect 85186 36758 85190 36814
rect 85126 36754 85190 36758
rect 2886 36270 2950 36274
rect 2886 36214 2890 36270
rect 2890 36214 2946 36270
rect 2946 36214 2950 36270
rect 2886 36210 2950 36214
rect 2966 36270 3030 36274
rect 2966 36214 2970 36270
rect 2970 36214 3026 36270
rect 3026 36214 3030 36270
rect 2966 36210 3030 36214
rect 3046 36270 3110 36274
rect 3046 36214 3050 36270
rect 3050 36214 3106 36270
rect 3106 36214 3110 36270
rect 3046 36210 3110 36214
rect 3126 36270 3190 36274
rect 3126 36214 3130 36270
rect 3130 36214 3186 36270
rect 3186 36214 3190 36270
rect 3126 36210 3190 36214
rect 86886 36270 86950 36274
rect 86886 36214 86890 36270
rect 86890 36214 86946 36270
rect 86946 36214 86950 36270
rect 86886 36210 86950 36214
rect 86966 36270 87030 36274
rect 86966 36214 86970 36270
rect 86970 36214 87026 36270
rect 87026 36214 87030 36270
rect 86966 36210 87030 36214
rect 87046 36270 87110 36274
rect 87046 36214 87050 36270
rect 87050 36214 87106 36270
rect 87106 36214 87110 36270
rect 87046 36210 87110 36214
rect 87126 36270 87190 36274
rect 87126 36214 87130 36270
rect 87130 36214 87186 36270
rect 87186 36214 87190 36270
rect 87126 36210 87190 36214
rect 886 35726 950 35730
rect 886 35670 890 35726
rect 890 35670 946 35726
rect 946 35670 950 35726
rect 886 35666 950 35670
rect 966 35726 1030 35730
rect 966 35670 970 35726
rect 970 35670 1026 35726
rect 1026 35670 1030 35726
rect 966 35666 1030 35670
rect 1046 35726 1110 35730
rect 1046 35670 1050 35726
rect 1050 35670 1106 35726
rect 1106 35670 1110 35726
rect 1046 35666 1110 35670
rect 1126 35726 1190 35730
rect 1126 35670 1130 35726
rect 1130 35670 1186 35726
rect 1186 35670 1190 35726
rect 1126 35666 1190 35670
rect 84886 35726 84950 35730
rect 84886 35670 84890 35726
rect 84890 35670 84946 35726
rect 84946 35670 84950 35726
rect 84886 35666 84950 35670
rect 84966 35726 85030 35730
rect 84966 35670 84970 35726
rect 84970 35670 85026 35726
rect 85026 35670 85030 35726
rect 84966 35666 85030 35670
rect 85046 35726 85110 35730
rect 85046 35670 85050 35726
rect 85050 35670 85106 35726
rect 85106 35670 85110 35726
rect 85046 35666 85110 35670
rect 85126 35726 85190 35730
rect 85126 35670 85130 35726
rect 85130 35670 85186 35726
rect 85186 35670 85190 35726
rect 85126 35666 85190 35670
rect 2886 35182 2950 35186
rect 2886 35126 2890 35182
rect 2890 35126 2946 35182
rect 2946 35126 2950 35182
rect 2886 35122 2950 35126
rect 2966 35182 3030 35186
rect 2966 35126 2970 35182
rect 2970 35126 3026 35182
rect 3026 35126 3030 35182
rect 2966 35122 3030 35126
rect 3046 35182 3110 35186
rect 3046 35126 3050 35182
rect 3050 35126 3106 35182
rect 3106 35126 3110 35182
rect 3046 35122 3110 35126
rect 3126 35182 3190 35186
rect 3126 35126 3130 35182
rect 3130 35126 3186 35182
rect 3186 35126 3190 35182
rect 3126 35122 3190 35126
rect 86886 35182 86950 35186
rect 86886 35126 86890 35182
rect 86890 35126 86946 35182
rect 86946 35126 86950 35182
rect 86886 35122 86950 35126
rect 86966 35182 87030 35186
rect 86966 35126 86970 35182
rect 86970 35126 87026 35182
rect 87026 35126 87030 35182
rect 86966 35122 87030 35126
rect 87046 35182 87110 35186
rect 87046 35126 87050 35182
rect 87050 35126 87106 35182
rect 87106 35126 87110 35182
rect 87046 35122 87110 35126
rect 87126 35182 87190 35186
rect 87126 35126 87130 35182
rect 87130 35126 87186 35182
rect 87186 35126 87190 35182
rect 87126 35122 87190 35126
rect 84738 34918 84802 34982
rect 886 34638 950 34642
rect 886 34582 890 34638
rect 890 34582 946 34638
rect 946 34582 950 34638
rect 886 34578 950 34582
rect 966 34638 1030 34642
rect 966 34582 970 34638
rect 970 34582 1026 34638
rect 1026 34582 1030 34638
rect 966 34578 1030 34582
rect 1046 34638 1110 34642
rect 1046 34582 1050 34638
rect 1050 34582 1106 34638
rect 1106 34582 1110 34638
rect 1046 34578 1110 34582
rect 1126 34638 1190 34642
rect 1126 34582 1130 34638
rect 1130 34582 1186 34638
rect 1186 34582 1190 34638
rect 1126 34578 1190 34582
rect 84886 34638 84950 34642
rect 84886 34582 84890 34638
rect 84890 34582 84946 34638
rect 84946 34582 84950 34638
rect 84886 34578 84950 34582
rect 84966 34638 85030 34642
rect 84966 34582 84970 34638
rect 84970 34582 85026 34638
rect 85026 34582 85030 34638
rect 84966 34578 85030 34582
rect 85046 34638 85110 34642
rect 85046 34582 85050 34638
rect 85050 34582 85106 34638
rect 85106 34582 85110 34638
rect 85046 34578 85110 34582
rect 85126 34638 85190 34642
rect 85126 34582 85130 34638
rect 85130 34582 85186 34638
rect 85186 34582 85190 34638
rect 85126 34578 85190 34582
rect 2886 34094 2950 34098
rect 2886 34038 2890 34094
rect 2890 34038 2946 34094
rect 2946 34038 2950 34094
rect 2886 34034 2950 34038
rect 2966 34094 3030 34098
rect 2966 34038 2970 34094
rect 2970 34038 3026 34094
rect 3026 34038 3030 34094
rect 2966 34034 3030 34038
rect 3046 34094 3110 34098
rect 3046 34038 3050 34094
rect 3050 34038 3106 34094
rect 3106 34038 3110 34094
rect 3046 34034 3110 34038
rect 3126 34094 3190 34098
rect 3126 34038 3130 34094
rect 3130 34038 3186 34094
rect 3186 34038 3190 34094
rect 3126 34034 3190 34038
rect 86886 34094 86950 34098
rect 86886 34038 86890 34094
rect 86890 34038 86946 34094
rect 86946 34038 86950 34094
rect 86886 34034 86950 34038
rect 86966 34094 87030 34098
rect 86966 34038 86970 34094
rect 86970 34038 87026 34094
rect 87026 34038 87030 34094
rect 86966 34034 87030 34038
rect 87046 34094 87110 34098
rect 87046 34038 87050 34094
rect 87050 34038 87106 34094
rect 87106 34038 87110 34094
rect 87046 34034 87110 34038
rect 87126 34094 87190 34098
rect 87126 34038 87130 34094
rect 87130 34038 87186 34094
rect 87186 34038 87190 34094
rect 87126 34034 87190 34038
rect 83634 33830 83698 33894
rect 886 33550 950 33554
rect 886 33494 890 33550
rect 890 33494 946 33550
rect 946 33494 950 33550
rect 886 33490 950 33494
rect 966 33550 1030 33554
rect 966 33494 970 33550
rect 970 33494 1026 33550
rect 1026 33494 1030 33550
rect 966 33490 1030 33494
rect 1046 33550 1110 33554
rect 1046 33494 1050 33550
rect 1050 33494 1106 33550
rect 1106 33494 1110 33550
rect 1046 33490 1110 33494
rect 1126 33550 1190 33554
rect 1126 33494 1130 33550
rect 1130 33494 1186 33550
rect 1186 33494 1190 33550
rect 1126 33490 1190 33494
rect 84886 33550 84950 33554
rect 84886 33494 84890 33550
rect 84890 33494 84946 33550
rect 84946 33494 84950 33550
rect 84886 33490 84950 33494
rect 84966 33550 85030 33554
rect 84966 33494 84970 33550
rect 84970 33494 85026 33550
rect 85026 33494 85030 33550
rect 84966 33490 85030 33494
rect 85046 33550 85110 33554
rect 85046 33494 85050 33550
rect 85050 33494 85106 33550
rect 85106 33494 85110 33550
rect 85046 33490 85110 33494
rect 85126 33550 85190 33554
rect 85126 33494 85130 33550
rect 85130 33494 85186 33550
rect 85186 33494 85190 33550
rect 85126 33490 85190 33494
rect 2886 33006 2950 33010
rect 2886 32950 2890 33006
rect 2890 32950 2946 33006
rect 2946 32950 2950 33006
rect 2886 32946 2950 32950
rect 2966 33006 3030 33010
rect 2966 32950 2970 33006
rect 2970 32950 3026 33006
rect 3026 32950 3030 33006
rect 2966 32946 3030 32950
rect 3046 33006 3110 33010
rect 3046 32950 3050 33006
rect 3050 32950 3106 33006
rect 3106 32950 3110 33006
rect 3046 32946 3110 32950
rect 3126 33006 3190 33010
rect 3126 32950 3130 33006
rect 3130 32950 3186 33006
rect 3186 32950 3190 33006
rect 3126 32946 3190 32950
rect 86886 33006 86950 33010
rect 86886 32950 86890 33006
rect 86890 32950 86946 33006
rect 86946 32950 86950 33006
rect 86886 32946 86950 32950
rect 86966 33006 87030 33010
rect 86966 32950 86970 33006
rect 86970 32950 87026 33006
rect 87026 32950 87030 33006
rect 86966 32946 87030 32950
rect 87046 33006 87110 33010
rect 87046 32950 87050 33006
rect 87050 32950 87106 33006
rect 87106 32950 87110 33006
rect 87046 32946 87110 32950
rect 87126 33006 87190 33010
rect 87126 32950 87130 33006
rect 87130 32950 87186 33006
rect 87186 32950 87190 33006
rect 87126 32946 87190 32950
rect 84370 32742 84434 32806
rect 886 32462 950 32466
rect 886 32406 890 32462
rect 890 32406 946 32462
rect 946 32406 950 32462
rect 886 32402 950 32406
rect 966 32462 1030 32466
rect 966 32406 970 32462
rect 970 32406 1026 32462
rect 1026 32406 1030 32462
rect 966 32402 1030 32406
rect 1046 32462 1110 32466
rect 1046 32406 1050 32462
rect 1050 32406 1106 32462
rect 1106 32406 1110 32462
rect 1046 32402 1110 32406
rect 1126 32462 1190 32466
rect 1126 32406 1130 32462
rect 1130 32406 1186 32462
rect 1186 32406 1190 32462
rect 1126 32402 1190 32406
rect 84886 32462 84950 32466
rect 84886 32406 84890 32462
rect 84890 32406 84946 32462
rect 84946 32406 84950 32462
rect 84886 32402 84950 32406
rect 84966 32462 85030 32466
rect 84966 32406 84970 32462
rect 84970 32406 85026 32462
rect 85026 32406 85030 32462
rect 84966 32402 85030 32406
rect 85046 32462 85110 32466
rect 85046 32406 85050 32462
rect 85050 32406 85106 32462
rect 85106 32406 85110 32462
rect 85046 32402 85110 32406
rect 85126 32462 85190 32466
rect 85126 32406 85130 32462
rect 85130 32406 85186 32462
rect 85186 32406 85190 32462
rect 85126 32402 85190 32406
rect 2886 31918 2950 31922
rect 2886 31862 2890 31918
rect 2890 31862 2946 31918
rect 2946 31862 2950 31918
rect 2886 31858 2950 31862
rect 2966 31918 3030 31922
rect 2966 31862 2970 31918
rect 2970 31862 3026 31918
rect 3026 31862 3030 31918
rect 2966 31858 3030 31862
rect 3046 31918 3110 31922
rect 3046 31862 3050 31918
rect 3050 31862 3106 31918
rect 3106 31862 3110 31918
rect 3046 31858 3110 31862
rect 3126 31918 3190 31922
rect 3126 31862 3130 31918
rect 3130 31862 3186 31918
rect 3186 31862 3190 31918
rect 3126 31858 3190 31862
rect 86886 31918 86950 31922
rect 86886 31862 86890 31918
rect 86890 31862 86946 31918
rect 86946 31862 86950 31918
rect 86886 31858 86950 31862
rect 86966 31918 87030 31922
rect 86966 31862 86970 31918
rect 86970 31862 87026 31918
rect 87026 31862 87030 31918
rect 86966 31858 87030 31862
rect 87046 31918 87110 31922
rect 87046 31862 87050 31918
rect 87050 31862 87106 31918
rect 87106 31862 87110 31918
rect 87046 31858 87110 31862
rect 87126 31918 87190 31922
rect 87126 31862 87130 31918
rect 87130 31862 87186 31918
rect 87186 31862 87190 31918
rect 87126 31858 87190 31862
rect 886 31374 950 31378
rect 886 31318 890 31374
rect 890 31318 946 31374
rect 946 31318 950 31374
rect 886 31314 950 31318
rect 966 31374 1030 31378
rect 966 31318 970 31374
rect 970 31318 1026 31374
rect 1026 31318 1030 31374
rect 966 31314 1030 31318
rect 1046 31374 1110 31378
rect 1046 31318 1050 31374
rect 1050 31318 1106 31374
rect 1106 31318 1110 31374
rect 1046 31314 1110 31318
rect 1126 31374 1190 31378
rect 1126 31318 1130 31374
rect 1130 31318 1186 31374
rect 1186 31318 1190 31374
rect 1126 31314 1190 31318
rect 84886 31374 84950 31378
rect 84886 31318 84890 31374
rect 84890 31318 84946 31374
rect 84946 31318 84950 31374
rect 84886 31314 84950 31318
rect 84966 31374 85030 31378
rect 84966 31318 84970 31374
rect 84970 31318 85026 31374
rect 85026 31318 85030 31374
rect 84966 31314 85030 31318
rect 85046 31374 85110 31378
rect 85046 31318 85050 31374
rect 85050 31318 85106 31374
rect 85106 31318 85110 31374
rect 85046 31314 85110 31318
rect 85126 31374 85190 31378
rect 85126 31318 85130 31374
rect 85130 31318 85186 31374
rect 85186 31318 85190 31374
rect 85126 31314 85190 31318
rect 2886 30830 2950 30834
rect 2886 30774 2890 30830
rect 2890 30774 2946 30830
rect 2946 30774 2950 30830
rect 2886 30770 2950 30774
rect 2966 30830 3030 30834
rect 2966 30774 2970 30830
rect 2970 30774 3026 30830
rect 3026 30774 3030 30830
rect 2966 30770 3030 30774
rect 3046 30830 3110 30834
rect 3046 30774 3050 30830
rect 3050 30774 3106 30830
rect 3106 30774 3110 30830
rect 3046 30770 3110 30774
rect 3126 30830 3190 30834
rect 3126 30774 3130 30830
rect 3130 30774 3186 30830
rect 3186 30774 3190 30830
rect 3126 30770 3190 30774
rect 86886 30830 86950 30834
rect 86886 30774 86890 30830
rect 86890 30774 86946 30830
rect 86946 30774 86950 30830
rect 86886 30770 86950 30774
rect 86966 30830 87030 30834
rect 86966 30774 86970 30830
rect 86970 30774 87026 30830
rect 87026 30774 87030 30830
rect 86966 30770 87030 30774
rect 87046 30830 87110 30834
rect 87046 30774 87050 30830
rect 87050 30774 87106 30830
rect 87106 30774 87110 30830
rect 87046 30770 87110 30774
rect 87126 30830 87190 30834
rect 87126 30774 87130 30830
rect 87130 30774 87186 30830
rect 87186 30774 87190 30830
rect 87126 30770 87190 30774
rect 886 30286 950 30290
rect 886 30230 890 30286
rect 890 30230 946 30286
rect 946 30230 950 30286
rect 886 30226 950 30230
rect 966 30286 1030 30290
rect 966 30230 970 30286
rect 970 30230 1026 30286
rect 1026 30230 1030 30286
rect 966 30226 1030 30230
rect 1046 30286 1110 30290
rect 1046 30230 1050 30286
rect 1050 30230 1106 30286
rect 1106 30230 1110 30286
rect 1046 30226 1110 30230
rect 1126 30286 1190 30290
rect 1126 30230 1130 30286
rect 1130 30230 1186 30286
rect 1186 30230 1190 30286
rect 1126 30226 1190 30230
rect 84886 30286 84950 30290
rect 84886 30230 84890 30286
rect 84890 30230 84946 30286
rect 84946 30230 84950 30286
rect 84886 30226 84950 30230
rect 84966 30286 85030 30290
rect 84966 30230 84970 30286
rect 84970 30230 85026 30286
rect 85026 30230 85030 30286
rect 84966 30226 85030 30230
rect 85046 30286 85110 30290
rect 85046 30230 85050 30286
rect 85050 30230 85106 30286
rect 85106 30230 85110 30286
rect 85046 30226 85110 30230
rect 85126 30286 85190 30290
rect 85126 30230 85130 30286
rect 85130 30230 85186 30286
rect 85186 30230 85190 30286
rect 85126 30226 85190 30230
rect 2886 29742 2950 29746
rect 2886 29686 2890 29742
rect 2890 29686 2946 29742
rect 2946 29686 2950 29742
rect 2886 29682 2950 29686
rect 2966 29742 3030 29746
rect 2966 29686 2970 29742
rect 2970 29686 3026 29742
rect 3026 29686 3030 29742
rect 2966 29682 3030 29686
rect 3046 29742 3110 29746
rect 3046 29686 3050 29742
rect 3050 29686 3106 29742
rect 3106 29686 3110 29742
rect 3046 29682 3110 29686
rect 3126 29742 3190 29746
rect 3126 29686 3130 29742
rect 3130 29686 3186 29742
rect 3186 29686 3190 29742
rect 3126 29682 3190 29686
rect 86886 29742 86950 29746
rect 86886 29686 86890 29742
rect 86890 29686 86946 29742
rect 86946 29686 86950 29742
rect 86886 29682 86950 29686
rect 86966 29742 87030 29746
rect 86966 29686 86970 29742
rect 86970 29686 87026 29742
rect 87026 29686 87030 29742
rect 86966 29682 87030 29686
rect 87046 29742 87110 29746
rect 87046 29686 87050 29742
rect 87050 29686 87106 29742
rect 87106 29686 87110 29742
rect 87046 29682 87110 29686
rect 87126 29742 87190 29746
rect 87126 29686 87130 29742
rect 87130 29686 87186 29742
rect 87186 29686 87190 29742
rect 87126 29682 87190 29686
rect 5618 29478 5682 29542
rect 85474 29342 85538 29406
rect 886 29198 950 29202
rect 886 29142 890 29198
rect 890 29142 946 29198
rect 946 29142 950 29198
rect 886 29138 950 29142
rect 966 29198 1030 29202
rect 966 29142 970 29198
rect 970 29142 1026 29198
rect 1026 29142 1030 29198
rect 966 29138 1030 29142
rect 1046 29198 1110 29202
rect 1046 29142 1050 29198
rect 1050 29142 1106 29198
rect 1106 29142 1110 29198
rect 1046 29138 1110 29142
rect 1126 29198 1190 29202
rect 1126 29142 1130 29198
rect 1130 29142 1186 29198
rect 1186 29142 1190 29198
rect 1126 29138 1190 29142
rect 84886 29198 84950 29202
rect 84886 29142 84890 29198
rect 84890 29142 84946 29198
rect 84946 29142 84950 29198
rect 84886 29138 84950 29142
rect 84966 29198 85030 29202
rect 84966 29142 84970 29198
rect 84970 29142 85026 29198
rect 85026 29142 85030 29198
rect 84966 29138 85030 29142
rect 85046 29198 85110 29202
rect 85046 29142 85050 29198
rect 85050 29142 85106 29198
rect 85106 29142 85110 29198
rect 85046 29138 85110 29142
rect 85126 29198 85190 29202
rect 85126 29142 85130 29198
rect 85130 29142 85186 29198
rect 85186 29142 85190 29198
rect 85126 29138 85190 29142
rect 2886 28654 2950 28658
rect 2886 28598 2890 28654
rect 2890 28598 2946 28654
rect 2946 28598 2950 28654
rect 2886 28594 2950 28598
rect 2966 28654 3030 28658
rect 2966 28598 2970 28654
rect 2970 28598 3026 28654
rect 3026 28598 3030 28654
rect 2966 28594 3030 28598
rect 3046 28654 3110 28658
rect 3046 28598 3050 28654
rect 3050 28598 3106 28654
rect 3106 28598 3110 28654
rect 3046 28594 3110 28598
rect 3126 28654 3190 28658
rect 3126 28598 3130 28654
rect 3130 28598 3186 28654
rect 3186 28598 3190 28654
rect 3126 28594 3190 28598
rect 86886 28654 86950 28658
rect 86886 28598 86890 28654
rect 86890 28598 86946 28654
rect 86946 28598 86950 28654
rect 86886 28594 86950 28598
rect 86966 28654 87030 28658
rect 86966 28598 86970 28654
rect 86970 28598 87026 28654
rect 87026 28598 87030 28654
rect 86966 28594 87030 28598
rect 87046 28654 87110 28658
rect 87046 28598 87050 28654
rect 87050 28598 87106 28654
rect 87106 28598 87110 28654
rect 87046 28594 87110 28598
rect 87126 28654 87190 28658
rect 87126 28598 87130 28654
rect 87130 28598 87186 28654
rect 87186 28598 87190 28654
rect 87126 28594 87190 28598
rect 85474 28254 85538 28318
rect 886 28110 950 28114
rect 886 28054 890 28110
rect 890 28054 946 28110
rect 946 28054 950 28110
rect 886 28050 950 28054
rect 966 28110 1030 28114
rect 966 28054 970 28110
rect 970 28054 1026 28110
rect 1026 28054 1030 28110
rect 966 28050 1030 28054
rect 1046 28110 1110 28114
rect 1046 28054 1050 28110
rect 1050 28054 1106 28110
rect 1106 28054 1110 28110
rect 1046 28050 1110 28054
rect 1126 28110 1190 28114
rect 1126 28054 1130 28110
rect 1130 28054 1186 28110
rect 1186 28054 1190 28110
rect 1126 28050 1190 28054
rect 84886 28110 84950 28114
rect 84886 28054 84890 28110
rect 84890 28054 84946 28110
rect 84946 28054 84950 28110
rect 84886 28050 84950 28054
rect 84966 28110 85030 28114
rect 84966 28054 84970 28110
rect 84970 28054 85026 28110
rect 85026 28054 85030 28110
rect 84966 28050 85030 28054
rect 85046 28110 85110 28114
rect 85046 28054 85050 28110
rect 85050 28054 85106 28110
rect 85106 28054 85110 28110
rect 85046 28050 85110 28054
rect 85126 28110 85190 28114
rect 85126 28054 85130 28110
rect 85130 28054 85186 28110
rect 85186 28054 85190 28110
rect 85126 28050 85190 28054
rect 5618 27982 5682 28046
rect 2886 27566 2950 27570
rect 2886 27510 2890 27566
rect 2890 27510 2946 27566
rect 2946 27510 2950 27566
rect 2886 27506 2950 27510
rect 2966 27566 3030 27570
rect 2966 27510 2970 27566
rect 2970 27510 3026 27566
rect 3026 27510 3030 27566
rect 2966 27506 3030 27510
rect 3046 27566 3110 27570
rect 3046 27510 3050 27566
rect 3050 27510 3106 27566
rect 3106 27510 3110 27566
rect 3046 27506 3110 27510
rect 3126 27566 3190 27570
rect 3126 27510 3130 27566
rect 3130 27510 3186 27566
rect 3186 27510 3190 27566
rect 3126 27506 3190 27510
rect 86886 27566 86950 27570
rect 86886 27510 86890 27566
rect 86890 27510 86946 27566
rect 86946 27510 86950 27566
rect 86886 27506 86950 27510
rect 86966 27566 87030 27570
rect 86966 27510 86970 27566
rect 86970 27510 87026 27566
rect 87026 27510 87030 27566
rect 86966 27506 87030 27510
rect 87046 27566 87110 27570
rect 87046 27510 87050 27566
rect 87050 27510 87106 27566
rect 87106 27510 87110 27566
rect 87046 27506 87110 27510
rect 87126 27566 87190 27570
rect 87126 27510 87130 27566
rect 87130 27510 87186 27566
rect 87186 27510 87190 27566
rect 87126 27506 87190 27510
rect 886 27022 950 27026
rect 886 26966 890 27022
rect 890 26966 946 27022
rect 946 26966 950 27022
rect 886 26962 950 26966
rect 966 27022 1030 27026
rect 966 26966 970 27022
rect 970 26966 1026 27022
rect 1026 26966 1030 27022
rect 966 26962 1030 26966
rect 1046 27022 1110 27026
rect 1046 26966 1050 27022
rect 1050 26966 1106 27022
rect 1106 26966 1110 27022
rect 1046 26962 1110 26966
rect 1126 27022 1190 27026
rect 1126 26966 1130 27022
rect 1130 26966 1186 27022
rect 1186 26966 1190 27022
rect 1126 26962 1190 26966
rect 84886 27022 84950 27026
rect 84886 26966 84890 27022
rect 84890 26966 84946 27022
rect 84946 26966 84950 27022
rect 84886 26962 84950 26966
rect 84966 27022 85030 27026
rect 84966 26966 84970 27022
rect 84970 26966 85026 27022
rect 85026 26966 85030 27022
rect 84966 26962 85030 26966
rect 85046 27022 85110 27026
rect 85046 26966 85050 27022
rect 85050 26966 85106 27022
rect 85106 26966 85110 27022
rect 85046 26962 85110 26966
rect 85126 27022 85190 27026
rect 85126 26966 85130 27022
rect 85130 26966 85186 27022
rect 85186 26966 85190 27022
rect 85126 26962 85190 26966
rect 2886 26478 2950 26482
rect 2886 26422 2890 26478
rect 2890 26422 2946 26478
rect 2946 26422 2950 26478
rect 2886 26418 2950 26422
rect 2966 26478 3030 26482
rect 2966 26422 2970 26478
rect 2970 26422 3026 26478
rect 3026 26422 3030 26478
rect 2966 26418 3030 26422
rect 3046 26478 3110 26482
rect 3046 26422 3050 26478
rect 3050 26422 3106 26478
rect 3106 26422 3110 26478
rect 3046 26418 3110 26422
rect 3126 26478 3190 26482
rect 3126 26422 3130 26478
rect 3130 26422 3186 26478
rect 3186 26422 3190 26478
rect 3126 26418 3190 26422
rect 86886 26478 86950 26482
rect 86886 26422 86890 26478
rect 86890 26422 86946 26478
rect 86946 26422 86950 26478
rect 86886 26418 86950 26422
rect 86966 26478 87030 26482
rect 86966 26422 86970 26478
rect 86970 26422 87026 26478
rect 87026 26422 87030 26478
rect 86966 26418 87030 26422
rect 87046 26478 87110 26482
rect 87046 26422 87050 26478
rect 87050 26422 87106 26478
rect 87106 26422 87110 26478
rect 87046 26418 87110 26422
rect 87126 26478 87190 26482
rect 87126 26422 87130 26478
rect 87130 26422 87186 26478
rect 87186 26422 87190 26478
rect 87126 26418 87190 26422
rect 886 25934 950 25938
rect 886 25878 890 25934
rect 890 25878 946 25934
rect 946 25878 950 25934
rect 886 25874 950 25878
rect 966 25934 1030 25938
rect 966 25878 970 25934
rect 970 25878 1026 25934
rect 1026 25878 1030 25934
rect 966 25874 1030 25878
rect 1046 25934 1110 25938
rect 1046 25878 1050 25934
rect 1050 25878 1106 25934
rect 1106 25878 1110 25934
rect 1046 25874 1110 25878
rect 1126 25934 1190 25938
rect 1126 25878 1130 25934
rect 1130 25878 1186 25934
rect 1186 25878 1190 25934
rect 1126 25874 1190 25878
rect 84886 25934 84950 25938
rect 84886 25878 84890 25934
rect 84890 25878 84946 25934
rect 84946 25878 84950 25934
rect 84886 25874 84950 25878
rect 84966 25934 85030 25938
rect 84966 25878 84970 25934
rect 84970 25878 85026 25934
rect 85026 25878 85030 25934
rect 84966 25874 85030 25878
rect 85046 25934 85110 25938
rect 85046 25878 85050 25934
rect 85050 25878 85106 25934
rect 85106 25878 85110 25934
rect 85046 25874 85110 25878
rect 85126 25934 85190 25938
rect 85126 25878 85130 25934
rect 85130 25878 85186 25934
rect 85186 25878 85190 25934
rect 85126 25874 85190 25878
rect 2886 25390 2950 25394
rect 2886 25334 2890 25390
rect 2890 25334 2946 25390
rect 2946 25334 2950 25390
rect 2886 25330 2950 25334
rect 2966 25390 3030 25394
rect 2966 25334 2970 25390
rect 2970 25334 3026 25390
rect 3026 25334 3030 25390
rect 2966 25330 3030 25334
rect 3046 25390 3110 25394
rect 3046 25334 3050 25390
rect 3050 25334 3106 25390
rect 3106 25334 3110 25390
rect 3046 25330 3110 25334
rect 3126 25390 3190 25394
rect 3126 25334 3130 25390
rect 3130 25334 3186 25390
rect 3186 25334 3190 25390
rect 3126 25330 3190 25334
rect 86886 25390 86950 25394
rect 86886 25334 86890 25390
rect 86890 25334 86946 25390
rect 86946 25334 86950 25390
rect 86886 25330 86950 25334
rect 86966 25390 87030 25394
rect 86966 25334 86970 25390
rect 86970 25334 87026 25390
rect 87026 25334 87030 25390
rect 86966 25330 87030 25334
rect 87046 25390 87110 25394
rect 87046 25334 87050 25390
rect 87050 25334 87106 25390
rect 87106 25334 87110 25390
rect 87046 25330 87110 25334
rect 87126 25390 87190 25394
rect 87126 25334 87130 25390
rect 87130 25334 87186 25390
rect 87186 25334 87190 25390
rect 87126 25330 87190 25334
rect 886 24846 950 24850
rect 886 24790 890 24846
rect 890 24790 946 24846
rect 946 24790 950 24846
rect 886 24786 950 24790
rect 966 24846 1030 24850
rect 966 24790 970 24846
rect 970 24790 1026 24846
rect 1026 24790 1030 24846
rect 966 24786 1030 24790
rect 1046 24846 1110 24850
rect 1046 24790 1050 24846
rect 1050 24790 1106 24846
rect 1106 24790 1110 24846
rect 1046 24786 1110 24790
rect 1126 24846 1190 24850
rect 1126 24790 1130 24846
rect 1130 24790 1186 24846
rect 1186 24790 1190 24846
rect 1126 24786 1190 24790
rect 84886 24846 84950 24850
rect 84886 24790 84890 24846
rect 84890 24790 84946 24846
rect 84946 24790 84950 24846
rect 84886 24786 84950 24790
rect 84966 24846 85030 24850
rect 84966 24790 84970 24846
rect 84970 24790 85026 24846
rect 85026 24790 85030 24846
rect 84966 24786 85030 24790
rect 85046 24846 85110 24850
rect 85046 24790 85050 24846
rect 85050 24790 85106 24846
rect 85106 24790 85110 24846
rect 85046 24786 85110 24790
rect 85126 24846 85190 24850
rect 85126 24790 85130 24846
rect 85130 24790 85186 24846
rect 85186 24790 85190 24846
rect 85126 24786 85190 24790
rect 82346 24446 82410 24510
rect 2886 24302 2950 24306
rect 2886 24246 2890 24302
rect 2890 24246 2946 24302
rect 2946 24246 2950 24302
rect 2886 24242 2950 24246
rect 2966 24302 3030 24306
rect 2966 24246 2970 24302
rect 2970 24246 3026 24302
rect 3026 24246 3030 24302
rect 2966 24242 3030 24246
rect 3046 24302 3110 24306
rect 3046 24246 3050 24302
rect 3050 24246 3106 24302
rect 3106 24246 3110 24302
rect 3046 24242 3110 24246
rect 3126 24302 3190 24306
rect 3126 24246 3130 24302
rect 3130 24246 3186 24302
rect 3186 24246 3190 24302
rect 3126 24242 3190 24246
rect 82346 24038 82410 24102
rect 86886 24302 86950 24306
rect 86886 24246 86890 24302
rect 86890 24246 86946 24302
rect 86946 24246 86950 24302
rect 86886 24242 86950 24246
rect 86966 24302 87030 24306
rect 86966 24246 86970 24302
rect 86970 24246 87026 24302
rect 87026 24246 87030 24302
rect 86966 24242 87030 24246
rect 87046 24302 87110 24306
rect 87046 24246 87050 24302
rect 87050 24246 87106 24302
rect 87106 24246 87110 24302
rect 87046 24242 87110 24246
rect 87126 24302 87190 24306
rect 87126 24246 87130 24302
rect 87130 24246 87186 24302
rect 87186 24246 87190 24302
rect 87126 24242 87190 24246
rect 84002 24174 84066 24238
rect 886 23758 950 23762
rect 886 23702 890 23758
rect 890 23702 946 23758
rect 946 23702 950 23758
rect 886 23698 950 23702
rect 966 23758 1030 23762
rect 966 23702 970 23758
rect 970 23702 1026 23758
rect 1026 23702 1030 23758
rect 966 23698 1030 23702
rect 1046 23758 1110 23762
rect 1046 23702 1050 23758
rect 1050 23702 1106 23758
rect 1106 23702 1110 23758
rect 1046 23698 1110 23702
rect 1126 23758 1190 23762
rect 1126 23702 1130 23758
rect 1130 23702 1186 23758
rect 1186 23702 1190 23758
rect 1126 23698 1190 23702
rect 84886 23758 84950 23762
rect 84886 23702 84890 23758
rect 84890 23702 84946 23758
rect 84946 23702 84950 23758
rect 84886 23698 84950 23702
rect 84966 23758 85030 23762
rect 84966 23702 84970 23758
rect 84970 23702 85026 23758
rect 85026 23702 85030 23758
rect 84966 23698 85030 23702
rect 85046 23758 85110 23762
rect 85046 23702 85050 23758
rect 85050 23702 85106 23758
rect 85106 23702 85110 23758
rect 85046 23698 85110 23702
rect 85126 23758 85190 23762
rect 85126 23702 85130 23758
rect 85130 23702 85186 23758
rect 85186 23702 85190 23758
rect 85126 23698 85190 23702
rect 2886 23214 2950 23218
rect 2886 23158 2890 23214
rect 2890 23158 2946 23214
rect 2946 23158 2950 23214
rect 2886 23154 2950 23158
rect 2966 23214 3030 23218
rect 2966 23158 2970 23214
rect 2970 23158 3026 23214
rect 3026 23158 3030 23214
rect 2966 23154 3030 23158
rect 3046 23214 3110 23218
rect 3046 23158 3050 23214
rect 3050 23158 3106 23214
rect 3106 23158 3110 23214
rect 3046 23154 3110 23158
rect 3126 23214 3190 23218
rect 3126 23158 3130 23214
rect 3130 23158 3186 23214
rect 3186 23158 3190 23214
rect 3126 23154 3190 23158
rect 86886 23214 86950 23218
rect 86886 23158 86890 23214
rect 86890 23158 86946 23214
rect 86946 23158 86950 23214
rect 86886 23154 86950 23158
rect 86966 23214 87030 23218
rect 86966 23158 86970 23214
rect 86970 23158 87026 23214
rect 87026 23158 87030 23214
rect 86966 23154 87030 23158
rect 87046 23214 87110 23218
rect 87046 23158 87050 23214
rect 87050 23158 87106 23214
rect 87106 23158 87110 23214
rect 87046 23154 87110 23158
rect 87126 23214 87190 23218
rect 87126 23158 87130 23214
rect 87130 23158 87186 23214
rect 87186 23158 87190 23214
rect 87126 23154 87190 23158
rect 4146 22814 4210 22878
rect 886 22670 950 22674
rect 886 22614 890 22670
rect 890 22614 946 22670
rect 946 22614 950 22670
rect 886 22610 950 22614
rect 966 22670 1030 22674
rect 966 22614 970 22670
rect 970 22614 1026 22670
rect 1026 22614 1030 22670
rect 966 22610 1030 22614
rect 1046 22670 1110 22674
rect 1046 22614 1050 22670
rect 1050 22614 1106 22670
rect 1106 22614 1110 22670
rect 1046 22610 1110 22614
rect 1126 22670 1190 22674
rect 1126 22614 1130 22670
rect 1130 22614 1186 22670
rect 1186 22614 1190 22670
rect 1126 22610 1190 22614
rect 84886 22670 84950 22674
rect 84886 22614 84890 22670
rect 84890 22614 84946 22670
rect 84946 22614 84950 22670
rect 84886 22610 84950 22614
rect 84966 22670 85030 22674
rect 84966 22614 84970 22670
rect 84970 22614 85026 22670
rect 85026 22614 85030 22670
rect 84966 22610 85030 22614
rect 85046 22670 85110 22674
rect 85046 22614 85050 22670
rect 85050 22614 85106 22670
rect 85106 22614 85110 22670
rect 85046 22610 85110 22614
rect 85126 22670 85190 22674
rect 85126 22614 85130 22670
rect 85130 22614 85186 22670
rect 85186 22614 85190 22670
rect 85126 22610 85190 22614
rect 2886 22126 2950 22130
rect 2886 22070 2890 22126
rect 2890 22070 2946 22126
rect 2946 22070 2950 22126
rect 2886 22066 2950 22070
rect 2966 22126 3030 22130
rect 2966 22070 2970 22126
rect 2970 22070 3026 22126
rect 3026 22070 3030 22126
rect 2966 22066 3030 22070
rect 3046 22126 3110 22130
rect 3046 22070 3050 22126
rect 3050 22070 3106 22126
rect 3106 22070 3110 22126
rect 3046 22066 3110 22070
rect 3126 22126 3190 22130
rect 3126 22070 3130 22126
rect 3130 22070 3186 22126
rect 3186 22070 3190 22126
rect 3126 22066 3190 22070
rect 86886 22126 86950 22130
rect 86886 22070 86890 22126
rect 86890 22070 86946 22126
rect 86946 22070 86950 22126
rect 86886 22066 86950 22070
rect 86966 22126 87030 22130
rect 86966 22070 86970 22126
rect 86970 22070 87026 22126
rect 87026 22070 87030 22126
rect 86966 22066 87030 22070
rect 87046 22126 87110 22130
rect 87046 22070 87050 22126
rect 87050 22070 87106 22126
rect 87106 22070 87110 22126
rect 87046 22066 87110 22070
rect 87126 22126 87190 22130
rect 87126 22070 87130 22126
rect 87130 22070 87186 22126
rect 87186 22070 87190 22126
rect 87126 22066 87190 22070
rect 84186 21862 84250 21926
rect 886 21582 950 21586
rect 886 21526 890 21582
rect 890 21526 946 21582
rect 946 21526 950 21582
rect 886 21522 950 21526
rect 966 21582 1030 21586
rect 966 21526 970 21582
rect 970 21526 1026 21582
rect 1026 21526 1030 21582
rect 966 21522 1030 21526
rect 1046 21582 1110 21586
rect 1046 21526 1050 21582
rect 1050 21526 1106 21582
rect 1106 21526 1110 21582
rect 1046 21522 1110 21526
rect 1126 21582 1190 21586
rect 1126 21526 1130 21582
rect 1130 21526 1186 21582
rect 1186 21526 1190 21582
rect 1126 21522 1190 21526
rect 84886 21582 84950 21586
rect 84886 21526 84890 21582
rect 84890 21526 84946 21582
rect 84946 21526 84950 21582
rect 84886 21522 84950 21526
rect 84966 21582 85030 21586
rect 84966 21526 84970 21582
rect 84970 21526 85026 21582
rect 85026 21526 85030 21582
rect 84966 21522 85030 21526
rect 85046 21582 85110 21586
rect 85046 21526 85050 21582
rect 85050 21526 85106 21582
rect 85106 21526 85110 21582
rect 85046 21522 85110 21526
rect 85126 21582 85190 21586
rect 85126 21526 85130 21582
rect 85130 21526 85186 21582
rect 85186 21526 85190 21582
rect 85126 21522 85190 21526
rect 2886 21038 2950 21042
rect 2886 20982 2890 21038
rect 2890 20982 2946 21038
rect 2946 20982 2950 21038
rect 2886 20978 2950 20982
rect 2966 21038 3030 21042
rect 2966 20982 2970 21038
rect 2970 20982 3026 21038
rect 3026 20982 3030 21038
rect 2966 20978 3030 20982
rect 3046 21038 3110 21042
rect 3046 20982 3050 21038
rect 3050 20982 3106 21038
rect 3106 20982 3110 21038
rect 3046 20978 3110 20982
rect 3126 21038 3190 21042
rect 3126 20982 3130 21038
rect 3130 20982 3186 21038
rect 3186 20982 3190 21038
rect 3126 20978 3190 20982
rect 86886 21038 86950 21042
rect 86886 20982 86890 21038
rect 86890 20982 86946 21038
rect 86946 20982 86950 21038
rect 86886 20978 86950 20982
rect 86966 21038 87030 21042
rect 86966 20982 86970 21038
rect 86970 20982 87026 21038
rect 87026 20982 87030 21038
rect 86966 20978 87030 20982
rect 87046 21038 87110 21042
rect 87046 20982 87050 21038
rect 87050 20982 87106 21038
rect 87106 20982 87110 21038
rect 87046 20978 87110 20982
rect 87126 21038 87190 21042
rect 87126 20982 87130 21038
rect 87130 20982 87186 21038
rect 87186 20982 87190 21038
rect 87126 20978 87190 20982
rect 886 20494 950 20498
rect 886 20438 890 20494
rect 890 20438 946 20494
rect 946 20438 950 20494
rect 886 20434 950 20438
rect 966 20494 1030 20498
rect 966 20438 970 20494
rect 970 20438 1026 20494
rect 1026 20438 1030 20494
rect 966 20434 1030 20438
rect 1046 20494 1110 20498
rect 1046 20438 1050 20494
rect 1050 20438 1106 20494
rect 1106 20438 1110 20494
rect 1046 20434 1110 20438
rect 1126 20494 1190 20498
rect 1126 20438 1130 20494
rect 1130 20438 1186 20494
rect 1186 20438 1190 20494
rect 1126 20434 1190 20438
rect 84886 20494 84950 20498
rect 84886 20438 84890 20494
rect 84890 20438 84946 20494
rect 84946 20438 84950 20494
rect 84886 20434 84950 20438
rect 84966 20494 85030 20498
rect 84966 20438 84970 20494
rect 84970 20438 85026 20494
rect 85026 20438 85030 20494
rect 84966 20434 85030 20438
rect 85046 20494 85110 20498
rect 85046 20438 85050 20494
rect 85050 20438 85106 20494
rect 85106 20438 85110 20494
rect 85046 20434 85110 20438
rect 85126 20494 85190 20498
rect 85126 20438 85130 20494
rect 85130 20438 85186 20494
rect 85186 20438 85190 20494
rect 85126 20434 85190 20438
rect 2886 19950 2950 19954
rect 2886 19894 2890 19950
rect 2890 19894 2946 19950
rect 2946 19894 2950 19950
rect 2886 19890 2950 19894
rect 2966 19950 3030 19954
rect 2966 19894 2970 19950
rect 2970 19894 3026 19950
rect 3026 19894 3030 19950
rect 2966 19890 3030 19894
rect 3046 19950 3110 19954
rect 3046 19894 3050 19950
rect 3050 19894 3106 19950
rect 3106 19894 3110 19950
rect 3046 19890 3110 19894
rect 3126 19950 3190 19954
rect 3126 19894 3130 19950
rect 3130 19894 3186 19950
rect 3186 19894 3190 19950
rect 3126 19890 3190 19894
rect 86886 19950 86950 19954
rect 86886 19894 86890 19950
rect 86890 19894 86946 19950
rect 86946 19894 86950 19950
rect 86886 19890 86950 19894
rect 86966 19950 87030 19954
rect 86966 19894 86970 19950
rect 86970 19894 87026 19950
rect 87026 19894 87030 19950
rect 86966 19890 87030 19894
rect 87046 19950 87110 19954
rect 87046 19894 87050 19950
rect 87050 19894 87106 19950
rect 87106 19894 87110 19950
rect 87046 19890 87110 19894
rect 87126 19950 87190 19954
rect 87126 19894 87130 19950
rect 87130 19894 87186 19950
rect 87186 19894 87190 19950
rect 87126 19890 87190 19894
rect 84002 19550 84066 19614
rect 886 19406 950 19410
rect 886 19350 890 19406
rect 890 19350 946 19406
rect 946 19350 950 19406
rect 886 19346 950 19350
rect 966 19406 1030 19410
rect 966 19350 970 19406
rect 970 19350 1026 19406
rect 1026 19350 1030 19406
rect 966 19346 1030 19350
rect 1046 19406 1110 19410
rect 1046 19350 1050 19406
rect 1050 19350 1106 19406
rect 1106 19350 1110 19406
rect 1046 19346 1110 19350
rect 1126 19406 1190 19410
rect 1126 19350 1130 19406
rect 1130 19350 1186 19406
rect 1186 19350 1190 19406
rect 1126 19346 1190 19350
rect 84886 19406 84950 19410
rect 84886 19350 84890 19406
rect 84890 19350 84946 19406
rect 84946 19350 84950 19406
rect 84886 19346 84950 19350
rect 84966 19406 85030 19410
rect 84966 19350 84970 19406
rect 84970 19350 85026 19406
rect 85026 19350 85030 19406
rect 84966 19346 85030 19350
rect 85046 19406 85110 19410
rect 85046 19350 85050 19406
rect 85050 19350 85106 19406
rect 85106 19350 85110 19406
rect 85046 19346 85110 19350
rect 85126 19406 85190 19410
rect 85126 19350 85130 19406
rect 85130 19350 85186 19406
rect 85186 19350 85190 19406
rect 85126 19346 85190 19350
rect 2886 18862 2950 18866
rect 2886 18806 2890 18862
rect 2890 18806 2946 18862
rect 2946 18806 2950 18862
rect 2886 18802 2950 18806
rect 2966 18862 3030 18866
rect 2966 18806 2970 18862
rect 2970 18806 3026 18862
rect 3026 18806 3030 18862
rect 2966 18802 3030 18806
rect 3046 18862 3110 18866
rect 3046 18806 3050 18862
rect 3050 18806 3106 18862
rect 3106 18806 3110 18862
rect 3046 18802 3110 18806
rect 3126 18862 3190 18866
rect 3126 18806 3130 18862
rect 3130 18806 3186 18862
rect 3186 18806 3190 18862
rect 3126 18802 3190 18806
rect 86886 18862 86950 18866
rect 86886 18806 86890 18862
rect 86890 18806 86946 18862
rect 86946 18806 86950 18862
rect 86886 18802 86950 18806
rect 86966 18862 87030 18866
rect 86966 18806 86970 18862
rect 86970 18806 87026 18862
rect 87026 18806 87030 18862
rect 86966 18802 87030 18806
rect 87046 18862 87110 18866
rect 87046 18806 87050 18862
rect 87050 18806 87106 18862
rect 87106 18806 87110 18862
rect 87046 18802 87110 18806
rect 87126 18862 87190 18866
rect 87126 18806 87130 18862
rect 87130 18806 87186 18862
rect 87186 18806 87190 18862
rect 87126 18802 87190 18806
rect 886 18318 950 18322
rect 886 18262 890 18318
rect 890 18262 946 18318
rect 946 18262 950 18318
rect 886 18258 950 18262
rect 966 18318 1030 18322
rect 966 18262 970 18318
rect 970 18262 1026 18318
rect 1026 18262 1030 18318
rect 966 18258 1030 18262
rect 1046 18318 1110 18322
rect 1046 18262 1050 18318
rect 1050 18262 1106 18318
rect 1106 18262 1110 18318
rect 1046 18258 1110 18262
rect 1126 18318 1190 18322
rect 1126 18262 1130 18318
rect 1130 18262 1186 18318
rect 1186 18262 1190 18318
rect 1126 18258 1190 18262
rect 84886 18318 84950 18322
rect 84886 18262 84890 18318
rect 84890 18262 84946 18318
rect 84946 18262 84950 18318
rect 84886 18258 84950 18262
rect 84966 18318 85030 18322
rect 84966 18262 84970 18318
rect 84970 18262 85026 18318
rect 85026 18262 85030 18318
rect 84966 18258 85030 18262
rect 85046 18318 85110 18322
rect 85046 18262 85050 18318
rect 85050 18262 85106 18318
rect 85106 18262 85110 18318
rect 85046 18258 85110 18262
rect 85126 18318 85190 18322
rect 85126 18262 85130 18318
rect 85130 18262 85186 18318
rect 85186 18262 85190 18318
rect 85126 18258 85190 18262
rect 2886 17774 2950 17778
rect 2886 17718 2890 17774
rect 2890 17718 2946 17774
rect 2946 17718 2950 17774
rect 2886 17714 2950 17718
rect 2966 17774 3030 17778
rect 2966 17718 2970 17774
rect 2970 17718 3026 17774
rect 3026 17718 3030 17774
rect 2966 17714 3030 17718
rect 3046 17774 3110 17778
rect 3046 17718 3050 17774
rect 3050 17718 3106 17774
rect 3106 17718 3110 17774
rect 3046 17714 3110 17718
rect 3126 17774 3190 17778
rect 3126 17718 3130 17774
rect 3130 17718 3186 17774
rect 3186 17718 3190 17774
rect 3126 17714 3190 17718
rect 86886 17774 86950 17778
rect 86886 17718 86890 17774
rect 86890 17718 86946 17774
rect 86946 17718 86950 17774
rect 86886 17714 86950 17718
rect 86966 17774 87030 17778
rect 86966 17718 86970 17774
rect 86970 17718 87026 17774
rect 87026 17718 87030 17774
rect 86966 17714 87030 17718
rect 87046 17774 87110 17778
rect 87046 17718 87050 17774
rect 87050 17718 87106 17774
rect 87106 17718 87110 17774
rect 87046 17714 87110 17718
rect 87126 17774 87190 17778
rect 87126 17718 87130 17774
rect 87130 17718 87186 17774
rect 87186 17718 87190 17774
rect 87126 17714 87190 17718
rect 886 17230 950 17234
rect 886 17174 890 17230
rect 890 17174 946 17230
rect 946 17174 950 17230
rect 886 17170 950 17174
rect 966 17230 1030 17234
rect 966 17174 970 17230
rect 970 17174 1026 17230
rect 1026 17174 1030 17230
rect 966 17170 1030 17174
rect 1046 17230 1110 17234
rect 1046 17174 1050 17230
rect 1050 17174 1106 17230
rect 1106 17174 1110 17230
rect 1046 17170 1110 17174
rect 1126 17230 1190 17234
rect 1126 17174 1130 17230
rect 1130 17174 1186 17230
rect 1186 17174 1190 17230
rect 1126 17170 1190 17174
rect 84886 17230 84950 17234
rect 84886 17174 84890 17230
rect 84890 17174 84946 17230
rect 84946 17174 84950 17230
rect 84886 17170 84950 17174
rect 84966 17230 85030 17234
rect 84966 17174 84970 17230
rect 84970 17174 85026 17230
rect 85026 17174 85030 17230
rect 84966 17170 85030 17174
rect 85046 17230 85110 17234
rect 85046 17174 85050 17230
rect 85050 17174 85106 17230
rect 85106 17174 85110 17230
rect 85046 17170 85110 17174
rect 85126 17230 85190 17234
rect 85126 17174 85130 17230
rect 85130 17174 85186 17230
rect 85186 17174 85190 17230
rect 85126 17170 85190 17174
rect 2886 16686 2950 16690
rect 2886 16630 2890 16686
rect 2890 16630 2946 16686
rect 2946 16630 2950 16686
rect 2886 16626 2950 16630
rect 2966 16686 3030 16690
rect 2966 16630 2970 16686
rect 2970 16630 3026 16686
rect 3026 16630 3030 16686
rect 2966 16626 3030 16630
rect 3046 16686 3110 16690
rect 3046 16630 3050 16686
rect 3050 16630 3106 16686
rect 3106 16630 3110 16686
rect 3046 16626 3110 16630
rect 3126 16686 3190 16690
rect 3126 16630 3130 16686
rect 3130 16630 3186 16686
rect 3186 16630 3190 16686
rect 3126 16626 3190 16630
rect 86886 16686 86950 16690
rect 86886 16630 86890 16686
rect 86890 16630 86946 16686
rect 86946 16630 86950 16686
rect 86886 16626 86950 16630
rect 86966 16686 87030 16690
rect 86966 16630 86970 16686
rect 86970 16630 87026 16686
rect 87026 16630 87030 16686
rect 86966 16626 87030 16630
rect 87046 16686 87110 16690
rect 87046 16630 87050 16686
rect 87050 16630 87106 16686
rect 87106 16630 87110 16686
rect 87046 16626 87110 16630
rect 87126 16686 87190 16690
rect 87126 16630 87130 16686
rect 87130 16630 87186 16686
rect 87186 16630 87190 16686
rect 87126 16626 87190 16630
rect 886 16142 950 16146
rect 886 16086 890 16142
rect 890 16086 946 16142
rect 946 16086 950 16142
rect 886 16082 950 16086
rect 966 16142 1030 16146
rect 966 16086 970 16142
rect 970 16086 1026 16142
rect 1026 16086 1030 16142
rect 966 16082 1030 16086
rect 1046 16142 1110 16146
rect 1046 16086 1050 16142
rect 1050 16086 1106 16142
rect 1106 16086 1110 16142
rect 1046 16082 1110 16086
rect 1126 16142 1190 16146
rect 1126 16086 1130 16142
rect 1130 16086 1186 16142
rect 1186 16086 1190 16142
rect 1126 16082 1190 16086
rect 84886 16142 84950 16146
rect 84886 16086 84890 16142
rect 84890 16086 84946 16142
rect 84946 16086 84950 16142
rect 84886 16082 84950 16086
rect 84966 16142 85030 16146
rect 84966 16086 84970 16142
rect 84970 16086 85026 16142
rect 85026 16086 85030 16142
rect 84966 16082 85030 16086
rect 85046 16142 85110 16146
rect 85046 16086 85050 16142
rect 85050 16086 85106 16142
rect 85106 16086 85110 16142
rect 85046 16082 85110 16086
rect 85126 16142 85190 16146
rect 85126 16086 85130 16142
rect 85130 16086 85186 16142
rect 85186 16086 85190 16142
rect 85126 16082 85190 16086
rect 2886 15598 2950 15602
rect 2886 15542 2890 15598
rect 2890 15542 2946 15598
rect 2946 15542 2950 15598
rect 2886 15538 2950 15542
rect 2966 15598 3030 15602
rect 2966 15542 2970 15598
rect 2970 15542 3026 15598
rect 3026 15542 3030 15598
rect 2966 15538 3030 15542
rect 3046 15598 3110 15602
rect 3046 15542 3050 15598
rect 3050 15542 3106 15598
rect 3106 15542 3110 15598
rect 3046 15538 3110 15542
rect 3126 15598 3190 15602
rect 3126 15542 3130 15598
rect 3130 15542 3186 15598
rect 3186 15542 3190 15598
rect 3126 15538 3190 15542
rect 86886 15598 86950 15602
rect 86886 15542 86890 15598
rect 86890 15542 86946 15598
rect 86946 15542 86950 15598
rect 86886 15538 86950 15542
rect 86966 15598 87030 15602
rect 86966 15542 86970 15598
rect 86970 15542 87026 15598
rect 87026 15542 87030 15598
rect 86966 15538 87030 15542
rect 87046 15598 87110 15602
rect 87046 15542 87050 15598
rect 87050 15542 87106 15598
rect 87106 15542 87110 15598
rect 87046 15538 87110 15542
rect 87126 15598 87190 15602
rect 87126 15542 87130 15598
rect 87130 15542 87186 15598
rect 87186 15542 87190 15598
rect 87126 15538 87190 15542
rect 82346 15470 82410 15534
rect 82898 15470 82962 15534
rect 82346 15334 82410 15398
rect 886 15054 950 15058
rect 886 14998 890 15054
rect 890 14998 946 15054
rect 946 14998 950 15054
rect 886 14994 950 14998
rect 966 15054 1030 15058
rect 966 14998 970 15054
rect 970 14998 1026 15054
rect 1026 14998 1030 15054
rect 966 14994 1030 14998
rect 1046 15054 1110 15058
rect 1046 14998 1050 15054
rect 1050 14998 1106 15054
rect 1106 14998 1110 15054
rect 1046 14994 1110 14998
rect 1126 15054 1190 15058
rect 1126 14998 1130 15054
rect 1130 14998 1186 15054
rect 1186 14998 1190 15054
rect 1126 14994 1190 14998
rect 84886 15054 84950 15058
rect 84886 14998 84890 15054
rect 84890 14998 84946 15054
rect 84946 14998 84950 15054
rect 84886 14994 84950 14998
rect 84966 15054 85030 15058
rect 84966 14998 84970 15054
rect 84970 14998 85026 15054
rect 85026 14998 85030 15054
rect 84966 14994 85030 14998
rect 85046 15054 85110 15058
rect 85046 14998 85050 15054
rect 85050 14998 85106 15054
rect 85106 14998 85110 15054
rect 85046 14994 85110 14998
rect 85126 15054 85190 15058
rect 85126 14998 85130 15054
rect 85130 14998 85186 15054
rect 85186 14998 85190 15054
rect 85126 14994 85190 14998
rect 2886 14510 2950 14514
rect 2886 14454 2890 14510
rect 2890 14454 2946 14510
rect 2946 14454 2950 14510
rect 2886 14450 2950 14454
rect 2966 14510 3030 14514
rect 2966 14454 2970 14510
rect 2970 14454 3026 14510
rect 3026 14454 3030 14510
rect 2966 14450 3030 14454
rect 3046 14510 3110 14514
rect 3046 14454 3050 14510
rect 3050 14454 3106 14510
rect 3106 14454 3110 14510
rect 3046 14450 3110 14454
rect 3126 14510 3190 14514
rect 3126 14454 3130 14510
rect 3130 14454 3186 14510
rect 3186 14454 3190 14510
rect 3126 14450 3190 14454
rect 86886 14510 86950 14514
rect 86886 14454 86890 14510
rect 86890 14454 86946 14510
rect 86946 14454 86950 14510
rect 86886 14450 86950 14454
rect 86966 14510 87030 14514
rect 86966 14454 86970 14510
rect 86970 14454 87026 14510
rect 87026 14454 87030 14510
rect 86966 14450 87030 14454
rect 87046 14510 87110 14514
rect 87046 14454 87050 14510
rect 87050 14454 87106 14510
rect 87106 14454 87110 14510
rect 87046 14450 87110 14454
rect 87126 14510 87190 14514
rect 87126 14454 87130 14510
rect 87130 14454 87186 14510
rect 87186 14454 87190 14510
rect 87126 14450 87190 14454
rect 886 13966 950 13970
rect 886 13910 890 13966
rect 890 13910 946 13966
rect 946 13910 950 13966
rect 886 13906 950 13910
rect 966 13966 1030 13970
rect 966 13910 970 13966
rect 970 13910 1026 13966
rect 1026 13910 1030 13966
rect 966 13906 1030 13910
rect 1046 13966 1110 13970
rect 1046 13910 1050 13966
rect 1050 13910 1106 13966
rect 1106 13910 1110 13966
rect 1046 13906 1110 13910
rect 1126 13966 1190 13970
rect 1126 13910 1130 13966
rect 1130 13910 1186 13966
rect 1186 13910 1190 13966
rect 1126 13906 1190 13910
rect 84886 13966 84950 13970
rect 84886 13910 84890 13966
rect 84890 13910 84946 13966
rect 84946 13910 84950 13966
rect 84886 13906 84950 13910
rect 84966 13966 85030 13970
rect 84966 13910 84970 13966
rect 84970 13910 85026 13966
rect 85026 13910 85030 13966
rect 84966 13906 85030 13910
rect 85046 13966 85110 13970
rect 85046 13910 85050 13966
rect 85050 13910 85106 13966
rect 85106 13910 85110 13966
rect 85046 13906 85110 13910
rect 85126 13966 85190 13970
rect 85126 13910 85130 13966
rect 85130 13910 85186 13966
rect 85186 13910 85190 13966
rect 85126 13906 85190 13910
rect 2886 13422 2950 13426
rect 2886 13366 2890 13422
rect 2890 13366 2946 13422
rect 2946 13366 2950 13422
rect 2886 13362 2950 13366
rect 2966 13422 3030 13426
rect 2966 13366 2970 13422
rect 2970 13366 3026 13422
rect 3026 13366 3030 13422
rect 2966 13362 3030 13366
rect 3046 13422 3110 13426
rect 3046 13366 3050 13422
rect 3050 13366 3106 13422
rect 3106 13366 3110 13422
rect 3046 13362 3110 13366
rect 3126 13422 3190 13426
rect 3126 13366 3130 13422
rect 3130 13366 3186 13422
rect 3186 13366 3190 13422
rect 3126 13362 3190 13366
rect 86886 13422 86950 13426
rect 86886 13366 86890 13422
rect 86890 13366 86946 13422
rect 86946 13366 86950 13422
rect 86886 13362 86950 13366
rect 86966 13422 87030 13426
rect 86966 13366 86970 13422
rect 86970 13366 87026 13422
rect 87026 13366 87030 13422
rect 86966 13362 87030 13366
rect 87046 13422 87110 13426
rect 87046 13366 87050 13422
rect 87050 13366 87106 13422
rect 87106 13366 87110 13422
rect 87046 13362 87110 13366
rect 87126 13422 87190 13426
rect 87126 13366 87130 13422
rect 87130 13366 87186 13422
rect 87186 13366 87190 13422
rect 87126 13362 87190 13366
rect 886 12878 950 12882
rect 886 12822 890 12878
rect 890 12822 946 12878
rect 946 12822 950 12878
rect 886 12818 950 12822
rect 966 12878 1030 12882
rect 966 12822 970 12878
rect 970 12822 1026 12878
rect 1026 12822 1030 12878
rect 966 12818 1030 12822
rect 1046 12878 1110 12882
rect 1046 12822 1050 12878
rect 1050 12822 1106 12878
rect 1106 12822 1110 12878
rect 1046 12818 1110 12822
rect 1126 12878 1190 12882
rect 1126 12822 1130 12878
rect 1130 12822 1186 12878
rect 1186 12822 1190 12878
rect 1126 12818 1190 12822
rect 84886 12878 84950 12882
rect 84886 12822 84890 12878
rect 84890 12822 84946 12878
rect 84946 12822 84950 12878
rect 84886 12818 84950 12822
rect 84966 12878 85030 12882
rect 84966 12822 84970 12878
rect 84970 12822 85026 12878
rect 85026 12822 85030 12878
rect 84966 12818 85030 12822
rect 85046 12878 85110 12882
rect 85046 12822 85050 12878
rect 85050 12822 85106 12878
rect 85106 12822 85110 12878
rect 85046 12818 85110 12822
rect 85126 12878 85190 12882
rect 85126 12822 85130 12878
rect 85130 12822 85186 12878
rect 85186 12822 85190 12878
rect 85126 12818 85190 12822
rect 2886 12334 2950 12338
rect 2886 12278 2890 12334
rect 2890 12278 2946 12334
rect 2946 12278 2950 12334
rect 2886 12274 2950 12278
rect 2966 12334 3030 12338
rect 2966 12278 2970 12334
rect 2970 12278 3026 12334
rect 3026 12278 3030 12334
rect 2966 12274 3030 12278
rect 3046 12334 3110 12338
rect 3046 12278 3050 12334
rect 3050 12278 3106 12334
rect 3106 12278 3110 12334
rect 3046 12274 3110 12278
rect 3126 12334 3190 12338
rect 3126 12278 3130 12334
rect 3130 12278 3186 12334
rect 3186 12278 3190 12334
rect 3126 12274 3190 12278
rect 86886 12334 86950 12338
rect 86886 12278 86890 12334
rect 86890 12278 86946 12334
rect 86946 12278 86950 12334
rect 86886 12274 86950 12278
rect 86966 12334 87030 12338
rect 86966 12278 86970 12334
rect 86970 12278 87026 12334
rect 87026 12278 87030 12334
rect 86966 12274 87030 12278
rect 87046 12334 87110 12338
rect 87046 12278 87050 12334
rect 87050 12278 87106 12334
rect 87106 12278 87110 12334
rect 87046 12274 87110 12278
rect 87126 12334 87190 12338
rect 87126 12278 87130 12334
rect 87130 12278 87186 12334
rect 87186 12278 87190 12334
rect 87126 12274 87190 12278
rect 886 11790 950 11794
rect 886 11734 890 11790
rect 890 11734 946 11790
rect 946 11734 950 11790
rect 886 11730 950 11734
rect 966 11790 1030 11794
rect 966 11734 970 11790
rect 970 11734 1026 11790
rect 1026 11734 1030 11790
rect 966 11730 1030 11734
rect 1046 11790 1110 11794
rect 1046 11734 1050 11790
rect 1050 11734 1106 11790
rect 1106 11734 1110 11790
rect 1046 11730 1110 11734
rect 1126 11790 1190 11794
rect 1126 11734 1130 11790
rect 1130 11734 1186 11790
rect 1186 11734 1190 11790
rect 1126 11730 1190 11734
rect 84886 11790 84950 11794
rect 84886 11734 84890 11790
rect 84890 11734 84946 11790
rect 84946 11734 84950 11790
rect 84886 11730 84950 11734
rect 84966 11790 85030 11794
rect 84966 11734 84970 11790
rect 84970 11734 85026 11790
rect 85026 11734 85030 11790
rect 84966 11730 85030 11734
rect 85046 11790 85110 11794
rect 85046 11734 85050 11790
rect 85050 11734 85106 11790
rect 85106 11734 85110 11790
rect 85046 11730 85110 11734
rect 85126 11790 85190 11794
rect 85126 11734 85130 11790
rect 85130 11734 85186 11790
rect 85186 11734 85190 11790
rect 85126 11730 85190 11734
rect 2886 11246 2950 11250
rect 2886 11190 2890 11246
rect 2890 11190 2946 11246
rect 2946 11190 2950 11246
rect 2886 11186 2950 11190
rect 2966 11246 3030 11250
rect 2966 11190 2970 11246
rect 2970 11190 3026 11246
rect 3026 11190 3030 11246
rect 2966 11186 3030 11190
rect 3046 11246 3110 11250
rect 3046 11190 3050 11246
rect 3050 11190 3106 11246
rect 3106 11190 3110 11246
rect 3046 11186 3110 11190
rect 3126 11246 3190 11250
rect 3126 11190 3130 11246
rect 3130 11190 3186 11246
rect 3186 11190 3190 11246
rect 3126 11186 3190 11190
rect 86886 11246 86950 11250
rect 86886 11190 86890 11246
rect 86890 11190 86946 11246
rect 86946 11190 86950 11246
rect 86886 11186 86950 11190
rect 86966 11246 87030 11250
rect 86966 11190 86970 11246
rect 86970 11190 87026 11246
rect 87026 11190 87030 11246
rect 86966 11186 87030 11190
rect 87046 11246 87110 11250
rect 87046 11190 87050 11246
rect 87050 11190 87106 11246
rect 87106 11190 87110 11246
rect 87046 11186 87110 11190
rect 87126 11246 87190 11250
rect 87126 11190 87130 11246
rect 87130 11190 87186 11246
rect 87186 11190 87190 11246
rect 87126 11186 87190 11190
rect 886 10702 950 10706
rect 886 10646 890 10702
rect 890 10646 946 10702
rect 946 10646 950 10702
rect 886 10642 950 10646
rect 966 10702 1030 10706
rect 966 10646 970 10702
rect 970 10646 1026 10702
rect 1026 10646 1030 10702
rect 966 10642 1030 10646
rect 1046 10702 1110 10706
rect 1046 10646 1050 10702
rect 1050 10646 1106 10702
rect 1106 10646 1110 10702
rect 1046 10642 1110 10646
rect 1126 10702 1190 10706
rect 1126 10646 1130 10702
rect 1130 10646 1186 10702
rect 1186 10646 1190 10702
rect 1126 10642 1190 10646
rect 84886 10702 84950 10706
rect 84886 10646 84890 10702
rect 84890 10646 84946 10702
rect 84946 10646 84950 10702
rect 84886 10642 84950 10646
rect 84966 10702 85030 10706
rect 84966 10646 84970 10702
rect 84970 10646 85026 10702
rect 85026 10646 85030 10702
rect 84966 10642 85030 10646
rect 85046 10702 85110 10706
rect 85046 10646 85050 10702
rect 85050 10646 85106 10702
rect 85106 10646 85110 10702
rect 85046 10642 85110 10646
rect 85126 10702 85190 10706
rect 85126 10646 85130 10702
rect 85130 10646 85186 10702
rect 85186 10646 85190 10702
rect 85126 10642 85190 10646
rect 2886 10158 2950 10162
rect 2886 10102 2890 10158
rect 2890 10102 2946 10158
rect 2946 10102 2950 10158
rect 2886 10098 2950 10102
rect 2966 10158 3030 10162
rect 2966 10102 2970 10158
rect 2970 10102 3026 10158
rect 3026 10102 3030 10158
rect 2966 10098 3030 10102
rect 3046 10158 3110 10162
rect 3046 10102 3050 10158
rect 3050 10102 3106 10158
rect 3106 10102 3110 10158
rect 3046 10098 3110 10102
rect 3126 10158 3190 10162
rect 3126 10102 3130 10158
rect 3130 10102 3186 10158
rect 3186 10102 3190 10158
rect 3126 10098 3190 10102
rect 86886 10158 86950 10162
rect 86886 10102 86890 10158
rect 86890 10102 86946 10158
rect 86946 10102 86950 10158
rect 86886 10098 86950 10102
rect 86966 10158 87030 10162
rect 86966 10102 86970 10158
rect 86970 10102 87026 10158
rect 87026 10102 87030 10158
rect 86966 10098 87030 10102
rect 87046 10158 87110 10162
rect 87046 10102 87050 10158
rect 87050 10102 87106 10158
rect 87106 10102 87110 10158
rect 87046 10098 87110 10102
rect 87126 10158 87190 10162
rect 87126 10102 87130 10158
rect 87130 10102 87186 10158
rect 87186 10102 87190 10158
rect 87126 10098 87190 10102
rect 886 9614 950 9618
rect 886 9558 890 9614
rect 890 9558 946 9614
rect 946 9558 950 9614
rect 886 9554 950 9558
rect 966 9614 1030 9618
rect 966 9558 970 9614
rect 970 9558 1026 9614
rect 1026 9558 1030 9614
rect 966 9554 1030 9558
rect 1046 9614 1110 9618
rect 1046 9558 1050 9614
rect 1050 9558 1106 9614
rect 1106 9558 1110 9614
rect 1046 9554 1110 9558
rect 1126 9614 1190 9618
rect 1126 9558 1130 9614
rect 1130 9558 1186 9614
rect 1186 9558 1190 9614
rect 1126 9554 1190 9558
rect 84886 9614 84950 9618
rect 84886 9558 84890 9614
rect 84890 9558 84946 9614
rect 84946 9558 84950 9614
rect 84886 9554 84950 9558
rect 84966 9614 85030 9618
rect 84966 9558 84970 9614
rect 84970 9558 85026 9614
rect 85026 9558 85030 9614
rect 84966 9554 85030 9558
rect 85046 9614 85110 9618
rect 85046 9558 85050 9614
rect 85050 9558 85106 9614
rect 85106 9558 85110 9614
rect 85046 9554 85110 9558
rect 85126 9614 85190 9618
rect 85126 9558 85130 9614
rect 85130 9558 85186 9614
rect 85186 9558 85190 9614
rect 85126 9554 85190 9558
rect 2886 9070 2950 9074
rect 2886 9014 2890 9070
rect 2890 9014 2946 9070
rect 2946 9014 2950 9070
rect 2886 9010 2950 9014
rect 2966 9070 3030 9074
rect 2966 9014 2970 9070
rect 2970 9014 3026 9070
rect 3026 9014 3030 9070
rect 2966 9010 3030 9014
rect 3046 9070 3110 9074
rect 3046 9014 3050 9070
rect 3050 9014 3106 9070
rect 3106 9014 3110 9070
rect 3046 9010 3110 9014
rect 3126 9070 3190 9074
rect 3126 9014 3130 9070
rect 3130 9014 3186 9070
rect 3186 9014 3190 9070
rect 3126 9010 3190 9014
rect 86886 9070 86950 9074
rect 86886 9014 86890 9070
rect 86890 9014 86946 9070
rect 86946 9014 86950 9070
rect 86886 9010 86950 9014
rect 86966 9070 87030 9074
rect 86966 9014 86970 9070
rect 86970 9014 87026 9070
rect 87026 9014 87030 9070
rect 86966 9010 87030 9014
rect 87046 9070 87110 9074
rect 87046 9014 87050 9070
rect 87050 9014 87106 9070
rect 87106 9014 87110 9070
rect 87046 9010 87110 9014
rect 87126 9070 87190 9074
rect 87126 9014 87130 9070
rect 87130 9014 87186 9070
rect 87186 9014 87190 9070
rect 87126 9010 87190 9014
rect 886 8526 950 8530
rect 886 8470 890 8526
rect 890 8470 946 8526
rect 946 8470 950 8526
rect 886 8466 950 8470
rect 966 8526 1030 8530
rect 966 8470 970 8526
rect 970 8470 1026 8526
rect 1026 8470 1030 8526
rect 966 8466 1030 8470
rect 1046 8526 1110 8530
rect 1046 8470 1050 8526
rect 1050 8470 1106 8526
rect 1106 8470 1110 8526
rect 1046 8466 1110 8470
rect 1126 8526 1190 8530
rect 1126 8470 1130 8526
rect 1130 8470 1186 8526
rect 1186 8470 1190 8526
rect 1126 8466 1190 8470
rect 84886 8526 84950 8530
rect 84886 8470 84890 8526
rect 84890 8470 84946 8526
rect 84946 8470 84950 8526
rect 84886 8466 84950 8470
rect 84966 8526 85030 8530
rect 84966 8470 84970 8526
rect 84970 8470 85026 8526
rect 85026 8470 85030 8526
rect 84966 8466 85030 8470
rect 85046 8526 85110 8530
rect 85046 8470 85050 8526
rect 85050 8470 85106 8526
rect 85106 8470 85110 8526
rect 85046 8466 85110 8470
rect 85126 8526 85190 8530
rect 85126 8470 85130 8526
rect 85130 8470 85186 8526
rect 85186 8470 85190 8526
rect 85126 8466 85190 8470
rect 2886 7982 2950 7986
rect 2886 7926 2890 7982
rect 2890 7926 2946 7982
rect 2946 7926 2950 7982
rect 2886 7922 2950 7926
rect 2966 7982 3030 7986
rect 2966 7926 2970 7982
rect 2970 7926 3026 7982
rect 3026 7926 3030 7982
rect 2966 7922 3030 7926
rect 3046 7982 3110 7986
rect 3046 7926 3050 7982
rect 3050 7926 3106 7982
rect 3106 7926 3110 7982
rect 3046 7922 3110 7926
rect 3126 7982 3190 7986
rect 3126 7926 3130 7982
rect 3130 7926 3186 7982
rect 3186 7926 3190 7982
rect 3126 7922 3190 7926
rect 86886 7982 86950 7986
rect 86886 7926 86890 7982
rect 86890 7926 86946 7982
rect 86946 7926 86950 7982
rect 86886 7922 86950 7926
rect 86966 7982 87030 7986
rect 86966 7926 86970 7982
rect 86970 7926 87026 7982
rect 87026 7926 87030 7982
rect 86966 7922 87030 7926
rect 87046 7982 87110 7986
rect 87046 7926 87050 7982
rect 87050 7926 87106 7982
rect 87106 7926 87110 7982
rect 87046 7922 87110 7926
rect 87126 7982 87190 7986
rect 87126 7926 87130 7982
rect 87130 7926 87186 7982
rect 87186 7926 87190 7982
rect 87126 7922 87190 7926
rect 886 7438 950 7442
rect 886 7382 890 7438
rect 890 7382 946 7438
rect 946 7382 950 7438
rect 886 7378 950 7382
rect 966 7438 1030 7442
rect 966 7382 970 7438
rect 970 7382 1026 7438
rect 1026 7382 1030 7438
rect 966 7378 1030 7382
rect 1046 7438 1110 7442
rect 1046 7382 1050 7438
rect 1050 7382 1106 7438
rect 1106 7382 1110 7438
rect 1046 7378 1110 7382
rect 1126 7438 1190 7442
rect 1126 7382 1130 7438
rect 1130 7382 1186 7438
rect 1186 7382 1190 7438
rect 1126 7378 1190 7382
rect 84886 7438 84950 7442
rect 84886 7382 84890 7438
rect 84890 7382 84946 7438
rect 84946 7382 84950 7438
rect 84886 7378 84950 7382
rect 84966 7438 85030 7442
rect 84966 7382 84970 7438
rect 84970 7382 85026 7438
rect 85026 7382 85030 7438
rect 84966 7378 85030 7382
rect 85046 7438 85110 7442
rect 85046 7382 85050 7438
rect 85050 7382 85106 7438
rect 85106 7382 85110 7438
rect 85046 7378 85110 7382
rect 85126 7438 85190 7442
rect 85126 7382 85130 7438
rect 85130 7382 85186 7438
rect 85186 7382 85190 7438
rect 85126 7378 85190 7382
rect 2886 6894 2950 6898
rect 2886 6838 2890 6894
rect 2890 6838 2946 6894
rect 2946 6838 2950 6894
rect 2886 6834 2950 6838
rect 2966 6894 3030 6898
rect 2966 6838 2970 6894
rect 2970 6838 3026 6894
rect 3026 6838 3030 6894
rect 2966 6834 3030 6838
rect 3046 6894 3110 6898
rect 3046 6838 3050 6894
rect 3050 6838 3106 6894
rect 3106 6838 3110 6894
rect 3046 6834 3110 6838
rect 3126 6894 3190 6898
rect 3126 6838 3130 6894
rect 3130 6838 3186 6894
rect 3186 6838 3190 6894
rect 3126 6834 3190 6838
rect 86886 6894 86950 6898
rect 86886 6838 86890 6894
rect 86890 6838 86946 6894
rect 86946 6838 86950 6894
rect 86886 6834 86950 6838
rect 86966 6894 87030 6898
rect 86966 6838 86970 6894
rect 86970 6838 87026 6894
rect 87026 6838 87030 6894
rect 86966 6834 87030 6838
rect 87046 6894 87110 6898
rect 87046 6838 87050 6894
rect 87050 6838 87106 6894
rect 87106 6838 87110 6894
rect 87046 6834 87110 6838
rect 87126 6894 87190 6898
rect 87126 6838 87130 6894
rect 87130 6838 87186 6894
rect 87186 6838 87190 6894
rect 87126 6834 87190 6838
rect 886 6350 950 6354
rect 886 6294 890 6350
rect 890 6294 946 6350
rect 946 6294 950 6350
rect 886 6290 950 6294
rect 966 6350 1030 6354
rect 966 6294 970 6350
rect 970 6294 1026 6350
rect 1026 6294 1030 6350
rect 966 6290 1030 6294
rect 1046 6350 1110 6354
rect 1046 6294 1050 6350
rect 1050 6294 1106 6350
rect 1106 6294 1110 6350
rect 1046 6290 1110 6294
rect 1126 6350 1190 6354
rect 1126 6294 1130 6350
rect 1130 6294 1186 6350
rect 1186 6294 1190 6350
rect 1126 6290 1190 6294
rect 84886 6350 84950 6354
rect 84886 6294 84890 6350
rect 84890 6294 84946 6350
rect 84946 6294 84950 6350
rect 84886 6290 84950 6294
rect 84966 6350 85030 6354
rect 84966 6294 84970 6350
rect 84970 6294 85026 6350
rect 85026 6294 85030 6350
rect 84966 6290 85030 6294
rect 85046 6350 85110 6354
rect 85046 6294 85050 6350
rect 85050 6294 85106 6350
rect 85106 6294 85110 6350
rect 85046 6290 85110 6294
rect 85126 6350 85190 6354
rect 85126 6294 85130 6350
rect 85130 6294 85186 6350
rect 85186 6294 85190 6350
rect 85126 6290 85190 6294
rect 82346 6086 82410 6150
rect 2886 5806 2950 5810
rect 2886 5750 2890 5806
rect 2890 5750 2946 5806
rect 2946 5750 2950 5806
rect 2886 5746 2950 5750
rect 2966 5806 3030 5810
rect 2966 5750 2970 5806
rect 2970 5750 3026 5806
rect 3026 5750 3030 5806
rect 2966 5746 3030 5750
rect 3046 5806 3110 5810
rect 3046 5750 3050 5806
rect 3050 5750 3106 5806
rect 3106 5750 3110 5806
rect 3046 5746 3110 5750
rect 3126 5806 3190 5810
rect 3126 5750 3130 5806
rect 3130 5750 3186 5806
rect 3186 5750 3190 5806
rect 3126 5746 3190 5750
rect 86886 5806 86950 5810
rect 86886 5750 86890 5806
rect 86890 5750 86946 5806
rect 86946 5750 86950 5806
rect 86886 5746 86950 5750
rect 86966 5806 87030 5810
rect 86966 5750 86970 5806
rect 86970 5750 87026 5806
rect 87026 5750 87030 5806
rect 86966 5746 87030 5750
rect 87046 5806 87110 5810
rect 87046 5750 87050 5806
rect 87050 5750 87106 5806
rect 87106 5750 87110 5806
rect 87046 5746 87110 5750
rect 87126 5806 87190 5810
rect 87126 5750 87130 5806
rect 87130 5750 87186 5806
rect 87186 5750 87190 5806
rect 87126 5746 87190 5750
rect 886 5262 950 5266
rect 886 5206 890 5262
rect 890 5206 946 5262
rect 946 5206 950 5262
rect 886 5202 950 5206
rect 966 5262 1030 5266
rect 966 5206 970 5262
rect 970 5206 1026 5262
rect 1026 5206 1030 5262
rect 966 5202 1030 5206
rect 1046 5262 1110 5266
rect 1046 5206 1050 5262
rect 1050 5206 1106 5262
rect 1106 5206 1110 5262
rect 1046 5202 1110 5206
rect 1126 5262 1190 5266
rect 1126 5206 1130 5262
rect 1130 5206 1186 5262
rect 1186 5206 1190 5262
rect 1126 5202 1190 5206
rect 84886 5262 84950 5266
rect 84886 5206 84890 5262
rect 84890 5206 84946 5262
rect 84946 5206 84950 5262
rect 84886 5202 84950 5206
rect 84966 5262 85030 5266
rect 84966 5206 84970 5262
rect 84970 5206 85026 5262
rect 85026 5206 85030 5262
rect 84966 5202 85030 5206
rect 85046 5262 85110 5266
rect 85046 5206 85050 5262
rect 85050 5206 85106 5262
rect 85106 5206 85110 5262
rect 85046 5202 85110 5206
rect 85126 5262 85190 5266
rect 85126 5206 85130 5262
rect 85130 5206 85186 5262
rect 85186 5206 85190 5262
rect 85126 5202 85190 5206
rect 3594 5194 3658 5198
rect 3594 5138 3644 5194
rect 3644 5138 3658 5194
rect 3594 5134 3658 5138
rect 2886 4718 2950 4722
rect 2886 4662 2890 4718
rect 2890 4662 2946 4718
rect 2946 4662 2950 4718
rect 2886 4658 2950 4662
rect 2966 4718 3030 4722
rect 2966 4662 2970 4718
rect 2970 4662 3026 4718
rect 3026 4662 3030 4718
rect 2966 4658 3030 4662
rect 3046 4718 3110 4722
rect 3046 4662 3050 4718
rect 3050 4662 3106 4718
rect 3106 4662 3110 4718
rect 3046 4658 3110 4662
rect 3126 4718 3190 4722
rect 3126 4662 3130 4718
rect 3130 4662 3186 4718
rect 3186 4662 3190 4718
rect 3126 4658 3190 4662
rect 86886 4718 86950 4722
rect 86886 4662 86890 4718
rect 86890 4662 86946 4718
rect 86946 4662 86950 4718
rect 86886 4658 86950 4662
rect 86966 4718 87030 4722
rect 86966 4662 86970 4718
rect 86970 4662 87026 4718
rect 87026 4662 87030 4718
rect 86966 4658 87030 4662
rect 87046 4718 87110 4722
rect 87046 4662 87050 4718
rect 87050 4662 87106 4718
rect 87106 4662 87110 4718
rect 87046 4658 87110 4662
rect 87126 4718 87190 4722
rect 87126 4662 87130 4718
rect 87130 4662 87186 4718
rect 87186 4662 87190 4718
rect 87126 4658 87190 4662
rect 4146 4590 4210 4654
rect 4514 4590 4578 4654
rect 4146 4182 4210 4246
rect 886 4174 950 4178
rect 886 4118 890 4174
rect 890 4118 946 4174
rect 946 4118 950 4174
rect 886 4114 950 4118
rect 966 4174 1030 4178
rect 966 4118 970 4174
rect 970 4118 1026 4174
rect 1026 4118 1030 4174
rect 966 4114 1030 4118
rect 1046 4174 1110 4178
rect 1046 4118 1050 4174
rect 1050 4118 1106 4174
rect 1106 4118 1110 4174
rect 1046 4114 1110 4118
rect 1126 4174 1190 4178
rect 1126 4118 1130 4174
rect 1130 4118 1186 4174
rect 1186 4118 1190 4174
rect 1126 4114 1190 4118
rect 84886 4174 84950 4178
rect 84886 4118 84890 4174
rect 84890 4118 84946 4174
rect 84946 4118 84950 4174
rect 84886 4114 84950 4118
rect 84966 4174 85030 4178
rect 84966 4118 84970 4174
rect 84970 4118 85026 4174
rect 85026 4118 85030 4174
rect 84966 4114 85030 4118
rect 85046 4174 85110 4178
rect 85046 4118 85050 4174
rect 85050 4118 85106 4174
rect 85106 4118 85110 4174
rect 85046 4114 85110 4118
rect 85126 4174 85190 4178
rect 85126 4118 85130 4174
rect 85130 4118 85186 4174
rect 85186 4118 85190 4174
rect 85126 4114 85190 4118
rect 83818 4106 83882 4110
rect 83818 4050 83832 4106
rect 83832 4050 83882 4106
rect 83818 4046 83882 4050
rect 82898 3774 82962 3838
rect 2886 3630 2950 3634
rect 2886 3574 2890 3630
rect 2890 3574 2946 3630
rect 2946 3574 2950 3630
rect 2886 3570 2950 3574
rect 2966 3630 3030 3634
rect 2966 3574 2970 3630
rect 2970 3574 3026 3630
rect 3026 3574 3030 3630
rect 2966 3570 3030 3574
rect 3046 3630 3110 3634
rect 3046 3574 3050 3630
rect 3050 3574 3106 3630
rect 3106 3574 3110 3630
rect 3046 3570 3110 3574
rect 3126 3630 3190 3634
rect 3126 3574 3130 3630
rect 3130 3574 3186 3630
rect 3186 3574 3190 3630
rect 3126 3570 3190 3574
rect 86886 3630 86950 3634
rect 86886 3574 86890 3630
rect 86890 3574 86946 3630
rect 86946 3574 86950 3630
rect 86886 3570 86950 3574
rect 86966 3630 87030 3634
rect 86966 3574 86970 3630
rect 86970 3574 87026 3630
rect 87026 3574 87030 3630
rect 86966 3570 87030 3574
rect 87046 3630 87110 3634
rect 87046 3574 87050 3630
rect 87050 3574 87106 3630
rect 87106 3574 87110 3630
rect 87046 3570 87110 3574
rect 87126 3630 87190 3634
rect 87126 3574 87130 3630
rect 87130 3574 87186 3630
rect 87186 3574 87190 3630
rect 87126 3570 87190 3574
rect 3410 3502 3474 3566
rect 84554 3230 84618 3294
rect 3778 3094 3842 3158
rect 84370 3094 84434 3158
rect 886 3086 950 3090
rect 886 3030 890 3086
rect 890 3030 946 3086
rect 946 3030 950 3086
rect 886 3026 950 3030
rect 966 3086 1030 3090
rect 966 3030 970 3086
rect 970 3030 1026 3086
rect 1026 3030 1030 3086
rect 966 3026 1030 3030
rect 1046 3086 1110 3090
rect 1046 3030 1050 3086
rect 1050 3030 1106 3086
rect 1106 3030 1110 3086
rect 1046 3026 1110 3030
rect 1126 3086 1190 3090
rect 1126 3030 1130 3086
rect 1130 3030 1186 3086
rect 1186 3030 1190 3086
rect 1126 3026 1190 3030
rect 84886 3086 84950 3090
rect 84886 3030 84890 3086
rect 84890 3030 84946 3086
rect 84946 3030 84950 3086
rect 84886 3026 84950 3030
rect 84966 3086 85030 3090
rect 84966 3030 84970 3086
rect 84970 3030 85026 3086
rect 85026 3030 85030 3086
rect 84966 3026 85030 3030
rect 85046 3086 85110 3090
rect 85046 3030 85050 3086
rect 85050 3030 85106 3086
rect 85106 3030 85110 3086
rect 85046 3026 85110 3030
rect 85126 3086 85190 3090
rect 85126 3030 85130 3086
rect 85130 3030 85186 3086
rect 85186 3030 85190 3086
rect 85126 3026 85190 3030
rect 39106 2958 39170 3022
rect 42970 2958 43034 3022
rect 13530 2822 13594 2886
rect 19786 2882 19850 2886
rect 19786 2826 19800 2882
rect 19800 2826 19850 2882
rect 19786 2822 19850 2826
rect 21994 2822 22058 2886
rect 24018 2882 24082 2886
rect 24018 2826 24032 2882
rect 24032 2826 24082 2882
rect 24018 2822 24082 2826
rect 25122 2882 25186 2886
rect 25122 2826 25136 2882
rect 25136 2826 25186 2882
rect 25122 2822 25186 2826
rect 27514 2882 27578 2886
rect 27514 2826 27528 2882
rect 27528 2826 27578 2882
rect 27514 2822 27578 2826
rect 31056 2882 31120 2886
rect 31056 2826 31060 2882
rect 31060 2826 31116 2882
rect 31116 2826 31120 2882
rect 31056 2822 31120 2826
rect 33724 2882 33788 2886
rect 33724 2826 33728 2882
rect 33728 2826 33784 2882
rect 33784 2826 33788 2882
rect 33724 2822 33788 2826
rect 36898 2882 36962 2886
rect 36898 2826 36948 2882
rect 36948 2826 36962 2882
rect 36898 2822 36962 2826
rect 38922 2822 38986 2886
rect 41314 2882 41378 2886
rect 41314 2826 41364 2882
rect 41364 2826 41378 2882
rect 41314 2822 41378 2826
rect 44258 2822 44322 2886
rect 82530 2822 82594 2886
rect 37082 2686 37146 2750
rect 45362 2686 45426 2750
rect 48858 2550 48922 2614
rect 50146 2610 50210 2614
rect 50146 2554 50196 2610
rect 50196 2554 50210 2610
rect 50146 2550 50210 2554
rect 53642 2610 53706 2614
rect 53642 2554 53692 2610
rect 53692 2554 53706 2610
rect 53642 2550 53706 2554
rect 2886 2542 2950 2546
rect 2886 2486 2890 2542
rect 2890 2486 2946 2542
rect 2946 2486 2950 2542
rect 2886 2482 2950 2486
rect 2966 2542 3030 2546
rect 2966 2486 2970 2542
rect 2970 2486 3026 2542
rect 3026 2486 3030 2542
rect 2966 2482 3030 2486
rect 3046 2542 3110 2546
rect 3046 2486 3050 2542
rect 3050 2486 3106 2542
rect 3106 2486 3110 2542
rect 3046 2482 3110 2486
rect 3126 2542 3190 2546
rect 3126 2486 3130 2542
rect 3130 2486 3186 2542
rect 3186 2486 3190 2542
rect 3126 2482 3190 2486
rect 18314 2338 18378 2342
rect 18314 2282 18328 2338
rect 18328 2282 18378 2338
rect 18314 2278 18378 2282
rect 26410 2202 26474 2206
rect 26410 2146 26424 2202
rect 26424 2146 26474 2202
rect 26410 2142 26474 2146
rect 34874 2278 34938 2342
rect 54194 2338 54258 2342
rect 86886 2542 86950 2546
rect 86886 2486 86890 2542
rect 86890 2486 86946 2542
rect 86946 2486 86950 2542
rect 86886 2482 86950 2486
rect 86966 2542 87030 2546
rect 86966 2486 86970 2542
rect 86970 2486 87026 2542
rect 87026 2486 87030 2542
rect 86966 2482 87030 2486
rect 87046 2542 87110 2546
rect 87046 2486 87050 2542
rect 87050 2486 87106 2542
rect 87106 2486 87110 2542
rect 87046 2482 87110 2486
rect 87126 2542 87190 2546
rect 87126 2486 87130 2542
rect 87130 2486 87186 2542
rect 87186 2486 87190 2542
rect 87126 2482 87190 2486
rect 84002 2474 84066 2478
rect 84002 2418 84016 2474
rect 84016 2418 84066 2474
rect 84002 2414 84066 2418
rect 54194 2282 54244 2338
rect 54244 2282 54258 2338
rect 54194 2278 54258 2282
rect 82714 2278 82778 2342
rect 41866 2202 41930 2206
rect 41866 2146 41880 2202
rect 41880 2146 41930 2202
rect 41866 2142 41930 2146
rect 45178 2202 45242 2206
rect 45178 2146 45228 2202
rect 45228 2146 45242 2202
rect 45178 2142 45242 2146
rect 46650 2202 46714 2206
rect 46650 2146 46700 2202
rect 46700 2146 46714 2202
rect 46650 2142 46714 2146
rect 47570 2142 47634 2206
rect 49778 2202 49842 2206
rect 49778 2146 49828 2202
rect 49828 2146 49842 2202
rect 49778 2142 49842 2146
rect 84002 2142 84066 2206
rect 886 1998 950 2002
rect 886 1942 890 1998
rect 890 1942 946 1998
rect 946 1942 950 1998
rect 886 1938 950 1942
rect 966 1998 1030 2002
rect 966 1942 970 1998
rect 970 1942 1026 1998
rect 1026 1942 1030 1998
rect 966 1938 1030 1942
rect 1046 1998 1110 2002
rect 1046 1942 1050 1998
rect 1050 1942 1106 1998
rect 1106 1942 1110 1998
rect 1046 1938 1110 1942
rect 1126 1998 1190 2002
rect 1126 1942 1130 1998
rect 1130 1942 1186 1998
rect 1186 1942 1190 1998
rect 1126 1938 1190 1942
rect 84886 1998 84950 2002
rect 84886 1942 84890 1998
rect 84890 1942 84946 1998
rect 84946 1942 84950 1998
rect 84886 1938 84950 1942
rect 84966 1998 85030 2002
rect 84966 1942 84970 1998
rect 84970 1942 85026 1998
rect 85026 1942 85030 1998
rect 84966 1938 85030 1942
rect 85046 1998 85110 2002
rect 85046 1942 85050 1998
rect 85050 1942 85106 1998
rect 85106 1942 85110 1998
rect 85046 1938 85110 1942
rect 85126 1998 85190 2002
rect 85126 1942 85130 1998
rect 85130 1942 85186 1998
rect 85186 1942 85190 1998
rect 85126 1938 85190 1942
rect 8735 1658 8799 1662
rect 8735 1602 8760 1658
rect 8760 1602 8799 1658
rect 8735 1598 8799 1602
rect 22370 1658 22434 1662
rect 22370 1602 22412 1658
rect 22412 1602 22434 1658
rect 22370 1598 22434 1602
rect 24706 1658 24770 1662
rect 24706 1602 24712 1658
rect 24712 1602 24768 1658
rect 24768 1602 24770 1658
rect 24706 1598 24770 1602
rect 29254 1658 29318 1662
rect 29254 1602 29276 1658
rect 29276 1602 29318 1658
rect 29254 1598 29318 1602
rect 36262 1658 36326 1662
rect 36262 1602 36304 1658
rect 36304 1602 36326 1658
rect 36262 1598 36326 1602
rect 84186 1598 84250 1662
rect 42234 1386 42298 1390
rect 42234 1330 42284 1386
rect 42284 1330 42298 1386
rect 42234 1326 42298 1330
rect 51434 1386 51498 1390
rect 51434 1330 51484 1386
rect 51484 1330 51498 1386
rect 51434 1326 51498 1330
rect 84738 1326 84802 1390
rect 27146 1054 27210 1118
rect 83634 1054 83698 1118
rect 11690 978 11754 982
rect 11690 922 11704 978
rect 11704 922 11754 978
rect 11690 918 11754 922
rect 12242 918 12306 982
rect 15186 918 15250 982
rect 17578 918 17642 982
rect 17762 918 17826 982
rect 18866 978 18930 982
rect 18866 922 18916 978
rect 18916 922 18930 978
rect 18866 918 18930 922
rect 21074 918 21138 982
rect 21258 978 21322 982
rect 21258 922 21308 978
rect 21308 922 21322 978
rect 21258 918 21322 922
rect 23466 978 23530 982
rect 23466 922 23480 978
rect 23480 922 23530 978
rect 23466 918 23530 922
rect 24202 978 24266 982
rect 24202 922 24252 978
rect 24252 922 24266 978
rect 24202 918 24266 922
rect 28250 978 28314 982
rect 28250 922 28300 978
rect 28300 922 28314 978
rect 28250 918 28314 922
rect 29354 978 29418 982
rect 29354 922 29404 978
rect 29404 922 29418 978
rect 29354 918 29418 922
rect 31010 978 31074 982
rect 31010 922 31060 978
rect 31060 922 31074 978
rect 31010 918 31074 922
rect 31746 918 31810 982
rect 32850 978 32914 982
rect 32850 922 32900 978
rect 32900 922 32914 978
rect 32850 918 32914 922
rect 34690 978 34754 982
rect 34690 922 34740 978
rect 34740 922 34754 978
rect 34690 918 34754 922
rect 35242 978 35306 982
rect 35242 922 35292 978
rect 35292 922 35306 978
rect 35242 918 35306 922
rect 38186 918 38250 982
rect 40026 978 40090 982
rect 40026 922 40076 978
rect 40076 922 40090 978
rect 40026 918 40090 922
rect 43890 978 43954 982
rect 43890 922 43940 978
rect 43940 922 43954 978
rect 43890 918 43954 922
rect 45730 918 45794 982
rect 47938 918 48002 982
rect 4514 782 4578 846
rect 40946 782 41010 846
rect 48122 782 48186 846
rect 4146 646 4210 710
rect 15738 646 15802 710
rect 20706 706 20770 710
rect 20706 650 20756 706
rect 20756 650 20770 706
rect 20706 646 20770 650
rect 29906 706 29970 710
rect 29906 650 29920 706
rect 29920 650 29970 706
rect 29906 646 29970 650
rect 51618 646 51682 710
rect 83266 646 83330 710
rect 32482 570 32546 574
rect 32482 514 32496 570
rect 32496 514 32546 570
rect 32482 510 32546 514
rect 52722 510 52786 574
rect 38554 374 38618 438
rect 52906 374 52970 438
rect 83450 374 83514 438
rect 50330 238 50394 302
rect 25858 102 25922 166
<< metal4 >>
rect 5249 187982 5315 187983
rect 5249 187918 5250 187982
rect 5314 187918 5315 187982
rect 5249 187917 5315 187918
rect 878 186962 1198 187522
rect 878 186898 886 186962
rect 950 186898 966 186962
rect 1030 186898 1046 186962
rect 1110 186898 1126 186962
rect 1190 186898 1198 186962
rect 878 185874 1198 186898
rect 878 185810 886 185874
rect 950 185810 966 185874
rect 1030 185810 1046 185874
rect 1110 185810 1126 185874
rect 1190 185810 1198 185874
rect 878 185370 1198 185810
rect 878 185134 920 185370
rect 1156 185134 1198 185370
rect 878 184786 1198 185134
rect 878 184722 886 184786
rect 950 184722 966 184786
rect 1030 184722 1046 184786
rect 1110 184722 1126 184786
rect 1190 184722 1198 184786
rect 878 183698 1198 184722
rect 878 183634 886 183698
rect 950 183634 966 183698
rect 1030 183634 1046 183698
rect 1110 183634 1126 183698
rect 1190 183634 1198 183698
rect 878 182610 1198 183634
rect 878 182546 886 182610
rect 950 182546 966 182610
rect 1030 182546 1046 182610
rect 1110 182546 1126 182610
rect 1190 182546 1198 182610
rect 878 181522 1198 182546
rect 878 181458 886 181522
rect 950 181458 966 181522
rect 1030 181458 1046 181522
rect 1110 181458 1126 181522
rect 1190 181458 1198 181522
rect 878 180434 1198 181458
rect 878 180370 886 180434
rect 950 180370 966 180434
rect 1030 180370 1046 180434
rect 1110 180370 1126 180434
rect 1190 180370 1198 180434
rect 878 179346 1198 180370
rect 878 179282 886 179346
rect 950 179282 966 179346
rect 1030 179282 1046 179346
rect 1110 179282 1126 179346
rect 1190 179282 1198 179346
rect 878 178258 1198 179282
rect 878 178194 886 178258
rect 950 178194 966 178258
rect 1030 178194 1046 178258
rect 1110 178194 1126 178258
rect 1190 178194 1198 178258
rect 878 177170 1198 178194
rect 878 177106 886 177170
rect 950 177106 966 177170
rect 1030 177106 1046 177170
rect 1110 177106 1126 177170
rect 1190 177106 1198 177170
rect 878 176082 1198 177106
rect 878 176018 886 176082
rect 950 176018 966 176082
rect 1030 176018 1046 176082
rect 1110 176018 1126 176082
rect 1190 176018 1198 176082
rect 878 175370 1198 176018
rect 878 175134 920 175370
rect 1156 175134 1198 175370
rect 878 174994 1198 175134
rect 878 174930 886 174994
rect 950 174930 966 174994
rect 1030 174930 1046 174994
rect 1110 174930 1126 174994
rect 1190 174930 1198 174994
rect 878 173906 1198 174930
rect 878 173842 886 173906
rect 950 173842 966 173906
rect 1030 173842 1046 173906
rect 1110 173842 1126 173906
rect 1190 173842 1198 173906
rect 878 172818 1198 173842
rect 878 172754 886 172818
rect 950 172754 966 172818
rect 1030 172754 1046 172818
rect 1110 172754 1126 172818
rect 1190 172754 1198 172818
rect 878 171730 1198 172754
rect 878 171666 886 171730
rect 950 171666 966 171730
rect 1030 171666 1046 171730
rect 1110 171666 1126 171730
rect 1190 171666 1198 171730
rect 878 170642 1198 171666
rect 878 170578 886 170642
rect 950 170578 966 170642
rect 1030 170578 1046 170642
rect 1110 170578 1126 170642
rect 1190 170578 1198 170642
rect 878 169554 1198 170578
rect 878 169490 886 169554
rect 950 169490 966 169554
rect 1030 169490 1046 169554
rect 1110 169490 1126 169554
rect 1190 169490 1198 169554
rect 878 168466 1198 169490
rect 878 168402 886 168466
rect 950 168402 966 168466
rect 1030 168402 1046 168466
rect 1110 168402 1126 168466
rect 1190 168402 1198 168466
rect 878 167378 1198 168402
rect 878 167314 886 167378
rect 950 167314 966 167378
rect 1030 167314 1046 167378
rect 1110 167314 1126 167378
rect 1190 167314 1198 167378
rect 878 166290 1198 167314
rect 878 166226 886 166290
rect 950 166226 966 166290
rect 1030 166226 1046 166290
rect 1110 166226 1126 166290
rect 1190 166226 1198 166290
rect 878 165370 1198 166226
rect 878 165202 920 165370
rect 1156 165202 1198 165370
rect 878 165138 886 165202
rect 1190 165138 1198 165202
rect 878 165134 920 165138
rect 1156 165134 1198 165138
rect 878 164114 1198 165134
rect 878 164050 886 164114
rect 950 164050 966 164114
rect 1030 164050 1046 164114
rect 1110 164050 1126 164114
rect 1190 164050 1198 164114
rect 878 163026 1198 164050
rect 878 162962 886 163026
rect 950 162962 966 163026
rect 1030 162962 1046 163026
rect 1110 162962 1126 163026
rect 1190 162962 1198 163026
rect 878 161938 1198 162962
rect 878 161874 886 161938
rect 950 161874 966 161938
rect 1030 161874 1046 161938
rect 1110 161874 1126 161938
rect 1190 161874 1198 161938
rect 878 160850 1198 161874
rect 878 160786 886 160850
rect 950 160786 966 160850
rect 1030 160786 1046 160850
rect 1110 160786 1126 160850
rect 1190 160786 1198 160850
rect 878 159762 1198 160786
rect 878 159698 886 159762
rect 950 159698 966 159762
rect 1030 159698 1046 159762
rect 1110 159698 1126 159762
rect 1190 159698 1198 159762
rect 878 158674 1198 159698
rect 878 158610 886 158674
rect 950 158610 966 158674
rect 1030 158610 1046 158674
rect 1110 158610 1126 158674
rect 1190 158610 1198 158674
rect 878 157586 1198 158610
rect 878 157522 886 157586
rect 950 157522 966 157586
rect 1030 157522 1046 157586
rect 1110 157522 1126 157586
rect 1190 157522 1198 157586
rect 878 156498 1198 157522
rect 878 156434 886 156498
rect 950 156434 966 156498
rect 1030 156434 1046 156498
rect 1110 156434 1126 156498
rect 1190 156434 1198 156498
rect 878 155410 1198 156434
rect 878 155346 886 155410
rect 950 155370 966 155410
rect 1030 155370 1046 155410
rect 1110 155370 1126 155410
rect 1190 155346 1198 155410
rect 878 155134 920 155346
rect 1156 155134 1198 155346
rect 878 154322 1198 155134
rect 878 154258 886 154322
rect 950 154258 966 154322
rect 1030 154258 1046 154322
rect 1110 154258 1126 154322
rect 1190 154258 1198 154322
rect 878 153234 1198 154258
rect 878 153170 886 153234
rect 950 153170 966 153234
rect 1030 153170 1046 153234
rect 1110 153170 1126 153234
rect 1190 153170 1198 153234
rect 878 152146 1198 153170
rect 878 152082 886 152146
rect 950 152082 966 152146
rect 1030 152082 1046 152146
rect 1110 152082 1126 152146
rect 1190 152082 1198 152146
rect 878 151058 1198 152082
rect 878 150994 886 151058
rect 950 150994 966 151058
rect 1030 150994 1046 151058
rect 1110 150994 1126 151058
rect 1190 150994 1198 151058
rect 878 149970 1198 150994
rect 878 149906 886 149970
rect 950 149906 966 149970
rect 1030 149906 1046 149970
rect 1110 149906 1126 149970
rect 1190 149906 1198 149970
rect 878 148882 1198 149906
rect 878 148818 886 148882
rect 950 148818 966 148882
rect 1030 148818 1046 148882
rect 1110 148818 1126 148882
rect 1190 148818 1198 148882
rect 878 147794 1198 148818
rect 878 147730 886 147794
rect 950 147730 966 147794
rect 1030 147730 1046 147794
rect 1110 147730 1126 147794
rect 1190 147730 1198 147794
rect 878 146706 1198 147730
rect 878 146642 886 146706
rect 950 146642 966 146706
rect 1030 146642 1046 146706
rect 1110 146642 1126 146706
rect 1190 146642 1198 146706
rect 878 145618 1198 146642
rect 878 145554 886 145618
rect 950 145554 966 145618
rect 1030 145554 1046 145618
rect 1110 145554 1126 145618
rect 1190 145554 1198 145618
rect 878 145370 1198 145554
rect 878 145134 920 145370
rect 1156 145134 1198 145370
rect 878 144530 1198 145134
rect 878 144466 886 144530
rect 950 144466 966 144530
rect 1030 144466 1046 144530
rect 1110 144466 1126 144530
rect 1190 144466 1198 144530
rect 878 143442 1198 144466
rect 878 143378 886 143442
rect 950 143378 966 143442
rect 1030 143378 1046 143442
rect 1110 143378 1126 143442
rect 1190 143378 1198 143442
rect 878 142354 1198 143378
rect 878 142290 886 142354
rect 950 142290 966 142354
rect 1030 142290 1046 142354
rect 1110 142290 1126 142354
rect 1190 142290 1198 142354
rect 878 141266 1198 142290
rect 878 141202 886 141266
rect 950 141202 966 141266
rect 1030 141202 1046 141266
rect 1110 141202 1126 141266
rect 1190 141202 1198 141266
rect 878 140178 1198 141202
rect 878 140114 886 140178
rect 950 140114 966 140178
rect 1030 140114 1046 140178
rect 1110 140114 1126 140178
rect 1190 140114 1198 140178
rect 878 139090 1198 140114
rect 878 139026 886 139090
rect 950 139026 966 139090
rect 1030 139026 1046 139090
rect 1110 139026 1126 139090
rect 1190 139026 1198 139090
rect 878 138002 1198 139026
rect 878 137938 886 138002
rect 950 137938 966 138002
rect 1030 137938 1046 138002
rect 1110 137938 1126 138002
rect 1190 137938 1198 138002
rect 878 136914 1198 137938
rect 878 136850 886 136914
rect 950 136850 966 136914
rect 1030 136850 1046 136914
rect 1110 136850 1126 136914
rect 1190 136850 1198 136914
rect 878 135826 1198 136850
rect 878 135762 886 135826
rect 950 135762 966 135826
rect 1030 135762 1046 135826
rect 1110 135762 1126 135826
rect 1190 135762 1198 135826
rect 878 135370 1198 135762
rect 878 135134 920 135370
rect 1156 135134 1198 135370
rect 878 134738 1198 135134
rect 878 134674 886 134738
rect 950 134674 966 134738
rect 1030 134674 1046 134738
rect 1110 134674 1126 134738
rect 1190 134674 1198 134738
rect 878 133650 1198 134674
rect 878 133586 886 133650
rect 950 133586 966 133650
rect 1030 133586 1046 133650
rect 1110 133586 1126 133650
rect 1190 133586 1198 133650
rect 878 132562 1198 133586
rect 878 132498 886 132562
rect 950 132498 966 132562
rect 1030 132498 1046 132562
rect 1110 132498 1126 132562
rect 1190 132498 1198 132562
rect 878 131474 1198 132498
rect 878 131410 886 131474
rect 950 131410 966 131474
rect 1030 131410 1046 131474
rect 1110 131410 1126 131474
rect 1190 131410 1198 131474
rect 878 130386 1198 131410
rect 878 130322 886 130386
rect 950 130322 966 130386
rect 1030 130322 1046 130386
rect 1110 130322 1126 130386
rect 1190 130322 1198 130386
rect 878 129298 1198 130322
rect 878 129234 886 129298
rect 950 129234 966 129298
rect 1030 129234 1046 129298
rect 1110 129234 1126 129298
rect 1190 129234 1198 129298
rect 878 128210 1198 129234
rect 878 128146 886 128210
rect 950 128146 966 128210
rect 1030 128146 1046 128210
rect 1110 128146 1126 128210
rect 1190 128146 1198 128210
rect 878 127122 1198 128146
rect 878 127058 886 127122
rect 950 127058 966 127122
rect 1030 127058 1046 127122
rect 1110 127058 1126 127122
rect 1190 127058 1198 127122
rect 878 126034 1198 127058
rect 878 125970 886 126034
rect 950 125970 966 126034
rect 1030 125970 1046 126034
rect 1110 125970 1126 126034
rect 1190 125970 1198 126034
rect 878 125370 1198 125970
rect 878 125134 920 125370
rect 1156 125134 1198 125370
rect 878 124946 1198 125134
rect 878 124882 886 124946
rect 950 124882 966 124946
rect 1030 124882 1046 124946
rect 1110 124882 1126 124946
rect 1190 124882 1198 124946
rect 878 123858 1198 124882
rect 2878 187506 3198 187522
rect 2878 187442 2886 187506
rect 2950 187442 2966 187506
rect 3030 187442 3046 187506
rect 3110 187442 3126 187506
rect 3190 187442 3198 187506
rect 2878 186418 3198 187442
rect 4145 187438 4211 187439
rect 4145 187374 4146 187438
rect 4210 187374 4211 187438
rect 4145 187373 4211 187374
rect 3593 187166 3659 187167
rect 3593 187102 3594 187166
rect 3658 187102 3659 187166
rect 3593 187101 3659 187102
rect 2878 186354 2886 186418
rect 2950 186354 2966 186418
rect 3030 186354 3046 186418
rect 3110 186354 3126 186418
rect 3190 186354 3198 186418
rect 2878 185330 3198 186354
rect 2878 185266 2886 185330
rect 2950 185266 2966 185330
rect 3030 185266 3046 185330
rect 3110 185266 3126 185330
rect 3190 185266 3198 185330
rect 2878 184242 3198 185266
rect 2878 184178 2886 184242
rect 2950 184178 2966 184242
rect 3030 184178 3046 184242
rect 3110 184178 3126 184242
rect 3190 184178 3198 184242
rect 2878 183154 3198 184178
rect 2878 183090 2886 183154
rect 2950 183090 2966 183154
rect 3030 183090 3046 183154
rect 3110 183090 3126 183154
rect 3190 183090 3198 183154
rect 2878 182066 3198 183090
rect 2878 182002 2886 182066
rect 2950 182002 2966 182066
rect 3030 182002 3046 182066
rect 3110 182002 3126 182066
rect 3190 182002 3198 182066
rect 2878 180978 3198 182002
rect 2878 180914 2886 180978
rect 2950 180914 2966 180978
rect 3030 180914 3046 180978
rect 3110 180914 3126 180978
rect 3190 180914 3198 180978
rect 2878 180370 3198 180914
rect 2878 180134 2920 180370
rect 3156 180134 3198 180370
rect 2878 179890 3198 180134
rect 2878 179826 2886 179890
rect 2950 179826 2966 179890
rect 3030 179826 3046 179890
rect 3110 179826 3126 179890
rect 3190 179826 3198 179890
rect 2878 178802 3198 179826
rect 2878 178738 2886 178802
rect 2950 178738 2966 178802
rect 3030 178738 3046 178802
rect 3110 178738 3126 178802
rect 3190 178738 3198 178802
rect 2878 177714 3198 178738
rect 2878 177650 2886 177714
rect 2950 177650 2966 177714
rect 3030 177650 3046 177714
rect 3110 177650 3126 177714
rect 3190 177650 3198 177714
rect 2878 176626 3198 177650
rect 2878 176562 2886 176626
rect 2950 176562 2966 176626
rect 3030 176562 3046 176626
rect 3110 176562 3126 176626
rect 3190 176562 3198 176626
rect 2878 175538 3198 176562
rect 2878 175474 2886 175538
rect 2950 175474 2966 175538
rect 3030 175474 3046 175538
rect 3110 175474 3126 175538
rect 3190 175474 3198 175538
rect 2878 174450 3198 175474
rect 2878 174386 2886 174450
rect 2950 174386 2966 174450
rect 3030 174386 3046 174450
rect 3110 174386 3126 174450
rect 3190 174386 3198 174450
rect 2878 173362 3198 174386
rect 2878 173298 2886 173362
rect 2950 173298 2966 173362
rect 3030 173298 3046 173362
rect 3110 173298 3126 173362
rect 3190 173298 3198 173362
rect 2878 172274 3198 173298
rect 2878 172210 2886 172274
rect 2950 172210 2966 172274
rect 3030 172210 3046 172274
rect 3110 172210 3126 172274
rect 3190 172210 3198 172274
rect 2878 171186 3198 172210
rect 2878 171122 2886 171186
rect 2950 171122 2966 171186
rect 3030 171122 3046 171186
rect 3110 171122 3126 171186
rect 3190 171122 3198 171186
rect 2878 170370 3198 171122
rect 2878 170134 2920 170370
rect 3156 170134 3198 170370
rect 2878 170098 3198 170134
rect 2878 170034 2886 170098
rect 2950 170034 2966 170098
rect 3030 170034 3046 170098
rect 3110 170034 3126 170098
rect 3190 170034 3198 170098
rect 2878 169010 3198 170034
rect 2878 168946 2886 169010
rect 2950 168946 2966 169010
rect 3030 168946 3046 169010
rect 3110 168946 3126 169010
rect 3190 168946 3198 169010
rect 2878 167922 3198 168946
rect 2878 167858 2886 167922
rect 2950 167858 2966 167922
rect 3030 167858 3046 167922
rect 3110 167858 3126 167922
rect 3190 167858 3198 167922
rect 2878 166834 3198 167858
rect 2878 166770 2886 166834
rect 2950 166770 2966 166834
rect 3030 166770 3046 166834
rect 3110 166770 3126 166834
rect 3190 166770 3198 166834
rect 2878 165746 3198 166770
rect 2878 165682 2886 165746
rect 2950 165682 2966 165746
rect 3030 165682 3046 165746
rect 3110 165682 3126 165746
rect 3190 165682 3198 165746
rect 2878 164658 3198 165682
rect 2878 164594 2886 164658
rect 2950 164594 2966 164658
rect 3030 164594 3046 164658
rect 3110 164594 3126 164658
rect 3190 164594 3198 164658
rect 2878 163570 3198 164594
rect 2878 163506 2886 163570
rect 2950 163506 2966 163570
rect 3030 163506 3046 163570
rect 3110 163506 3126 163570
rect 3190 163506 3198 163570
rect 2878 162482 3198 163506
rect 2878 162418 2886 162482
rect 2950 162418 2966 162482
rect 3030 162418 3046 162482
rect 3110 162418 3126 162482
rect 3190 162418 3198 162482
rect 2878 161394 3198 162418
rect 2878 161330 2886 161394
rect 2950 161330 2966 161394
rect 3030 161330 3046 161394
rect 3110 161330 3126 161394
rect 3190 161330 3198 161394
rect 2878 160370 3198 161330
rect 2878 160306 2920 160370
rect 3156 160306 3198 160370
rect 2878 160242 2886 160306
rect 3190 160242 3198 160306
rect 2878 160134 2920 160242
rect 3156 160134 3198 160242
rect 2878 159218 3198 160134
rect 2878 159154 2886 159218
rect 2950 159154 2966 159218
rect 3030 159154 3046 159218
rect 3110 159154 3126 159218
rect 3190 159154 3198 159218
rect 2878 158130 3198 159154
rect 2878 158066 2886 158130
rect 2950 158066 2966 158130
rect 3030 158066 3046 158130
rect 3110 158066 3126 158130
rect 3190 158066 3198 158130
rect 2878 157042 3198 158066
rect 2878 156978 2886 157042
rect 2950 156978 2966 157042
rect 3030 156978 3046 157042
rect 3110 156978 3126 157042
rect 3190 156978 3198 157042
rect 2878 155954 3198 156978
rect 2878 155890 2886 155954
rect 2950 155890 2966 155954
rect 3030 155890 3046 155954
rect 3110 155890 3126 155954
rect 3190 155890 3198 155954
rect 2878 154866 3198 155890
rect 2878 154802 2886 154866
rect 2950 154802 2966 154866
rect 3030 154802 3046 154866
rect 3110 154802 3126 154866
rect 3190 154802 3198 154866
rect 2878 153778 3198 154802
rect 2878 153714 2886 153778
rect 2950 153714 2966 153778
rect 3030 153714 3046 153778
rect 3110 153714 3126 153778
rect 3190 153714 3198 153778
rect 2878 152690 3198 153714
rect 2878 152626 2886 152690
rect 2950 152626 2966 152690
rect 3030 152626 3046 152690
rect 3110 152626 3126 152690
rect 3190 152626 3198 152690
rect 2878 151602 3198 152626
rect 2878 151538 2886 151602
rect 2950 151538 2966 151602
rect 3030 151538 3046 151602
rect 3110 151538 3126 151602
rect 3190 151538 3198 151602
rect 2878 150514 3198 151538
rect 2878 150450 2886 150514
rect 2950 150450 2966 150514
rect 3030 150450 3046 150514
rect 3110 150450 3126 150514
rect 3190 150450 3198 150514
rect 2878 150370 3198 150450
rect 2878 150134 2920 150370
rect 3156 150134 3198 150370
rect 2878 149426 3198 150134
rect 2878 149362 2886 149426
rect 2950 149362 2966 149426
rect 3030 149362 3046 149426
rect 3110 149362 3126 149426
rect 3190 149362 3198 149426
rect 2878 148338 3198 149362
rect 2878 148274 2886 148338
rect 2950 148274 2966 148338
rect 3030 148274 3046 148338
rect 3110 148274 3126 148338
rect 3190 148274 3198 148338
rect 2878 147250 3198 148274
rect 2878 147186 2886 147250
rect 2950 147186 2966 147250
rect 3030 147186 3046 147250
rect 3110 147186 3126 147250
rect 3190 147186 3198 147250
rect 2878 146162 3198 147186
rect 2878 146098 2886 146162
rect 2950 146098 2966 146162
rect 3030 146098 3046 146162
rect 3110 146098 3126 146162
rect 3190 146098 3198 146162
rect 2878 145074 3198 146098
rect 2878 145010 2886 145074
rect 2950 145010 2966 145074
rect 3030 145010 3046 145074
rect 3110 145010 3126 145074
rect 3190 145010 3198 145074
rect 2878 143986 3198 145010
rect 2878 143922 2886 143986
rect 2950 143922 2966 143986
rect 3030 143922 3046 143986
rect 3110 143922 3126 143986
rect 3190 143922 3198 143986
rect 2878 142898 3198 143922
rect 2878 142834 2886 142898
rect 2950 142834 2966 142898
rect 3030 142834 3046 142898
rect 3110 142834 3126 142898
rect 3190 142834 3198 142898
rect 2878 141810 3198 142834
rect 2878 141746 2886 141810
rect 2950 141746 2966 141810
rect 3030 141746 3046 141810
rect 3110 141746 3126 141810
rect 3190 141746 3198 141810
rect 2878 140722 3198 141746
rect 2878 140658 2886 140722
rect 2950 140658 2966 140722
rect 3030 140658 3046 140722
rect 3110 140658 3126 140722
rect 3190 140658 3198 140722
rect 2878 140370 3198 140658
rect 2878 140134 2920 140370
rect 3156 140134 3198 140370
rect 2878 139634 3198 140134
rect 2878 139570 2886 139634
rect 2950 139570 2966 139634
rect 3030 139570 3046 139634
rect 3110 139570 3126 139634
rect 3190 139570 3198 139634
rect 2878 138546 3198 139570
rect 2878 138482 2886 138546
rect 2950 138482 2966 138546
rect 3030 138482 3046 138546
rect 3110 138482 3126 138546
rect 3190 138482 3198 138546
rect 2878 137458 3198 138482
rect 2878 137394 2886 137458
rect 2950 137394 2966 137458
rect 3030 137394 3046 137458
rect 3110 137394 3126 137458
rect 3190 137394 3198 137458
rect 2878 136370 3198 137394
rect 2878 136306 2886 136370
rect 2950 136306 2966 136370
rect 3030 136306 3046 136370
rect 3110 136306 3126 136370
rect 3190 136306 3198 136370
rect 2878 135282 3198 136306
rect 2878 135218 2886 135282
rect 2950 135218 2966 135282
rect 3030 135218 3046 135282
rect 3110 135218 3126 135282
rect 3190 135218 3198 135282
rect 2878 134194 3198 135218
rect 2878 134130 2886 134194
rect 2950 134130 2966 134194
rect 3030 134130 3046 134194
rect 3110 134130 3126 134194
rect 3190 134130 3198 134194
rect 2878 133106 3198 134130
rect 2878 133042 2886 133106
rect 2950 133042 2966 133106
rect 3030 133042 3046 133106
rect 3110 133042 3126 133106
rect 3190 133042 3198 133106
rect 2878 132018 3198 133042
rect 2878 131954 2886 132018
rect 2950 131954 2966 132018
rect 3030 131954 3046 132018
rect 3110 131954 3126 132018
rect 3190 131954 3198 132018
rect 2878 130930 3198 131954
rect 2878 130866 2886 130930
rect 2950 130866 2966 130930
rect 3030 130866 3046 130930
rect 3110 130866 3126 130930
rect 3190 130866 3198 130930
rect 2878 130370 3198 130866
rect 2878 130134 2920 130370
rect 3156 130134 3198 130370
rect 2878 129842 3198 130134
rect 2878 129778 2886 129842
rect 2950 129778 2966 129842
rect 3030 129778 3046 129842
rect 3110 129778 3126 129842
rect 3190 129778 3198 129842
rect 2878 128754 3198 129778
rect 2878 128690 2886 128754
rect 2950 128690 2966 128754
rect 3030 128690 3046 128754
rect 3110 128690 3126 128754
rect 3190 128690 3198 128754
rect 2878 127666 3198 128690
rect 2878 127602 2886 127666
rect 2950 127602 2966 127666
rect 3030 127602 3046 127666
rect 3110 127602 3126 127666
rect 3190 127602 3198 127666
rect 2878 126578 3198 127602
rect 2878 126514 2886 126578
rect 2950 126514 2966 126578
rect 3030 126514 3046 126578
rect 3110 126514 3126 126578
rect 3190 126514 3198 126578
rect 2878 125490 3198 126514
rect 2878 125426 2886 125490
rect 2950 125426 2966 125490
rect 3030 125426 3046 125490
rect 3110 125426 3126 125490
rect 3190 125426 3198 125490
rect 2305 124742 2371 124743
rect 2305 124678 2306 124742
rect 2370 124678 2371 124742
rect 2305 124677 2371 124678
rect 878 123794 886 123858
rect 950 123794 966 123858
rect 1030 123794 1046 123858
rect 1110 123794 1126 123858
rect 1190 123794 1198 123858
rect 878 122770 1198 123794
rect 878 122706 886 122770
rect 950 122706 966 122770
rect 1030 122706 1046 122770
rect 1110 122706 1126 122770
rect 1190 122706 1198 122770
rect 878 121682 1198 122706
rect 878 121618 886 121682
rect 950 121618 966 121682
rect 1030 121618 1046 121682
rect 1110 121618 1126 121682
rect 1190 121618 1198 121682
rect 878 120594 1198 121618
rect 878 120530 886 120594
rect 950 120530 966 120594
rect 1030 120530 1046 120594
rect 1110 120530 1126 120594
rect 1190 120530 1198 120594
rect 878 119506 1198 120530
rect 878 119442 886 119506
rect 950 119442 966 119506
rect 1030 119442 1046 119506
rect 1110 119442 1126 119506
rect 1190 119442 1198 119506
rect 878 118418 1198 119442
rect 878 118354 886 118418
rect 950 118354 966 118418
rect 1030 118354 1046 118418
rect 1110 118354 1126 118418
rect 1190 118354 1198 118418
rect 878 117330 1198 118354
rect 878 117266 886 117330
rect 950 117266 966 117330
rect 1030 117266 1046 117330
rect 1110 117266 1126 117330
rect 1190 117266 1198 117330
rect 878 116242 1198 117266
rect 878 116178 886 116242
rect 950 116178 966 116242
rect 1030 116178 1046 116242
rect 1110 116178 1126 116242
rect 1190 116178 1198 116242
rect 878 115370 1198 116178
rect 878 115154 920 115370
rect 1156 115154 1198 115370
rect 878 115090 886 115154
rect 950 115090 966 115134
rect 1030 115090 1046 115134
rect 1110 115090 1126 115134
rect 1190 115090 1198 115154
rect 878 114066 1198 115090
rect 878 114002 886 114066
rect 950 114002 966 114066
rect 1030 114002 1046 114066
rect 1110 114002 1126 114066
rect 1190 114002 1198 114066
rect 878 112978 1198 114002
rect 878 112914 886 112978
rect 950 112914 966 112978
rect 1030 112914 1046 112978
rect 1110 112914 1126 112978
rect 1190 112914 1198 112978
rect 878 111890 1198 112914
rect 878 111826 886 111890
rect 950 111826 966 111890
rect 1030 111826 1046 111890
rect 1110 111826 1126 111890
rect 1190 111826 1198 111890
rect 878 110802 1198 111826
rect 878 110738 886 110802
rect 950 110738 966 110802
rect 1030 110738 1046 110802
rect 1110 110738 1126 110802
rect 1190 110738 1198 110802
rect 878 109714 1198 110738
rect 878 109650 886 109714
rect 950 109650 966 109714
rect 1030 109650 1046 109714
rect 1110 109650 1126 109714
rect 1190 109650 1198 109714
rect 878 108626 1198 109650
rect 878 108562 886 108626
rect 950 108562 966 108626
rect 1030 108562 1046 108626
rect 1110 108562 1126 108626
rect 1190 108562 1198 108626
rect 878 107538 1198 108562
rect 2308 108151 2368 124677
rect 2878 124402 3198 125426
rect 2878 124338 2886 124402
rect 2950 124338 2966 124402
rect 3030 124338 3046 124402
rect 3110 124338 3126 124402
rect 3190 124338 3198 124402
rect 2878 123314 3198 124338
rect 2878 123250 2886 123314
rect 2950 123250 2966 123314
rect 3030 123250 3046 123314
rect 3110 123250 3126 123314
rect 3190 123250 3198 123314
rect 2878 122226 3198 123250
rect 2878 122162 2886 122226
rect 2950 122162 2966 122226
rect 3030 122162 3046 122226
rect 3110 122162 3126 122226
rect 3190 122162 3198 122226
rect 2878 121138 3198 122162
rect 2878 121074 2886 121138
rect 2950 121074 2966 121138
rect 3030 121074 3046 121138
rect 3110 121074 3126 121138
rect 3190 121074 3198 121138
rect 2878 120370 3198 121074
rect 2878 120134 2920 120370
rect 3156 120134 3198 120370
rect 2878 120050 3198 120134
rect 2878 119986 2886 120050
rect 2950 119986 2966 120050
rect 3030 119986 3046 120050
rect 3110 119986 3126 120050
rect 3190 119986 3198 120050
rect 2878 118962 3198 119986
rect 2878 118898 2886 118962
rect 2950 118898 2966 118962
rect 3030 118898 3046 118962
rect 3110 118898 3126 118962
rect 3190 118898 3198 118962
rect 2878 117874 3198 118898
rect 2878 117810 2886 117874
rect 2950 117810 2966 117874
rect 3030 117810 3046 117874
rect 3110 117810 3126 117874
rect 3190 117810 3198 117874
rect 2878 116786 3198 117810
rect 2878 116722 2886 116786
rect 2950 116722 2966 116786
rect 3030 116722 3046 116786
rect 3110 116722 3126 116786
rect 3190 116722 3198 116786
rect 2878 115698 3198 116722
rect 2878 115634 2886 115698
rect 2950 115634 2966 115698
rect 3030 115634 3046 115698
rect 3110 115634 3126 115698
rect 3190 115634 3198 115698
rect 2878 114610 3198 115634
rect 2878 114546 2886 114610
rect 2950 114546 2966 114610
rect 3030 114546 3046 114610
rect 3110 114546 3126 114610
rect 3190 114546 3198 114610
rect 2878 113522 3198 114546
rect 2878 113458 2886 113522
rect 2950 113458 2966 113522
rect 3030 113458 3046 113522
rect 3110 113458 3126 113522
rect 3190 113458 3198 113522
rect 2878 112434 3198 113458
rect 2878 112370 2886 112434
rect 2950 112370 2966 112434
rect 3030 112370 3046 112434
rect 3110 112370 3126 112434
rect 3190 112370 3198 112434
rect 2878 111346 3198 112370
rect 2878 111282 2886 111346
rect 2950 111282 2966 111346
rect 3030 111282 3046 111346
rect 3110 111282 3126 111346
rect 3190 111282 3198 111346
rect 2878 110370 3198 111282
rect 2878 110258 2920 110370
rect 3156 110258 3198 110370
rect 2878 110194 2886 110258
rect 3190 110194 3198 110258
rect 2878 110134 2920 110194
rect 3156 110134 3198 110194
rect 2878 109170 3198 110134
rect 2878 109106 2886 109170
rect 2950 109106 2966 109170
rect 3030 109106 3046 109170
rect 3110 109106 3126 109170
rect 3190 109106 3198 109170
rect 2305 108150 2371 108151
rect 2305 108086 2306 108150
rect 2370 108086 2371 108150
rect 2305 108085 2371 108086
rect 878 107474 886 107538
rect 950 107474 966 107538
rect 1030 107474 1046 107538
rect 1110 107474 1126 107538
rect 1190 107474 1198 107538
rect 878 106450 1198 107474
rect 878 106386 886 106450
rect 950 106386 966 106450
rect 1030 106386 1046 106450
rect 1110 106386 1126 106450
rect 1190 106386 1198 106450
rect 878 105370 1198 106386
rect 878 105362 920 105370
rect 1156 105362 1198 105370
rect 878 105298 886 105362
rect 1190 105298 1198 105362
rect 878 105134 920 105298
rect 1156 105134 1198 105298
rect 878 104274 1198 105134
rect 878 104210 886 104274
rect 950 104210 966 104274
rect 1030 104210 1046 104274
rect 1110 104210 1126 104274
rect 1190 104210 1198 104274
rect 878 103186 1198 104210
rect 878 103122 886 103186
rect 950 103122 966 103186
rect 1030 103122 1046 103186
rect 1110 103122 1126 103186
rect 1190 103122 1198 103186
rect 878 102098 1198 103122
rect 878 102034 886 102098
rect 950 102034 966 102098
rect 1030 102034 1046 102098
rect 1110 102034 1126 102098
rect 1190 102034 1198 102098
rect 878 101010 1198 102034
rect 878 100946 886 101010
rect 950 100946 966 101010
rect 1030 100946 1046 101010
rect 1110 100946 1126 101010
rect 1190 100946 1198 101010
rect 878 99922 1198 100946
rect 878 99858 886 99922
rect 950 99858 966 99922
rect 1030 99858 1046 99922
rect 1110 99858 1126 99922
rect 1190 99858 1198 99922
rect 878 98834 1198 99858
rect 878 98770 886 98834
rect 950 98770 966 98834
rect 1030 98770 1046 98834
rect 1110 98770 1126 98834
rect 1190 98770 1198 98834
rect 878 97746 1198 98770
rect 878 97682 886 97746
rect 950 97682 966 97746
rect 1030 97682 1046 97746
rect 1110 97682 1126 97746
rect 1190 97682 1198 97746
rect 878 96658 1198 97682
rect 878 96594 886 96658
rect 950 96594 966 96658
rect 1030 96594 1046 96658
rect 1110 96594 1126 96658
rect 1190 96594 1198 96658
rect 878 95570 1198 96594
rect 878 95506 886 95570
rect 950 95506 966 95570
rect 1030 95506 1046 95570
rect 1110 95506 1126 95570
rect 1190 95506 1198 95570
rect 878 95370 1198 95506
rect 878 95134 920 95370
rect 1156 95134 1198 95370
rect 878 94482 1198 95134
rect 878 94418 886 94482
rect 950 94418 966 94482
rect 1030 94418 1046 94482
rect 1110 94418 1126 94482
rect 1190 94418 1198 94482
rect 878 93394 1198 94418
rect 878 93330 886 93394
rect 950 93330 966 93394
rect 1030 93330 1046 93394
rect 1110 93330 1126 93394
rect 1190 93330 1198 93394
rect 878 92306 1198 93330
rect 878 92242 886 92306
rect 950 92242 966 92306
rect 1030 92242 1046 92306
rect 1110 92242 1126 92306
rect 1190 92242 1198 92306
rect 878 91218 1198 92242
rect 878 91154 886 91218
rect 950 91154 966 91218
rect 1030 91154 1046 91218
rect 1110 91154 1126 91218
rect 1190 91154 1198 91218
rect 878 90130 1198 91154
rect 878 90066 886 90130
rect 950 90066 966 90130
rect 1030 90066 1046 90130
rect 1110 90066 1126 90130
rect 1190 90066 1198 90130
rect 878 89042 1198 90066
rect 878 88978 886 89042
rect 950 88978 966 89042
rect 1030 88978 1046 89042
rect 1110 88978 1126 89042
rect 1190 88978 1198 89042
rect 878 87954 1198 88978
rect 878 87890 886 87954
rect 950 87890 966 87954
rect 1030 87890 1046 87954
rect 1110 87890 1126 87954
rect 1190 87890 1198 87954
rect 878 86866 1198 87890
rect 878 86802 886 86866
rect 950 86802 966 86866
rect 1030 86802 1046 86866
rect 1110 86802 1126 86866
rect 1190 86802 1198 86866
rect 878 85778 1198 86802
rect 878 85714 886 85778
rect 950 85714 966 85778
rect 1030 85714 1046 85778
rect 1110 85714 1126 85778
rect 1190 85714 1198 85778
rect 878 85370 1198 85714
rect 878 85134 920 85370
rect 1156 85134 1198 85370
rect 878 84690 1198 85134
rect 878 84626 886 84690
rect 950 84626 966 84690
rect 1030 84626 1046 84690
rect 1110 84626 1126 84690
rect 1190 84626 1198 84690
rect 878 83602 1198 84626
rect 878 83538 886 83602
rect 950 83538 966 83602
rect 1030 83538 1046 83602
rect 1110 83538 1126 83602
rect 1190 83538 1198 83602
rect 878 82514 1198 83538
rect 878 82450 886 82514
rect 950 82450 966 82514
rect 1030 82450 1046 82514
rect 1110 82450 1126 82514
rect 1190 82450 1198 82514
rect 878 81426 1198 82450
rect 878 81362 886 81426
rect 950 81362 966 81426
rect 1030 81362 1046 81426
rect 1110 81362 1126 81426
rect 1190 81362 1198 81426
rect 878 80338 1198 81362
rect 878 80274 886 80338
rect 950 80274 966 80338
rect 1030 80274 1046 80338
rect 1110 80274 1126 80338
rect 1190 80274 1198 80338
rect 878 79250 1198 80274
rect 878 79186 886 79250
rect 950 79186 966 79250
rect 1030 79186 1046 79250
rect 1110 79186 1126 79250
rect 1190 79186 1198 79250
rect 878 78162 1198 79186
rect 878 78098 886 78162
rect 950 78098 966 78162
rect 1030 78098 1046 78162
rect 1110 78098 1126 78162
rect 1190 78098 1198 78162
rect 878 77074 1198 78098
rect 878 77010 886 77074
rect 950 77010 966 77074
rect 1030 77010 1046 77074
rect 1110 77010 1126 77074
rect 1190 77010 1198 77074
rect 878 75986 1198 77010
rect 878 75922 886 75986
rect 950 75922 966 75986
rect 1030 75922 1046 75986
rect 1110 75922 1126 75986
rect 1190 75922 1198 75986
rect 878 75370 1198 75922
rect 878 75134 920 75370
rect 1156 75134 1198 75370
rect 878 74898 1198 75134
rect 878 74834 886 74898
rect 950 74834 966 74898
rect 1030 74834 1046 74898
rect 1110 74834 1126 74898
rect 1190 74834 1198 74898
rect 878 73810 1198 74834
rect 878 73746 886 73810
rect 950 73746 966 73810
rect 1030 73746 1046 73810
rect 1110 73746 1126 73810
rect 1190 73746 1198 73810
rect 878 72722 1198 73746
rect 878 72658 886 72722
rect 950 72658 966 72722
rect 1030 72658 1046 72722
rect 1110 72658 1126 72722
rect 1190 72658 1198 72722
rect 878 71634 1198 72658
rect 878 71570 886 71634
rect 950 71570 966 71634
rect 1030 71570 1046 71634
rect 1110 71570 1126 71634
rect 1190 71570 1198 71634
rect 878 70546 1198 71570
rect 878 70482 886 70546
rect 950 70482 966 70546
rect 1030 70482 1046 70546
rect 1110 70482 1126 70546
rect 1190 70482 1198 70546
rect 878 69458 1198 70482
rect 878 69394 886 69458
rect 950 69394 966 69458
rect 1030 69394 1046 69458
rect 1110 69394 1126 69458
rect 1190 69394 1198 69458
rect 878 68370 1198 69394
rect 878 68306 886 68370
rect 950 68306 966 68370
rect 1030 68306 1046 68370
rect 1110 68306 1126 68370
rect 1190 68306 1198 68370
rect 878 67282 1198 68306
rect 878 67218 886 67282
rect 950 67218 966 67282
rect 1030 67218 1046 67282
rect 1110 67218 1126 67282
rect 1190 67218 1198 67282
rect 878 66194 1198 67218
rect 878 66130 886 66194
rect 950 66130 966 66194
rect 1030 66130 1046 66194
rect 1110 66130 1126 66194
rect 1190 66130 1198 66194
rect 878 65370 1198 66130
rect 878 65134 920 65370
rect 1156 65134 1198 65370
rect 878 65106 1198 65134
rect 878 65042 886 65106
rect 950 65042 966 65106
rect 1030 65042 1046 65106
rect 1110 65042 1126 65106
rect 1190 65042 1198 65106
rect 878 64018 1198 65042
rect 878 63954 886 64018
rect 950 63954 966 64018
rect 1030 63954 1046 64018
rect 1110 63954 1126 64018
rect 1190 63954 1198 64018
rect 878 62930 1198 63954
rect 878 62866 886 62930
rect 950 62866 966 62930
rect 1030 62866 1046 62930
rect 1110 62866 1126 62930
rect 1190 62866 1198 62930
rect 878 61842 1198 62866
rect 878 61778 886 61842
rect 950 61778 966 61842
rect 1030 61778 1046 61842
rect 1110 61778 1126 61842
rect 1190 61778 1198 61842
rect 878 60754 1198 61778
rect 878 60690 886 60754
rect 950 60690 966 60754
rect 1030 60690 1046 60754
rect 1110 60690 1126 60754
rect 1190 60690 1198 60754
rect 878 59666 1198 60690
rect 878 59602 886 59666
rect 950 59602 966 59666
rect 1030 59602 1046 59666
rect 1110 59602 1126 59666
rect 1190 59602 1198 59666
rect 878 58578 1198 59602
rect 878 58514 886 58578
rect 950 58514 966 58578
rect 1030 58514 1046 58578
rect 1110 58514 1126 58578
rect 1190 58514 1198 58578
rect 878 57490 1198 58514
rect 878 57426 886 57490
rect 950 57426 966 57490
rect 1030 57426 1046 57490
rect 1110 57426 1126 57490
rect 1190 57426 1198 57490
rect 878 56402 1198 57426
rect 878 56338 886 56402
rect 950 56338 966 56402
rect 1030 56338 1046 56402
rect 1110 56338 1126 56402
rect 1190 56338 1198 56402
rect 878 55370 1198 56338
rect 878 55314 920 55370
rect 1156 55314 1198 55370
rect 878 55250 886 55314
rect 1190 55250 1198 55314
rect 878 55134 920 55250
rect 1156 55134 1198 55250
rect 878 54226 1198 55134
rect 878 54162 886 54226
rect 950 54162 966 54226
rect 1030 54162 1046 54226
rect 1110 54162 1126 54226
rect 1190 54162 1198 54226
rect 878 53138 1198 54162
rect 878 53074 886 53138
rect 950 53074 966 53138
rect 1030 53074 1046 53138
rect 1110 53074 1126 53138
rect 1190 53074 1198 53138
rect 878 52050 1198 53074
rect 878 51986 886 52050
rect 950 51986 966 52050
rect 1030 51986 1046 52050
rect 1110 51986 1126 52050
rect 1190 51986 1198 52050
rect 878 50962 1198 51986
rect 878 50898 886 50962
rect 950 50898 966 50962
rect 1030 50898 1046 50962
rect 1110 50898 1126 50962
rect 1190 50898 1198 50962
rect 878 49874 1198 50898
rect 878 49810 886 49874
rect 950 49810 966 49874
rect 1030 49810 1046 49874
rect 1110 49810 1126 49874
rect 1190 49810 1198 49874
rect 878 48786 1198 49810
rect 878 48722 886 48786
rect 950 48722 966 48786
rect 1030 48722 1046 48786
rect 1110 48722 1126 48786
rect 1190 48722 1198 48786
rect 878 47698 1198 48722
rect 878 47634 886 47698
rect 950 47634 966 47698
rect 1030 47634 1046 47698
rect 1110 47634 1126 47698
rect 1190 47634 1198 47698
rect 878 46610 1198 47634
rect 878 46546 886 46610
rect 950 46546 966 46610
rect 1030 46546 1046 46610
rect 1110 46546 1126 46610
rect 1190 46546 1198 46610
rect 878 45522 1198 46546
rect 878 45458 886 45522
rect 950 45458 966 45522
rect 1030 45458 1046 45522
rect 1110 45458 1126 45522
rect 1190 45458 1198 45522
rect 878 45370 1198 45458
rect 878 45134 920 45370
rect 1156 45134 1198 45370
rect 878 44434 1198 45134
rect 878 44370 886 44434
rect 950 44370 966 44434
rect 1030 44370 1046 44434
rect 1110 44370 1126 44434
rect 1190 44370 1198 44434
rect 878 43346 1198 44370
rect 878 43282 886 43346
rect 950 43282 966 43346
rect 1030 43282 1046 43346
rect 1110 43282 1126 43346
rect 1190 43282 1198 43346
rect 878 42258 1198 43282
rect 878 42194 886 42258
rect 950 42194 966 42258
rect 1030 42194 1046 42258
rect 1110 42194 1126 42258
rect 1190 42194 1198 42258
rect 878 41170 1198 42194
rect 878 41106 886 41170
rect 950 41106 966 41170
rect 1030 41106 1046 41170
rect 1110 41106 1126 41170
rect 1190 41106 1198 41170
rect 878 40082 1198 41106
rect 878 40018 886 40082
rect 950 40018 966 40082
rect 1030 40018 1046 40082
rect 1110 40018 1126 40082
rect 1190 40018 1198 40082
rect 878 38994 1198 40018
rect 878 38930 886 38994
rect 950 38930 966 38994
rect 1030 38930 1046 38994
rect 1110 38930 1126 38994
rect 1190 38930 1198 38994
rect 878 37906 1198 38930
rect 878 37842 886 37906
rect 950 37842 966 37906
rect 1030 37842 1046 37906
rect 1110 37842 1126 37906
rect 1190 37842 1198 37906
rect 878 36818 1198 37842
rect 878 36754 886 36818
rect 950 36754 966 36818
rect 1030 36754 1046 36818
rect 1110 36754 1126 36818
rect 1190 36754 1198 36818
rect 878 35730 1198 36754
rect 878 35666 886 35730
rect 950 35666 966 35730
rect 1030 35666 1046 35730
rect 1110 35666 1126 35730
rect 1190 35666 1198 35730
rect 878 35370 1198 35666
rect 878 35134 920 35370
rect 1156 35134 1198 35370
rect 878 34642 1198 35134
rect 878 34578 886 34642
rect 950 34578 966 34642
rect 1030 34578 1046 34642
rect 1110 34578 1126 34642
rect 1190 34578 1198 34642
rect 878 33554 1198 34578
rect 878 33490 886 33554
rect 950 33490 966 33554
rect 1030 33490 1046 33554
rect 1110 33490 1126 33554
rect 1190 33490 1198 33554
rect 878 32466 1198 33490
rect 878 32402 886 32466
rect 950 32402 966 32466
rect 1030 32402 1046 32466
rect 1110 32402 1126 32466
rect 1190 32402 1198 32466
rect 878 31378 1198 32402
rect 878 31314 886 31378
rect 950 31314 966 31378
rect 1030 31314 1046 31378
rect 1110 31314 1126 31378
rect 1190 31314 1198 31378
rect 878 30290 1198 31314
rect 878 30226 886 30290
rect 950 30226 966 30290
rect 1030 30226 1046 30290
rect 1110 30226 1126 30290
rect 1190 30226 1198 30290
rect 878 29202 1198 30226
rect 878 29138 886 29202
rect 950 29138 966 29202
rect 1030 29138 1046 29202
rect 1110 29138 1126 29202
rect 1190 29138 1198 29202
rect 878 28114 1198 29138
rect 878 28050 886 28114
rect 950 28050 966 28114
rect 1030 28050 1046 28114
rect 1110 28050 1126 28114
rect 1190 28050 1198 28114
rect 878 27026 1198 28050
rect 878 26962 886 27026
rect 950 26962 966 27026
rect 1030 26962 1046 27026
rect 1110 26962 1126 27026
rect 1190 26962 1198 27026
rect 878 25938 1198 26962
rect 878 25874 886 25938
rect 950 25874 966 25938
rect 1030 25874 1046 25938
rect 1110 25874 1126 25938
rect 1190 25874 1198 25938
rect 878 25370 1198 25874
rect 878 25134 920 25370
rect 1156 25134 1198 25370
rect 878 24850 1198 25134
rect 878 24786 886 24850
rect 950 24786 966 24850
rect 1030 24786 1046 24850
rect 1110 24786 1126 24850
rect 1190 24786 1198 24850
rect 878 23762 1198 24786
rect 878 23698 886 23762
rect 950 23698 966 23762
rect 1030 23698 1046 23762
rect 1110 23698 1126 23762
rect 1190 23698 1198 23762
rect 878 22674 1198 23698
rect 878 22610 886 22674
rect 950 22610 966 22674
rect 1030 22610 1046 22674
rect 1110 22610 1126 22674
rect 1190 22610 1198 22674
rect 878 21586 1198 22610
rect 878 21522 886 21586
rect 950 21522 966 21586
rect 1030 21522 1046 21586
rect 1110 21522 1126 21586
rect 1190 21522 1198 21586
rect 878 20498 1198 21522
rect 878 20434 886 20498
rect 950 20434 966 20498
rect 1030 20434 1046 20498
rect 1110 20434 1126 20498
rect 1190 20434 1198 20498
rect 878 19410 1198 20434
rect 878 19346 886 19410
rect 950 19346 966 19410
rect 1030 19346 1046 19410
rect 1110 19346 1126 19410
rect 1190 19346 1198 19410
rect 878 18322 1198 19346
rect 878 18258 886 18322
rect 950 18258 966 18322
rect 1030 18258 1046 18322
rect 1110 18258 1126 18322
rect 1190 18258 1198 18322
rect 878 17234 1198 18258
rect 878 17170 886 17234
rect 950 17170 966 17234
rect 1030 17170 1046 17234
rect 1110 17170 1126 17234
rect 1190 17170 1198 17234
rect 878 16146 1198 17170
rect 878 16082 886 16146
rect 950 16082 966 16146
rect 1030 16082 1046 16146
rect 1110 16082 1126 16146
rect 1190 16082 1198 16146
rect 878 15370 1198 16082
rect 878 15134 920 15370
rect 1156 15134 1198 15370
rect 878 15058 1198 15134
rect 878 14994 886 15058
rect 950 14994 966 15058
rect 1030 14994 1046 15058
rect 1110 14994 1126 15058
rect 1190 14994 1198 15058
rect 878 13970 1198 14994
rect 878 13906 886 13970
rect 950 13906 966 13970
rect 1030 13906 1046 13970
rect 1110 13906 1126 13970
rect 1190 13906 1198 13970
rect 878 12882 1198 13906
rect 878 12818 886 12882
rect 950 12818 966 12882
rect 1030 12818 1046 12882
rect 1110 12818 1126 12882
rect 1190 12818 1198 12882
rect 878 11794 1198 12818
rect 878 11730 886 11794
rect 950 11730 966 11794
rect 1030 11730 1046 11794
rect 1110 11730 1126 11794
rect 1190 11730 1198 11794
rect 878 10706 1198 11730
rect 878 10642 886 10706
rect 950 10642 966 10706
rect 1030 10642 1046 10706
rect 1110 10642 1126 10706
rect 1190 10642 1198 10706
rect 878 9618 1198 10642
rect 878 9554 886 9618
rect 950 9554 966 9618
rect 1030 9554 1046 9618
rect 1110 9554 1126 9618
rect 1190 9554 1198 9618
rect 878 8530 1198 9554
rect 878 8466 886 8530
rect 950 8466 966 8530
rect 1030 8466 1046 8530
rect 1110 8466 1126 8530
rect 1190 8466 1198 8530
rect 878 7442 1198 8466
rect 878 7378 886 7442
rect 950 7378 966 7442
rect 1030 7378 1046 7442
rect 1110 7378 1126 7442
rect 1190 7378 1198 7442
rect 878 6354 1198 7378
rect 878 6290 886 6354
rect 950 6290 966 6354
rect 1030 6290 1046 6354
rect 1110 6290 1126 6354
rect 1190 6290 1198 6354
rect 878 5370 1198 6290
rect 878 5266 920 5370
rect 1156 5266 1198 5370
rect 878 5202 886 5266
rect 1190 5202 1198 5266
rect 878 5134 920 5202
rect 1156 5134 1198 5202
rect 878 4178 1198 5134
rect 878 4114 886 4178
rect 950 4114 966 4178
rect 1030 4114 1046 4178
rect 1110 4114 1126 4178
rect 1190 4114 1198 4178
rect 878 3090 1198 4114
rect 878 3026 886 3090
rect 950 3026 966 3090
rect 1030 3026 1046 3090
rect 1110 3026 1126 3090
rect 1190 3026 1198 3090
rect 878 2002 1198 3026
rect 878 1938 886 2002
rect 950 1938 966 2002
rect 1030 1938 1046 2002
rect 1110 1938 1126 2002
rect 1190 1938 1198 2002
rect 878 1922 1198 1938
rect 2878 108082 3198 109106
rect 2878 108018 2886 108082
rect 2950 108018 2966 108082
rect 3030 108018 3046 108082
rect 3110 108018 3126 108082
rect 3190 108018 3198 108082
rect 2878 106994 3198 108018
rect 2878 106930 2886 106994
rect 2950 106930 2966 106994
rect 3030 106930 3046 106994
rect 3110 106930 3126 106994
rect 3190 106930 3198 106994
rect 2878 105906 3198 106930
rect 2878 105842 2886 105906
rect 2950 105842 2966 105906
rect 3030 105842 3046 105906
rect 3110 105842 3126 105906
rect 3190 105842 3198 105906
rect 2878 104818 3198 105842
rect 2878 104754 2886 104818
rect 2950 104754 2966 104818
rect 3030 104754 3046 104818
rect 3110 104754 3126 104818
rect 3190 104754 3198 104818
rect 2878 103730 3198 104754
rect 2878 103666 2886 103730
rect 2950 103666 2966 103730
rect 3030 103666 3046 103730
rect 3110 103666 3126 103730
rect 3190 103666 3198 103730
rect 2878 102642 3198 103666
rect 2878 102578 2886 102642
rect 2950 102578 2966 102642
rect 3030 102578 3046 102642
rect 3110 102578 3126 102642
rect 3190 102578 3198 102642
rect 2878 101554 3198 102578
rect 2878 101490 2886 101554
rect 2950 101490 2966 101554
rect 3030 101490 3046 101554
rect 3110 101490 3126 101554
rect 3190 101490 3198 101554
rect 2878 100466 3198 101490
rect 2878 100402 2886 100466
rect 2950 100402 2966 100466
rect 3030 100402 3046 100466
rect 3110 100402 3126 100466
rect 3190 100402 3198 100466
rect 2878 100370 3198 100402
rect 2878 100134 2920 100370
rect 3156 100134 3198 100370
rect 2878 99378 3198 100134
rect 2878 99314 2886 99378
rect 2950 99314 2966 99378
rect 3030 99314 3046 99378
rect 3110 99314 3126 99378
rect 3190 99314 3198 99378
rect 2878 98290 3198 99314
rect 2878 98226 2886 98290
rect 2950 98226 2966 98290
rect 3030 98226 3046 98290
rect 3110 98226 3126 98290
rect 3190 98226 3198 98290
rect 2878 97202 3198 98226
rect 2878 97138 2886 97202
rect 2950 97138 2966 97202
rect 3030 97138 3046 97202
rect 3110 97138 3126 97202
rect 3190 97138 3198 97202
rect 2878 96114 3198 97138
rect 3409 96726 3475 96727
rect 3409 96662 3410 96726
rect 3474 96662 3475 96726
rect 3409 96661 3475 96662
rect 2878 96050 2886 96114
rect 2950 96050 2966 96114
rect 3030 96050 3046 96114
rect 3110 96050 3126 96114
rect 3190 96050 3198 96114
rect 2878 95026 3198 96050
rect 2878 94962 2886 95026
rect 2950 94962 2966 95026
rect 3030 94962 3046 95026
rect 3110 94962 3126 95026
rect 3190 94962 3198 95026
rect 2878 93938 3198 94962
rect 2878 93874 2886 93938
rect 2950 93874 2966 93938
rect 3030 93874 3046 93938
rect 3110 93874 3126 93938
rect 3190 93874 3198 93938
rect 2878 92850 3198 93874
rect 2878 92786 2886 92850
rect 2950 92786 2966 92850
rect 3030 92786 3046 92850
rect 3110 92786 3126 92850
rect 3190 92786 3198 92850
rect 2878 91762 3198 92786
rect 2878 91698 2886 91762
rect 2950 91698 2966 91762
rect 3030 91698 3046 91762
rect 3110 91698 3126 91762
rect 3190 91698 3198 91762
rect 2878 90674 3198 91698
rect 2878 90610 2886 90674
rect 2950 90610 2966 90674
rect 3030 90610 3046 90674
rect 3110 90610 3126 90674
rect 3190 90610 3198 90674
rect 2878 90370 3198 90610
rect 2878 90134 2920 90370
rect 3156 90134 3198 90370
rect 2878 89586 3198 90134
rect 2878 89522 2886 89586
rect 2950 89522 2966 89586
rect 3030 89522 3046 89586
rect 3110 89522 3126 89586
rect 3190 89522 3198 89586
rect 2878 88498 3198 89522
rect 2878 88434 2886 88498
rect 2950 88434 2966 88498
rect 3030 88434 3046 88498
rect 3110 88434 3126 88498
rect 3190 88434 3198 88498
rect 2878 87410 3198 88434
rect 2878 87346 2886 87410
rect 2950 87346 2966 87410
rect 3030 87346 3046 87410
rect 3110 87346 3126 87410
rect 3190 87346 3198 87410
rect 2878 86322 3198 87346
rect 2878 86258 2886 86322
rect 2950 86258 2966 86322
rect 3030 86258 3046 86322
rect 3110 86258 3126 86322
rect 3190 86258 3198 86322
rect 2878 85234 3198 86258
rect 2878 85170 2886 85234
rect 2950 85170 2966 85234
rect 3030 85170 3046 85234
rect 3110 85170 3126 85234
rect 3190 85170 3198 85234
rect 2878 84146 3198 85170
rect 2878 84082 2886 84146
rect 2950 84082 2966 84146
rect 3030 84082 3046 84146
rect 3110 84082 3126 84146
rect 3190 84082 3198 84146
rect 2878 83058 3198 84082
rect 2878 82994 2886 83058
rect 2950 82994 2966 83058
rect 3030 82994 3046 83058
rect 3110 82994 3126 83058
rect 3190 82994 3198 83058
rect 2878 81970 3198 82994
rect 2878 81906 2886 81970
rect 2950 81906 2966 81970
rect 3030 81906 3046 81970
rect 3110 81906 3126 81970
rect 3190 81906 3198 81970
rect 2878 80882 3198 81906
rect 2878 80818 2886 80882
rect 2950 80818 2966 80882
rect 3030 80818 3046 80882
rect 3110 80818 3126 80882
rect 3190 80818 3198 80882
rect 2878 80370 3198 80818
rect 2878 80134 2920 80370
rect 3156 80134 3198 80370
rect 2878 79794 3198 80134
rect 2878 79730 2886 79794
rect 2950 79730 2966 79794
rect 3030 79730 3046 79794
rect 3110 79730 3126 79794
rect 3190 79730 3198 79794
rect 2878 78706 3198 79730
rect 2878 78642 2886 78706
rect 2950 78642 2966 78706
rect 3030 78642 3046 78706
rect 3110 78642 3126 78706
rect 3190 78642 3198 78706
rect 2878 77618 3198 78642
rect 2878 77554 2886 77618
rect 2950 77554 2966 77618
rect 3030 77554 3046 77618
rect 3110 77554 3126 77618
rect 3190 77554 3198 77618
rect 2878 76530 3198 77554
rect 2878 76466 2886 76530
rect 2950 76466 2966 76530
rect 3030 76466 3046 76530
rect 3110 76466 3126 76530
rect 3190 76466 3198 76530
rect 2878 75442 3198 76466
rect 2878 75378 2886 75442
rect 2950 75378 2966 75442
rect 3030 75378 3046 75442
rect 3110 75378 3126 75442
rect 3190 75378 3198 75442
rect 2878 74354 3198 75378
rect 2878 74290 2886 74354
rect 2950 74290 2966 74354
rect 3030 74290 3046 74354
rect 3110 74290 3126 74354
rect 3190 74290 3198 74354
rect 2878 73266 3198 74290
rect 2878 73202 2886 73266
rect 2950 73202 2966 73266
rect 3030 73202 3046 73266
rect 3110 73202 3126 73266
rect 3190 73202 3198 73266
rect 2878 72178 3198 73202
rect 2878 72114 2886 72178
rect 2950 72114 2966 72178
rect 3030 72114 3046 72178
rect 3110 72114 3126 72178
rect 3190 72114 3198 72178
rect 2878 71090 3198 72114
rect 2878 71026 2886 71090
rect 2950 71026 2966 71090
rect 3030 71026 3046 71090
rect 3110 71026 3126 71090
rect 3190 71026 3198 71090
rect 2878 70370 3198 71026
rect 2878 70134 2920 70370
rect 3156 70134 3198 70370
rect 2878 70002 3198 70134
rect 2878 69938 2886 70002
rect 2950 69938 2966 70002
rect 3030 69938 3046 70002
rect 3110 69938 3126 70002
rect 3190 69938 3198 70002
rect 2878 68914 3198 69938
rect 2878 68850 2886 68914
rect 2950 68850 2966 68914
rect 3030 68850 3046 68914
rect 3110 68850 3126 68914
rect 3190 68850 3198 68914
rect 2878 67826 3198 68850
rect 2878 67762 2886 67826
rect 2950 67762 2966 67826
rect 3030 67762 3046 67826
rect 3110 67762 3126 67826
rect 3190 67762 3198 67826
rect 2878 66738 3198 67762
rect 2878 66674 2886 66738
rect 2950 66674 2966 66738
rect 3030 66674 3046 66738
rect 3110 66674 3126 66738
rect 3190 66674 3198 66738
rect 2878 65650 3198 66674
rect 2878 65586 2886 65650
rect 2950 65586 2966 65650
rect 3030 65586 3046 65650
rect 3110 65586 3126 65650
rect 3190 65586 3198 65650
rect 2878 64562 3198 65586
rect 2878 64498 2886 64562
rect 2950 64498 2966 64562
rect 3030 64498 3046 64562
rect 3110 64498 3126 64562
rect 3190 64498 3198 64562
rect 2878 63474 3198 64498
rect 2878 63410 2886 63474
rect 2950 63410 2966 63474
rect 3030 63410 3046 63474
rect 3110 63410 3126 63474
rect 3190 63410 3198 63474
rect 2878 62386 3198 63410
rect 2878 62322 2886 62386
rect 2950 62322 2966 62386
rect 3030 62322 3046 62386
rect 3110 62322 3126 62386
rect 3190 62322 3198 62386
rect 2878 61298 3198 62322
rect 2878 61234 2886 61298
rect 2950 61234 2966 61298
rect 3030 61234 3046 61298
rect 3110 61234 3126 61298
rect 3190 61234 3198 61298
rect 2878 60370 3198 61234
rect 2878 60210 2920 60370
rect 3156 60210 3198 60370
rect 2878 60146 2886 60210
rect 3190 60146 3198 60210
rect 2878 60134 2920 60146
rect 3156 60134 3198 60146
rect 2878 59122 3198 60134
rect 2878 59058 2886 59122
rect 2950 59058 2966 59122
rect 3030 59058 3046 59122
rect 3110 59058 3126 59122
rect 3190 59058 3198 59122
rect 2878 58034 3198 59058
rect 2878 57970 2886 58034
rect 2950 57970 2966 58034
rect 3030 57970 3046 58034
rect 3110 57970 3126 58034
rect 3190 57970 3198 58034
rect 2878 56946 3198 57970
rect 2878 56882 2886 56946
rect 2950 56882 2966 56946
rect 3030 56882 3046 56946
rect 3110 56882 3126 56946
rect 3190 56882 3198 56946
rect 2878 55858 3198 56882
rect 2878 55794 2886 55858
rect 2950 55794 2966 55858
rect 3030 55794 3046 55858
rect 3110 55794 3126 55858
rect 3190 55794 3198 55858
rect 2878 54770 3198 55794
rect 2878 54706 2886 54770
rect 2950 54706 2966 54770
rect 3030 54706 3046 54770
rect 3110 54706 3126 54770
rect 3190 54706 3198 54770
rect 2878 53682 3198 54706
rect 2878 53618 2886 53682
rect 2950 53618 2966 53682
rect 3030 53618 3046 53682
rect 3110 53618 3126 53682
rect 3190 53618 3198 53682
rect 2878 52594 3198 53618
rect 2878 52530 2886 52594
rect 2950 52530 2966 52594
rect 3030 52530 3046 52594
rect 3110 52530 3126 52594
rect 3190 52530 3198 52594
rect 2878 51506 3198 52530
rect 2878 51442 2886 51506
rect 2950 51442 2966 51506
rect 3030 51442 3046 51506
rect 3110 51442 3126 51506
rect 3190 51442 3198 51506
rect 2878 50418 3198 51442
rect 2878 50354 2886 50418
rect 2950 50370 2966 50418
rect 3030 50370 3046 50418
rect 3110 50370 3126 50418
rect 3190 50354 3198 50418
rect 2878 50134 2920 50354
rect 3156 50134 3198 50354
rect 2878 49330 3198 50134
rect 2878 49266 2886 49330
rect 2950 49266 2966 49330
rect 3030 49266 3046 49330
rect 3110 49266 3126 49330
rect 3190 49266 3198 49330
rect 2878 48242 3198 49266
rect 2878 48178 2886 48242
rect 2950 48178 2966 48242
rect 3030 48178 3046 48242
rect 3110 48178 3126 48242
rect 3190 48178 3198 48242
rect 2878 47154 3198 48178
rect 2878 47090 2886 47154
rect 2950 47090 2966 47154
rect 3030 47090 3046 47154
rect 3110 47090 3126 47154
rect 3190 47090 3198 47154
rect 2878 46066 3198 47090
rect 2878 46002 2886 46066
rect 2950 46002 2966 46066
rect 3030 46002 3046 46066
rect 3110 46002 3126 46066
rect 3190 46002 3198 46066
rect 2878 44978 3198 46002
rect 2878 44914 2886 44978
rect 2950 44914 2966 44978
rect 3030 44914 3046 44978
rect 3110 44914 3126 44978
rect 3190 44914 3198 44978
rect 2878 43890 3198 44914
rect 2878 43826 2886 43890
rect 2950 43826 2966 43890
rect 3030 43826 3046 43890
rect 3110 43826 3126 43890
rect 3190 43826 3198 43890
rect 2878 42802 3198 43826
rect 2878 42738 2886 42802
rect 2950 42738 2966 42802
rect 3030 42738 3046 42802
rect 3110 42738 3126 42802
rect 3190 42738 3198 42802
rect 2878 41714 3198 42738
rect 2878 41650 2886 41714
rect 2950 41650 2966 41714
rect 3030 41650 3046 41714
rect 3110 41650 3126 41714
rect 3190 41650 3198 41714
rect 2878 40626 3198 41650
rect 2878 40562 2886 40626
rect 2950 40562 2966 40626
rect 3030 40562 3046 40626
rect 3110 40562 3126 40626
rect 3190 40562 3198 40626
rect 2878 40370 3198 40562
rect 2878 40134 2920 40370
rect 3156 40134 3198 40370
rect 2878 39538 3198 40134
rect 2878 39474 2886 39538
rect 2950 39474 2966 39538
rect 3030 39474 3046 39538
rect 3110 39474 3126 39538
rect 3190 39474 3198 39538
rect 2878 38450 3198 39474
rect 2878 38386 2886 38450
rect 2950 38386 2966 38450
rect 3030 38386 3046 38450
rect 3110 38386 3126 38450
rect 3190 38386 3198 38450
rect 2878 37362 3198 38386
rect 2878 37298 2886 37362
rect 2950 37298 2966 37362
rect 3030 37298 3046 37362
rect 3110 37298 3126 37362
rect 3190 37298 3198 37362
rect 2878 36274 3198 37298
rect 2878 36210 2886 36274
rect 2950 36210 2966 36274
rect 3030 36210 3046 36274
rect 3110 36210 3126 36274
rect 3190 36210 3198 36274
rect 2878 35186 3198 36210
rect 2878 35122 2886 35186
rect 2950 35122 2966 35186
rect 3030 35122 3046 35186
rect 3110 35122 3126 35186
rect 3190 35122 3198 35186
rect 2878 34098 3198 35122
rect 2878 34034 2886 34098
rect 2950 34034 2966 34098
rect 3030 34034 3046 34098
rect 3110 34034 3126 34098
rect 3190 34034 3198 34098
rect 2878 33010 3198 34034
rect 2878 32946 2886 33010
rect 2950 32946 2966 33010
rect 3030 32946 3046 33010
rect 3110 32946 3126 33010
rect 3190 32946 3198 33010
rect 2878 31922 3198 32946
rect 2878 31858 2886 31922
rect 2950 31858 2966 31922
rect 3030 31858 3046 31922
rect 3110 31858 3126 31922
rect 3190 31858 3198 31922
rect 2878 30834 3198 31858
rect 2878 30770 2886 30834
rect 2950 30770 2966 30834
rect 3030 30770 3046 30834
rect 3110 30770 3126 30834
rect 3190 30770 3198 30834
rect 2878 30370 3198 30770
rect 2878 30134 2920 30370
rect 3156 30134 3198 30370
rect 2878 29746 3198 30134
rect 2878 29682 2886 29746
rect 2950 29682 2966 29746
rect 3030 29682 3046 29746
rect 3110 29682 3126 29746
rect 3190 29682 3198 29746
rect 2878 28658 3198 29682
rect 2878 28594 2886 28658
rect 2950 28594 2966 28658
rect 3030 28594 3046 28658
rect 3110 28594 3126 28658
rect 3190 28594 3198 28658
rect 2878 27570 3198 28594
rect 2878 27506 2886 27570
rect 2950 27506 2966 27570
rect 3030 27506 3046 27570
rect 3110 27506 3126 27570
rect 3190 27506 3198 27570
rect 2878 26482 3198 27506
rect 2878 26418 2886 26482
rect 2950 26418 2966 26482
rect 3030 26418 3046 26482
rect 3110 26418 3126 26482
rect 3190 26418 3198 26482
rect 2878 25394 3198 26418
rect 2878 25330 2886 25394
rect 2950 25330 2966 25394
rect 3030 25330 3046 25394
rect 3110 25330 3126 25394
rect 3190 25330 3198 25394
rect 2878 24306 3198 25330
rect 2878 24242 2886 24306
rect 2950 24242 2966 24306
rect 3030 24242 3046 24306
rect 3110 24242 3126 24306
rect 3190 24242 3198 24306
rect 2878 23218 3198 24242
rect 2878 23154 2886 23218
rect 2950 23154 2966 23218
rect 3030 23154 3046 23218
rect 3110 23154 3126 23218
rect 3190 23154 3198 23218
rect 2878 22130 3198 23154
rect 2878 22066 2886 22130
rect 2950 22066 2966 22130
rect 3030 22066 3046 22130
rect 3110 22066 3126 22130
rect 3190 22066 3198 22130
rect 2878 21042 3198 22066
rect 2878 20978 2886 21042
rect 2950 20978 2966 21042
rect 3030 20978 3046 21042
rect 3110 20978 3126 21042
rect 3190 20978 3198 21042
rect 2878 20370 3198 20978
rect 2878 20134 2920 20370
rect 3156 20134 3198 20370
rect 2878 19954 3198 20134
rect 2878 19890 2886 19954
rect 2950 19890 2966 19954
rect 3030 19890 3046 19954
rect 3110 19890 3126 19954
rect 3190 19890 3198 19954
rect 2878 18866 3198 19890
rect 2878 18802 2886 18866
rect 2950 18802 2966 18866
rect 3030 18802 3046 18866
rect 3110 18802 3126 18866
rect 3190 18802 3198 18866
rect 2878 17778 3198 18802
rect 2878 17714 2886 17778
rect 2950 17714 2966 17778
rect 3030 17714 3046 17778
rect 3110 17714 3126 17778
rect 3190 17714 3198 17778
rect 2878 16690 3198 17714
rect 2878 16626 2886 16690
rect 2950 16626 2966 16690
rect 3030 16626 3046 16690
rect 3110 16626 3126 16690
rect 3190 16626 3198 16690
rect 2878 15602 3198 16626
rect 2878 15538 2886 15602
rect 2950 15538 2966 15602
rect 3030 15538 3046 15602
rect 3110 15538 3126 15602
rect 3190 15538 3198 15602
rect 2878 14514 3198 15538
rect 2878 14450 2886 14514
rect 2950 14450 2966 14514
rect 3030 14450 3046 14514
rect 3110 14450 3126 14514
rect 3190 14450 3198 14514
rect 2878 13426 3198 14450
rect 2878 13362 2886 13426
rect 2950 13362 2966 13426
rect 3030 13362 3046 13426
rect 3110 13362 3126 13426
rect 3190 13362 3198 13426
rect 2878 12338 3198 13362
rect 2878 12274 2886 12338
rect 2950 12274 2966 12338
rect 3030 12274 3046 12338
rect 3110 12274 3126 12338
rect 3190 12274 3198 12338
rect 2878 11250 3198 12274
rect 2878 11186 2886 11250
rect 2950 11186 2966 11250
rect 3030 11186 3046 11250
rect 3110 11186 3126 11250
rect 3190 11186 3198 11250
rect 2878 10370 3198 11186
rect 2878 10162 2920 10370
rect 3156 10162 3198 10370
rect 2878 10098 2886 10162
rect 2950 10098 2966 10134
rect 3030 10098 3046 10134
rect 3110 10098 3126 10134
rect 3190 10098 3198 10162
rect 2878 9074 3198 10098
rect 2878 9010 2886 9074
rect 2950 9010 2966 9074
rect 3030 9010 3046 9074
rect 3110 9010 3126 9074
rect 3190 9010 3198 9074
rect 2878 7986 3198 9010
rect 2878 7922 2886 7986
rect 2950 7922 2966 7986
rect 3030 7922 3046 7986
rect 3110 7922 3126 7986
rect 3190 7922 3198 7986
rect 2878 6898 3198 7922
rect 2878 6834 2886 6898
rect 2950 6834 2966 6898
rect 3030 6834 3046 6898
rect 3110 6834 3126 6898
rect 3190 6834 3198 6898
rect 2878 5810 3198 6834
rect 2878 5746 2886 5810
rect 2950 5746 2966 5810
rect 3030 5746 3046 5810
rect 3110 5746 3126 5810
rect 3190 5746 3198 5810
rect 2878 4722 3198 5746
rect 2878 4658 2886 4722
rect 2950 4658 2966 4722
rect 3030 4658 3046 4722
rect 3110 4658 3126 4722
rect 3190 4658 3198 4722
rect 2878 3634 3198 4658
rect 2878 3570 2886 3634
rect 2950 3570 2966 3634
rect 3030 3570 3046 3634
rect 3110 3570 3126 3634
rect 3190 3570 3198 3634
rect 2878 2546 3198 3570
rect 3412 3567 3472 96661
rect 3596 5199 3656 187101
rect 3777 187030 3843 187031
rect 3777 186966 3778 187030
rect 3842 186966 3843 187030
rect 3777 186965 3843 186966
rect 3780 98223 3840 186965
rect 3777 98222 3843 98223
rect 3777 98158 3778 98222
rect 3842 98158 3843 98222
rect 3777 98157 3843 98158
rect 3777 96318 3843 96319
rect 3777 96254 3778 96318
rect 3842 96254 3843 96318
rect 3777 96253 3843 96254
rect 3593 5198 3659 5199
rect 3593 5134 3594 5198
rect 3658 5134 3659 5198
rect 3593 5133 3659 5134
rect 3409 3566 3475 3567
rect 3409 3502 3410 3566
rect 3474 3502 3475 3566
rect 3409 3501 3475 3502
rect 3780 3159 3840 96253
rect 4148 22879 4208 187373
rect 4329 98358 4395 98359
rect 4329 98294 4330 98358
rect 4394 98294 4395 98358
rect 4329 98293 4395 98294
rect 4332 95095 4392 98293
rect 5252 96591 5312 187917
rect 84185 187302 84251 187303
rect 84185 187238 84186 187302
rect 84250 187238 84251 187302
rect 84185 187237 84251 187238
rect 84188 183084 84248 187237
rect 84553 187166 84619 187167
rect 84553 187102 84554 187166
rect 84618 187102 84619 187166
rect 84553 187101 84619 187102
rect 84556 183359 84616 187101
rect 84878 186962 85198 187522
rect 84878 186898 84886 186962
rect 84950 186898 84966 186962
rect 85030 186898 85046 186962
rect 85110 186898 85126 186962
rect 85190 186898 85198 186962
rect 84737 186622 84803 186623
rect 84737 186558 84738 186622
rect 84802 186558 84803 186622
rect 84737 186557 84803 186558
rect 84740 184447 84800 186557
rect 84878 185874 85198 186898
rect 84878 185810 84886 185874
rect 84950 185810 84966 185874
rect 85030 185810 85046 185874
rect 85110 185810 85126 185874
rect 85190 185810 85198 185874
rect 84878 185370 85198 185810
rect 84878 185134 84920 185370
rect 85156 185134 85198 185370
rect 84878 184786 85198 185134
rect 84878 184722 84886 184786
rect 84950 184722 84966 184786
rect 85030 184722 85046 184786
rect 85110 184722 85126 184786
rect 85190 184722 85198 184786
rect 84737 184446 84803 184447
rect 84737 184382 84738 184446
rect 84802 184382 84803 184446
rect 84737 184381 84803 184382
rect 84878 183698 85198 184722
rect 84878 183634 84886 183698
rect 84950 183634 84966 183698
rect 85030 183634 85046 183698
rect 85110 183634 85126 183698
rect 85190 183634 85198 183698
rect 84553 183358 84619 183359
rect 84553 183294 84554 183358
rect 84618 183294 84619 183358
rect 84553 183293 84619 183294
rect 84188 183024 84616 183084
rect 84556 182271 84616 183024
rect 84878 182610 85198 183634
rect 84878 182546 84886 182610
rect 84950 182546 84966 182610
rect 85030 182546 85046 182610
rect 85110 182546 85126 182610
rect 85190 182546 85198 182610
rect 84553 182270 84619 182271
rect 84553 182206 84554 182270
rect 84618 182206 84619 182270
rect 84553 182205 84619 182206
rect 84878 181522 85198 182546
rect 84878 181458 84886 181522
rect 84950 181458 84966 181522
rect 85030 181458 85046 181522
rect 85110 181458 85126 181522
rect 85190 181458 85198 181522
rect 84878 180434 85198 181458
rect 81872 180370 82196 180412
rect 81872 180134 81916 180370
rect 82152 180134 82196 180370
rect 81872 180092 82196 180134
rect 84878 180370 84886 180434
rect 84950 180370 84966 180434
rect 85030 180370 85046 180434
rect 85110 180370 85126 180434
rect 85190 180370 85198 180434
rect 84878 179346 85198 180370
rect 84878 179282 84886 179346
rect 84950 179282 84966 179346
rect 85030 179282 85046 179346
rect 85110 179282 85126 179346
rect 85190 179282 85198 179346
rect 84878 178258 85198 179282
rect 84878 178194 84886 178258
rect 84950 178194 84966 178258
rect 85030 178194 85046 178258
rect 85110 178194 85126 178258
rect 85190 178194 85198 178258
rect 84878 177170 85198 178194
rect 84878 177106 84886 177170
rect 84950 177106 84966 177170
rect 85030 177106 85046 177170
rect 85110 177106 85126 177170
rect 85190 177106 85198 177170
rect 84878 176082 85198 177106
rect 84878 176018 84886 176082
rect 84950 176018 84966 176082
rect 85030 176018 85046 176082
rect 85110 176018 85126 176082
rect 85190 176018 85198 176082
rect 81428 175370 81748 175412
rect 81428 175134 81470 175370
rect 81706 175134 81748 175370
rect 81428 175092 81748 175134
rect 84878 175370 85198 176018
rect 84878 175134 84920 175370
rect 85156 175134 85198 175370
rect 84878 174994 85198 175134
rect 84878 174930 84886 174994
rect 84950 174930 84966 174994
rect 85030 174930 85046 174994
rect 85110 174930 85126 174994
rect 85190 174930 85198 174994
rect 84878 173906 85198 174930
rect 84878 173842 84886 173906
rect 84950 173842 84966 173906
rect 85030 173842 85046 173906
rect 85110 173842 85126 173906
rect 85190 173842 85198 173906
rect 84878 172818 85198 173842
rect 84878 172754 84886 172818
rect 84950 172754 84966 172818
rect 85030 172754 85046 172818
rect 85110 172754 85126 172818
rect 85190 172754 85198 172818
rect 84737 172070 84803 172071
rect 84737 172006 84738 172070
rect 84802 172006 84803 172070
rect 84737 172005 84803 172006
rect 81872 170370 82196 170412
rect 81872 170134 81916 170370
rect 82152 170134 82196 170370
rect 81872 170092 82196 170134
rect 83817 169894 83883 169895
rect 83817 169830 83818 169894
rect 83882 169830 83883 169894
rect 83817 169829 83883 169830
rect 83633 168670 83699 168671
rect 83633 168606 83634 168670
rect 83698 168606 83699 168670
rect 83633 168605 83699 168606
rect 83449 166086 83515 166087
rect 83449 166022 83450 166086
rect 83514 166022 83515 166086
rect 83449 166021 83515 166022
rect 81428 165370 81748 165412
rect 81428 165134 81470 165370
rect 81706 165134 81748 165370
rect 81428 165092 81748 165134
rect 81872 160370 82196 160412
rect 81872 160134 81916 160370
rect 82152 160134 82196 160370
rect 81872 160092 82196 160134
rect 81428 155370 81748 155412
rect 81428 155134 81470 155370
rect 81706 155134 81748 155370
rect 81428 155092 81748 155134
rect 81872 150370 82196 150412
rect 81872 150134 81916 150370
rect 82152 150134 82196 150370
rect 81872 150092 82196 150134
rect 81428 145370 81748 145412
rect 81428 145134 81470 145370
rect 81706 145134 81748 145370
rect 81428 145092 81748 145134
rect 82345 141062 82411 141063
rect 82345 140998 82346 141062
rect 82410 140998 82411 141062
rect 82345 140997 82411 140998
rect 81872 140370 82196 140412
rect 81872 140134 81916 140370
rect 82152 140134 82196 140370
rect 81872 140092 82196 140134
rect 81428 135370 81748 135412
rect 81428 135134 81470 135370
rect 81706 135134 81748 135370
rect 81428 135092 81748 135134
rect 81872 130370 82196 130412
rect 81872 130134 81916 130370
rect 82152 130134 82196 130370
rect 81872 130092 82196 130134
rect 81428 125370 81748 125412
rect 81428 125134 81470 125370
rect 81706 125134 81748 125370
rect 81428 125092 81748 125134
rect 81872 120370 82196 120412
rect 81872 120134 81916 120370
rect 82152 120134 82196 120370
rect 81872 120092 82196 120134
rect 81428 115370 81748 115412
rect 81428 115134 81470 115370
rect 81706 115134 81748 115370
rect 81428 115092 81748 115134
rect 81872 110370 82196 110412
rect 81872 110134 81916 110370
rect 82152 110134 82196 110370
rect 81872 110092 82196 110134
rect 81428 105370 81748 105412
rect 81428 105134 81470 105370
rect 81706 105134 81748 105370
rect 81428 105092 81748 105134
rect 81872 100370 82196 100412
rect 81872 100134 81916 100370
rect 82152 100134 82196 100370
rect 81872 100092 82196 100134
rect 82348 96999 82408 140997
rect 39105 96998 39171 96999
rect 39105 96934 39106 96998
rect 39170 96934 39171 96998
rect 39105 96933 39171 96934
rect 82345 96998 82411 96999
rect 82345 96934 82346 96998
rect 82410 96934 82411 96998
rect 82345 96933 82411 96934
rect 14633 96862 14699 96863
rect 14633 96798 14634 96862
rect 14698 96798 14699 96862
rect 14633 96797 14699 96798
rect 33401 96862 33467 96863
rect 33401 96798 33402 96862
rect 33466 96798 33467 96862
rect 33401 96797 33467 96798
rect 14636 96724 14696 96797
rect 15737 96726 15803 96727
rect 14636 96664 15270 96724
rect 15737 96662 15738 96726
rect 15802 96724 15803 96726
rect 21993 96726 22059 96727
rect 15802 96664 16438 96724
rect 15802 96662 15803 96664
rect 15737 96661 15803 96662
rect 21993 96662 21994 96726
rect 22058 96724 22059 96726
rect 25305 96726 25371 96727
rect 22058 96664 22278 96724
rect 22058 96662 22059 96664
rect 21993 96661 22059 96662
rect 25305 96662 25306 96726
rect 25370 96724 25371 96726
rect 28985 96726 29051 96727
rect 25370 96664 25782 96724
rect 25370 96662 25371 96664
rect 25305 96661 25371 96662
rect 28985 96662 28986 96726
rect 29050 96724 29051 96726
rect 29976 96726 30042 96727
rect 29050 96664 29286 96724
rect 29050 96662 29051 96664
rect 28985 96661 29051 96662
rect 29976 96662 29977 96726
rect 30041 96724 30042 96726
rect 33404 96724 33464 96797
rect 34968 96726 35034 96727
rect 30041 96664 30454 96724
rect 33404 96664 33958 96724
rect 30041 96662 30042 96664
rect 29976 96661 30042 96662
rect 34968 96662 34969 96726
rect 35033 96724 35034 96726
rect 36897 96726 36963 96727
rect 35033 96664 35126 96724
rect 35033 96662 35034 96664
rect 34968 96661 35034 96662
rect 36897 96662 36898 96726
rect 36962 96724 36963 96726
rect 39108 96724 39168 96933
rect 83452 96863 83512 166021
rect 83636 97679 83696 168605
rect 83633 97678 83699 97679
rect 83633 97614 83634 97678
rect 83698 97614 83699 97678
rect 83633 97613 83699 97614
rect 45361 96862 45427 96863
rect 45361 96798 45362 96862
rect 45426 96798 45427 96862
rect 45361 96797 45427 96798
rect 83449 96862 83515 96863
rect 83449 96798 83450 96862
rect 83514 96798 83515 96862
rect 83449 96797 83515 96798
rect 44257 96726 44323 96727
rect 36962 96664 37462 96724
rect 39108 96664 39798 96724
rect 40396 96664 40966 96724
rect 36962 96662 36963 96664
rect 36897 96661 36963 96662
rect 5249 96590 5315 96591
rect 5249 96526 5250 96590
rect 5314 96526 5315 96590
rect 5249 96525 5315 96526
rect 40396 96455 40456 96664
rect 44257 96662 44258 96726
rect 44322 96724 44323 96726
rect 45364 96724 45424 96797
rect 48857 96726 48923 96727
rect 44322 96664 44470 96724
rect 45364 96664 45638 96724
rect 44322 96662 44323 96664
rect 44257 96661 44323 96662
rect 48857 96662 48858 96726
rect 48922 96724 48923 96726
rect 50145 96726 50211 96727
rect 48922 96664 49142 96724
rect 48922 96662 48923 96664
rect 48857 96661 48923 96662
rect 50145 96662 50146 96726
rect 50210 96724 50211 96726
rect 82161 96726 82227 96727
rect 50210 96664 50310 96724
rect 52356 96664 52646 96724
rect 50210 96662 50211 96664
rect 50145 96661 50211 96662
rect 4513 96454 4579 96455
rect 4513 96390 4514 96454
rect 4578 96390 4579 96454
rect 4513 96389 4579 96390
rect 40393 96454 40459 96455
rect 40393 96390 40394 96454
rect 40458 96390 40459 96454
rect 40393 96389 40459 96390
rect 4329 95094 4395 95095
rect 4329 95030 4330 95094
rect 4394 95030 4395 95094
rect 4329 95029 4395 95030
rect 4516 89924 4576 96389
rect 8196 96324 8767 96384
rect 11324 96324 11766 96384
rect 12244 96324 12934 96384
rect 4878 94354 5198 95250
rect 6878 94354 7198 95250
rect 8196 95095 8256 96324
rect 8193 95094 8259 95095
rect 8193 95030 8194 95094
rect 8258 95030 8259 95094
rect 8193 95029 8259 95030
rect 8878 94354 9198 95250
rect 10878 94354 11198 95250
rect 11324 94959 11384 96324
rect 12244 95095 12304 96324
rect 14072 95911 14132 96354
rect 17576 95911 17636 96354
rect 17730 96324 18192 96384
rect 14069 95910 14135 95911
rect 14069 95846 14070 95910
rect 14134 95846 14135 95910
rect 14069 95845 14135 95846
rect 17573 95910 17639 95911
rect 17573 95846 17574 95910
rect 17638 95846 17639 95910
rect 17573 95845 17639 95846
rect 12241 95094 12307 95095
rect 12241 95030 12242 95094
rect 12306 95030 12307 95094
rect 12241 95029 12307 95030
rect 11321 94958 11387 94959
rect 11321 94894 11322 94958
rect 11386 94894 11387 94958
rect 11321 94893 11387 94894
rect 12878 94354 13198 95250
rect 14878 94354 15198 95250
rect 16878 94354 17198 95250
rect 18132 94823 18192 96324
rect 18500 96324 18774 96384
rect 18500 96047 18560 96324
rect 18497 96046 18563 96047
rect 18497 95982 18498 96046
rect 18562 95982 18563 96046
rect 18497 95981 18563 95982
rect 18868 95908 18928 96354
rect 18684 95848 18928 95908
rect 19788 96324 19942 96384
rect 18129 94822 18195 94823
rect 18129 94758 18130 94822
rect 18194 94758 18195 94822
rect 18129 94757 18195 94758
rect 18684 94415 18744 95848
rect 19788 95775 19848 96324
rect 20036 96044 20096 96354
rect 19972 95984 20096 96044
rect 21080 96044 21140 96354
rect 21234 96324 21872 96384
rect 22402 96324 22792 96384
rect 21080 95984 21504 96044
rect 19785 95774 19851 95775
rect 19785 95710 19786 95774
rect 19850 95710 19851 95774
rect 19785 95709 19851 95710
rect 18681 94414 18747 94415
rect 18681 94350 18682 94414
rect 18746 94350 18747 94414
rect 18878 94354 19198 95250
rect 19972 94823 20032 95984
rect 19969 94822 20035 94823
rect 19969 94758 19970 94822
rect 20034 94758 20035 94822
rect 19969 94757 20035 94758
rect 20878 94354 21198 95250
rect 21444 94823 21504 95984
rect 21441 94822 21507 94823
rect 21441 94758 21442 94822
rect 21506 94758 21507 94822
rect 21441 94757 21507 94758
rect 18681 94349 18747 94350
rect 21812 94279 21872 96324
rect 22732 94959 22792 96324
rect 23416 96047 23476 96354
rect 23570 96324 23896 96384
rect 23413 96046 23479 96047
rect 23413 95982 23414 96046
rect 23478 95982 23479 96046
rect 23413 95981 23479 95982
rect 22729 94958 22795 94959
rect 22729 94894 22730 94958
rect 22794 94894 22795 94958
rect 22729 94893 22795 94894
rect 22878 94354 23198 95250
rect 21809 94278 21875 94279
rect 21809 94214 21810 94278
rect 21874 94214 21875 94278
rect 21809 94213 21875 94214
rect 23836 94143 23896 96324
rect 24020 96324 24614 96384
rect 24738 96324 25368 96384
rect 24020 95911 24080 96324
rect 24017 95910 24083 95911
rect 24017 95846 24018 95910
rect 24082 95846 24083 95910
rect 24017 95845 24083 95846
rect 24385 95230 24451 95231
rect 24385 95166 24386 95230
rect 24450 95166 24451 95230
rect 24385 95165 24451 95166
rect 23833 94142 23899 94143
rect 23833 94078 23834 94142
rect 23898 94078 23899 94142
rect 23833 94077 23899 94078
rect 24388 93324 24448 95165
rect 24878 94354 25198 95250
rect 25308 94959 25368 96324
rect 25876 96044 25936 96354
rect 25860 95984 25936 96044
rect 26412 96324 26950 96384
rect 25673 95230 25739 95231
rect 25673 95166 25674 95230
rect 25738 95166 25739 95230
rect 25673 95165 25739 95166
rect 25305 94958 25371 94959
rect 25305 94894 25306 94958
rect 25370 94894 25371 94958
rect 25305 94893 25371 94894
rect 25676 93324 25736 95165
rect 23769 93264 24448 93324
rect 25017 93264 25736 93324
rect 25860 93191 25920 95984
rect 26412 94823 26472 96324
rect 27044 96044 27104 96354
rect 27516 96324 28118 96384
rect 28242 96324 28312 96384
rect 29410 96324 29784 96384
rect 27044 95984 27208 96044
rect 27148 95639 27208 95984
rect 27145 95638 27211 95639
rect 27145 95574 27146 95638
rect 27210 95574 27211 95638
rect 27145 95573 27211 95574
rect 26593 95230 26659 95231
rect 26593 95166 26594 95230
rect 26658 95166 26659 95230
rect 26593 95165 26659 95166
rect 26409 94822 26475 94823
rect 26409 94758 26410 94822
rect 26474 94758 26475 94822
rect 26409 94757 26475 94758
rect 26596 93324 26656 95165
rect 26878 94354 27198 95250
rect 27516 94687 27576 96324
rect 27513 94686 27579 94687
rect 27513 94622 27514 94686
rect 27578 94622 27579 94686
rect 27513 94621 27579 94622
rect 28252 94143 28312 96324
rect 29353 95774 29419 95775
rect 29353 95710 29354 95774
rect 29418 95710 29419 95774
rect 29353 95709 29419 95710
rect 28878 94354 29198 95250
rect 28249 94142 28315 94143
rect 28249 94078 28250 94142
rect 28314 94078 28315 94142
rect 28249 94077 28315 94078
rect 27480 93598 27546 93599
rect 27480 93534 27481 93598
rect 27545 93534 27546 93598
rect 27480 93533 27546 93534
rect 26265 93264 26656 93324
rect 27483 93294 27543 93533
rect 29356 93324 29416 95709
rect 29724 94415 29784 96324
rect 30548 96044 30608 96354
rect 31380 96324 31622 96384
rect 31746 96324 32360 96384
rect 30548 95984 30704 96044
rect 29721 94414 29787 94415
rect 29721 94350 29722 94414
rect 29786 94350 29787 94414
rect 29721 94349 29787 94350
rect 30644 94007 30704 95984
rect 30878 94354 31198 95250
rect 31380 95095 31440 96324
rect 31745 95910 31811 95911
rect 31745 95846 31746 95910
rect 31810 95846 31811 95910
rect 31745 95845 31811 95846
rect 31377 95094 31443 95095
rect 31377 95030 31378 95094
rect 31442 95030 31443 95094
rect 31377 95029 31443 95030
rect 30641 94006 30707 94007
rect 30641 93942 30642 94006
rect 30706 93942 30707 94006
rect 30641 93941 30707 93942
rect 30641 93870 30707 93871
rect 30641 93806 30642 93870
rect 30706 93806 30707 93870
rect 30641 93805 30707 93806
rect 30644 93324 30704 93805
rect 31748 93324 31808 95845
rect 32300 93871 32360 96324
rect 32484 96324 32790 96384
rect 32914 96324 33464 96384
rect 34082 96324 34752 96384
rect 35250 96324 35856 96384
rect 32484 94687 32544 96324
rect 32665 96046 32731 96047
rect 32665 95982 32666 96046
rect 32730 95982 32731 96046
rect 32665 95981 32731 95982
rect 32481 94686 32547 94687
rect 32481 94622 32482 94686
rect 32546 94622 32547 94686
rect 32481 94621 32547 94622
rect 32297 93870 32363 93871
rect 32297 93806 32298 93870
rect 32362 93806 32363 93870
rect 32297 93805 32363 93806
rect 32668 93324 32728 95981
rect 32878 94354 33198 95250
rect 33404 93871 33464 96324
rect 34321 95230 34387 95231
rect 34321 95166 34322 95230
rect 34386 95166 34387 95230
rect 34321 95165 34387 95166
rect 33401 93870 33467 93871
rect 33401 93806 33402 93870
rect 33466 93806 33467 93870
rect 33401 93805 33467 93806
rect 34324 93324 34384 95165
rect 34692 93871 34752 96324
rect 34878 94354 35198 95250
rect 35609 95230 35675 95231
rect 35609 95166 35610 95230
rect 35674 95166 35675 95230
rect 35609 95165 35675 95166
rect 34689 93870 34755 93871
rect 34689 93806 34690 93870
rect 34754 93806 34755 93870
rect 34689 93805 34755 93806
rect 35612 93324 35672 95165
rect 35796 93871 35856 96324
rect 36264 96044 36324 96354
rect 36418 96324 36776 96384
rect 37586 96324 38064 96384
rect 36264 95984 36408 96044
rect 36161 95230 36227 95231
rect 36161 95166 36162 95230
rect 36226 95166 36227 95230
rect 36161 95165 36227 95166
rect 35793 93870 35859 93871
rect 35793 93806 35794 93870
rect 35858 93806 35859 93870
rect 35793 93805 35859 93806
rect 28761 93264 29416 93324
rect 30009 93264 30704 93324
rect 31257 93264 31808 93324
rect 32505 93264 32728 93324
rect 33753 93264 34384 93324
rect 35001 93264 35672 93324
rect 36164 93324 36224 95165
rect 36348 95095 36408 95984
rect 36716 95095 36776 96324
rect 36345 95094 36411 95095
rect 36345 95030 36346 95094
rect 36410 95030 36411 95094
rect 36345 95029 36411 95030
rect 36713 95094 36779 95095
rect 36713 95030 36714 95094
rect 36778 95030 36779 95094
rect 36713 95029 36779 95030
rect 36878 94354 37198 95250
rect 37449 95230 37515 95231
rect 37449 95166 37450 95230
rect 37514 95166 37515 95230
rect 37449 95165 37515 95166
rect 36164 93264 36249 93324
rect 37452 93264 37512 95165
rect 38004 93871 38064 96324
rect 38188 96324 38630 96384
rect 38188 96183 38248 96324
rect 38185 96182 38251 96183
rect 38185 96118 38186 96182
rect 38250 96118 38251 96182
rect 38185 96117 38251 96118
rect 38553 95230 38619 95231
rect 38553 95166 38554 95230
rect 38618 95166 38619 95230
rect 38553 95165 38619 95166
rect 38001 93870 38067 93871
rect 38001 93806 38002 93870
rect 38066 93806 38067 93870
rect 38001 93805 38067 93806
rect 38556 93324 38616 95165
rect 38740 95095 38800 96384
rect 39922 96324 40088 96384
rect 41090 96324 41376 96384
rect 38737 95094 38803 95095
rect 38737 95030 38738 95094
rect 38802 95030 38803 95094
rect 38737 95029 38803 95030
rect 38878 94354 39198 95250
rect 40028 94551 40088 96324
rect 40025 94550 40091 94551
rect 40025 94486 40026 94550
rect 40090 94486 40091 94550
rect 40025 94485 40091 94486
rect 40878 94354 41198 95250
rect 41316 94415 41376 96324
rect 41500 96324 42134 96384
rect 42258 96324 42664 96384
rect 41500 94551 41560 96324
rect 41865 95230 41931 95231
rect 41865 95166 41866 95230
rect 41930 95166 41931 95230
rect 41865 95165 41931 95166
rect 41497 94550 41563 94551
rect 41497 94486 41498 94550
rect 41562 94486 41563 94550
rect 41497 94485 41563 94486
rect 41313 94414 41379 94415
rect 41313 94350 41314 94414
rect 41378 94350 41379 94414
rect 41313 94349 41379 94350
rect 41681 94414 41747 94415
rect 41681 94350 41682 94414
rect 41746 94350 41747 94414
rect 41681 94349 41747 94350
rect 39960 93870 40026 93871
rect 39960 93806 39961 93870
rect 40025 93806 40026 93870
rect 39960 93805 40026 93806
rect 38556 93264 38745 93324
rect 39963 93294 40023 93805
rect 25857 93190 25923 93191
rect 25857 93126 25858 93190
rect 25922 93126 25923 93190
rect 25857 93125 25923 93126
rect 41684 92984 41744 94349
rect 41868 93324 41928 95165
rect 42604 94551 42664 96324
rect 43272 96044 43332 96354
rect 43426 96324 43952 96384
rect 43272 95984 43400 96044
rect 42601 94550 42667 94551
rect 42601 94486 42602 94550
rect 42666 94486 42667 94550
rect 42601 94485 42667 94486
rect 42878 94354 43198 95250
rect 43340 95095 43400 95984
rect 43705 95230 43771 95231
rect 43705 95166 43706 95230
rect 43770 95166 43771 95230
rect 43705 95165 43771 95166
rect 43337 95094 43403 95095
rect 43337 95030 43338 95094
rect 43402 95030 43403 95094
rect 43337 95029 43403 95030
rect 41868 93264 42489 93324
rect 43708 93264 43768 95165
rect 43892 94415 43952 96324
rect 44564 96044 44624 96354
rect 44564 95984 44688 96044
rect 44441 95230 44507 95231
rect 44441 95166 44442 95230
rect 44506 95166 44507 95230
rect 44441 95165 44507 95166
rect 43889 94414 43955 94415
rect 43889 94350 43890 94414
rect 43954 94350 43955 94414
rect 43889 94349 43955 94350
rect 44444 93324 44504 95165
rect 44628 94415 44688 95984
rect 44625 94414 44691 94415
rect 44625 94350 44626 94414
rect 44690 94350 44691 94414
rect 44878 94354 45198 95250
rect 44625 94349 44691 94350
rect 45732 94007 45792 96354
rect 46776 96044 46836 96354
rect 46930 96324 47632 96384
rect 47572 96183 47632 96324
rect 47017 96182 47083 96183
rect 47017 96118 47018 96182
rect 47082 96118 47083 96182
rect 47017 96117 47083 96118
rect 47569 96182 47635 96183
rect 47569 96118 47570 96182
rect 47634 96118 47635 96182
rect 47569 96117 47635 96118
rect 47020 96044 47080 96117
rect 46776 95984 47080 96044
rect 46465 95230 46531 95231
rect 46465 95166 46466 95230
rect 46530 95166 46531 95230
rect 46465 95165 46531 95166
rect 45729 94006 45795 94007
rect 45729 93942 45730 94006
rect 45794 93942 45795 94006
rect 45729 93941 45795 93942
rect 46468 93324 46528 95165
rect 46878 94354 47198 95250
rect 47753 95230 47819 95231
rect 47753 95166 47754 95230
rect 47818 95166 47819 95230
rect 47753 95165 47819 95166
rect 47756 93324 47816 95165
rect 47940 95095 48000 96384
rect 48098 96324 48552 96384
rect 49266 96324 49840 96384
rect 47937 95094 48003 95095
rect 47937 95030 47938 95094
rect 48002 95030 48003 95094
rect 47937 95029 48003 95030
rect 48492 94687 48552 96324
rect 48673 95230 48739 95231
rect 48673 95166 48674 95230
rect 48738 95166 48739 95230
rect 48673 95165 48739 95166
rect 48489 94686 48555 94687
rect 48489 94622 48490 94686
rect 48554 94622 48555 94686
rect 48489 94621 48555 94622
rect 44444 93264 44985 93324
rect 46233 93264 46528 93324
rect 47481 93264 47816 93324
rect 48676 93264 48736 95165
rect 48878 94354 49198 95250
rect 49780 94823 49840 96324
rect 50404 96044 50464 96354
rect 50332 95984 50464 96044
rect 50145 95230 50211 95231
rect 50145 95166 50146 95230
rect 50210 95166 50211 95230
rect 50145 95165 50211 95166
rect 49777 94822 49843 94823
rect 49777 94758 49778 94822
rect 49842 94758 49843 94822
rect 49777 94757 49843 94758
rect 50148 93324 50208 95165
rect 50332 95095 50392 95984
rect 51436 95639 51496 96384
rect 51602 96324 51680 96384
rect 51433 95638 51499 95639
rect 51433 95574 51434 95638
rect 51498 95574 51499 95638
rect 51433 95573 51499 95574
rect 50329 95094 50395 95095
rect 50329 95030 50330 95094
rect 50394 95030 50395 95094
rect 50329 95029 50395 95030
rect 50878 94354 51198 95250
rect 51433 95230 51499 95231
rect 51433 95166 51434 95230
rect 51498 95166 51499 95230
rect 51433 95165 51499 95166
rect 51436 93324 51496 95165
rect 51620 94415 51680 96324
rect 52356 94823 52416 96664
rect 82161 96662 82162 96726
rect 82226 96662 82227 96726
rect 82161 96661 82227 96662
rect 52740 96044 52800 96354
rect 52724 95984 52800 96044
rect 53784 96044 53844 96354
rect 53938 96324 54256 96384
rect 53784 95984 53888 96044
rect 52353 94822 52419 94823
rect 52353 94758 52354 94822
rect 52418 94758 52419 94822
rect 52353 94757 52419 94758
rect 52724 94687 52784 95984
rect 52721 94686 52787 94687
rect 52721 94622 52722 94686
rect 52786 94622 52787 94686
rect 52721 94621 52787 94622
rect 51617 94414 51683 94415
rect 51617 94350 51618 94414
rect 51682 94350 51683 94414
rect 52878 94354 53198 95250
rect 53828 94551 53888 95984
rect 54196 95095 54256 96324
rect 82164 95364 82224 96661
rect 82529 96590 82595 96591
rect 82529 96526 82530 96590
rect 82594 96526 82595 96590
rect 82529 96525 82595 96526
rect 82164 95304 82408 95364
rect 54193 95094 54259 95095
rect 54193 95030 54194 95094
rect 54258 95030 54259 95094
rect 54193 95029 54259 95030
rect 53825 94550 53891 94551
rect 53825 94486 53826 94550
rect 53890 94486 53891 94550
rect 53825 94485 53891 94486
rect 54878 94354 55198 95250
rect 56585 95230 56651 95231
rect 56585 95166 56586 95230
rect 56650 95166 56651 95230
rect 56585 95165 56651 95166
rect 51617 94349 51683 94350
rect 52905 94006 52971 94007
rect 52905 93942 52906 94006
rect 52970 93942 52971 94006
rect 52905 93941 52971 93942
rect 52908 93324 52968 93941
rect 53688 93870 53754 93871
rect 53688 93806 53689 93870
rect 53753 93806 53754 93870
rect 53688 93805 53754 93806
rect 49977 93264 50208 93324
rect 51225 93264 51496 93324
rect 52473 93264 52968 93324
rect 53691 93294 53751 93805
rect 56588 93324 56648 95165
rect 56878 94354 57198 95250
rect 57873 95230 57939 95231
rect 57873 95166 57874 95230
rect 57938 95166 57939 95230
rect 57873 95165 57939 95166
rect 57876 93324 57936 95165
rect 58878 94354 59198 95250
rect 59345 95230 59411 95231
rect 59345 95166 59346 95230
rect 59410 95166 59411 95230
rect 59345 95165 59411 95166
rect 59348 93324 59408 95165
rect 60878 94354 61198 95250
rect 61737 95230 61803 95231
rect 61737 95166 61738 95230
rect 61802 95166 61803 95230
rect 61737 95165 61803 95166
rect 62657 95230 62723 95231
rect 62657 95166 62658 95230
rect 62722 95166 62723 95230
rect 62657 95165 62723 95166
rect 61740 93324 61800 95165
rect 62660 93324 62720 95165
rect 62878 94354 63198 95250
rect 64878 94354 65198 95250
rect 66878 94354 67198 95250
rect 68878 94354 69198 95250
rect 69833 94414 69899 94415
rect 69833 94350 69834 94414
rect 69898 94350 69899 94414
rect 70878 94354 71198 95250
rect 72878 94354 73198 95250
rect 74878 94354 75198 95250
rect 76878 94354 77198 95250
rect 78878 94354 79198 95250
rect 80878 94354 81198 95250
rect 69833 94349 69899 94350
rect 69836 93871 69896 94349
rect 69833 93870 69899 93871
rect 69833 93806 69834 93870
rect 69898 93806 69899 93870
rect 69833 93805 69899 93806
rect 78481 93870 78547 93871
rect 78481 93806 78482 93870
rect 78546 93806 78547 93870
rect 78481 93805 78547 93806
rect 56217 93264 56648 93324
rect 57465 93264 57936 93324
rect 58713 93264 59408 93324
rect 61209 93264 61800 93324
rect 62457 93264 62720 93324
rect 78484 93264 78544 93805
rect 41241 92924 41744 92984
rect 55297 92646 55363 92647
rect 55297 92644 55298 92646
rect 54969 92584 55298 92644
rect 55297 92582 55298 92584
rect 55362 92582 55363 92646
rect 60449 92646 60515 92647
rect 60449 92644 60450 92646
rect 59961 92584 60450 92644
rect 55297 92581 55363 92582
rect 60449 92582 60450 92584
rect 60514 92582 60515 92646
rect 73697 92646 73763 92647
rect 73697 92644 73698 92646
rect 73542 92584 73698 92644
rect 60449 92581 60515 92582
rect 73697 92582 73698 92584
rect 73762 92582 73763 92646
rect 73697 92581 73763 92582
rect 81872 90370 82196 90412
rect 81872 90134 81916 90370
rect 82152 90134 82196 90370
rect 81872 90092 82196 90134
rect 4516 89864 4760 89924
rect 4700 83671 4760 89864
rect 81428 85370 81748 85412
rect 81428 85134 81470 85370
rect 81706 85134 81748 85370
rect 81428 85092 81748 85134
rect 4697 83670 4763 83671
rect 4697 83606 4698 83670
rect 4762 83606 4763 83670
rect 4697 83605 4763 83606
rect 4697 83398 4763 83399
rect 4697 83334 4698 83398
rect 4762 83334 4763 83398
rect 4697 83333 4763 83334
rect 4700 74695 4760 83333
rect 81872 80370 82196 80412
rect 81872 80134 81916 80370
rect 82152 80134 82196 80370
rect 81872 80092 82196 80134
rect 81428 75370 81748 75412
rect 81428 75134 81470 75370
rect 81706 75134 81748 75370
rect 81428 75092 81748 75134
rect 4697 74694 4763 74695
rect 4697 74630 4698 74694
rect 4762 74630 4763 74694
rect 4697 74629 4763 74630
rect 4513 74422 4579 74423
rect 4513 74358 4514 74422
rect 4578 74358 4579 74422
rect 4513 74357 4579 74358
rect 4516 65583 4576 74357
rect 81872 70370 82196 70412
rect 81872 70134 81916 70370
rect 82152 70134 82196 70370
rect 81872 70092 82196 70134
rect 4513 65582 4579 65583
rect 4513 65518 4514 65582
rect 4578 65518 4579 65582
rect 4513 65517 4579 65518
rect 81428 65370 81748 65412
rect 4697 65310 4763 65311
rect 4697 65246 4698 65310
rect 4762 65246 4763 65310
rect 4697 65245 4763 65246
rect 4700 56604 4760 65245
rect 81428 65134 81470 65370
rect 81706 65134 81748 65370
rect 81428 65092 81748 65134
rect 81872 60370 82196 60412
rect 81872 60134 81916 60370
rect 82152 60134 82196 60370
rect 81872 60092 82196 60134
rect 4332 56544 4760 56604
rect 4332 55924 4392 56544
rect 4332 55864 4760 55924
rect 4145 22878 4211 22879
rect 4145 22814 4146 22878
rect 4210 22814 4211 22878
rect 4145 22813 4211 22814
rect 4700 20564 4760 55864
rect 81428 55370 81748 55412
rect 81428 55134 81470 55370
rect 81706 55134 81748 55370
rect 81428 55092 81748 55134
rect 81872 50370 82196 50412
rect 81872 50134 81916 50370
rect 82152 50134 82196 50370
rect 81872 50092 82196 50134
rect 81428 45370 81748 45412
rect 81428 45134 81470 45370
rect 81706 45134 81748 45370
rect 81428 45092 81748 45134
rect 81872 40370 82196 40412
rect 81872 40134 81916 40370
rect 82152 40134 82196 40370
rect 81872 40092 82196 40134
rect 81428 35370 81748 35412
rect 81428 35134 81470 35370
rect 81706 35134 81748 35370
rect 81428 35092 81748 35134
rect 81872 30370 82196 30412
rect 81872 30134 81916 30370
rect 82152 30134 82196 30370
rect 81872 30092 82196 30134
rect 5617 29542 5683 29543
rect 5617 29492 5618 29542
rect 5682 29492 5683 29542
rect 81428 25370 81748 25412
rect 81428 25134 81470 25370
rect 81706 25134 81748 25370
rect 81428 25092 81748 25134
rect 82348 24511 82408 95304
rect 82345 24510 82411 24511
rect 82345 24446 82346 24510
rect 82410 24446 82411 24510
rect 82345 24445 82411 24446
rect 82345 24102 82411 24103
rect 82345 24038 82346 24102
rect 82410 24038 82411 24102
rect 82345 24037 82411 24038
rect 4516 20504 4760 20564
rect 4516 11724 4576 20504
rect 81872 20370 82196 20412
rect 81872 20134 81916 20370
rect 82152 20134 82196 20370
rect 81872 20092 82196 20134
rect 82348 15535 82408 24037
rect 82345 15534 82411 15535
rect 82345 15470 82346 15534
rect 82410 15470 82411 15534
rect 82345 15469 82411 15470
rect 81428 15370 81748 15412
rect 81428 15134 81470 15370
rect 81706 15134 81748 15370
rect 82345 15398 82411 15399
rect 82345 15334 82346 15398
rect 82410 15334 82411 15398
rect 82345 15333 82411 15334
rect 81428 15092 81748 15134
rect 4148 11664 4576 11724
rect 4148 4655 4208 11664
rect 81872 10370 82196 10412
rect 81872 10134 81916 10370
rect 82152 10134 82196 10370
rect 81872 10092 82196 10134
rect 82348 6151 82408 15333
rect 82345 6150 82411 6151
rect 82345 6086 82346 6150
rect 82410 6086 82411 6150
rect 82345 6085 82411 6086
rect 81428 5370 81748 5412
rect 81428 5134 81470 5370
rect 81706 5134 81748 5370
rect 81428 5092 81748 5134
rect 4145 4654 4211 4655
rect 4145 4590 4146 4654
rect 4210 4590 4211 4654
rect 4145 4589 4211 4590
rect 4513 4654 4579 4655
rect 4513 4590 4514 4654
rect 4578 4590 4579 4654
rect 4513 4589 4579 4590
rect 4145 4246 4211 4247
rect 4145 4182 4146 4246
rect 4210 4182 4211 4246
rect 4145 4181 4211 4182
rect 3777 3158 3843 3159
rect 3777 3094 3778 3158
rect 3842 3094 3843 3158
rect 3777 3093 3843 3094
rect 2878 2482 2886 2546
rect 2950 2482 2966 2546
rect 3030 2482 3046 2546
rect 3110 2482 3126 2546
rect 3190 2482 3198 2546
rect 2878 1922 3198 2482
rect 4148 711 4208 4181
rect 4516 847 4576 4589
rect 39105 3022 39171 3023
rect 39105 2958 39106 3022
rect 39170 2958 39171 3022
rect 39105 2957 39171 2958
rect 42969 3022 43035 3023
rect 42969 2958 42970 3022
rect 43034 2958 43035 3022
rect 42969 2957 43035 2958
rect 13529 2886 13595 2887
rect 13529 2822 13530 2886
rect 13594 2884 13595 2886
rect 19785 2886 19851 2887
rect 13594 2824 14102 2884
rect 13594 2822 13595 2824
rect 13529 2821 13595 2822
rect 19785 2822 19786 2886
rect 19850 2884 19851 2886
rect 21993 2886 22059 2887
rect 19850 2824 19942 2884
rect 19850 2822 19851 2824
rect 19785 2821 19851 2822
rect 21993 2822 21994 2886
rect 22058 2884 22059 2886
rect 24017 2886 24083 2887
rect 22058 2824 22278 2884
rect 22058 2822 22059 2824
rect 21993 2821 22059 2822
rect 24017 2822 24018 2886
rect 24082 2884 24083 2886
rect 25121 2886 25187 2887
rect 24082 2824 24614 2884
rect 24082 2822 24083 2824
rect 24017 2821 24083 2822
rect 25121 2822 25122 2886
rect 25186 2884 25187 2886
rect 27513 2886 27579 2887
rect 25186 2824 25782 2884
rect 25186 2822 25187 2824
rect 25121 2821 25187 2822
rect 27513 2822 27514 2886
rect 27578 2884 27579 2886
rect 31055 2886 31121 2887
rect 27578 2824 28118 2884
rect 27578 2822 27579 2824
rect 27513 2821 27579 2822
rect 31055 2822 31056 2886
rect 31120 2884 31121 2886
rect 33723 2886 33789 2887
rect 31120 2824 31622 2884
rect 31120 2822 31121 2824
rect 31055 2821 31121 2822
rect 33723 2822 33724 2886
rect 33788 2884 33789 2886
rect 36897 2886 36963 2887
rect 36897 2884 36898 2886
rect 33788 2824 33958 2884
rect 36418 2824 36898 2884
rect 33788 2822 33789 2824
rect 33723 2821 33789 2822
rect 36897 2822 36898 2824
rect 36962 2822 36963 2886
rect 38921 2886 38987 2887
rect 38921 2884 38922 2886
rect 36897 2821 36963 2822
rect 37084 2824 37462 2884
rect 38754 2824 38922 2884
rect 37084 2751 37144 2824
rect 38921 2822 38922 2824
rect 38986 2822 38987 2886
rect 39108 2884 39168 2957
rect 41313 2886 41379 2887
rect 41313 2884 41314 2886
rect 39108 2824 39798 2884
rect 41090 2824 41314 2884
rect 38921 2821 38987 2822
rect 41313 2822 41314 2824
rect 41378 2822 41379 2886
rect 42972 2884 43032 2957
rect 82532 2887 82592 96525
rect 83820 96319 83880 169829
rect 84185 167582 84251 167583
rect 84185 167518 84186 167582
rect 84250 167518 84251 167582
rect 84185 167517 84251 167518
rect 84188 97135 84248 167517
rect 84369 164998 84435 164999
rect 84369 164934 84370 164998
rect 84434 164934 84435 164998
rect 84369 164933 84435 164934
rect 84372 164455 84432 164933
rect 84553 164862 84619 164863
rect 84553 164798 84554 164862
rect 84618 164798 84619 164862
rect 84553 164797 84619 164798
rect 84369 164454 84435 164455
rect 84369 164390 84370 164454
rect 84434 164390 84435 164454
rect 84369 164389 84435 164390
rect 84556 164319 84616 164797
rect 84553 164318 84619 164319
rect 84553 164254 84554 164318
rect 84618 164254 84619 164318
rect 84553 164253 84619 164254
rect 84185 97134 84251 97135
rect 84185 97070 84186 97134
rect 84250 97070 84251 97134
rect 84185 97069 84251 97070
rect 84740 96863 84800 172005
rect 84878 171730 85198 172754
rect 84878 171666 84886 171730
rect 84950 171666 84966 171730
rect 85030 171666 85046 171730
rect 85110 171666 85126 171730
rect 85190 171666 85198 171730
rect 84878 170642 85198 171666
rect 84878 170578 84886 170642
rect 84950 170578 84966 170642
rect 85030 170578 85046 170642
rect 85110 170578 85126 170642
rect 85190 170578 85198 170642
rect 84878 169554 85198 170578
rect 84878 169490 84886 169554
rect 84950 169490 84966 169554
rect 85030 169490 85046 169554
rect 85110 169490 85126 169554
rect 85190 169490 85198 169554
rect 84878 168466 85198 169490
rect 84878 168402 84886 168466
rect 84950 168402 84966 168466
rect 85030 168402 85046 168466
rect 85110 168402 85126 168466
rect 85190 168402 85198 168466
rect 84878 167378 85198 168402
rect 84878 167314 84886 167378
rect 84950 167314 84966 167378
rect 85030 167314 85046 167378
rect 85110 167314 85126 167378
rect 85190 167314 85198 167378
rect 84878 166290 85198 167314
rect 84878 166226 84886 166290
rect 84950 166226 84966 166290
rect 85030 166226 85046 166290
rect 85110 166226 85126 166290
rect 85190 166226 85198 166290
rect 84878 165370 85198 166226
rect 84878 165202 84920 165370
rect 85156 165202 85198 165370
rect 84878 165138 84886 165202
rect 85190 165138 85198 165202
rect 84878 165134 84920 165138
rect 85156 165134 85198 165138
rect 84878 164114 85198 165134
rect 84878 164050 84886 164114
rect 84950 164050 84966 164114
rect 85030 164050 85046 164114
rect 85110 164050 85126 164114
rect 85190 164050 85198 164114
rect 84878 163026 85198 164050
rect 84878 162962 84886 163026
rect 84950 162962 84966 163026
rect 85030 162962 85046 163026
rect 85110 162962 85126 163026
rect 85190 162962 85198 163026
rect 84878 161938 85198 162962
rect 84878 161874 84886 161938
rect 84950 161874 84966 161938
rect 85030 161874 85046 161938
rect 85110 161874 85126 161938
rect 85190 161874 85198 161938
rect 84878 160850 85198 161874
rect 84878 160786 84886 160850
rect 84950 160786 84966 160850
rect 85030 160786 85046 160850
rect 85110 160786 85126 160850
rect 85190 160786 85198 160850
rect 84878 159762 85198 160786
rect 84878 159698 84886 159762
rect 84950 159698 84966 159762
rect 85030 159698 85046 159762
rect 85110 159698 85126 159762
rect 85190 159698 85198 159762
rect 84878 158674 85198 159698
rect 84878 158610 84886 158674
rect 84950 158610 84966 158674
rect 85030 158610 85046 158674
rect 85110 158610 85126 158674
rect 85190 158610 85198 158674
rect 84878 157586 85198 158610
rect 84878 157522 84886 157586
rect 84950 157522 84966 157586
rect 85030 157522 85046 157586
rect 85110 157522 85126 157586
rect 85190 157522 85198 157586
rect 84878 156498 85198 157522
rect 84878 156434 84886 156498
rect 84950 156434 84966 156498
rect 85030 156434 85046 156498
rect 85110 156434 85126 156498
rect 85190 156434 85198 156498
rect 84878 155410 85198 156434
rect 84878 155346 84886 155410
rect 84950 155370 84966 155410
rect 85030 155370 85046 155410
rect 85110 155370 85126 155410
rect 85190 155346 85198 155410
rect 84878 155134 84920 155346
rect 85156 155134 85198 155346
rect 84878 154322 85198 155134
rect 84878 154258 84886 154322
rect 84950 154258 84966 154322
rect 85030 154258 85046 154322
rect 85110 154258 85126 154322
rect 85190 154258 85198 154322
rect 84878 153234 85198 154258
rect 84878 153170 84886 153234
rect 84950 153170 84966 153234
rect 85030 153170 85046 153234
rect 85110 153170 85126 153234
rect 85190 153170 85198 153234
rect 84878 152146 85198 153170
rect 84878 152082 84886 152146
rect 84950 152082 84966 152146
rect 85030 152082 85046 152146
rect 85110 152082 85126 152146
rect 85190 152082 85198 152146
rect 84878 151058 85198 152082
rect 84878 150994 84886 151058
rect 84950 150994 84966 151058
rect 85030 150994 85046 151058
rect 85110 150994 85126 151058
rect 85190 150994 85198 151058
rect 84878 149970 85198 150994
rect 84878 149906 84886 149970
rect 84950 149906 84966 149970
rect 85030 149906 85046 149970
rect 85110 149906 85126 149970
rect 85190 149906 85198 149970
rect 84878 148882 85198 149906
rect 84878 148818 84886 148882
rect 84950 148818 84966 148882
rect 85030 148818 85046 148882
rect 85110 148818 85126 148882
rect 85190 148818 85198 148882
rect 84878 147794 85198 148818
rect 84878 147730 84886 147794
rect 84950 147730 84966 147794
rect 85030 147730 85046 147794
rect 85110 147730 85126 147794
rect 85190 147730 85198 147794
rect 84878 146706 85198 147730
rect 84878 146642 84886 146706
rect 84950 146642 84966 146706
rect 85030 146642 85046 146706
rect 85110 146642 85126 146706
rect 85190 146642 85198 146706
rect 84878 145618 85198 146642
rect 84878 145554 84886 145618
rect 84950 145554 84966 145618
rect 85030 145554 85046 145618
rect 85110 145554 85126 145618
rect 85190 145554 85198 145618
rect 84878 145370 85198 145554
rect 84878 145134 84920 145370
rect 85156 145134 85198 145370
rect 84878 144530 85198 145134
rect 84878 144466 84886 144530
rect 84950 144466 84966 144530
rect 85030 144466 85046 144530
rect 85110 144466 85126 144530
rect 85190 144466 85198 144530
rect 84878 143442 85198 144466
rect 84878 143378 84886 143442
rect 84950 143378 84966 143442
rect 85030 143378 85046 143442
rect 85110 143378 85126 143442
rect 85190 143378 85198 143442
rect 84878 142354 85198 143378
rect 84878 142290 84886 142354
rect 84950 142290 84966 142354
rect 85030 142290 85046 142354
rect 85110 142290 85126 142354
rect 85190 142290 85198 142354
rect 84878 141266 85198 142290
rect 84878 141202 84886 141266
rect 84950 141202 84966 141266
rect 85030 141202 85046 141266
rect 85110 141202 85126 141266
rect 85190 141202 85198 141266
rect 84878 140178 85198 141202
rect 84878 140114 84886 140178
rect 84950 140114 84966 140178
rect 85030 140114 85046 140178
rect 85110 140114 85126 140178
rect 85190 140114 85198 140178
rect 84878 139090 85198 140114
rect 84878 139026 84886 139090
rect 84950 139026 84966 139090
rect 85030 139026 85046 139090
rect 85110 139026 85126 139090
rect 85190 139026 85198 139090
rect 84878 138002 85198 139026
rect 84878 137938 84886 138002
rect 84950 137938 84966 138002
rect 85030 137938 85046 138002
rect 85110 137938 85126 138002
rect 85190 137938 85198 138002
rect 84878 136914 85198 137938
rect 84878 136850 84886 136914
rect 84950 136850 84966 136914
rect 85030 136850 85046 136914
rect 85110 136850 85126 136914
rect 85190 136850 85198 136914
rect 84878 135826 85198 136850
rect 84878 135762 84886 135826
rect 84950 135762 84966 135826
rect 85030 135762 85046 135826
rect 85110 135762 85126 135826
rect 85190 135762 85198 135826
rect 84878 135370 85198 135762
rect 84878 135134 84920 135370
rect 85156 135134 85198 135370
rect 84878 134738 85198 135134
rect 84878 134674 84886 134738
rect 84950 134674 84966 134738
rect 85030 134674 85046 134738
rect 85110 134674 85126 134738
rect 85190 134674 85198 134738
rect 84878 133650 85198 134674
rect 84878 133586 84886 133650
rect 84950 133586 84966 133650
rect 85030 133586 85046 133650
rect 85110 133586 85126 133650
rect 85190 133586 85198 133650
rect 84878 132562 85198 133586
rect 84878 132498 84886 132562
rect 84950 132498 84966 132562
rect 85030 132498 85046 132562
rect 85110 132498 85126 132562
rect 85190 132498 85198 132562
rect 84878 131474 85198 132498
rect 84878 131410 84886 131474
rect 84950 131410 84966 131474
rect 85030 131410 85046 131474
rect 85110 131410 85126 131474
rect 85190 131410 85198 131474
rect 84878 130386 85198 131410
rect 84878 130322 84886 130386
rect 84950 130322 84966 130386
rect 85030 130322 85046 130386
rect 85110 130322 85126 130386
rect 85190 130322 85198 130386
rect 84878 129298 85198 130322
rect 84878 129234 84886 129298
rect 84950 129234 84966 129298
rect 85030 129234 85046 129298
rect 85110 129234 85126 129298
rect 85190 129234 85198 129298
rect 84878 128210 85198 129234
rect 84878 128146 84886 128210
rect 84950 128146 84966 128210
rect 85030 128146 85046 128210
rect 85110 128146 85126 128210
rect 85190 128146 85198 128210
rect 84878 127122 85198 128146
rect 84878 127058 84886 127122
rect 84950 127058 84966 127122
rect 85030 127058 85046 127122
rect 85110 127058 85126 127122
rect 85190 127058 85198 127122
rect 84878 126034 85198 127058
rect 84878 125970 84886 126034
rect 84950 125970 84966 126034
rect 85030 125970 85046 126034
rect 85110 125970 85126 126034
rect 85190 125970 85198 126034
rect 84878 125370 85198 125970
rect 84878 125134 84920 125370
rect 85156 125134 85198 125370
rect 84878 124946 85198 125134
rect 84878 124882 84886 124946
rect 84950 124882 84966 124946
rect 85030 124882 85046 124946
rect 85110 124882 85126 124946
rect 85190 124882 85198 124946
rect 84878 123858 85198 124882
rect 84878 123794 84886 123858
rect 84950 123794 84966 123858
rect 85030 123794 85046 123858
rect 85110 123794 85126 123858
rect 85190 123794 85198 123858
rect 84878 122770 85198 123794
rect 84878 122706 84886 122770
rect 84950 122706 84966 122770
rect 85030 122706 85046 122770
rect 85110 122706 85126 122770
rect 85190 122706 85198 122770
rect 84878 121682 85198 122706
rect 84878 121618 84886 121682
rect 84950 121618 84966 121682
rect 85030 121618 85046 121682
rect 85110 121618 85126 121682
rect 85190 121618 85198 121682
rect 84878 120594 85198 121618
rect 84878 120530 84886 120594
rect 84950 120530 84966 120594
rect 85030 120530 85046 120594
rect 85110 120530 85126 120594
rect 85190 120530 85198 120594
rect 84878 119506 85198 120530
rect 84878 119442 84886 119506
rect 84950 119442 84966 119506
rect 85030 119442 85046 119506
rect 85110 119442 85126 119506
rect 85190 119442 85198 119506
rect 84878 118418 85198 119442
rect 84878 118354 84886 118418
rect 84950 118354 84966 118418
rect 85030 118354 85046 118418
rect 85110 118354 85126 118418
rect 85190 118354 85198 118418
rect 84878 117330 85198 118354
rect 84878 117266 84886 117330
rect 84950 117266 84966 117330
rect 85030 117266 85046 117330
rect 85110 117266 85126 117330
rect 85190 117266 85198 117330
rect 84878 116242 85198 117266
rect 84878 116178 84886 116242
rect 84950 116178 84966 116242
rect 85030 116178 85046 116242
rect 85110 116178 85126 116242
rect 85190 116178 85198 116242
rect 84878 115370 85198 116178
rect 84878 115154 84920 115370
rect 85156 115154 85198 115370
rect 84878 115090 84886 115154
rect 84950 115090 84966 115134
rect 85030 115090 85046 115134
rect 85110 115090 85126 115134
rect 85190 115090 85198 115154
rect 84878 114066 85198 115090
rect 84878 114002 84886 114066
rect 84950 114002 84966 114066
rect 85030 114002 85046 114066
rect 85110 114002 85126 114066
rect 85190 114002 85198 114066
rect 84878 112978 85198 114002
rect 84878 112914 84886 112978
rect 84950 112914 84966 112978
rect 85030 112914 85046 112978
rect 85110 112914 85126 112978
rect 85190 112914 85198 112978
rect 84878 111890 85198 112914
rect 84878 111826 84886 111890
rect 84950 111826 84966 111890
rect 85030 111826 85046 111890
rect 85110 111826 85126 111890
rect 85190 111826 85198 111890
rect 84878 110802 85198 111826
rect 84878 110738 84886 110802
rect 84950 110738 84966 110802
rect 85030 110738 85046 110802
rect 85110 110738 85126 110802
rect 85190 110738 85198 110802
rect 84878 109714 85198 110738
rect 84878 109650 84886 109714
rect 84950 109650 84966 109714
rect 85030 109650 85046 109714
rect 85110 109650 85126 109714
rect 85190 109650 85198 109714
rect 84878 108626 85198 109650
rect 84878 108562 84886 108626
rect 84950 108562 84966 108626
rect 85030 108562 85046 108626
rect 85110 108562 85126 108626
rect 85190 108562 85198 108626
rect 84878 107538 85198 108562
rect 84878 107474 84886 107538
rect 84950 107474 84966 107538
rect 85030 107474 85046 107538
rect 85110 107474 85126 107538
rect 85190 107474 85198 107538
rect 84878 106450 85198 107474
rect 84878 106386 84886 106450
rect 84950 106386 84966 106450
rect 85030 106386 85046 106450
rect 85110 106386 85126 106450
rect 85190 106386 85198 106450
rect 84878 105370 85198 106386
rect 84878 105362 84920 105370
rect 85156 105362 85198 105370
rect 84878 105298 84886 105362
rect 85190 105298 85198 105362
rect 84878 105134 84920 105298
rect 85156 105134 85198 105298
rect 84878 104274 85198 105134
rect 84878 104210 84886 104274
rect 84950 104210 84966 104274
rect 85030 104210 85046 104274
rect 85110 104210 85126 104274
rect 85190 104210 85198 104274
rect 84878 103186 85198 104210
rect 84878 103122 84886 103186
rect 84950 103122 84966 103186
rect 85030 103122 85046 103186
rect 85110 103122 85126 103186
rect 85190 103122 85198 103186
rect 84878 102098 85198 103122
rect 84878 102034 84886 102098
rect 84950 102034 84966 102098
rect 85030 102034 85046 102098
rect 85110 102034 85126 102098
rect 85190 102034 85198 102098
rect 84878 101010 85198 102034
rect 84878 100946 84886 101010
rect 84950 100946 84966 101010
rect 85030 100946 85046 101010
rect 85110 100946 85126 101010
rect 85190 100946 85198 101010
rect 84878 99922 85198 100946
rect 84878 99858 84886 99922
rect 84950 99858 84966 99922
rect 85030 99858 85046 99922
rect 85110 99858 85126 99922
rect 85190 99858 85198 99922
rect 84878 98834 85198 99858
rect 84878 98770 84886 98834
rect 84950 98770 84966 98834
rect 85030 98770 85046 98834
rect 85110 98770 85126 98834
rect 85190 98770 85198 98834
rect 84878 97746 85198 98770
rect 84878 97682 84886 97746
rect 84950 97682 84966 97746
rect 85030 97682 85046 97746
rect 85110 97682 85126 97746
rect 85190 97682 85198 97746
rect 84737 96862 84803 96863
rect 84737 96798 84738 96862
rect 84802 96798 84803 96862
rect 84737 96797 84803 96798
rect 84878 96658 85198 97682
rect 84878 96594 84886 96658
rect 84950 96594 84966 96658
rect 85030 96594 85046 96658
rect 85110 96594 85126 96658
rect 85190 96594 85198 96658
rect 83817 96318 83883 96319
rect 83817 96254 83818 96318
rect 83882 96254 83883 96318
rect 83817 96253 83883 96254
rect 84878 95570 85198 96594
rect 84878 95506 84886 95570
rect 84950 95506 84966 95570
rect 85030 95506 85046 95570
rect 85110 95506 85126 95570
rect 85190 95506 85198 95570
rect 84878 95370 85198 95506
rect 82878 94354 83198 95250
rect 84878 95134 84920 95370
rect 85156 95134 85198 95370
rect 83817 94686 83883 94687
rect 83817 94622 83818 94686
rect 83882 94622 83883 94686
rect 83817 94621 83883 94622
rect 82713 94006 82779 94007
rect 82713 93942 82714 94006
rect 82778 93942 82779 94006
rect 82713 93941 82779 93942
rect 44257 2886 44323 2887
rect 42972 2824 43302 2884
rect 41313 2821 41379 2822
rect 44257 2822 44258 2886
rect 44322 2884 44323 2886
rect 82529 2886 82595 2887
rect 44322 2824 44470 2884
rect 45364 2824 45638 2884
rect 48860 2824 49142 2884
rect 50148 2824 50310 2884
rect 53644 2824 53814 2884
rect 44322 2822 44323 2824
rect 44257 2821 44323 2822
rect 45364 2751 45424 2824
rect 37081 2750 37147 2751
rect 37081 2686 37082 2750
rect 37146 2686 37147 2750
rect 37081 2685 37147 2686
rect 45361 2750 45427 2751
rect 45361 2686 45362 2750
rect 45426 2686 45427 2750
rect 45361 2685 45427 2686
rect 48860 2615 48920 2824
rect 50148 2615 50208 2824
rect 53644 2615 53704 2824
rect 82529 2822 82530 2886
rect 82594 2822 82595 2886
rect 82529 2821 82595 2822
rect 48857 2614 48923 2615
rect 48857 2550 48858 2614
rect 48922 2550 48923 2614
rect 48857 2549 48923 2550
rect 50145 2614 50211 2615
rect 50145 2550 50146 2614
rect 50210 2550 50211 2614
rect 50145 2549 50211 2550
rect 53641 2614 53707 2615
rect 53641 2550 53642 2614
rect 53706 2550 53707 2614
rect 53641 2549 53707 2550
rect 12244 2484 12934 2544
rect 15740 2484 16438 2544
rect 18316 2484 18774 2544
rect 20066 2484 20768 2544
rect 23570 2484 24264 2544
rect 8737 1663 8797 2174
rect 8734 1662 8800 1663
rect 8734 1598 8735 1662
rect 8799 1598 8800 1662
rect 8734 1597 8800 1598
rect 11736 1524 11796 2174
rect 11692 1464 11796 1524
rect 11692 983 11752 1464
rect 12244 983 12304 2484
rect 15240 1524 15300 2174
rect 15188 1464 15300 1524
rect 15188 983 15248 1464
rect 11689 982 11755 983
rect 11689 918 11690 982
rect 11754 918 11755 982
rect 11689 917 11755 918
rect 12241 982 12307 983
rect 12241 918 12242 982
rect 12306 918 12307 982
rect 12241 917 12307 918
rect 15185 982 15251 983
rect 15185 918 15186 982
rect 15250 918 15251 982
rect 15185 917 15251 918
rect 4513 846 4579 847
rect 4513 782 4514 846
rect 4578 782 4579 846
rect 4513 781 4579 782
rect 15740 711 15800 2484
rect 18316 2343 18376 2484
rect 18313 2342 18379 2343
rect 18313 2278 18314 2342
rect 18378 2278 18379 2342
rect 18313 2277 18379 2278
rect 17576 1524 17636 2174
rect 17700 1524 17760 2174
rect 17576 1464 17640 1524
rect 17700 1464 17824 1524
rect 17580 983 17640 1464
rect 17764 983 17824 1464
rect 18868 983 18928 2174
rect 17577 982 17643 983
rect 17577 918 17578 982
rect 17642 918 17643 982
rect 17577 917 17643 918
rect 17761 982 17827 983
rect 17761 918 17762 982
rect 17826 918 17827 982
rect 17761 917 17827 918
rect 18865 982 18931 983
rect 18865 918 18866 982
rect 18930 918 18931 982
rect 18865 917 18931 918
rect 20708 711 20768 2484
rect 21080 1524 21140 2174
rect 21076 1464 21140 1524
rect 21204 1524 21264 2174
rect 22372 1663 22432 2174
rect 22369 1662 22435 1663
rect 22369 1598 22370 1662
rect 22434 1598 22435 1662
rect 22369 1597 22435 1598
rect 23416 1524 23476 2174
rect 21204 1464 21320 1524
rect 23416 1464 23528 1524
rect 21076 983 21136 1464
rect 21260 983 21320 1464
rect 23468 983 23528 1464
rect 24204 983 24264 2484
rect 26412 2484 26950 2544
rect 29908 2484 30454 2544
rect 30578 2484 31072 2544
rect 26412 2207 26472 2484
rect 26409 2206 26475 2207
rect 24708 1663 24768 2174
rect 24705 1662 24771 1663
rect 24705 1598 24706 1662
rect 24770 1598 24771 1662
rect 24705 1597 24771 1598
rect 25876 1524 25936 2174
rect 26409 2142 26410 2206
rect 26474 2142 26475 2206
rect 26409 2141 26475 2142
rect 25860 1464 25936 1524
rect 27044 1524 27104 2174
rect 28212 1524 28272 2174
rect 29256 1663 29316 2174
rect 29253 1662 29319 1663
rect 29253 1598 29254 1662
rect 29318 1598 29319 1662
rect 29253 1597 29319 1598
rect 29380 1524 29440 2174
rect 27044 1464 27208 1524
rect 28212 1464 28312 1524
rect 21073 982 21139 983
rect 21073 918 21074 982
rect 21138 918 21139 982
rect 21073 917 21139 918
rect 21257 982 21323 983
rect 21257 918 21258 982
rect 21322 918 21323 982
rect 21257 917 21323 918
rect 23465 982 23531 983
rect 23465 918 23466 982
rect 23530 918 23531 982
rect 23465 917 23531 918
rect 24201 982 24267 983
rect 24201 918 24202 982
rect 24266 918 24267 982
rect 24201 917 24267 918
rect 4145 710 4211 711
rect 4145 646 4146 710
rect 4210 646 4211 710
rect 4145 645 4211 646
rect 15737 710 15803 711
rect 15737 646 15738 710
rect 15802 646 15803 710
rect 15737 645 15803 646
rect 20705 710 20771 711
rect 20705 646 20706 710
rect 20770 646 20771 710
rect 20705 645 20771 646
rect 25860 167 25920 1464
rect 27148 1119 27208 1464
rect 27145 1118 27211 1119
rect 27145 1054 27146 1118
rect 27210 1054 27211 1118
rect 27145 1053 27211 1054
rect 28252 983 28312 1464
rect 29356 1464 29440 1524
rect 29356 983 29416 1464
rect 28249 982 28315 983
rect 28249 918 28250 982
rect 28314 918 28315 982
rect 28249 917 28315 918
rect 29353 982 29419 983
rect 29353 918 29354 982
rect 29418 918 29419 982
rect 29353 917 29419 918
rect 29908 711 29968 2484
rect 31012 983 31072 2484
rect 32484 2484 32790 2544
rect 34082 2484 34752 2544
rect 31716 1524 31776 2174
rect 31716 1464 31808 1524
rect 31748 983 31808 1464
rect 31009 982 31075 983
rect 31009 918 31010 982
rect 31074 918 31075 982
rect 31009 917 31075 918
rect 31745 982 31811 983
rect 31745 918 31746 982
rect 31810 918 31811 982
rect 31745 917 31811 918
rect 29905 710 29971 711
rect 29905 646 29906 710
rect 29970 646 29971 710
rect 29905 645 29971 646
rect 32484 575 32544 2484
rect 32884 1524 32944 2174
rect 32852 1464 32944 1524
rect 32852 983 32912 1464
rect 34692 983 34752 2484
rect 35060 2484 35126 2544
rect 37586 2484 38248 2544
rect 39922 2484 40088 2544
rect 34873 2342 34939 2343
rect 34873 2278 34874 2342
rect 34938 2278 34939 2342
rect 34873 2277 34939 2278
rect 34876 2204 34936 2277
rect 35060 2204 35120 2484
rect 34876 2144 35120 2204
rect 35220 1524 35280 2174
rect 36264 1663 36324 2174
rect 36261 1662 36327 1663
rect 36261 1598 36262 1662
rect 36326 1598 36327 1662
rect 36261 1597 36327 1598
rect 35220 1464 35304 1524
rect 35244 983 35304 1464
rect 38188 983 38248 2484
rect 38600 1524 38660 2174
rect 38556 1464 38660 1524
rect 32849 982 32915 983
rect 32849 918 32850 982
rect 32914 918 32915 982
rect 32849 917 32915 918
rect 34689 982 34755 983
rect 34689 918 34690 982
rect 34754 918 34755 982
rect 34689 917 34755 918
rect 35241 982 35307 983
rect 35241 918 35242 982
rect 35306 918 35307 982
rect 35241 917 35307 918
rect 38185 982 38251 983
rect 38185 918 38186 982
rect 38250 918 38251 982
rect 38185 917 38251 918
rect 32481 574 32547 575
rect 32481 510 32482 574
rect 32546 510 32547 574
rect 32481 509 32547 510
rect 38556 439 38616 1464
rect 40028 983 40088 2484
rect 41868 2484 42134 2544
rect 43426 2484 43952 2544
rect 44594 2484 45240 2544
rect 41868 2207 41928 2484
rect 41865 2206 41931 2207
rect 40936 1524 40996 2174
rect 41865 2142 41866 2206
rect 41930 2142 41931 2206
rect 41865 2141 41931 2142
rect 42228 1524 42288 2174
rect 40936 1464 41008 1524
rect 42228 1464 42296 1524
rect 40025 982 40091 983
rect 40025 918 40026 982
rect 40090 918 40091 982
rect 40025 917 40091 918
rect 40948 847 41008 1464
rect 42236 1391 42296 1464
rect 42233 1390 42299 1391
rect 42233 1326 42234 1390
rect 42298 1326 42299 1390
rect 42233 1325 42299 1326
rect 43892 983 43952 2484
rect 45180 2207 45240 2484
rect 46652 2484 46806 2544
rect 46930 2484 47632 2544
rect 49266 2484 49840 2544
rect 52770 2484 52968 2544
rect 53938 2484 54256 2544
rect 46652 2207 46712 2484
rect 47572 2207 47632 2484
rect 49780 2207 49840 2484
rect 45177 2206 45243 2207
rect 45177 2142 45178 2206
rect 45242 2142 45243 2206
rect 46649 2206 46715 2207
rect 45177 2141 45243 2142
rect 45732 983 45792 2174
rect 46649 2142 46650 2206
rect 46714 2142 46715 2206
rect 46649 2141 46715 2142
rect 47569 2206 47635 2207
rect 47569 2142 47570 2206
rect 47634 2142 47635 2206
rect 49777 2206 49843 2207
rect 47569 2141 47635 2142
rect 47944 1524 48004 2174
rect 47940 1464 48004 1524
rect 48068 1524 48128 2174
rect 49777 2142 49778 2206
rect 49842 2142 49843 2206
rect 49777 2141 49843 2142
rect 50404 1524 50464 2174
rect 51448 1524 51508 2174
rect 48068 1464 48184 1524
rect 47940 983 48000 1464
rect 43889 982 43955 983
rect 43889 918 43890 982
rect 43954 918 43955 982
rect 43889 917 43955 918
rect 45729 982 45795 983
rect 45729 918 45730 982
rect 45794 918 45795 982
rect 45729 917 45795 918
rect 47937 982 48003 983
rect 47937 918 47938 982
rect 48002 918 48003 982
rect 47937 917 48003 918
rect 48124 847 48184 1464
rect 50332 1464 50464 1524
rect 51436 1464 51508 1524
rect 51572 1524 51632 2174
rect 52616 1524 52676 2174
rect 51572 1464 51680 1524
rect 52616 1464 52784 1524
rect 40945 846 41011 847
rect 40945 782 40946 846
rect 41010 782 41011 846
rect 40945 781 41011 782
rect 48121 846 48187 847
rect 48121 782 48122 846
rect 48186 782 48187 846
rect 48121 781 48187 782
rect 38553 438 38619 439
rect 38553 374 38554 438
rect 38618 374 38619 438
rect 38553 373 38619 374
rect 50332 303 50392 1464
rect 51436 1391 51496 1464
rect 51433 1390 51499 1391
rect 51433 1326 51434 1390
rect 51498 1326 51499 1390
rect 51433 1325 51499 1326
rect 51620 711 51680 1464
rect 51617 710 51683 711
rect 51617 646 51618 710
rect 51682 646 51683 710
rect 51617 645 51683 646
rect 52724 575 52784 1464
rect 52721 574 52787 575
rect 52721 510 52722 574
rect 52786 510 52787 574
rect 52721 509 52787 510
rect 52908 439 52968 2484
rect 54196 2343 54256 2484
rect 82716 2343 82776 93941
rect 83265 59326 83331 59327
rect 83265 59262 83266 59326
rect 83330 59262 83331 59326
rect 83265 59261 83331 59262
rect 82897 15534 82963 15535
rect 82897 15470 82898 15534
rect 82962 15470 82963 15534
rect 82897 15469 82963 15470
rect 82900 3839 82960 15469
rect 82897 3838 82963 3839
rect 82897 3774 82898 3838
rect 82962 3774 82963 3838
rect 82897 3773 82963 3774
rect 54193 2342 54259 2343
rect 54193 2278 54194 2342
rect 54258 2278 54259 2342
rect 54193 2277 54259 2278
rect 82713 2342 82779 2343
rect 82713 2278 82714 2342
rect 82778 2278 82779 2342
rect 82713 2277 82779 2278
rect 83268 711 83328 59261
rect 83449 55246 83515 55247
rect 83449 55182 83450 55246
rect 83514 55182 83515 55246
rect 83449 55181 83515 55182
rect 83265 710 83331 711
rect 83265 646 83266 710
rect 83330 646 83331 710
rect 83265 645 83331 646
rect 83452 439 83512 55181
rect 83633 33894 83699 33895
rect 83633 33830 83634 33894
rect 83698 33830 83699 33894
rect 83633 33829 83699 33830
rect 83636 1119 83696 33829
rect 83820 4111 83880 94621
rect 84878 94482 85198 95134
rect 84878 94418 84886 94482
rect 84950 94418 84966 94482
rect 85030 94418 85046 94482
rect 85110 94418 85126 94482
rect 85190 94418 85198 94482
rect 84878 93394 85198 94418
rect 84878 93330 84886 93394
rect 84950 93330 84966 93394
rect 85030 93330 85046 93394
rect 85110 93330 85126 93394
rect 85190 93330 85198 93394
rect 84878 92306 85198 93330
rect 84878 92242 84886 92306
rect 84950 92242 84966 92306
rect 85030 92242 85046 92306
rect 85110 92242 85126 92306
rect 85190 92242 85198 92306
rect 84878 91218 85198 92242
rect 84878 91154 84886 91218
rect 84950 91154 84966 91218
rect 85030 91154 85046 91218
rect 85110 91154 85126 91218
rect 85190 91154 85198 91218
rect 84878 90130 85198 91154
rect 84878 90066 84886 90130
rect 84950 90066 84966 90130
rect 85030 90066 85046 90130
rect 85110 90066 85126 90130
rect 85190 90066 85198 90130
rect 84878 89042 85198 90066
rect 84878 88978 84886 89042
rect 84950 88978 84966 89042
rect 85030 88978 85046 89042
rect 85110 88978 85126 89042
rect 85190 88978 85198 89042
rect 84878 87954 85198 88978
rect 84878 87890 84886 87954
rect 84950 87890 84966 87954
rect 85030 87890 85046 87954
rect 85110 87890 85126 87954
rect 85190 87890 85198 87954
rect 84878 86866 85198 87890
rect 84878 86802 84886 86866
rect 84950 86802 84966 86866
rect 85030 86802 85046 86866
rect 85110 86802 85126 86866
rect 85190 86802 85198 86866
rect 84878 85778 85198 86802
rect 84878 85714 84886 85778
rect 84950 85714 84966 85778
rect 85030 85714 85046 85778
rect 85110 85714 85126 85778
rect 85190 85714 85198 85778
rect 84878 85370 85198 85714
rect 84878 85134 84920 85370
rect 85156 85134 85198 85370
rect 84878 84690 85198 85134
rect 84878 84626 84886 84690
rect 84950 84626 84966 84690
rect 85030 84626 85046 84690
rect 85110 84626 85126 84690
rect 85190 84626 85198 84690
rect 84878 83602 85198 84626
rect 84878 83538 84886 83602
rect 84950 83538 84966 83602
rect 85030 83538 85046 83602
rect 85110 83538 85126 83602
rect 85190 83538 85198 83602
rect 84878 82514 85198 83538
rect 84878 82450 84886 82514
rect 84950 82450 84966 82514
rect 85030 82450 85046 82514
rect 85110 82450 85126 82514
rect 85190 82450 85198 82514
rect 84878 81426 85198 82450
rect 84878 81362 84886 81426
rect 84950 81362 84966 81426
rect 85030 81362 85046 81426
rect 85110 81362 85126 81426
rect 85190 81362 85198 81426
rect 84878 80338 85198 81362
rect 84878 80274 84886 80338
rect 84950 80274 84966 80338
rect 85030 80274 85046 80338
rect 85110 80274 85126 80338
rect 85190 80274 85198 80338
rect 84878 79250 85198 80274
rect 84878 79186 84886 79250
rect 84950 79186 84966 79250
rect 85030 79186 85046 79250
rect 85110 79186 85126 79250
rect 85190 79186 85198 79250
rect 84878 78162 85198 79186
rect 84878 78098 84886 78162
rect 84950 78098 84966 78162
rect 85030 78098 85046 78162
rect 85110 78098 85126 78162
rect 85190 78098 85198 78162
rect 84878 77074 85198 78098
rect 84878 77010 84886 77074
rect 84950 77010 84966 77074
rect 85030 77010 85046 77074
rect 85110 77010 85126 77074
rect 85190 77010 85198 77074
rect 84878 75986 85198 77010
rect 84878 75922 84886 75986
rect 84950 75922 84966 75986
rect 85030 75922 85046 75986
rect 85110 75922 85126 75986
rect 85190 75922 85198 75986
rect 84878 75370 85198 75922
rect 84878 75134 84920 75370
rect 85156 75134 85198 75370
rect 84878 74898 85198 75134
rect 84878 74834 84886 74898
rect 84950 74834 84966 74898
rect 85030 74834 85046 74898
rect 85110 74834 85126 74898
rect 85190 74834 85198 74898
rect 84878 73810 85198 74834
rect 84878 73746 84886 73810
rect 84950 73746 84966 73810
rect 85030 73746 85046 73810
rect 85110 73746 85126 73810
rect 85190 73746 85198 73810
rect 84878 72722 85198 73746
rect 84878 72658 84886 72722
rect 84950 72658 84966 72722
rect 85030 72658 85046 72722
rect 85110 72658 85126 72722
rect 85190 72658 85198 72722
rect 84878 71634 85198 72658
rect 84878 71570 84886 71634
rect 84950 71570 84966 71634
rect 85030 71570 85046 71634
rect 85110 71570 85126 71634
rect 85190 71570 85198 71634
rect 84878 70546 85198 71570
rect 84878 70482 84886 70546
rect 84950 70482 84966 70546
rect 85030 70482 85046 70546
rect 85110 70482 85126 70546
rect 85190 70482 85198 70546
rect 84878 69458 85198 70482
rect 84878 69394 84886 69458
rect 84950 69394 84966 69458
rect 85030 69394 85046 69458
rect 85110 69394 85126 69458
rect 85190 69394 85198 69458
rect 84878 68370 85198 69394
rect 84878 68306 84886 68370
rect 84950 68306 84966 68370
rect 85030 68306 85046 68370
rect 85110 68306 85126 68370
rect 85190 68306 85198 68370
rect 84878 67282 85198 68306
rect 84878 67218 84886 67282
rect 84950 67218 84966 67282
rect 85030 67218 85046 67282
rect 85110 67218 85126 67282
rect 85190 67218 85198 67282
rect 84878 66194 85198 67218
rect 84878 66130 84886 66194
rect 84950 66130 84966 66194
rect 85030 66130 85046 66194
rect 85110 66130 85126 66194
rect 85190 66130 85198 66194
rect 84878 65370 85198 66130
rect 84878 65134 84920 65370
rect 85156 65134 85198 65370
rect 84878 65106 85198 65134
rect 84878 65042 84886 65106
rect 84950 65042 84966 65106
rect 85030 65042 85046 65106
rect 85110 65042 85126 65106
rect 85190 65042 85198 65106
rect 84878 64018 85198 65042
rect 84878 63954 84886 64018
rect 84950 63954 84966 64018
rect 85030 63954 85046 64018
rect 85110 63954 85126 64018
rect 85190 63954 85198 64018
rect 84878 62930 85198 63954
rect 84878 62866 84886 62930
rect 84950 62866 84966 62930
rect 85030 62866 85046 62930
rect 85110 62866 85126 62930
rect 85190 62866 85198 62930
rect 84878 61842 85198 62866
rect 84878 61778 84886 61842
rect 84950 61778 84966 61842
rect 85030 61778 85046 61842
rect 85110 61778 85126 61842
rect 85190 61778 85198 61842
rect 84878 60754 85198 61778
rect 84878 60690 84886 60754
rect 84950 60690 84966 60754
rect 85030 60690 85046 60754
rect 85110 60690 85126 60754
rect 85190 60690 85198 60754
rect 84878 59666 85198 60690
rect 84878 59602 84886 59666
rect 84950 59602 84966 59666
rect 85030 59602 85046 59666
rect 85110 59602 85126 59666
rect 85190 59602 85198 59666
rect 84878 58578 85198 59602
rect 84878 58514 84886 58578
rect 84950 58514 84966 58578
rect 85030 58514 85046 58578
rect 85110 58514 85126 58578
rect 85190 58514 85198 58578
rect 84553 57830 84619 57831
rect 84553 57766 84554 57830
rect 84618 57766 84619 57830
rect 84553 57765 84619 57766
rect 84369 32806 84435 32807
rect 84369 32742 84370 32806
rect 84434 32742 84435 32806
rect 84369 32741 84435 32742
rect 84001 24238 84067 24239
rect 84001 24174 84002 24238
rect 84066 24174 84067 24238
rect 84001 24173 84067 24174
rect 84004 19615 84064 24173
rect 84185 21926 84251 21927
rect 84185 21862 84186 21926
rect 84250 21862 84251 21926
rect 84185 21861 84251 21862
rect 84001 19614 84067 19615
rect 84001 19550 84002 19614
rect 84066 19550 84067 19614
rect 84001 19549 84067 19550
rect 83817 4110 83883 4111
rect 83817 4046 83818 4110
rect 83882 4046 83883 4110
rect 83817 4045 83883 4046
rect 84001 2478 84067 2479
rect 84001 2414 84002 2478
rect 84066 2414 84067 2478
rect 84001 2413 84067 2414
rect 84004 2207 84064 2413
rect 84001 2206 84067 2207
rect 84001 2142 84002 2206
rect 84066 2142 84067 2206
rect 84001 2141 84067 2142
rect 84188 1663 84248 21861
rect 84372 3159 84432 32741
rect 84556 3295 84616 57765
rect 84878 57490 85198 58514
rect 84878 57426 84886 57490
rect 84950 57426 84966 57490
rect 85030 57426 85046 57490
rect 85110 57426 85126 57490
rect 85190 57426 85198 57490
rect 84878 56402 85198 57426
rect 84878 56338 84886 56402
rect 84950 56338 84966 56402
rect 85030 56338 85046 56402
rect 85110 56338 85126 56402
rect 85190 56338 85198 56402
rect 84878 55370 85198 56338
rect 84878 55314 84920 55370
rect 85156 55314 85198 55370
rect 84878 55250 84886 55314
rect 85190 55250 85198 55314
rect 84878 55134 84920 55250
rect 85156 55134 85198 55250
rect 84878 54226 85198 55134
rect 84878 54162 84886 54226
rect 84950 54162 84966 54226
rect 85030 54162 85046 54226
rect 85110 54162 85126 54226
rect 85190 54162 85198 54226
rect 84878 53138 85198 54162
rect 84878 53074 84886 53138
rect 84950 53074 84966 53138
rect 85030 53074 85046 53138
rect 85110 53074 85126 53138
rect 85190 53074 85198 53138
rect 84878 52050 85198 53074
rect 84878 51986 84886 52050
rect 84950 51986 84966 52050
rect 85030 51986 85046 52050
rect 85110 51986 85126 52050
rect 85190 51986 85198 52050
rect 84878 50962 85198 51986
rect 84878 50898 84886 50962
rect 84950 50898 84966 50962
rect 85030 50898 85046 50962
rect 85110 50898 85126 50962
rect 85190 50898 85198 50962
rect 84878 49874 85198 50898
rect 84878 49810 84886 49874
rect 84950 49810 84966 49874
rect 85030 49810 85046 49874
rect 85110 49810 85126 49874
rect 85190 49810 85198 49874
rect 84878 48786 85198 49810
rect 84878 48722 84886 48786
rect 84950 48722 84966 48786
rect 85030 48722 85046 48786
rect 85110 48722 85126 48786
rect 85190 48722 85198 48786
rect 84878 47698 85198 48722
rect 84878 47634 84886 47698
rect 84950 47634 84966 47698
rect 85030 47634 85046 47698
rect 85110 47634 85126 47698
rect 85190 47634 85198 47698
rect 84878 46610 85198 47634
rect 84878 46546 84886 46610
rect 84950 46546 84966 46610
rect 85030 46546 85046 46610
rect 85110 46546 85126 46610
rect 85190 46546 85198 46610
rect 84878 45522 85198 46546
rect 84878 45458 84886 45522
rect 84950 45458 84966 45522
rect 85030 45458 85046 45522
rect 85110 45458 85126 45522
rect 85190 45458 85198 45522
rect 84878 45370 85198 45458
rect 84878 45134 84920 45370
rect 85156 45134 85198 45370
rect 84878 44434 85198 45134
rect 84878 44370 84886 44434
rect 84950 44370 84966 44434
rect 85030 44370 85046 44434
rect 85110 44370 85126 44434
rect 85190 44370 85198 44434
rect 84878 43346 85198 44370
rect 84878 43282 84886 43346
rect 84950 43282 84966 43346
rect 85030 43282 85046 43346
rect 85110 43282 85126 43346
rect 85190 43282 85198 43346
rect 84878 42258 85198 43282
rect 84878 42194 84886 42258
rect 84950 42194 84966 42258
rect 85030 42194 85046 42258
rect 85110 42194 85126 42258
rect 85190 42194 85198 42258
rect 84878 41170 85198 42194
rect 84878 41106 84886 41170
rect 84950 41106 84966 41170
rect 85030 41106 85046 41170
rect 85110 41106 85126 41170
rect 85190 41106 85198 41170
rect 84878 40082 85198 41106
rect 84878 40018 84886 40082
rect 84950 40018 84966 40082
rect 85030 40018 85046 40082
rect 85110 40018 85126 40082
rect 85190 40018 85198 40082
rect 84878 38994 85198 40018
rect 84878 38930 84886 38994
rect 84950 38930 84966 38994
rect 85030 38930 85046 38994
rect 85110 38930 85126 38994
rect 85190 38930 85198 38994
rect 84878 37906 85198 38930
rect 84878 37842 84886 37906
rect 84950 37842 84966 37906
rect 85030 37842 85046 37906
rect 85110 37842 85126 37906
rect 85190 37842 85198 37906
rect 84878 36818 85198 37842
rect 84878 36754 84886 36818
rect 84950 36754 84966 36818
rect 85030 36754 85046 36818
rect 85110 36754 85126 36818
rect 85190 36754 85198 36818
rect 84878 35730 85198 36754
rect 84878 35666 84886 35730
rect 84950 35666 84966 35730
rect 85030 35666 85046 35730
rect 85110 35666 85126 35730
rect 85190 35666 85198 35730
rect 84878 35370 85198 35666
rect 84878 35134 84920 35370
rect 85156 35134 85198 35370
rect 84737 34982 84803 34983
rect 84737 34918 84738 34982
rect 84802 34918 84803 34982
rect 84737 34917 84803 34918
rect 84553 3294 84619 3295
rect 84553 3230 84554 3294
rect 84618 3230 84619 3294
rect 84553 3229 84619 3230
rect 84369 3158 84435 3159
rect 84369 3094 84370 3158
rect 84434 3094 84435 3158
rect 84369 3093 84435 3094
rect 84185 1662 84251 1663
rect 84185 1598 84186 1662
rect 84250 1598 84251 1662
rect 84185 1597 84251 1598
rect 84740 1391 84800 34917
rect 84878 34642 85198 35134
rect 84878 34578 84886 34642
rect 84950 34578 84966 34642
rect 85030 34578 85046 34642
rect 85110 34578 85126 34642
rect 85190 34578 85198 34642
rect 84878 33554 85198 34578
rect 84878 33490 84886 33554
rect 84950 33490 84966 33554
rect 85030 33490 85046 33554
rect 85110 33490 85126 33554
rect 85190 33490 85198 33554
rect 84878 32466 85198 33490
rect 84878 32402 84886 32466
rect 84950 32402 84966 32466
rect 85030 32402 85046 32466
rect 85110 32402 85126 32466
rect 85190 32402 85198 32466
rect 84878 31378 85198 32402
rect 84878 31314 84886 31378
rect 84950 31314 84966 31378
rect 85030 31314 85046 31378
rect 85110 31314 85126 31378
rect 85190 31314 85198 31378
rect 84878 30290 85198 31314
rect 84878 30226 84886 30290
rect 84950 30226 84966 30290
rect 85030 30226 85046 30290
rect 85110 30226 85126 30290
rect 85190 30226 85198 30290
rect 84878 29202 85198 30226
rect 86878 187506 87198 187522
rect 86878 187442 86886 187506
rect 86950 187442 86966 187506
rect 87030 187442 87046 187506
rect 87110 187442 87126 187506
rect 87190 187442 87198 187506
rect 86878 186418 87198 187442
rect 86878 186354 86886 186418
rect 86950 186354 86966 186418
rect 87030 186354 87046 186418
rect 87110 186354 87126 186418
rect 87190 186354 87198 186418
rect 86878 185330 87198 186354
rect 86878 185266 86886 185330
rect 86950 185266 86966 185330
rect 87030 185266 87046 185330
rect 87110 185266 87126 185330
rect 87190 185266 87198 185330
rect 86878 184242 87198 185266
rect 86878 184178 86886 184242
rect 86950 184178 86966 184242
rect 87030 184178 87046 184242
rect 87110 184178 87126 184242
rect 87190 184178 87198 184242
rect 86878 183154 87198 184178
rect 86878 183090 86886 183154
rect 86950 183090 86966 183154
rect 87030 183090 87046 183154
rect 87110 183090 87126 183154
rect 87190 183090 87198 183154
rect 86878 182066 87198 183090
rect 86878 182002 86886 182066
rect 86950 182002 86966 182066
rect 87030 182002 87046 182066
rect 87110 182002 87126 182066
rect 87190 182002 87198 182066
rect 86878 180978 87198 182002
rect 86878 180914 86886 180978
rect 86950 180914 86966 180978
rect 87030 180914 87046 180978
rect 87110 180914 87126 180978
rect 87190 180914 87198 180978
rect 86878 180370 87198 180914
rect 86878 180134 86920 180370
rect 87156 180134 87198 180370
rect 86878 179890 87198 180134
rect 86878 179826 86886 179890
rect 86950 179826 86966 179890
rect 87030 179826 87046 179890
rect 87110 179826 87126 179890
rect 87190 179826 87198 179890
rect 86878 178802 87198 179826
rect 86878 178738 86886 178802
rect 86950 178738 86966 178802
rect 87030 178738 87046 178802
rect 87110 178738 87126 178802
rect 87190 178738 87198 178802
rect 86878 177714 87198 178738
rect 86878 177650 86886 177714
rect 86950 177650 86966 177714
rect 87030 177650 87046 177714
rect 87110 177650 87126 177714
rect 87190 177650 87198 177714
rect 86878 176626 87198 177650
rect 86878 176562 86886 176626
rect 86950 176562 86966 176626
rect 87030 176562 87046 176626
rect 87110 176562 87126 176626
rect 87190 176562 87198 176626
rect 86878 175538 87198 176562
rect 86878 175474 86886 175538
rect 86950 175474 86966 175538
rect 87030 175474 87046 175538
rect 87110 175474 87126 175538
rect 87190 175474 87198 175538
rect 86878 174450 87198 175474
rect 86878 174386 86886 174450
rect 86950 174386 86966 174450
rect 87030 174386 87046 174450
rect 87110 174386 87126 174450
rect 87190 174386 87198 174450
rect 86878 173362 87198 174386
rect 86878 173298 86886 173362
rect 86950 173298 86966 173362
rect 87030 173298 87046 173362
rect 87110 173298 87126 173362
rect 87190 173298 87198 173362
rect 86878 172274 87198 173298
rect 86878 172210 86886 172274
rect 86950 172210 86966 172274
rect 87030 172210 87046 172274
rect 87110 172210 87126 172274
rect 87190 172210 87198 172274
rect 86878 171186 87198 172210
rect 86878 171122 86886 171186
rect 86950 171122 86966 171186
rect 87030 171122 87046 171186
rect 87110 171122 87126 171186
rect 87190 171122 87198 171186
rect 86878 170370 87198 171122
rect 86878 170134 86920 170370
rect 87156 170134 87198 170370
rect 86878 170098 87198 170134
rect 86878 170034 86886 170098
rect 86950 170034 86966 170098
rect 87030 170034 87046 170098
rect 87110 170034 87126 170098
rect 87190 170034 87198 170098
rect 86878 169010 87198 170034
rect 86878 168946 86886 169010
rect 86950 168946 86966 169010
rect 87030 168946 87046 169010
rect 87110 168946 87126 169010
rect 87190 168946 87198 169010
rect 86878 167922 87198 168946
rect 86878 167858 86886 167922
rect 86950 167858 86966 167922
rect 87030 167858 87046 167922
rect 87110 167858 87126 167922
rect 87190 167858 87198 167922
rect 86878 166834 87198 167858
rect 86878 166770 86886 166834
rect 86950 166770 86966 166834
rect 87030 166770 87046 166834
rect 87110 166770 87126 166834
rect 87190 166770 87198 166834
rect 86878 165746 87198 166770
rect 86878 165682 86886 165746
rect 86950 165682 86966 165746
rect 87030 165682 87046 165746
rect 87110 165682 87126 165746
rect 87190 165682 87198 165746
rect 86878 164658 87198 165682
rect 86878 164594 86886 164658
rect 86950 164594 86966 164658
rect 87030 164594 87046 164658
rect 87110 164594 87126 164658
rect 87190 164594 87198 164658
rect 86878 163570 87198 164594
rect 86878 163506 86886 163570
rect 86950 163506 86966 163570
rect 87030 163506 87046 163570
rect 87110 163506 87126 163570
rect 87190 163506 87198 163570
rect 86878 162482 87198 163506
rect 86878 162418 86886 162482
rect 86950 162418 86966 162482
rect 87030 162418 87046 162482
rect 87110 162418 87126 162482
rect 87190 162418 87198 162482
rect 86878 161394 87198 162418
rect 86878 161330 86886 161394
rect 86950 161330 86966 161394
rect 87030 161330 87046 161394
rect 87110 161330 87126 161394
rect 87190 161330 87198 161394
rect 86878 160370 87198 161330
rect 86878 160306 86920 160370
rect 87156 160306 87198 160370
rect 86878 160242 86886 160306
rect 87190 160242 87198 160306
rect 86878 160134 86920 160242
rect 87156 160134 87198 160242
rect 86878 159218 87198 160134
rect 86878 159154 86886 159218
rect 86950 159154 86966 159218
rect 87030 159154 87046 159218
rect 87110 159154 87126 159218
rect 87190 159154 87198 159218
rect 86878 158130 87198 159154
rect 86878 158066 86886 158130
rect 86950 158066 86966 158130
rect 87030 158066 87046 158130
rect 87110 158066 87126 158130
rect 87190 158066 87198 158130
rect 86878 157042 87198 158066
rect 86878 156978 86886 157042
rect 86950 156978 86966 157042
rect 87030 156978 87046 157042
rect 87110 156978 87126 157042
rect 87190 156978 87198 157042
rect 86878 155954 87198 156978
rect 86878 155890 86886 155954
rect 86950 155890 86966 155954
rect 87030 155890 87046 155954
rect 87110 155890 87126 155954
rect 87190 155890 87198 155954
rect 86878 154866 87198 155890
rect 86878 154802 86886 154866
rect 86950 154802 86966 154866
rect 87030 154802 87046 154866
rect 87110 154802 87126 154866
rect 87190 154802 87198 154866
rect 86878 153778 87198 154802
rect 86878 153714 86886 153778
rect 86950 153714 86966 153778
rect 87030 153714 87046 153778
rect 87110 153714 87126 153778
rect 87190 153714 87198 153778
rect 86878 152690 87198 153714
rect 86878 152626 86886 152690
rect 86950 152626 86966 152690
rect 87030 152626 87046 152690
rect 87110 152626 87126 152690
rect 87190 152626 87198 152690
rect 86878 151602 87198 152626
rect 86878 151538 86886 151602
rect 86950 151538 86966 151602
rect 87030 151538 87046 151602
rect 87110 151538 87126 151602
rect 87190 151538 87198 151602
rect 86878 150514 87198 151538
rect 86878 150450 86886 150514
rect 86950 150450 86966 150514
rect 87030 150450 87046 150514
rect 87110 150450 87126 150514
rect 87190 150450 87198 150514
rect 86878 150370 87198 150450
rect 86878 150134 86920 150370
rect 87156 150134 87198 150370
rect 86878 149426 87198 150134
rect 86878 149362 86886 149426
rect 86950 149362 86966 149426
rect 87030 149362 87046 149426
rect 87110 149362 87126 149426
rect 87190 149362 87198 149426
rect 86878 148338 87198 149362
rect 86878 148274 86886 148338
rect 86950 148274 86966 148338
rect 87030 148274 87046 148338
rect 87110 148274 87126 148338
rect 87190 148274 87198 148338
rect 86878 147250 87198 148274
rect 86878 147186 86886 147250
rect 86950 147186 86966 147250
rect 87030 147186 87046 147250
rect 87110 147186 87126 147250
rect 87190 147186 87198 147250
rect 86878 146162 87198 147186
rect 86878 146098 86886 146162
rect 86950 146098 86966 146162
rect 87030 146098 87046 146162
rect 87110 146098 87126 146162
rect 87190 146098 87198 146162
rect 86878 145074 87198 146098
rect 86878 145010 86886 145074
rect 86950 145010 86966 145074
rect 87030 145010 87046 145074
rect 87110 145010 87126 145074
rect 87190 145010 87198 145074
rect 86878 143986 87198 145010
rect 86878 143922 86886 143986
rect 86950 143922 86966 143986
rect 87030 143922 87046 143986
rect 87110 143922 87126 143986
rect 87190 143922 87198 143986
rect 86878 142898 87198 143922
rect 86878 142834 86886 142898
rect 86950 142834 86966 142898
rect 87030 142834 87046 142898
rect 87110 142834 87126 142898
rect 87190 142834 87198 142898
rect 86878 141810 87198 142834
rect 86878 141746 86886 141810
rect 86950 141746 86966 141810
rect 87030 141746 87046 141810
rect 87110 141746 87126 141810
rect 87190 141746 87198 141810
rect 86878 140722 87198 141746
rect 86878 140658 86886 140722
rect 86950 140658 86966 140722
rect 87030 140658 87046 140722
rect 87110 140658 87126 140722
rect 87190 140658 87198 140722
rect 86878 140370 87198 140658
rect 86878 140134 86920 140370
rect 87156 140134 87198 140370
rect 86878 139634 87198 140134
rect 86878 139570 86886 139634
rect 86950 139570 86966 139634
rect 87030 139570 87046 139634
rect 87110 139570 87126 139634
rect 87190 139570 87198 139634
rect 86878 138546 87198 139570
rect 86878 138482 86886 138546
rect 86950 138482 86966 138546
rect 87030 138482 87046 138546
rect 87110 138482 87126 138546
rect 87190 138482 87198 138546
rect 86878 137458 87198 138482
rect 86878 137394 86886 137458
rect 86950 137394 86966 137458
rect 87030 137394 87046 137458
rect 87110 137394 87126 137458
rect 87190 137394 87198 137458
rect 86878 136370 87198 137394
rect 86878 136306 86886 136370
rect 86950 136306 86966 136370
rect 87030 136306 87046 136370
rect 87110 136306 87126 136370
rect 87190 136306 87198 136370
rect 86878 135282 87198 136306
rect 86878 135218 86886 135282
rect 86950 135218 86966 135282
rect 87030 135218 87046 135282
rect 87110 135218 87126 135282
rect 87190 135218 87198 135282
rect 86878 134194 87198 135218
rect 86878 134130 86886 134194
rect 86950 134130 86966 134194
rect 87030 134130 87046 134194
rect 87110 134130 87126 134194
rect 87190 134130 87198 134194
rect 86878 133106 87198 134130
rect 86878 133042 86886 133106
rect 86950 133042 86966 133106
rect 87030 133042 87046 133106
rect 87110 133042 87126 133106
rect 87190 133042 87198 133106
rect 86878 132018 87198 133042
rect 86878 131954 86886 132018
rect 86950 131954 86966 132018
rect 87030 131954 87046 132018
rect 87110 131954 87126 132018
rect 87190 131954 87198 132018
rect 86878 130930 87198 131954
rect 86878 130866 86886 130930
rect 86950 130866 86966 130930
rect 87030 130866 87046 130930
rect 87110 130866 87126 130930
rect 87190 130866 87198 130930
rect 86878 130370 87198 130866
rect 86878 130134 86920 130370
rect 87156 130134 87198 130370
rect 86878 129842 87198 130134
rect 86878 129778 86886 129842
rect 86950 129778 86966 129842
rect 87030 129778 87046 129842
rect 87110 129778 87126 129842
rect 87190 129778 87198 129842
rect 86878 128754 87198 129778
rect 86878 128690 86886 128754
rect 86950 128690 86966 128754
rect 87030 128690 87046 128754
rect 87110 128690 87126 128754
rect 87190 128690 87198 128754
rect 86878 127666 87198 128690
rect 86878 127602 86886 127666
rect 86950 127602 86966 127666
rect 87030 127602 87046 127666
rect 87110 127602 87126 127666
rect 87190 127602 87198 127666
rect 86878 126578 87198 127602
rect 86878 126514 86886 126578
rect 86950 126514 86966 126578
rect 87030 126514 87046 126578
rect 87110 126514 87126 126578
rect 87190 126514 87198 126578
rect 86878 125490 87198 126514
rect 86878 125426 86886 125490
rect 86950 125426 86966 125490
rect 87030 125426 87046 125490
rect 87110 125426 87126 125490
rect 87190 125426 87198 125490
rect 86878 124402 87198 125426
rect 86878 124338 86886 124402
rect 86950 124338 86966 124402
rect 87030 124338 87046 124402
rect 87110 124338 87126 124402
rect 87190 124338 87198 124402
rect 86878 123314 87198 124338
rect 86878 123250 86886 123314
rect 86950 123250 86966 123314
rect 87030 123250 87046 123314
rect 87110 123250 87126 123314
rect 87190 123250 87198 123314
rect 86878 122226 87198 123250
rect 86878 122162 86886 122226
rect 86950 122162 86966 122226
rect 87030 122162 87046 122226
rect 87110 122162 87126 122226
rect 87190 122162 87198 122226
rect 86878 121138 87198 122162
rect 86878 121074 86886 121138
rect 86950 121074 86966 121138
rect 87030 121074 87046 121138
rect 87110 121074 87126 121138
rect 87190 121074 87198 121138
rect 86878 120370 87198 121074
rect 86878 120134 86920 120370
rect 87156 120134 87198 120370
rect 86878 120050 87198 120134
rect 86878 119986 86886 120050
rect 86950 119986 86966 120050
rect 87030 119986 87046 120050
rect 87110 119986 87126 120050
rect 87190 119986 87198 120050
rect 86878 118962 87198 119986
rect 86878 118898 86886 118962
rect 86950 118898 86966 118962
rect 87030 118898 87046 118962
rect 87110 118898 87126 118962
rect 87190 118898 87198 118962
rect 86878 117874 87198 118898
rect 86878 117810 86886 117874
rect 86950 117810 86966 117874
rect 87030 117810 87046 117874
rect 87110 117810 87126 117874
rect 87190 117810 87198 117874
rect 86878 116786 87198 117810
rect 86878 116722 86886 116786
rect 86950 116722 86966 116786
rect 87030 116722 87046 116786
rect 87110 116722 87126 116786
rect 87190 116722 87198 116786
rect 86878 115698 87198 116722
rect 86878 115634 86886 115698
rect 86950 115634 86966 115698
rect 87030 115634 87046 115698
rect 87110 115634 87126 115698
rect 87190 115634 87198 115698
rect 86878 114610 87198 115634
rect 86878 114546 86886 114610
rect 86950 114546 86966 114610
rect 87030 114546 87046 114610
rect 87110 114546 87126 114610
rect 87190 114546 87198 114610
rect 86878 113522 87198 114546
rect 86878 113458 86886 113522
rect 86950 113458 86966 113522
rect 87030 113458 87046 113522
rect 87110 113458 87126 113522
rect 87190 113458 87198 113522
rect 86878 112434 87198 113458
rect 86878 112370 86886 112434
rect 86950 112370 86966 112434
rect 87030 112370 87046 112434
rect 87110 112370 87126 112434
rect 87190 112370 87198 112434
rect 86878 111346 87198 112370
rect 86878 111282 86886 111346
rect 86950 111282 86966 111346
rect 87030 111282 87046 111346
rect 87110 111282 87126 111346
rect 87190 111282 87198 111346
rect 86878 110370 87198 111282
rect 86878 110258 86920 110370
rect 87156 110258 87198 110370
rect 86878 110194 86886 110258
rect 87190 110194 87198 110258
rect 86878 110134 86920 110194
rect 87156 110134 87198 110194
rect 86878 109170 87198 110134
rect 86878 109106 86886 109170
rect 86950 109106 86966 109170
rect 87030 109106 87046 109170
rect 87110 109106 87126 109170
rect 87190 109106 87198 109170
rect 86878 108082 87198 109106
rect 86878 108018 86886 108082
rect 86950 108018 86966 108082
rect 87030 108018 87046 108082
rect 87110 108018 87126 108082
rect 87190 108018 87198 108082
rect 86878 106994 87198 108018
rect 86878 106930 86886 106994
rect 86950 106930 86966 106994
rect 87030 106930 87046 106994
rect 87110 106930 87126 106994
rect 87190 106930 87198 106994
rect 86878 105906 87198 106930
rect 86878 105842 86886 105906
rect 86950 105842 86966 105906
rect 87030 105842 87046 105906
rect 87110 105842 87126 105906
rect 87190 105842 87198 105906
rect 86878 104818 87198 105842
rect 86878 104754 86886 104818
rect 86950 104754 86966 104818
rect 87030 104754 87046 104818
rect 87110 104754 87126 104818
rect 87190 104754 87198 104818
rect 86878 103730 87198 104754
rect 86878 103666 86886 103730
rect 86950 103666 86966 103730
rect 87030 103666 87046 103730
rect 87110 103666 87126 103730
rect 87190 103666 87198 103730
rect 86878 102642 87198 103666
rect 86878 102578 86886 102642
rect 86950 102578 86966 102642
rect 87030 102578 87046 102642
rect 87110 102578 87126 102642
rect 87190 102578 87198 102642
rect 86878 101554 87198 102578
rect 86878 101490 86886 101554
rect 86950 101490 86966 101554
rect 87030 101490 87046 101554
rect 87110 101490 87126 101554
rect 87190 101490 87198 101554
rect 86878 100466 87198 101490
rect 86878 100402 86886 100466
rect 86950 100402 86966 100466
rect 87030 100402 87046 100466
rect 87110 100402 87126 100466
rect 87190 100402 87198 100466
rect 86878 100370 87198 100402
rect 86878 100134 86920 100370
rect 87156 100134 87198 100370
rect 86878 99378 87198 100134
rect 86878 99314 86886 99378
rect 86950 99314 86966 99378
rect 87030 99314 87046 99378
rect 87110 99314 87126 99378
rect 87190 99314 87198 99378
rect 86878 98290 87198 99314
rect 86878 98226 86886 98290
rect 86950 98226 86966 98290
rect 87030 98226 87046 98290
rect 87110 98226 87126 98290
rect 87190 98226 87198 98290
rect 86878 97202 87198 98226
rect 86878 97138 86886 97202
rect 86950 97138 86966 97202
rect 87030 97138 87046 97202
rect 87110 97138 87126 97202
rect 87190 97138 87198 97202
rect 86878 96114 87198 97138
rect 86878 96050 86886 96114
rect 86950 96050 86966 96114
rect 87030 96050 87046 96114
rect 87110 96050 87126 96114
rect 87190 96050 87198 96114
rect 86878 95026 87198 96050
rect 86878 94962 86886 95026
rect 86950 94962 86966 95026
rect 87030 94962 87046 95026
rect 87110 94962 87126 95026
rect 87190 94962 87198 95026
rect 86878 93938 87198 94962
rect 86878 93874 86886 93938
rect 86950 93874 86966 93938
rect 87030 93874 87046 93938
rect 87110 93874 87126 93938
rect 87190 93874 87198 93938
rect 86878 92850 87198 93874
rect 86878 92786 86886 92850
rect 86950 92786 86966 92850
rect 87030 92786 87046 92850
rect 87110 92786 87126 92850
rect 87190 92786 87198 92850
rect 86878 91762 87198 92786
rect 86878 91698 86886 91762
rect 86950 91698 86966 91762
rect 87030 91698 87046 91762
rect 87110 91698 87126 91762
rect 87190 91698 87198 91762
rect 86878 90674 87198 91698
rect 86878 90610 86886 90674
rect 86950 90610 86966 90674
rect 87030 90610 87046 90674
rect 87110 90610 87126 90674
rect 87190 90610 87198 90674
rect 86878 90370 87198 90610
rect 86878 90134 86920 90370
rect 87156 90134 87198 90370
rect 86878 89586 87198 90134
rect 86878 89522 86886 89586
rect 86950 89522 86966 89586
rect 87030 89522 87046 89586
rect 87110 89522 87126 89586
rect 87190 89522 87198 89586
rect 86878 88498 87198 89522
rect 86878 88434 86886 88498
rect 86950 88434 86966 88498
rect 87030 88434 87046 88498
rect 87110 88434 87126 88498
rect 87190 88434 87198 88498
rect 86878 87410 87198 88434
rect 86878 87346 86886 87410
rect 86950 87346 86966 87410
rect 87030 87346 87046 87410
rect 87110 87346 87126 87410
rect 87190 87346 87198 87410
rect 86878 86322 87198 87346
rect 86878 86258 86886 86322
rect 86950 86258 86966 86322
rect 87030 86258 87046 86322
rect 87110 86258 87126 86322
rect 87190 86258 87198 86322
rect 86878 85234 87198 86258
rect 86878 85170 86886 85234
rect 86950 85170 86966 85234
rect 87030 85170 87046 85234
rect 87110 85170 87126 85234
rect 87190 85170 87198 85234
rect 86878 84146 87198 85170
rect 86878 84082 86886 84146
rect 86950 84082 86966 84146
rect 87030 84082 87046 84146
rect 87110 84082 87126 84146
rect 87190 84082 87198 84146
rect 86878 83058 87198 84082
rect 86878 82994 86886 83058
rect 86950 82994 86966 83058
rect 87030 82994 87046 83058
rect 87110 82994 87126 83058
rect 87190 82994 87198 83058
rect 86878 81970 87198 82994
rect 86878 81906 86886 81970
rect 86950 81906 86966 81970
rect 87030 81906 87046 81970
rect 87110 81906 87126 81970
rect 87190 81906 87198 81970
rect 86878 80882 87198 81906
rect 86878 80818 86886 80882
rect 86950 80818 86966 80882
rect 87030 80818 87046 80882
rect 87110 80818 87126 80882
rect 87190 80818 87198 80882
rect 86878 80370 87198 80818
rect 86878 80134 86920 80370
rect 87156 80134 87198 80370
rect 86878 79794 87198 80134
rect 86878 79730 86886 79794
rect 86950 79730 86966 79794
rect 87030 79730 87046 79794
rect 87110 79730 87126 79794
rect 87190 79730 87198 79794
rect 86878 78706 87198 79730
rect 86878 78642 86886 78706
rect 86950 78642 86966 78706
rect 87030 78642 87046 78706
rect 87110 78642 87126 78706
rect 87190 78642 87198 78706
rect 86878 77618 87198 78642
rect 86878 77554 86886 77618
rect 86950 77554 86966 77618
rect 87030 77554 87046 77618
rect 87110 77554 87126 77618
rect 87190 77554 87198 77618
rect 86878 76530 87198 77554
rect 86878 76466 86886 76530
rect 86950 76466 86966 76530
rect 87030 76466 87046 76530
rect 87110 76466 87126 76530
rect 87190 76466 87198 76530
rect 86878 75442 87198 76466
rect 86878 75378 86886 75442
rect 86950 75378 86966 75442
rect 87030 75378 87046 75442
rect 87110 75378 87126 75442
rect 87190 75378 87198 75442
rect 86878 74354 87198 75378
rect 86878 74290 86886 74354
rect 86950 74290 86966 74354
rect 87030 74290 87046 74354
rect 87110 74290 87126 74354
rect 87190 74290 87198 74354
rect 86878 73266 87198 74290
rect 86878 73202 86886 73266
rect 86950 73202 86966 73266
rect 87030 73202 87046 73266
rect 87110 73202 87126 73266
rect 87190 73202 87198 73266
rect 86878 72178 87198 73202
rect 86878 72114 86886 72178
rect 86950 72114 86966 72178
rect 87030 72114 87046 72178
rect 87110 72114 87126 72178
rect 87190 72114 87198 72178
rect 86878 71090 87198 72114
rect 86878 71026 86886 71090
rect 86950 71026 86966 71090
rect 87030 71026 87046 71090
rect 87110 71026 87126 71090
rect 87190 71026 87198 71090
rect 86878 70370 87198 71026
rect 86878 70134 86920 70370
rect 87156 70134 87198 70370
rect 86878 70002 87198 70134
rect 86878 69938 86886 70002
rect 86950 69938 86966 70002
rect 87030 69938 87046 70002
rect 87110 69938 87126 70002
rect 87190 69938 87198 70002
rect 86878 68914 87198 69938
rect 86878 68850 86886 68914
rect 86950 68850 86966 68914
rect 87030 68850 87046 68914
rect 87110 68850 87126 68914
rect 87190 68850 87198 68914
rect 86878 67826 87198 68850
rect 86878 67762 86886 67826
rect 86950 67762 86966 67826
rect 87030 67762 87046 67826
rect 87110 67762 87126 67826
rect 87190 67762 87198 67826
rect 86878 66738 87198 67762
rect 86878 66674 86886 66738
rect 86950 66674 86966 66738
rect 87030 66674 87046 66738
rect 87110 66674 87126 66738
rect 87190 66674 87198 66738
rect 86878 65650 87198 66674
rect 86878 65586 86886 65650
rect 86950 65586 86966 65650
rect 87030 65586 87046 65650
rect 87110 65586 87126 65650
rect 87190 65586 87198 65650
rect 86878 64562 87198 65586
rect 86878 64498 86886 64562
rect 86950 64498 86966 64562
rect 87030 64498 87046 64562
rect 87110 64498 87126 64562
rect 87190 64498 87198 64562
rect 86878 63474 87198 64498
rect 86878 63410 86886 63474
rect 86950 63410 86966 63474
rect 87030 63410 87046 63474
rect 87110 63410 87126 63474
rect 87190 63410 87198 63474
rect 86878 62386 87198 63410
rect 86878 62322 86886 62386
rect 86950 62322 86966 62386
rect 87030 62322 87046 62386
rect 87110 62322 87126 62386
rect 87190 62322 87198 62386
rect 86878 61298 87198 62322
rect 86878 61234 86886 61298
rect 86950 61234 86966 61298
rect 87030 61234 87046 61298
rect 87110 61234 87126 61298
rect 87190 61234 87198 61298
rect 86878 60370 87198 61234
rect 86878 60210 86920 60370
rect 87156 60210 87198 60370
rect 86878 60146 86886 60210
rect 87190 60146 87198 60210
rect 86878 60134 86920 60146
rect 87156 60134 87198 60146
rect 86878 59122 87198 60134
rect 86878 59058 86886 59122
rect 86950 59058 86966 59122
rect 87030 59058 87046 59122
rect 87110 59058 87126 59122
rect 87190 59058 87198 59122
rect 86878 58034 87198 59058
rect 86878 57970 86886 58034
rect 86950 57970 86966 58034
rect 87030 57970 87046 58034
rect 87110 57970 87126 58034
rect 87190 57970 87198 58034
rect 86878 56946 87198 57970
rect 86878 56882 86886 56946
rect 86950 56882 86966 56946
rect 87030 56882 87046 56946
rect 87110 56882 87126 56946
rect 87190 56882 87198 56946
rect 86878 55858 87198 56882
rect 86878 55794 86886 55858
rect 86950 55794 86966 55858
rect 87030 55794 87046 55858
rect 87110 55794 87126 55858
rect 87190 55794 87198 55858
rect 86878 54770 87198 55794
rect 86878 54706 86886 54770
rect 86950 54706 86966 54770
rect 87030 54706 87046 54770
rect 87110 54706 87126 54770
rect 87190 54706 87198 54770
rect 86878 53682 87198 54706
rect 86878 53618 86886 53682
rect 86950 53618 86966 53682
rect 87030 53618 87046 53682
rect 87110 53618 87126 53682
rect 87190 53618 87198 53682
rect 86878 52594 87198 53618
rect 86878 52530 86886 52594
rect 86950 52530 86966 52594
rect 87030 52530 87046 52594
rect 87110 52530 87126 52594
rect 87190 52530 87198 52594
rect 86878 51506 87198 52530
rect 86878 51442 86886 51506
rect 86950 51442 86966 51506
rect 87030 51442 87046 51506
rect 87110 51442 87126 51506
rect 87190 51442 87198 51506
rect 86878 50418 87198 51442
rect 86878 50354 86886 50418
rect 86950 50370 86966 50418
rect 87030 50370 87046 50418
rect 87110 50370 87126 50418
rect 87190 50354 87198 50418
rect 86878 50134 86920 50354
rect 87156 50134 87198 50354
rect 86878 49330 87198 50134
rect 86878 49266 86886 49330
rect 86950 49266 86966 49330
rect 87030 49266 87046 49330
rect 87110 49266 87126 49330
rect 87190 49266 87198 49330
rect 86878 48242 87198 49266
rect 86878 48178 86886 48242
rect 86950 48178 86966 48242
rect 87030 48178 87046 48242
rect 87110 48178 87126 48242
rect 87190 48178 87198 48242
rect 86878 47154 87198 48178
rect 86878 47090 86886 47154
rect 86950 47090 86966 47154
rect 87030 47090 87046 47154
rect 87110 47090 87126 47154
rect 87190 47090 87198 47154
rect 86878 46066 87198 47090
rect 86878 46002 86886 46066
rect 86950 46002 86966 46066
rect 87030 46002 87046 46066
rect 87110 46002 87126 46066
rect 87190 46002 87198 46066
rect 86878 44978 87198 46002
rect 86878 44914 86886 44978
rect 86950 44914 86966 44978
rect 87030 44914 87046 44978
rect 87110 44914 87126 44978
rect 87190 44914 87198 44978
rect 86878 43890 87198 44914
rect 86878 43826 86886 43890
rect 86950 43826 86966 43890
rect 87030 43826 87046 43890
rect 87110 43826 87126 43890
rect 87190 43826 87198 43890
rect 86878 42802 87198 43826
rect 86878 42738 86886 42802
rect 86950 42738 86966 42802
rect 87030 42738 87046 42802
rect 87110 42738 87126 42802
rect 87190 42738 87198 42802
rect 86878 41714 87198 42738
rect 86878 41650 86886 41714
rect 86950 41650 86966 41714
rect 87030 41650 87046 41714
rect 87110 41650 87126 41714
rect 87190 41650 87198 41714
rect 86878 40626 87198 41650
rect 86878 40562 86886 40626
rect 86950 40562 86966 40626
rect 87030 40562 87046 40626
rect 87110 40562 87126 40626
rect 87190 40562 87198 40626
rect 86878 40370 87198 40562
rect 86878 40134 86920 40370
rect 87156 40134 87198 40370
rect 86878 39538 87198 40134
rect 86878 39474 86886 39538
rect 86950 39474 86966 39538
rect 87030 39474 87046 39538
rect 87110 39474 87126 39538
rect 87190 39474 87198 39538
rect 86878 38450 87198 39474
rect 86878 38386 86886 38450
rect 86950 38386 86966 38450
rect 87030 38386 87046 38450
rect 87110 38386 87126 38450
rect 87190 38386 87198 38450
rect 86878 37362 87198 38386
rect 86878 37298 86886 37362
rect 86950 37298 86966 37362
rect 87030 37298 87046 37362
rect 87110 37298 87126 37362
rect 87190 37298 87198 37362
rect 86878 36274 87198 37298
rect 86878 36210 86886 36274
rect 86950 36210 86966 36274
rect 87030 36210 87046 36274
rect 87110 36210 87126 36274
rect 87190 36210 87198 36274
rect 86878 35186 87198 36210
rect 86878 35122 86886 35186
rect 86950 35122 86966 35186
rect 87030 35122 87046 35186
rect 87110 35122 87126 35186
rect 87190 35122 87198 35186
rect 86878 34098 87198 35122
rect 86878 34034 86886 34098
rect 86950 34034 86966 34098
rect 87030 34034 87046 34098
rect 87110 34034 87126 34098
rect 87190 34034 87198 34098
rect 86878 33010 87198 34034
rect 86878 32946 86886 33010
rect 86950 32946 86966 33010
rect 87030 32946 87046 33010
rect 87110 32946 87126 33010
rect 87190 32946 87198 33010
rect 86878 31922 87198 32946
rect 86878 31858 86886 31922
rect 86950 31858 86966 31922
rect 87030 31858 87046 31922
rect 87110 31858 87126 31922
rect 87190 31858 87198 31922
rect 86878 30834 87198 31858
rect 86878 30770 86886 30834
rect 86950 30770 86966 30834
rect 87030 30770 87046 30834
rect 87110 30770 87126 30834
rect 87190 30770 87198 30834
rect 86878 30370 87198 30770
rect 86878 30134 86920 30370
rect 87156 30134 87198 30370
rect 86878 29746 87198 30134
rect 86878 29682 86886 29746
rect 86950 29682 86966 29746
rect 87030 29682 87046 29746
rect 87110 29682 87126 29746
rect 87190 29682 87198 29746
rect 84878 29138 84886 29202
rect 84950 29138 84966 29202
rect 85030 29138 85046 29202
rect 85110 29138 85126 29202
rect 85190 29138 85198 29202
rect 84878 28114 85198 29138
rect 86878 28658 87198 29682
rect 86878 28594 86886 28658
rect 86950 28594 86966 28658
rect 87030 28594 87046 28658
rect 87110 28594 87126 28658
rect 87190 28594 87198 28658
rect 85473 28318 85539 28319
rect 85473 28254 85474 28318
rect 85538 28254 85539 28318
rect 85473 28253 85539 28254
rect 85476 28132 85536 28253
rect 84878 28050 84886 28114
rect 84950 28050 84966 28114
rect 85030 28050 85046 28114
rect 85110 28050 85126 28114
rect 85190 28050 85198 28114
rect 84878 27026 85198 28050
rect 84878 26962 84886 27026
rect 84950 26962 84966 27026
rect 85030 26962 85046 27026
rect 85110 26962 85126 27026
rect 85190 26962 85198 27026
rect 84878 25938 85198 26962
rect 84878 25874 84886 25938
rect 84950 25874 84966 25938
rect 85030 25874 85046 25938
rect 85110 25874 85126 25938
rect 85190 25874 85198 25938
rect 84878 25370 85198 25874
rect 84878 25134 84920 25370
rect 85156 25134 85198 25370
rect 84878 24850 85198 25134
rect 84878 24786 84886 24850
rect 84950 24786 84966 24850
rect 85030 24786 85046 24850
rect 85110 24786 85126 24850
rect 85190 24786 85198 24850
rect 84878 23762 85198 24786
rect 84878 23698 84886 23762
rect 84950 23698 84966 23762
rect 85030 23698 85046 23762
rect 85110 23698 85126 23762
rect 85190 23698 85198 23762
rect 84878 22674 85198 23698
rect 84878 22610 84886 22674
rect 84950 22610 84966 22674
rect 85030 22610 85046 22674
rect 85110 22610 85126 22674
rect 85190 22610 85198 22674
rect 84878 21586 85198 22610
rect 84878 21522 84886 21586
rect 84950 21522 84966 21586
rect 85030 21522 85046 21586
rect 85110 21522 85126 21586
rect 85190 21522 85198 21586
rect 84878 20498 85198 21522
rect 84878 20434 84886 20498
rect 84950 20434 84966 20498
rect 85030 20434 85046 20498
rect 85110 20434 85126 20498
rect 85190 20434 85198 20498
rect 84878 19410 85198 20434
rect 84878 19346 84886 19410
rect 84950 19346 84966 19410
rect 85030 19346 85046 19410
rect 85110 19346 85126 19410
rect 85190 19346 85198 19410
rect 84878 18322 85198 19346
rect 84878 18258 84886 18322
rect 84950 18258 84966 18322
rect 85030 18258 85046 18322
rect 85110 18258 85126 18322
rect 85190 18258 85198 18322
rect 84878 17234 85198 18258
rect 84878 17170 84886 17234
rect 84950 17170 84966 17234
rect 85030 17170 85046 17234
rect 85110 17170 85126 17234
rect 85190 17170 85198 17234
rect 84878 16146 85198 17170
rect 84878 16082 84886 16146
rect 84950 16082 84966 16146
rect 85030 16082 85046 16146
rect 85110 16082 85126 16146
rect 85190 16082 85198 16146
rect 84878 15370 85198 16082
rect 84878 15134 84920 15370
rect 85156 15134 85198 15370
rect 84878 15058 85198 15134
rect 84878 14994 84886 15058
rect 84950 14994 84966 15058
rect 85030 14994 85046 15058
rect 85110 14994 85126 15058
rect 85190 14994 85198 15058
rect 84878 13970 85198 14994
rect 84878 13906 84886 13970
rect 84950 13906 84966 13970
rect 85030 13906 85046 13970
rect 85110 13906 85126 13970
rect 85190 13906 85198 13970
rect 84878 12882 85198 13906
rect 84878 12818 84886 12882
rect 84950 12818 84966 12882
rect 85030 12818 85046 12882
rect 85110 12818 85126 12882
rect 85190 12818 85198 12882
rect 84878 11794 85198 12818
rect 84878 11730 84886 11794
rect 84950 11730 84966 11794
rect 85030 11730 85046 11794
rect 85110 11730 85126 11794
rect 85190 11730 85198 11794
rect 84878 10706 85198 11730
rect 84878 10642 84886 10706
rect 84950 10642 84966 10706
rect 85030 10642 85046 10706
rect 85110 10642 85126 10706
rect 85190 10642 85198 10706
rect 84878 9618 85198 10642
rect 84878 9554 84886 9618
rect 84950 9554 84966 9618
rect 85030 9554 85046 9618
rect 85110 9554 85126 9618
rect 85190 9554 85198 9618
rect 84878 8530 85198 9554
rect 84878 8466 84886 8530
rect 84950 8466 84966 8530
rect 85030 8466 85046 8530
rect 85110 8466 85126 8530
rect 85190 8466 85198 8530
rect 84878 7442 85198 8466
rect 84878 7378 84886 7442
rect 84950 7378 84966 7442
rect 85030 7378 85046 7442
rect 85110 7378 85126 7442
rect 85190 7378 85198 7442
rect 84878 6354 85198 7378
rect 84878 6290 84886 6354
rect 84950 6290 84966 6354
rect 85030 6290 85046 6354
rect 85110 6290 85126 6354
rect 85190 6290 85198 6354
rect 84878 5370 85198 6290
rect 84878 5266 84920 5370
rect 85156 5266 85198 5370
rect 84878 5202 84886 5266
rect 85190 5202 85198 5266
rect 84878 5134 84920 5202
rect 85156 5134 85198 5202
rect 84878 4178 85198 5134
rect 84878 4114 84886 4178
rect 84950 4114 84966 4178
rect 85030 4114 85046 4178
rect 85110 4114 85126 4178
rect 85190 4114 85198 4178
rect 84878 3090 85198 4114
rect 84878 3026 84886 3090
rect 84950 3026 84966 3090
rect 85030 3026 85046 3090
rect 85110 3026 85126 3090
rect 85190 3026 85198 3090
rect 84878 2002 85198 3026
rect 84878 1938 84886 2002
rect 84950 1938 84966 2002
rect 85030 1938 85046 2002
rect 85110 1938 85126 2002
rect 85190 1938 85198 2002
rect 84878 1922 85198 1938
rect 86878 27570 87198 28594
rect 86878 27506 86886 27570
rect 86950 27506 86966 27570
rect 87030 27506 87046 27570
rect 87110 27506 87126 27570
rect 87190 27506 87198 27570
rect 86878 26482 87198 27506
rect 86878 26418 86886 26482
rect 86950 26418 86966 26482
rect 87030 26418 87046 26482
rect 87110 26418 87126 26482
rect 87190 26418 87198 26482
rect 86878 25394 87198 26418
rect 86878 25330 86886 25394
rect 86950 25330 86966 25394
rect 87030 25330 87046 25394
rect 87110 25330 87126 25394
rect 87190 25330 87198 25394
rect 86878 24306 87198 25330
rect 86878 24242 86886 24306
rect 86950 24242 86966 24306
rect 87030 24242 87046 24306
rect 87110 24242 87126 24306
rect 87190 24242 87198 24306
rect 86878 23218 87198 24242
rect 86878 23154 86886 23218
rect 86950 23154 86966 23218
rect 87030 23154 87046 23218
rect 87110 23154 87126 23218
rect 87190 23154 87198 23218
rect 86878 22130 87198 23154
rect 86878 22066 86886 22130
rect 86950 22066 86966 22130
rect 87030 22066 87046 22130
rect 87110 22066 87126 22130
rect 87190 22066 87198 22130
rect 86878 21042 87198 22066
rect 86878 20978 86886 21042
rect 86950 20978 86966 21042
rect 87030 20978 87046 21042
rect 87110 20978 87126 21042
rect 87190 20978 87198 21042
rect 86878 20370 87198 20978
rect 86878 20134 86920 20370
rect 87156 20134 87198 20370
rect 86878 19954 87198 20134
rect 86878 19890 86886 19954
rect 86950 19890 86966 19954
rect 87030 19890 87046 19954
rect 87110 19890 87126 19954
rect 87190 19890 87198 19954
rect 86878 18866 87198 19890
rect 86878 18802 86886 18866
rect 86950 18802 86966 18866
rect 87030 18802 87046 18866
rect 87110 18802 87126 18866
rect 87190 18802 87198 18866
rect 86878 17778 87198 18802
rect 86878 17714 86886 17778
rect 86950 17714 86966 17778
rect 87030 17714 87046 17778
rect 87110 17714 87126 17778
rect 87190 17714 87198 17778
rect 86878 16690 87198 17714
rect 86878 16626 86886 16690
rect 86950 16626 86966 16690
rect 87030 16626 87046 16690
rect 87110 16626 87126 16690
rect 87190 16626 87198 16690
rect 86878 15602 87198 16626
rect 86878 15538 86886 15602
rect 86950 15538 86966 15602
rect 87030 15538 87046 15602
rect 87110 15538 87126 15602
rect 87190 15538 87198 15602
rect 86878 14514 87198 15538
rect 86878 14450 86886 14514
rect 86950 14450 86966 14514
rect 87030 14450 87046 14514
rect 87110 14450 87126 14514
rect 87190 14450 87198 14514
rect 86878 13426 87198 14450
rect 86878 13362 86886 13426
rect 86950 13362 86966 13426
rect 87030 13362 87046 13426
rect 87110 13362 87126 13426
rect 87190 13362 87198 13426
rect 86878 12338 87198 13362
rect 86878 12274 86886 12338
rect 86950 12274 86966 12338
rect 87030 12274 87046 12338
rect 87110 12274 87126 12338
rect 87190 12274 87198 12338
rect 86878 11250 87198 12274
rect 86878 11186 86886 11250
rect 86950 11186 86966 11250
rect 87030 11186 87046 11250
rect 87110 11186 87126 11250
rect 87190 11186 87198 11250
rect 86878 10370 87198 11186
rect 86878 10162 86920 10370
rect 87156 10162 87198 10370
rect 86878 10098 86886 10162
rect 86950 10098 86966 10134
rect 87030 10098 87046 10134
rect 87110 10098 87126 10134
rect 87190 10098 87198 10162
rect 86878 9074 87198 10098
rect 86878 9010 86886 9074
rect 86950 9010 86966 9074
rect 87030 9010 87046 9074
rect 87110 9010 87126 9074
rect 87190 9010 87198 9074
rect 86878 7986 87198 9010
rect 86878 7922 86886 7986
rect 86950 7922 86966 7986
rect 87030 7922 87046 7986
rect 87110 7922 87126 7986
rect 87190 7922 87198 7986
rect 86878 6898 87198 7922
rect 86878 6834 86886 6898
rect 86950 6834 86966 6898
rect 87030 6834 87046 6898
rect 87110 6834 87126 6898
rect 87190 6834 87198 6898
rect 86878 5810 87198 6834
rect 86878 5746 86886 5810
rect 86950 5746 86966 5810
rect 87030 5746 87046 5810
rect 87110 5746 87126 5810
rect 87190 5746 87198 5810
rect 86878 4722 87198 5746
rect 86878 4658 86886 4722
rect 86950 4658 86966 4722
rect 87030 4658 87046 4722
rect 87110 4658 87126 4722
rect 87190 4658 87198 4722
rect 86878 3634 87198 4658
rect 86878 3570 86886 3634
rect 86950 3570 86966 3634
rect 87030 3570 87046 3634
rect 87110 3570 87126 3634
rect 87190 3570 87198 3634
rect 86878 2546 87198 3570
rect 86878 2482 86886 2546
rect 86950 2482 86966 2546
rect 87030 2482 87046 2546
rect 87110 2482 87126 2546
rect 87190 2482 87198 2546
rect 86878 1922 87198 2482
rect 84737 1390 84803 1391
rect 84737 1326 84738 1390
rect 84802 1326 84803 1390
rect 84737 1325 84803 1326
rect 83633 1118 83699 1119
rect 83633 1054 83634 1118
rect 83698 1054 83699 1118
rect 83633 1053 83699 1054
rect 52905 438 52971 439
rect 52905 374 52906 438
rect 52970 374 52971 438
rect 52905 373 52971 374
rect 83449 438 83515 439
rect 83449 374 83450 438
rect 83514 374 83515 438
rect 83449 373 83515 374
rect 50329 302 50395 303
rect 50329 238 50330 302
rect 50394 238 50395 302
rect 50329 237 50395 238
rect 25857 166 25923 167
rect 25857 102 25858 166
rect 25922 102 25923 166
rect 25857 101 25923 102
<< via4 >>
rect 920 185134 1156 185370
rect 920 175134 1156 175370
rect 920 165202 1156 165370
rect 920 165138 950 165202
rect 950 165138 966 165202
rect 966 165138 1030 165202
rect 1030 165138 1046 165202
rect 1046 165138 1110 165202
rect 1110 165138 1126 165202
rect 1126 165138 1156 165202
rect 920 165134 1156 165138
rect 920 155346 950 155370
rect 950 155346 966 155370
rect 966 155346 1030 155370
rect 1030 155346 1046 155370
rect 1046 155346 1110 155370
rect 1110 155346 1126 155370
rect 1126 155346 1156 155370
rect 920 155134 1156 155346
rect 920 145134 1156 145370
rect 920 135134 1156 135370
rect 920 125134 1156 125370
rect 2920 180134 3156 180370
rect 2920 170134 3156 170370
rect 2920 160306 3156 160370
rect 2920 160242 2950 160306
rect 2950 160242 2966 160306
rect 2966 160242 3030 160306
rect 3030 160242 3046 160306
rect 3046 160242 3110 160306
rect 3110 160242 3126 160306
rect 3126 160242 3156 160306
rect 2920 160134 3156 160242
rect 2920 150134 3156 150370
rect 2920 140134 3156 140370
rect 2920 130134 3156 130370
rect 920 115154 1156 115370
rect 920 115134 950 115154
rect 950 115134 966 115154
rect 966 115134 1030 115154
rect 1030 115134 1046 115154
rect 1046 115134 1110 115154
rect 1110 115134 1126 115154
rect 1126 115134 1156 115154
rect 2920 120134 3156 120370
rect 2920 110258 3156 110370
rect 2920 110194 2950 110258
rect 2950 110194 2966 110258
rect 2966 110194 3030 110258
rect 3030 110194 3046 110258
rect 3046 110194 3110 110258
rect 3110 110194 3126 110258
rect 3126 110194 3156 110258
rect 2920 110134 3156 110194
rect 920 105362 1156 105370
rect 920 105298 950 105362
rect 950 105298 966 105362
rect 966 105298 1030 105362
rect 1030 105298 1046 105362
rect 1046 105298 1110 105362
rect 1110 105298 1126 105362
rect 1126 105298 1156 105362
rect 920 105134 1156 105298
rect 920 95134 1156 95370
rect 920 85134 1156 85370
rect 920 75134 1156 75370
rect 920 65134 1156 65370
rect 920 55314 1156 55370
rect 920 55250 950 55314
rect 950 55250 966 55314
rect 966 55250 1030 55314
rect 1030 55250 1046 55314
rect 1046 55250 1110 55314
rect 1110 55250 1126 55314
rect 1126 55250 1156 55314
rect 920 55134 1156 55250
rect 920 45134 1156 45370
rect 920 35134 1156 35370
rect 920 25134 1156 25370
rect 920 15134 1156 15370
rect 920 5266 1156 5370
rect 920 5202 950 5266
rect 950 5202 966 5266
rect 966 5202 1030 5266
rect 1030 5202 1046 5266
rect 1046 5202 1110 5266
rect 1110 5202 1126 5266
rect 1126 5202 1156 5266
rect 920 5134 1156 5202
rect 2920 100134 3156 100370
rect 2920 90134 3156 90370
rect 2920 80134 3156 80370
rect 2920 70134 3156 70370
rect 2920 60210 3156 60370
rect 2920 60146 2950 60210
rect 2950 60146 2966 60210
rect 2966 60146 3030 60210
rect 3030 60146 3046 60210
rect 3046 60146 3110 60210
rect 3110 60146 3126 60210
rect 3126 60146 3156 60210
rect 2920 60134 3156 60146
rect 2920 50354 2950 50370
rect 2950 50354 2966 50370
rect 2966 50354 3030 50370
rect 3030 50354 3046 50370
rect 3046 50354 3110 50370
rect 3110 50354 3126 50370
rect 3126 50354 3156 50370
rect 2920 50134 3156 50354
rect 2920 40134 3156 40370
rect 2920 30134 3156 30370
rect 2920 20134 3156 20370
rect 2920 10162 3156 10370
rect 2920 10134 2950 10162
rect 2950 10134 2966 10162
rect 2966 10134 3030 10162
rect 3030 10134 3046 10162
rect 3046 10134 3110 10162
rect 3110 10134 3126 10162
rect 3126 10134 3156 10162
rect 84920 185134 85156 185370
rect 81916 180134 82152 180370
rect 81470 175134 81706 175370
rect 84920 175134 85156 175370
rect 81916 170134 82152 170370
rect 81470 165134 81706 165370
rect 81916 160134 82152 160370
rect 81470 155134 81706 155370
rect 5532 151806 5768 151892
rect 5532 151742 5618 151806
rect 5618 151742 5682 151806
rect 5682 151742 5768 151806
rect 5532 151656 5768 151742
rect 82260 151806 82496 151892
rect 82260 151742 82346 151806
rect 82346 151742 82410 151806
rect 82410 151742 82496 151806
rect 82260 151656 82496 151742
rect 81916 150134 82152 150370
rect 81470 145134 81706 145370
rect 81916 140134 82152 140370
rect 81470 135134 81706 135370
rect 81916 130134 82152 130370
rect 81470 125134 81706 125370
rect 81916 120134 82152 120370
rect 81470 115134 81706 115370
rect 81916 110134 82152 110370
rect 81470 105134 81706 105370
rect 81916 100134 82152 100370
rect 81916 90134 82152 90370
rect 81470 85134 81706 85370
rect 81916 80134 82152 80370
rect 81470 75134 81706 75370
rect 81916 70134 82152 70370
rect 81470 65134 81706 65370
rect 81916 60134 82152 60370
rect 81470 55134 81706 55370
rect 81916 50134 82152 50370
rect 81470 45134 81706 45370
rect 81916 40134 82152 40370
rect 81470 35134 81706 35370
rect 81916 30134 82152 30370
rect 5532 29478 5618 29492
rect 5618 29478 5682 29492
rect 5682 29478 5768 29492
rect 5532 29256 5768 29478
rect 5532 28046 5768 28132
rect 5532 27982 5618 28046
rect 5618 27982 5682 28046
rect 5682 27982 5768 28046
rect 5532 27896 5768 27982
rect 81470 25134 81706 25370
rect 81916 20134 82152 20370
rect 81470 15134 81706 15370
rect 81916 10134 82152 10370
rect 81470 5134 81706 5370
rect 84920 165202 85156 165370
rect 84920 165138 84950 165202
rect 84950 165138 84966 165202
rect 84966 165138 85030 165202
rect 85030 165138 85046 165202
rect 85046 165138 85110 165202
rect 85110 165138 85126 165202
rect 85126 165138 85156 165202
rect 84920 165134 85156 165138
rect 84920 155346 84950 155370
rect 84950 155346 84966 155370
rect 84966 155346 85030 155370
rect 85030 155346 85046 155370
rect 85046 155346 85110 155370
rect 85110 155346 85126 155370
rect 85126 155346 85156 155370
rect 84920 155134 85156 155346
rect 84920 145134 85156 145370
rect 84920 135134 85156 135370
rect 84920 125134 85156 125370
rect 84920 115154 85156 115370
rect 84920 115134 84950 115154
rect 84950 115134 84966 115154
rect 84966 115134 85030 115154
rect 85030 115134 85046 115154
rect 85046 115134 85110 115154
rect 85110 115134 85126 115154
rect 85126 115134 85156 115154
rect 84920 105362 85156 105370
rect 84920 105298 84950 105362
rect 84950 105298 84966 105362
rect 84966 105298 85030 105362
rect 85030 105298 85046 105362
rect 85046 105298 85110 105362
rect 85110 105298 85126 105362
rect 85126 105298 85156 105362
rect 84920 105134 85156 105298
rect 84920 95134 85156 95370
rect 84920 85134 85156 85370
rect 84920 75134 85156 75370
rect 84920 65134 85156 65370
rect 84920 55314 85156 55370
rect 84920 55250 84950 55314
rect 84950 55250 84966 55314
rect 84966 55250 85030 55314
rect 85030 55250 85046 55314
rect 85046 55250 85110 55314
rect 85110 55250 85126 55314
rect 85126 55250 85156 55314
rect 84920 55134 85156 55250
rect 84920 45134 85156 45370
rect 84920 35134 85156 35370
rect 86920 180134 87156 180370
rect 86920 170134 87156 170370
rect 86920 160306 87156 160370
rect 86920 160242 86950 160306
rect 86950 160242 86966 160306
rect 86966 160242 87030 160306
rect 87030 160242 87046 160306
rect 87046 160242 87110 160306
rect 87110 160242 87126 160306
rect 87126 160242 87156 160306
rect 86920 160134 87156 160242
rect 86920 150134 87156 150370
rect 86920 140134 87156 140370
rect 86920 130134 87156 130370
rect 86920 120134 87156 120370
rect 86920 110258 87156 110370
rect 86920 110194 86950 110258
rect 86950 110194 86966 110258
rect 86966 110194 87030 110258
rect 87030 110194 87046 110258
rect 87046 110194 87110 110258
rect 87110 110194 87126 110258
rect 87126 110194 87156 110258
rect 86920 110134 87156 110194
rect 86920 100134 87156 100370
rect 86920 90134 87156 90370
rect 86920 80134 87156 80370
rect 86920 70134 87156 70370
rect 86920 60210 87156 60370
rect 86920 60146 86950 60210
rect 86950 60146 86966 60210
rect 86966 60146 87030 60210
rect 87030 60146 87046 60210
rect 87046 60146 87110 60210
rect 87110 60146 87126 60210
rect 87126 60146 87156 60210
rect 86920 60134 87156 60146
rect 86920 50354 86950 50370
rect 86950 50354 86966 50370
rect 86966 50354 87030 50370
rect 87030 50354 87046 50370
rect 87046 50354 87110 50370
rect 87110 50354 87126 50370
rect 87126 50354 87156 50370
rect 86920 50134 87156 50354
rect 86920 40134 87156 40370
rect 86920 30134 87156 30370
rect 85388 29406 85624 29492
rect 85388 29342 85474 29406
rect 85474 29342 85538 29406
rect 85538 29342 85624 29406
rect 85388 29256 85624 29342
rect 85388 27896 85624 28132
rect 84920 25134 85156 25370
rect 84920 15134 85156 15370
rect 84920 5266 85156 5370
rect 84920 5202 84950 5266
rect 84950 5202 84966 5266
rect 84966 5202 85030 5266
rect 85030 5202 85046 5266
rect 85046 5202 85110 5266
rect 85110 5202 85126 5266
rect 85126 5202 85156 5266
rect 84920 5134 85156 5202
rect 86920 20134 87156 20370
rect 86920 10162 87156 10370
rect 86920 10134 86950 10162
rect 86950 10134 86966 10162
rect 86966 10134 87030 10162
rect 87030 10134 87046 10162
rect 87046 10134 87110 10162
rect 87110 10134 87126 10162
rect 87126 10134 87156 10162
<< metal5 >>
rect 38 185370 87806 185412
rect 38 185134 920 185370
rect 1156 185134 84920 185370
rect 85156 185134 87806 185370
rect 38 185092 87806 185134
rect 38 180370 87806 180412
rect 38 180134 2920 180370
rect 3156 180134 81916 180370
rect 82152 180134 86920 180370
rect 87156 180134 87806 180370
rect 38 180092 87806 180134
rect 38 175370 87806 175412
rect 38 175134 920 175370
rect 1156 175134 81470 175370
rect 81706 175134 84920 175370
rect 85156 175134 87806 175370
rect 38 175092 87806 175134
rect 38 170370 87806 170412
rect 38 170134 2920 170370
rect 3156 170134 81916 170370
rect 82152 170134 86920 170370
rect 87156 170134 87806 170370
rect 38 170092 87806 170134
rect 38 165370 87806 165412
rect 38 165134 920 165370
rect 1156 165134 81470 165370
rect 81706 165134 84920 165370
rect 85156 165134 87806 165370
rect 38 165092 87806 165134
rect 38 160370 87806 160412
rect 38 160134 2920 160370
rect 3156 160134 81916 160370
rect 82152 160134 86920 160370
rect 87156 160134 87806 160370
rect 38 160092 87806 160134
rect 38 155370 87806 155412
rect 38 155134 920 155370
rect 1156 155134 81470 155370
rect 81706 155134 84920 155370
rect 85156 155134 87806 155370
rect 38 155092 87806 155134
rect 5490 151892 82538 151934
rect 5490 151656 5532 151892
rect 5768 151656 82260 151892
rect 82496 151656 82538 151892
rect 5490 151614 82538 151656
rect 38 150370 87806 150412
rect 38 150134 2920 150370
rect 3156 150134 81916 150370
rect 82152 150134 86920 150370
rect 87156 150134 87806 150370
rect 38 150092 87806 150134
rect 38 145370 87806 145412
rect 38 145134 920 145370
rect 1156 145134 81470 145370
rect 81706 145134 84920 145370
rect 85156 145134 87806 145370
rect 38 145092 87806 145134
rect 38 140370 87806 140412
rect 38 140134 2920 140370
rect 3156 140134 81916 140370
rect 82152 140134 86920 140370
rect 87156 140134 87806 140370
rect 38 140092 87806 140134
rect 38 135370 87806 135412
rect 38 135134 920 135370
rect 1156 135134 81470 135370
rect 81706 135134 84920 135370
rect 85156 135134 87806 135370
rect 38 135092 87806 135134
rect 38 130370 87806 130412
rect 38 130134 2920 130370
rect 3156 130134 81916 130370
rect 82152 130134 86920 130370
rect 87156 130134 87806 130370
rect 38 130092 87806 130134
rect 38 125370 87806 125412
rect 38 125134 920 125370
rect 1156 125134 81470 125370
rect 81706 125134 84920 125370
rect 85156 125134 87806 125370
rect 38 125092 87806 125134
rect 38 120370 87806 120412
rect 38 120134 2920 120370
rect 3156 120134 81916 120370
rect 82152 120134 86920 120370
rect 87156 120134 87806 120370
rect 38 120092 87806 120134
rect 38 115370 87806 115412
rect 38 115134 920 115370
rect 1156 115134 81470 115370
rect 81706 115134 84920 115370
rect 85156 115134 87806 115370
rect 38 115092 87806 115134
rect 38 110370 87806 110412
rect 38 110134 2920 110370
rect 3156 110134 81916 110370
rect 82152 110134 86920 110370
rect 87156 110134 87806 110370
rect 38 110092 87806 110134
rect 38 105370 87806 105412
rect 38 105134 920 105370
rect 1156 105134 81470 105370
rect 81706 105134 84920 105370
rect 85156 105134 87806 105370
rect 38 105092 87806 105134
rect 38 100370 87806 100412
rect 38 100134 2920 100370
rect 3156 100134 81916 100370
rect 82152 100134 86920 100370
rect 87156 100134 87806 100370
rect 38 100092 87806 100134
rect 38 95370 87806 95412
rect 38 95134 920 95370
rect 1156 95134 84920 95370
rect 85156 95134 87806 95370
rect 38 95092 87806 95134
rect 38 90370 87806 90412
rect 38 90134 2920 90370
rect 3156 90134 81916 90370
rect 82152 90134 86920 90370
rect 87156 90134 87806 90370
rect 38 90092 87806 90134
rect 38 85370 87806 85412
rect 38 85134 920 85370
rect 1156 85134 81470 85370
rect 81706 85134 84920 85370
rect 85156 85134 87806 85370
rect 38 85092 87806 85134
rect 38 80370 87806 80412
rect 38 80134 2920 80370
rect 3156 80134 81916 80370
rect 82152 80134 86920 80370
rect 87156 80134 87806 80370
rect 38 80092 87806 80134
rect 38 75370 87806 75412
rect 38 75134 920 75370
rect 1156 75134 81470 75370
rect 81706 75134 84920 75370
rect 85156 75134 87806 75370
rect 38 75092 87806 75134
rect 38 70370 87806 70412
rect 38 70134 2920 70370
rect 3156 70134 81916 70370
rect 82152 70134 86920 70370
rect 87156 70134 87806 70370
rect 38 70092 87806 70134
rect 38 65370 87806 65412
rect 38 65134 920 65370
rect 1156 65134 81470 65370
rect 81706 65134 84920 65370
rect 85156 65134 87806 65370
rect 38 65092 87806 65134
rect 38 60370 87806 60412
rect 38 60134 2920 60370
rect 3156 60134 81916 60370
rect 82152 60134 86920 60370
rect 87156 60134 87806 60370
rect 38 60092 87806 60134
rect 38 55370 87806 55412
rect 38 55134 920 55370
rect 1156 55134 81470 55370
rect 81706 55134 84920 55370
rect 85156 55134 87806 55370
rect 38 55092 87806 55134
rect 38 50370 87806 50412
rect 38 50134 2920 50370
rect 3156 50134 81916 50370
rect 82152 50134 86920 50370
rect 87156 50134 87806 50370
rect 38 50092 87806 50134
rect 38 45370 87806 45412
rect 38 45134 920 45370
rect 1156 45134 81470 45370
rect 81706 45134 84920 45370
rect 85156 45134 87806 45370
rect 38 45092 87806 45134
rect 38 40370 87806 40412
rect 38 40134 2920 40370
rect 3156 40134 81916 40370
rect 82152 40134 86920 40370
rect 87156 40134 87806 40370
rect 38 40092 87806 40134
rect 38 35370 87806 35412
rect 38 35134 920 35370
rect 1156 35134 81470 35370
rect 81706 35134 84920 35370
rect 85156 35134 87806 35370
rect 38 35092 87806 35134
rect 38 30370 87806 30412
rect 38 30134 2920 30370
rect 3156 30134 81916 30370
rect 82152 30134 86920 30370
rect 87156 30134 87806 30370
rect 38 30092 87806 30134
rect 5490 29492 85666 29534
rect 5490 29256 5532 29492
rect 5768 29256 85388 29492
rect 85624 29256 85666 29492
rect 5490 29214 85666 29256
rect 5490 28132 85666 28174
rect 5490 27896 5532 28132
rect 5768 27896 85388 28132
rect 85624 27896 85666 28132
rect 5490 27854 85666 27896
rect 38 25370 87806 25412
rect 38 25134 920 25370
rect 1156 25134 81470 25370
rect 81706 25134 84920 25370
rect 85156 25134 87806 25370
rect 38 25092 87806 25134
rect 38 20370 87806 20412
rect 38 20134 2920 20370
rect 3156 20134 81916 20370
rect 82152 20134 86920 20370
rect 87156 20134 87806 20370
rect 38 20092 87806 20134
rect 38 15370 87806 15412
rect 38 15134 920 15370
rect 1156 15134 81470 15370
rect 81706 15134 84920 15370
rect 85156 15134 87806 15370
rect 38 15092 87806 15134
rect 38 10370 87806 10412
rect 38 10134 2920 10370
rect 3156 10134 81916 10370
rect 82152 10134 86920 10370
rect 87156 10134 87806 10370
rect 38 10092 87806 10134
rect 38 5370 87806 5412
rect 38 5134 920 5370
rect 1156 5134 81470 5370
rect 81706 5134 84920 5370
rect 85156 5134 87806 5370
rect 38 5092 87806 5134
use sky130_fd_sc_hd__decap_3  PHY_0 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 38 0 1 2514
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_680
timestamp 1604489732
transform 1 0 38 0 -1 2514
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[7] /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 866 0 1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[9]
timestamp 1604489732
transform 1 0 498 0 1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 314 0 1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_7
timestamp 1604489732
transform 1 0 682 0 1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[17]
timestamp 1604489732
transform 1 0 1602 0 1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[4]
timestamp 1604489732
transform 1 0 1234 0 1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[8]
timestamp 1604489732
transform 1 0 1602 0 -1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15
timestamp 1604489732
transform 1 0 1418 0 -1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19
timestamp 1604489732
transform 1 0 1786 0 -1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_11
timestamp 1604489732
transform 1 0 1050 0 1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_15
timestamp 1604489732
transform 1 0 1418 0 1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_19
timestamp 1604489732
transform 1 0 1786 0 1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 314 0 -1 2514
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_19
timestamp 1604489732
transform 1 0 1786 0 -1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_15
timestamp 1604489732
transform 1 0 1418 0 -1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_11
timestamp 1604489732
transform 1 0 1050 0 -1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 314 0 -1 3602
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_wmask0[1]
timestamp 1604489732
transform 1 0 1234 0 -1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[6]
timestamp 1604489732
transform 1 0 1602 0 -1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604489732
transform 1 0 38 0 -1 3602
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_15 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 1418 0 1 3602
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604489732
transform 1 0 314 0 1 3602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604489732
transform 1 0 38 0 1 3602
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_23
timestamp 1604489732
transform 1 0 2154 0 1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23
timestamp 1604489732
transform 1 0 2154 0 -1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[3]
timestamp 1604489732
transform 1 0 1970 0 -1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[15]
timestamp 1604489732
transform 1 0 1970 0 1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_27
timestamp 1604489732
transform 1 0 2522 0 1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27
timestamp 1604489732
transform 1 0 2522 0 -1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[1]
timestamp 1604489732
transform 1 0 2338 0 -1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[16]
timestamp 1604489732
transform 1 0 2706 0 -1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[12]
timestamp 1604489732
transform 1 0 2338 0 1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[11]
timestamp 1604489732
transform 1 0 2706 0 1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_31
timestamp 1604489732
transform 1 0 2890 0 1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 2982 0 -1 2514
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[0]
timestamp 1604489732
transform 1 0 3074 0 1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1534 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 2890 0 -1 2514
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_35
timestamp 1604489732
transform 1 0 3258 0 1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 3350 0 -1 2514
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[10]
timestamp 1604489732
transform 1 0 3442 0 -1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr0[0]
timestamp 1604489732
transform 1 0 3442 0 1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_23
timestamp 1604489732
transform 1 0 2154 0 -1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[2]
timestamp 1604489732
transform 1 0 1970 0 -1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1604489732
transform 1 0 2522 0 -1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[19]
timestamp 1604489732
transform 1 0 2338 0 -1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[14]
timestamp 1604489732
transform 1 0 2706 0 -1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_32
timestamp 1604489732
transform 1 0 2982 0 -1 3602
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1364
timestamp 1604489732
transform 1 0 2890 0 -1 3602
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_36
timestamp 1604489732
transform 1 0 3350 0 -1 3602
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_clk0
timestamp 1604489732
transform 1 0 3442 0 -1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_23
timestamp 1604489732
transform 1 0 2154 0 1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_wmask0[0]
timestamp 1604489732
transform 1 0 1970 0 1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_27
timestamp 1604489732
transform 1 0 2522 0 1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[5]
timestamp 1604489732
transform 1 0 2338 0 1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[21]
timestamp 1604489732
transform 1 0 2706 0 1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_31
timestamp 1604489732
transform 1 0 2890 0 1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[18]
timestamp 1604489732
transform 1 0 3074 0 1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_35
timestamp 1604489732
transform 1 0 3258 0 1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[13]
timestamp 1604489732
transform 1 0 3442 0 1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604489732
transform -1 0 3902 0 1 2514
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604489732
transform -1 0 3902 0 -1 3602
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604489732
transform -1 0 3902 0 1 3602
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_681
timestamp 1604489732
transform -1 0 3902 0 -1 2514
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_682
timestamp 1604489732
transform 1 0 83298 0 -1 2514
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_684
timestamp 1604489732
transform 1 0 83298 0 1 2514
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[22]
timestamp 1604489732
transform 1 0 83758 0 1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[24]
timestamp 1604489732
transform 1 0 84126 0 1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[25]
timestamp 1604489732
transform 1 0 83758 0 -1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[29]
timestamp 1604489732
transform 1 0 84126 0 -1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_908
timestamp 1604489732
transform 1 0 83574 0 -1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_912
timestamp 1604489732
transform 1 0 83942 0 -1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_908
timestamp 1604489732
transform 1 0 83574 0 1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_912
timestamp 1604489732
transform 1 0 83942 0 1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_916
timestamp 1604489732
transform 1 0 84310 0 1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_916
timestamp 1604489732
transform 1 0 84310 0 -1 2514
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_916
timestamp 1604489732
transform 1 0 84310 0 -1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_912
timestamp 1604489732
transform 1 0 83942 0 -1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_908
timestamp 1604489732
transform 1 0 83574 0 -1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[28]
timestamp 1604489732
transform 1 0 84126 0 -1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[23]
timestamp 1604489732
transform 1 0 83758 0 -1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_686
timestamp 1604489732
transform 1 0 83298 0 -1 3602
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_912
timestamp 1604489732
transform 1 0 83942 0 1 3602
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_908
timestamp 1604489732
transform 1 0 83574 0 1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[30]
timestamp 1604489732
transform 1 0 83758 0 1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_688
timestamp 1604489732
transform 1 0 83298 0 1 3602
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[26]
timestamp 1604489732
transform 1 0 84494 0 1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[27]
timestamp 1604489732
transform 1 0 84862 0 1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[31]
timestamp 1604489732
transform 1 0 84494 0 -1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_928
timestamp 1604489732
transform 1 0 85414 0 -1 2514
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_920
timestamp 1604489732
transform 1 0 84678 0 1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_924
timestamp 1604489732
transform 1 0 85046 0 1 2514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_920
timestamp 1604489732
transform 1 0 84678 0 -1 3602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_932
timestamp 1604489732
transform 1 0 85782 0 -1 3602
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_924
timestamp 1604489732
transform 1 0 85046 0 1 3602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_948
timestamp 1604489732
transform 1 0 87254 0 1 2514
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_936
timestamp 1604489732
transform 1 0 86150 0 1 2514
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_949
timestamp 1604489732
transform 1 0 87346 0 -1 2514
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_937
timestamp 1604489732
transform 1 0 86242 0 -1 2514
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1535
timestamp 1604489732
transform 1 0 86150 0 -1 2514
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_685
timestamp 1604489732
transform -1 0 87806 0 1 2514
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_683
timestamp 1604489732
transform -1 0 87806 0 -1 2514
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_949
timestamp 1604489732
transform 1 0 87346 0 -1 3602
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_937
timestamp 1604489732
transform 1 0 86242 0 -1 3602
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1536
timestamp 1604489732
transform 1 0 86150 0 -1 3602
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_687
timestamp 1604489732
transform -1 0 87806 0 -1 3602
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_948
timestamp 1604489732
transform 1 0 87254 0 1 3602
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_936
timestamp 1604489732
transform 1 0 86150 0 1 3602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_689
timestamp 1604489732
transform -1 0 87806 0 1 3602
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604489732
transform 1 0 38 0 -1 4690
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604489732
transform 1 0 38 0 1 4690
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604489732
transform 1 0 38 0 -1 5778
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604489732
transform 1 0 314 0 -1 4690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604489732
transform 1 0 1418 0 -1 4690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604489732
transform 1 0 314 0 1 4690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604489732
transform 1 0 1418 0 1 4690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604489732
transform 1 0 314 0 -1 5778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1604489732
transform 1 0 1418 0 -1 5778
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1604489732
transform 1 0 2522 0 -1 4690
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_36
timestamp 1604489732
transform 1 0 3350 0 -1 4690
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_32
timestamp 1604489732
transform 1 0 2982 0 -1 4690
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_wmask0[3]
timestamp 1604489732
transform 1 0 2706 0 -1 4690
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[20]
timestamp 1604489732
transform 1 0 3442 0 -1 4690
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1365
timestamp 1604489732
transform 1 0 2890 0 -1 4690
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_27
timestamp 1604489732
transform 1 0 2522 0 1 4690
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_35
timestamp 1604489732
transform 1 0 3258 0 1 4690
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_wmask0[2]
timestamp 1604489732
transform 1 0 3442 0 1 4690
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1604489732
transform 1 0 2522 0 -1 5778
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_32
timestamp 1604489732
transform 1 0 2982 0 -1 5778
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1366
timestamp 1604489732
transform 1 0 2890 0 -1 5778
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_38
timestamp 1604489732
transform 1 0 3534 0 -1 5778
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604489732
transform -1 0 3902 0 -1 4690
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604489732
transform -1 0 3902 0 1 4690
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604489732
transform -1 0 3902 0 -1 5778
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_690
timestamp 1604489732
transform 1 0 83298 0 -1 4690
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_692
timestamp 1604489732
transform 1 0 83298 0 1 4690
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_694
timestamp 1604489732
transform 1 0 83298 0 -1 5778
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_908
timestamp 1604489732
transform 1 0 83574 0 -1 4690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_908
timestamp 1604489732
transform 1 0 83574 0 1 4690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_908
timestamp 1604489732
transform 1 0 83574 0 -1 5778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_920
timestamp 1604489732
transform 1 0 84678 0 -1 4690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_932
timestamp 1604489732
transform 1 0 85782 0 -1 4690
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_920
timestamp 1604489732
transform 1 0 84678 0 1 4690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_932
timestamp 1604489732
transform 1 0 85782 0 1 4690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_920
timestamp 1604489732
transform 1 0 84678 0 -1 5778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_932
timestamp 1604489732
transform 1 0 85782 0 -1 5778
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_949
timestamp 1604489732
transform 1 0 87346 0 -1 4690
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_937
timestamp 1604489732
transform 1 0 86242 0 -1 4690
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1537
timestamp 1604489732
transform 1 0 86150 0 -1 4690
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_691
timestamp 1604489732
transform -1 0 87806 0 -1 4690
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_950
timestamp 1604489732
transform 1 0 87438 0 1 4690
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_944
timestamp 1604489732
transform 1 0 86886 0 1 4690
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_693
timestamp 1604489732
transform -1 0 87806 0 1 4690
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_949
timestamp 1604489732
transform 1 0 87346 0 -1 5778
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_937
timestamp 1604489732
transform 1 0 86242 0 -1 5778
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1538
timestamp 1604489732
transform 1 0 86150 0 -1 5778
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_695
timestamp 1604489732
transform -1 0 87806 0 -1 5778
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604489732
transform 1 0 38 0 1 5778
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604489732
transform 1 0 38 0 -1 6866
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604489732
transform 1 0 38 0 1 6866
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604489732
transform 1 0 314 0 1 5778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604489732
transform 1 0 1418 0 1 5778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604489732
transform 1 0 314 0 -1 6866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604489732
transform 1 0 1418 0 -1 6866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1604489732
transform 1 0 314 0 1 6866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1604489732
transform 1 0 1418 0 1 6866
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1367
timestamp 1604489732
transform 1 0 2890 0 -1 6866
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1604489732
transform 1 0 2522 0 1 5778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1604489732
transform 1 0 2522 0 -1 6866
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_32
timestamp 1604489732
transform 1 0 2982 0 -1 6866
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_38
timestamp 1604489732
transform 1 0 3534 0 -1 6866
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1604489732
transform 1 0 2522 0 1 6866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604489732
transform -1 0 3902 0 1 5778
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604489732
transform -1 0 3902 0 -1 6866
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604489732
transform -1 0 3902 0 1 6866
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_696
timestamp 1604489732
transform 1 0 83298 0 1 5778
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_698
timestamp 1604489732
transform 1 0 83298 0 -1 6866
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_700
timestamp 1604489732
transform 1 0 83298 0 1 6866
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_908
timestamp 1604489732
transform 1 0 83574 0 1 5778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_908
timestamp 1604489732
transform 1 0 83574 0 -1 6866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_908
timestamp 1604489732
transform 1 0 83574 0 1 6866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_920
timestamp 1604489732
transform 1 0 84678 0 1 5778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_932
timestamp 1604489732
transform 1 0 85782 0 1 5778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_920
timestamp 1604489732
transform 1 0 84678 0 -1 6866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_932
timestamp 1604489732
transform 1 0 85782 0 -1 6866
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_920
timestamp 1604489732
transform 1 0 84678 0 1 6866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_932
timestamp 1604489732
transform 1 0 85782 0 1 6866
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_950
timestamp 1604489732
transform 1 0 87438 0 1 5778
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_944
timestamp 1604489732
transform 1 0 86886 0 1 5778
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_697
timestamp 1604489732
transform -1 0 87806 0 1 5778
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_949
timestamp 1604489732
transform 1 0 87346 0 -1 6866
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_937
timestamp 1604489732
transform 1 0 86242 0 -1 6866
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1539
timestamp 1604489732
transform 1 0 86150 0 -1 6866
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_699
timestamp 1604489732
transform -1 0 87806 0 -1 6866
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_950
timestamp 1604489732
transform 1 0 87438 0 1 6866
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_944
timestamp 1604489732
transform 1 0 86886 0 1 6866
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_701
timestamp 1604489732
transform -1 0 87806 0 1 6866
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1604489732
transform 1 0 1418 0 1 7954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1604489732
transform 1 0 314 0 1 7954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1604489732
transform 1 0 1418 0 -1 7954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604489732
transform 1 0 314 0 -1 7954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604489732
transform 1 0 38 0 1 7954
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604489732
transform 1 0 38 0 -1 7954
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1604489732
transform 1 0 1418 0 -1 9042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1604489732
transform 1 0 314 0 -1 9042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604489732
transform 1 0 38 0 -1 9042
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1604489732
transform 1 0 1418 0 1 9042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1604489732
transform 1 0 314 0 1 9042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604489732
transform 1 0 38 0 1 9042
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1604489732
transform 1 0 2522 0 1 7954
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_38
timestamp 1604489732
transform 1 0 3534 0 -1 7954
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_32
timestamp 1604489732
transform 1 0 2982 0 -1 7954
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1604489732
transform 1 0 2522 0 -1 7954
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1368
timestamp 1604489732
transform 1 0 2890 0 -1 7954
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_38
timestamp 1604489732
transform 1 0 3534 0 -1 9042
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_32
timestamp 1604489732
transform 1 0 2982 0 -1 9042
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1604489732
transform 1 0 2522 0 -1 9042
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1369
timestamp 1604489732
transform 1 0 2890 0 -1 9042
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1604489732
transform 1 0 2522 0 1 9042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604489732
transform -1 0 3902 0 -1 7954
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604489732
transform -1 0 3902 0 1 7954
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604489732
transform -1 0 3902 0 -1 9042
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604489732
transform -1 0 3902 0 1 9042
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_702
timestamp 1604489732
transform 1 0 83298 0 -1 7954
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_704
timestamp 1604489732
transform 1 0 83298 0 1 7954
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_706
timestamp 1604489732
transform 1 0 83298 0 -1 9042
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_708
timestamp 1604489732
transform 1 0 83298 0 1 9042
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_908
timestamp 1604489732
transform 1 0 83574 0 -1 7954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_908
timestamp 1604489732
transform 1 0 83574 0 1 7954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_908
timestamp 1604489732
transform 1 0 83574 0 -1 9042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_908
timestamp 1604489732
transform 1 0 83574 0 1 9042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_920
timestamp 1604489732
transform 1 0 84678 0 -1 7954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_932
timestamp 1604489732
transform 1 0 85782 0 -1 7954
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_920
timestamp 1604489732
transform 1 0 84678 0 1 7954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_932
timestamp 1604489732
transform 1 0 85782 0 1 7954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_920
timestamp 1604489732
transform 1 0 84678 0 -1 9042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_932
timestamp 1604489732
transform 1 0 85782 0 -1 9042
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_920
timestamp 1604489732
transform 1 0 84678 0 1 9042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_932
timestamp 1604489732
transform 1 0 85782 0 1 9042
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_950
timestamp 1604489732
transform 1 0 87438 0 1 7954
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_944
timestamp 1604489732
transform 1 0 86886 0 1 7954
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_949
timestamp 1604489732
transform 1 0 87346 0 -1 7954
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_937
timestamp 1604489732
transform 1 0 86242 0 -1 7954
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1540
timestamp 1604489732
transform 1 0 86150 0 -1 7954
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_705
timestamp 1604489732
transform -1 0 87806 0 1 7954
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_703
timestamp 1604489732
transform -1 0 87806 0 -1 7954
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_949
timestamp 1604489732
transform 1 0 87346 0 -1 9042
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_937
timestamp 1604489732
transform 1 0 86242 0 -1 9042
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1541
timestamp 1604489732
transform 1 0 86150 0 -1 9042
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_707
timestamp 1604489732
transform -1 0 87806 0 -1 9042
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_950
timestamp 1604489732
transform 1 0 87438 0 1 9042
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_944
timestamp 1604489732
transform 1 0 86886 0 1 9042
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_709
timestamp 1604489732
transform -1 0 87806 0 1 9042
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604489732
transform 1 0 38 0 -1 10130
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604489732
transform 1 0 38 0 1 10130
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604489732
transform 1 0 38 0 -1 11218
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1604489732
transform 1 0 314 0 -1 10130
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1604489732
transform 1 0 1418 0 -1 10130
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1604489732
transform 1 0 314 0 1 10130
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1604489732
transform 1 0 1418 0 1 10130
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1604489732
transform 1 0 314 0 -1 11218
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1604489732
transform 1 0 1418 0 -1 11218
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1370
timestamp 1604489732
transform 1 0 2890 0 -1 10130
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1371
timestamp 1604489732
transform 1 0 2890 0 -1 11218
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1604489732
transform 1 0 2522 0 -1 10130
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_32
timestamp 1604489732
transform 1 0 2982 0 -1 10130
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_38
timestamp 1604489732
transform 1 0 3534 0 -1 10130
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1604489732
transform 1 0 2522 0 1 10130
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1604489732
transform 1 0 2522 0 -1 11218
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_32
timestamp 1604489732
transform 1 0 2982 0 -1 11218
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_38
timestamp 1604489732
transform 1 0 3534 0 -1 11218
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604489732
transform -1 0 3902 0 -1 10130
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604489732
transform -1 0 3902 0 1 10130
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604489732
transform -1 0 3902 0 -1 11218
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_710
timestamp 1604489732
transform 1 0 83298 0 -1 10130
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_712
timestamp 1604489732
transform 1 0 83298 0 1 10130
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_714
timestamp 1604489732
transform 1 0 83298 0 -1 11218
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_908
timestamp 1604489732
transform 1 0 83574 0 -1 10130
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_908
timestamp 1604489732
transform 1 0 83574 0 1 10130
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_908
timestamp 1604489732
transform 1 0 83574 0 -1 11218
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_920
timestamp 1604489732
transform 1 0 84678 0 -1 10130
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_932
timestamp 1604489732
transform 1 0 85782 0 -1 10130
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_920
timestamp 1604489732
transform 1 0 84678 0 1 10130
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_932
timestamp 1604489732
transform 1 0 85782 0 1 10130
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_920
timestamp 1604489732
transform 1 0 84678 0 -1 11218
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_932
timestamp 1604489732
transform 1 0 85782 0 -1 11218
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_949
timestamp 1604489732
transform 1 0 87346 0 -1 10130
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_937
timestamp 1604489732
transform 1 0 86242 0 -1 10130
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1542
timestamp 1604489732
transform 1 0 86150 0 -1 10130
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_711
timestamp 1604489732
transform -1 0 87806 0 -1 10130
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_950
timestamp 1604489732
transform 1 0 87438 0 1 10130
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_944
timestamp 1604489732
transform 1 0 86886 0 1 10130
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_713
timestamp 1604489732
transform -1 0 87806 0 1 10130
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_949
timestamp 1604489732
transform 1 0 87346 0 -1 11218
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_937
timestamp 1604489732
transform 1 0 86242 0 -1 11218
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1543
timestamp 1604489732
transform 1 0 86150 0 -1 11218
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_715
timestamp 1604489732
transform -1 0 87806 0 -1 11218
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604489732
transform 1 0 38 0 1 11218
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604489732
transform 1 0 38 0 -1 12306
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604489732
transform 1 0 38 0 1 12306
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1604489732
transform 1 0 314 0 1 11218
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1604489732
transform 1 0 1418 0 1 11218
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1604489732
transform 1 0 314 0 -1 12306
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1604489732
transform 1 0 1418 0 -1 12306
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1604489732
transform 1 0 314 0 1 12306
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1604489732
transform 1 0 1418 0 1 12306
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1372
timestamp 1604489732
transform 1 0 2890 0 -1 12306
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1604489732
transform 1 0 2522 0 1 11218
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1604489732
transform 1 0 2522 0 -1 12306
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_32
timestamp 1604489732
transform 1 0 2982 0 -1 12306
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_38
timestamp 1604489732
transform 1 0 3534 0 -1 12306
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1604489732
transform 1 0 2522 0 1 12306
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604489732
transform -1 0 3902 0 1 11218
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604489732
transform -1 0 3902 0 -1 12306
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604489732
transform -1 0 3902 0 1 12306
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_716
timestamp 1604489732
transform 1 0 83298 0 1 11218
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_718
timestamp 1604489732
transform 1 0 83298 0 -1 12306
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_720
timestamp 1604489732
transform 1 0 83298 0 1 12306
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_908
timestamp 1604489732
transform 1 0 83574 0 1 11218
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_908
timestamp 1604489732
transform 1 0 83574 0 -1 12306
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_908
timestamp 1604489732
transform 1 0 83574 0 1 12306
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_920
timestamp 1604489732
transform 1 0 84678 0 1 11218
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_932
timestamp 1604489732
transform 1 0 85782 0 1 11218
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_920
timestamp 1604489732
transform 1 0 84678 0 -1 12306
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_932
timestamp 1604489732
transform 1 0 85782 0 -1 12306
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_920
timestamp 1604489732
transform 1 0 84678 0 1 12306
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_932
timestamp 1604489732
transform 1 0 85782 0 1 12306
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_950
timestamp 1604489732
transform 1 0 87438 0 1 11218
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_944
timestamp 1604489732
transform 1 0 86886 0 1 11218
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_717
timestamp 1604489732
transform -1 0 87806 0 1 11218
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_949
timestamp 1604489732
transform 1 0 87346 0 -1 12306
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_937
timestamp 1604489732
transform 1 0 86242 0 -1 12306
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1544
timestamp 1604489732
transform 1 0 86150 0 -1 12306
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_719
timestamp 1604489732
transform -1 0 87806 0 -1 12306
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_950
timestamp 1604489732
transform 1 0 87438 0 1 12306
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_944
timestamp 1604489732
transform 1 0 86886 0 1 12306
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_721
timestamp 1604489732
transform -1 0 87806 0 1 12306
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1604489732
transform 1 0 1418 0 -1 13394
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1604489732
transform 1 0 314 0 -1 13394
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604489732
transform 1 0 38 0 -1 13394
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1604489732
transform 1 0 1418 0 -1 14482
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1604489732
transform 1 0 314 0 -1 14482
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1604489732
transform 1 0 1418 0 1 13394
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1604489732
transform 1 0 314 0 1 13394
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604489732
transform 1 0 38 0 -1 14482
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604489732
transform 1 0 38 0 1 13394
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1604489732
transform 1 0 1418 0 1 14482
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1604489732
transform 1 0 314 0 1 14482
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604489732
transform 1 0 38 0 1 14482
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_38
timestamp 1604489732
transform 1 0 3534 0 -1 13394
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_32
timestamp 1604489732
transform 1 0 2982 0 -1 13394
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1604489732
transform 1 0 2522 0 -1 13394
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1373
timestamp 1604489732
transform 1 0 2890 0 -1 13394
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_38
timestamp 1604489732
transform 1 0 3534 0 -1 14482
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_32
timestamp 1604489732
transform 1 0 2982 0 -1 14482
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1604489732
transform 1 0 2522 0 -1 14482
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1604489732
transform 1 0 2522 0 1 13394
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1374
timestamp 1604489732
transform 1 0 2890 0 -1 14482
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1604489732
transform 1 0 2522 0 1 14482
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604489732
transform -1 0 3902 0 -1 13394
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604489732
transform -1 0 3902 0 1 13394
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604489732
transform -1 0 3902 0 -1 14482
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604489732
transform -1 0 3902 0 1 14482
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_722
timestamp 1604489732
transform 1 0 83298 0 -1 13394
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_724
timestamp 1604489732
transform 1 0 83298 0 1 13394
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_726
timestamp 1604489732
transform 1 0 83298 0 -1 14482
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_728
timestamp 1604489732
transform 1 0 83298 0 1 14482
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_908
timestamp 1604489732
transform 1 0 83574 0 -1 13394
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_908
timestamp 1604489732
transform 1 0 83574 0 1 13394
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_908
timestamp 1604489732
transform 1 0 83574 0 -1 14482
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_908
timestamp 1604489732
transform 1 0 83574 0 1 14482
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_920
timestamp 1604489732
transform 1 0 84678 0 -1 13394
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_932
timestamp 1604489732
transform 1 0 85782 0 -1 13394
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_920
timestamp 1604489732
transform 1 0 84678 0 1 13394
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_932
timestamp 1604489732
transform 1 0 85782 0 1 13394
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_920
timestamp 1604489732
transform 1 0 84678 0 -1 14482
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_932
timestamp 1604489732
transform 1 0 85782 0 -1 14482
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_920
timestamp 1604489732
transform 1 0 84678 0 1 14482
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_932
timestamp 1604489732
transform 1 0 85782 0 1 14482
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_949
timestamp 1604489732
transform 1 0 87346 0 -1 13394
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_937
timestamp 1604489732
transform 1 0 86242 0 -1 13394
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1545
timestamp 1604489732
transform 1 0 86150 0 -1 13394
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_723
timestamp 1604489732
transform -1 0 87806 0 -1 13394
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_949
timestamp 1604489732
transform 1 0 87346 0 -1 14482
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_937
timestamp 1604489732
transform 1 0 86242 0 -1 14482
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_950
timestamp 1604489732
transform 1 0 87438 0 1 13394
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_944
timestamp 1604489732
transform 1 0 86886 0 1 13394
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1546
timestamp 1604489732
transform 1 0 86150 0 -1 14482
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_727
timestamp 1604489732
transform -1 0 87806 0 -1 14482
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_725
timestamp 1604489732
transform -1 0 87806 0 1 13394
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_950
timestamp 1604489732
transform 1 0 87438 0 1 14482
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_944
timestamp 1604489732
transform 1 0 86886 0 1 14482
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_729
timestamp 1604489732
transform -1 0 87806 0 1 14482
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604489732
transform 1 0 38 0 -1 15570
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604489732
transform 1 0 38 0 1 15570
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604489732
transform 1 0 38 0 -1 16658
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1604489732
transform 1 0 314 0 -1 15570
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604489732
transform 1 0 1418 0 -1 15570
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1604489732
transform 1 0 314 0 1 15570
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1604489732
transform 1 0 1418 0 1 15570
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1604489732
transform 1 0 314 0 -1 16658
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1604489732
transform 1 0 1418 0 -1 16658
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1375
timestamp 1604489732
transform 1 0 2890 0 -1 15570
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1376
timestamp 1604489732
transform 1 0 2890 0 -1 16658
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1604489732
transform 1 0 2522 0 -1 15570
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_32
timestamp 1604489732
transform 1 0 2982 0 -1 15570
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_38
timestamp 1604489732
transform 1 0 3534 0 -1 15570
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1604489732
transform 1 0 2522 0 1 15570
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1604489732
transform 1 0 2522 0 -1 16658
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_32
timestamp 1604489732
transform 1 0 2982 0 -1 16658
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_38
timestamp 1604489732
transform 1 0 3534 0 -1 16658
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604489732
transform -1 0 3902 0 -1 15570
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604489732
transform -1 0 3902 0 1 15570
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604489732
transform -1 0 3902 0 -1 16658
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_730
timestamp 1604489732
transform 1 0 83298 0 -1 15570
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_732
timestamp 1604489732
transform 1 0 83298 0 1 15570
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_734
timestamp 1604489732
transform 1 0 83298 0 -1 16658
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_908
timestamp 1604489732
transform 1 0 83574 0 -1 15570
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_908
timestamp 1604489732
transform 1 0 83574 0 1 15570
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_908
timestamp 1604489732
transform 1 0 83574 0 -1 16658
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_920
timestamp 1604489732
transform 1 0 84678 0 -1 15570
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_932
timestamp 1604489732
transform 1 0 85782 0 -1 15570
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_920
timestamp 1604489732
transform 1 0 84678 0 1 15570
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_932
timestamp 1604489732
transform 1 0 85782 0 1 15570
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_920
timestamp 1604489732
transform 1 0 84678 0 -1 16658
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_932
timestamp 1604489732
transform 1 0 85782 0 -1 16658
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_949
timestamp 1604489732
transform 1 0 87346 0 -1 15570
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_937
timestamp 1604489732
transform 1 0 86242 0 -1 15570
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1547
timestamp 1604489732
transform 1 0 86150 0 -1 15570
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_731
timestamp 1604489732
transform -1 0 87806 0 -1 15570
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_950
timestamp 1604489732
transform 1 0 87438 0 1 15570
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_944
timestamp 1604489732
transform 1 0 86886 0 1 15570
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_733
timestamp 1604489732
transform -1 0 87806 0 1 15570
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_949
timestamp 1604489732
transform 1 0 87346 0 -1 16658
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_937
timestamp 1604489732
transform 1 0 86242 0 -1 16658
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1548
timestamp 1604489732
transform 1 0 86150 0 -1 16658
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_735
timestamp 1604489732
transform -1 0 87806 0 -1 16658
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604489732
transform 1 0 38 0 1 16658
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604489732
transform 1 0 38 0 -1 17746
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604489732
transform 1 0 38 0 1 17746
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1604489732
transform 1 0 314 0 1 16658
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1604489732
transform 1 0 1418 0 1 16658
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1604489732
transform 1 0 314 0 -1 17746
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1604489732
transform 1 0 1418 0 -1 17746
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1604489732
transform 1 0 314 0 1 17746
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1604489732
transform 1 0 1418 0 1 17746
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1377
timestamp 1604489732
transform 1 0 2890 0 -1 17746
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1604489732
transform 1 0 2522 0 1 16658
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1604489732
transform 1 0 2522 0 -1 17746
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_32
timestamp 1604489732
transform 1 0 2982 0 -1 17746
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_38
timestamp 1604489732
transform 1 0 3534 0 -1 17746
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1604489732
transform 1 0 2522 0 1 17746
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604489732
transform -1 0 3902 0 1 16658
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604489732
transform -1 0 3902 0 -1 17746
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604489732
transform -1 0 3902 0 1 17746
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_736
timestamp 1604489732
transform 1 0 83298 0 1 16658
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_738
timestamp 1604489732
transform 1 0 83298 0 -1 17746
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_740
timestamp 1604489732
transform 1 0 83298 0 1 17746
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_908
timestamp 1604489732
transform 1 0 83574 0 1 16658
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_908
timestamp 1604489732
transform 1 0 83574 0 -1 17746
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_908
timestamp 1604489732
transform 1 0 83574 0 1 17746
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_920
timestamp 1604489732
transform 1 0 84678 0 1 16658
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_932
timestamp 1604489732
transform 1 0 85782 0 1 16658
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_920
timestamp 1604489732
transform 1 0 84678 0 -1 17746
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_932
timestamp 1604489732
transform 1 0 85782 0 -1 17746
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_920
timestamp 1604489732
transform 1 0 84678 0 1 17746
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_932
timestamp 1604489732
transform 1 0 85782 0 1 17746
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_950
timestamp 1604489732
transform 1 0 87438 0 1 16658
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_944
timestamp 1604489732
transform 1 0 86886 0 1 16658
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_737
timestamp 1604489732
transform -1 0 87806 0 1 16658
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_949
timestamp 1604489732
transform 1 0 87346 0 -1 17746
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_937
timestamp 1604489732
transform 1 0 86242 0 -1 17746
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1549
timestamp 1604489732
transform 1 0 86150 0 -1 17746
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_739
timestamp 1604489732
transform -1 0 87806 0 -1 17746
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_950
timestamp 1604489732
transform 1 0 87438 0 1 17746
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_944
timestamp 1604489732
transform 1 0 86886 0 1 17746
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_741
timestamp 1604489732
transform -1 0 87806 0 1 17746
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604489732
transform 1 0 38 0 -1 18834
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604489732
transform 1 0 38 0 1 18834
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604489732
transform 1 0 38 0 -1 19922
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1604489732
transform 1 0 314 0 -1 18834
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1604489732
transform 1 0 1418 0 -1 18834
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604489732
transform 1 0 314 0 1 18834
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1604489732
transform 1 0 1418 0 1 18834
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604489732
transform 1 0 314 0 -1 19922
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1604489732
transform 1 0 1418 0 -1 19922
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1378
timestamp 1604489732
transform 1 0 2890 0 -1 18834
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1379
timestamp 1604489732
transform 1 0 2890 0 -1 19922
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1604489732
transform 1 0 2522 0 -1 18834
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_32
timestamp 1604489732
transform 1 0 2982 0 -1 18834
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_38
timestamp 1604489732
transform 1 0 3534 0 -1 18834
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1604489732
transform 1 0 2522 0 1 18834
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1604489732
transform 1 0 2522 0 -1 19922
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_32
timestamp 1604489732
transform 1 0 2982 0 -1 19922
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_38
timestamp 1604489732
transform 1 0 3534 0 -1 19922
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604489732
transform -1 0 3902 0 -1 18834
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604489732
transform -1 0 3902 0 1 18834
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604489732
transform -1 0 3902 0 -1 19922
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_742
timestamp 1604489732
transform 1 0 83298 0 -1 18834
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_744
timestamp 1604489732
transform 1 0 83298 0 1 18834
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_746
timestamp 1604489732
transform 1 0 83298 0 -1 19922
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_908
timestamp 1604489732
transform 1 0 83574 0 -1 18834
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_908
timestamp 1604489732
transform 1 0 83574 0 1 18834
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_908
timestamp 1604489732
transform 1 0 83574 0 -1 19922
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_920
timestamp 1604489732
transform 1 0 84678 0 -1 18834
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_932
timestamp 1604489732
transform 1 0 85782 0 -1 18834
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_920
timestamp 1604489732
transform 1 0 84678 0 1 18834
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_932
timestamp 1604489732
transform 1 0 85782 0 1 18834
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_920
timestamp 1604489732
transform 1 0 84678 0 -1 19922
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_932
timestamp 1604489732
transform 1 0 85782 0 -1 19922
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_949
timestamp 1604489732
transform 1 0 87346 0 -1 18834
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_937
timestamp 1604489732
transform 1 0 86242 0 -1 18834
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1550
timestamp 1604489732
transform 1 0 86150 0 -1 18834
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_743
timestamp 1604489732
transform -1 0 87806 0 -1 18834
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_949
timestamp 1604489732
transform 1 0 87346 0 -1 19922
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_937
timestamp 1604489732
transform 1 0 86242 0 -1 19922
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_950
timestamp 1604489732
transform 1 0 87438 0 1 18834
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_944
timestamp 1604489732
transform 1 0 86886 0 1 18834
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1551
timestamp 1604489732
transform 1 0 86150 0 -1 19922
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_747
timestamp 1604489732
transform -1 0 87806 0 -1 19922
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_745
timestamp 1604489732
transform -1 0 87806 0 1 18834
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604489732
transform 1 0 1418 0 -1 21010
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604489732
transform 1 0 314 0 -1 21010
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604489732
transform 1 0 1418 0 1 19922
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604489732
transform 1 0 314 0 1 19922
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604489732
transform 1 0 38 0 -1 21010
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604489732
transform 1 0 38 0 1 19922
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604489732
transform 1 0 1418 0 1 21010
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604489732
transform 1 0 314 0 1 21010
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604489732
transform 1 0 38 0 1 21010
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1604489732
transform 1 0 1418 0 -1 22098
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1604489732
transform 1 0 314 0 -1 22098
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604489732
transform 1 0 38 0 -1 22098
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_36
timestamp 1604489732
transform 1 0 3350 0 -1 21010
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_32
timestamp 1604489732
transform 1 0 2982 0 -1 21010
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1604489732
transform 1 0 2522 0 -1 21010
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1604489732
transform 1 0 2522 0 1 19922
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_csb0
timestamp 1604489732
transform 1 0 3442 0 -1 21010
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1380
timestamp 1604489732
transform 1 0 2890 0 -1 21010
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1604489732
transform 1 0 2522 0 1 21010
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_38
timestamp 1604489732
transform 1 0 3534 0 -1 22098
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_32
timestamp 1604489732
transform 1 0 2982 0 -1 22098
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1604489732
transform 1 0 2522 0 -1 22098
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1381
timestamp 1604489732
transform 1 0 2890 0 -1 22098
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604489732
transform -1 0 3902 0 1 19922
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604489732
transform -1 0 3902 0 -1 21010
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604489732
transform -1 0 3902 0 1 21010
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604489732
transform -1 0 3902 0 -1 22098
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_748
timestamp 1604489732
transform 1 0 83298 0 1 19922
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_750
timestamp 1604489732
transform 1 0 83298 0 -1 21010
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_752
timestamp 1604489732
transform 1 0 83298 0 1 21010
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_754
timestamp 1604489732
transform 1 0 83298 0 -1 22098
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_908
timestamp 1604489732
transform 1 0 83574 0 1 19922
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_908
timestamp 1604489732
transform 1 0 83574 0 -1 21010
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_908
timestamp 1604489732
transform 1 0 83574 0 1 21010
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_908
timestamp 1604489732
transform 1 0 83574 0 -1 22098
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_920
timestamp 1604489732
transform 1 0 84678 0 1 19922
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_932
timestamp 1604489732
transform 1 0 85782 0 1 19922
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_920
timestamp 1604489732
transform 1 0 84678 0 -1 21010
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_932
timestamp 1604489732
transform 1 0 85782 0 -1 21010
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_920
timestamp 1604489732
transform 1 0 84678 0 1 21010
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_932
timestamp 1604489732
transform 1 0 85782 0 1 21010
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_920
timestamp 1604489732
transform 1 0 84678 0 -1 22098
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_932
timestamp 1604489732
transform 1 0 85782 0 -1 22098
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_949
timestamp 1604489732
transform 1 0 87346 0 -1 21010
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_937
timestamp 1604489732
transform 1 0 86242 0 -1 21010
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_950
timestamp 1604489732
transform 1 0 87438 0 1 19922
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_944
timestamp 1604489732
transform 1 0 86886 0 1 19922
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1552
timestamp 1604489732
transform 1 0 86150 0 -1 21010
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_751
timestamp 1604489732
transform -1 0 87806 0 -1 21010
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_749
timestamp 1604489732
transform -1 0 87806 0 1 19922
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_950
timestamp 1604489732
transform 1 0 87438 0 1 21010
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_944
timestamp 1604489732
transform 1 0 86886 0 1 21010
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_753
timestamp 1604489732
transform -1 0 87806 0 1 21010
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_949
timestamp 1604489732
transform 1 0 87346 0 -1 22098
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_937
timestamp 1604489732
transform 1 0 86242 0 -1 22098
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1553
timestamp 1604489732
transform 1 0 86150 0 -1 22098
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_755
timestamp 1604489732
transform -1 0 87806 0 -1 22098
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604489732
transform 1 0 38 0 1 22098
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604489732
transform 1 0 38 0 -1 23186
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604489732
transform 1 0 38 0 1 23186
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1604489732
transform 1 0 314 0 1 22098
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1604489732
transform 1 0 1418 0 1 22098
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1604489732
transform 1 0 314 0 -1 23186
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1604489732
transform 1 0 1418 0 -1 23186
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1604489732
transform 1 0 314 0 1 23186
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1604489732
transform 1 0 1418 0 1 23186
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1382
timestamp 1604489732
transform 1 0 2890 0 -1 23186
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_web0
timestamp 1604489732
transform 1 0 3442 0 1 22098
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_27
timestamp 1604489732
transform 1 0 2522 0 1 22098
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_35
timestamp 1604489732
transform 1 0 3258 0 1 22098
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1604489732
transform 1 0 2522 0 -1 23186
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_32
timestamp 1604489732
transform 1 0 2982 0 -1 23186
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_38
timestamp 1604489732
transform 1 0 3534 0 -1 23186
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1604489732
transform 1 0 2522 0 1 23186
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604489732
transform -1 0 3902 0 1 22098
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604489732
transform -1 0 3902 0 -1 23186
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604489732
transform -1 0 3902 0 1 23186
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_756
timestamp 1604489732
transform 1 0 83298 0 1 22098
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_758
timestamp 1604489732
transform 1 0 83298 0 -1 23186
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_760
timestamp 1604489732
transform 1 0 83298 0 1 23186
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr1[7]
timestamp 1604489732
transform 1 0 83758 0 -1 23186
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_908
timestamp 1604489732
transform 1 0 83574 0 1 22098
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_908
timestamp 1604489732
transform 1 0 83574 0 -1 23186
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_912
timestamp 1604489732
transform 1 0 83942 0 -1 23186
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_908
timestamp 1604489732
transform 1 0 83574 0 1 23186
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_920
timestamp 1604489732
transform 1 0 84678 0 1 22098
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_932
timestamp 1604489732
transform 1 0 85782 0 1 22098
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_924
timestamp 1604489732
transform 1 0 85046 0 -1 23186
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_920
timestamp 1604489732
transform 1 0 84678 0 1 23186
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_932
timestamp 1604489732
transform 1 0 85782 0 1 23186
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_950
timestamp 1604489732
transform 1 0 87438 0 1 22098
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_944
timestamp 1604489732
transform 1 0 86886 0 1 22098
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_757
timestamp 1604489732
transform -1 0 87806 0 1 22098
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_949
timestamp 1604489732
transform 1 0 87346 0 -1 23186
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_937
timestamp 1604489732
transform 1 0 86242 0 -1 23186
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1554
timestamp 1604489732
transform 1 0 86150 0 -1 23186
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_759
timestamp 1604489732
transform -1 0 87806 0 -1 23186
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_39_950
timestamp 1604489732
transform 1 0 87438 0 1 23186
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_944
timestamp 1604489732
transform 1 0 86886 0 1 23186
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_761
timestamp 1604489732
transform -1 0 87806 0 1 23186
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604489732
transform 1 0 38 0 -1 24274
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604489732
transform 1 0 38 0 1 24274
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604489732
transform 1 0 38 0 -1 25362
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1604489732
transform 1 0 314 0 -1 24274
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1604489732
transform 1 0 1418 0 -1 24274
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1604489732
transform 1 0 314 0 1 24274
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1604489732
transform 1 0 1418 0 1 24274
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1604489732
transform 1 0 314 0 -1 25362
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1604489732
transform 1 0 1418 0 -1 25362
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1383
timestamp 1604489732
transform 1 0 2890 0 -1 24274
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1384
timestamp 1604489732
transform 1 0 2890 0 -1 25362
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1604489732
transform 1 0 2522 0 -1 24274
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_32
timestamp 1604489732
transform 1 0 2982 0 -1 24274
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_38
timestamp 1604489732
transform 1 0 3534 0 -1 24274
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1604489732
transform 1 0 2522 0 1 24274
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1604489732
transform 1 0 2522 0 -1 25362
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_32
timestamp 1604489732
transform 1 0 2982 0 -1 25362
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_38
timestamp 1604489732
transform 1 0 3534 0 -1 25362
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604489732
transform -1 0 3902 0 -1 24274
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604489732
transform -1 0 3902 0 1 24274
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604489732
transform -1 0 3902 0 -1 25362
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_762
timestamp 1604489732
transform 1 0 83298 0 -1 24274
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_764
timestamp 1604489732
transform 1 0 83298 0 1 24274
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_766
timestamp 1604489732
transform 1 0 83298 0 -1 25362
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr1[6]
timestamp 1604489732
transform 1 0 83758 0 -1 24274
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_908
timestamp 1604489732
transform 1 0 83574 0 -1 24274
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_912
timestamp 1604489732
transform 1 0 83942 0 -1 24274
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_908
timestamp 1604489732
transform 1 0 83574 0 1 24274
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_908
timestamp 1604489732
transform 1 0 83574 0 -1 25362
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_924
timestamp 1604489732
transform 1 0 85046 0 -1 24274
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_920
timestamp 1604489732
transform 1 0 84678 0 1 24274
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_932
timestamp 1604489732
transform 1 0 85782 0 1 24274
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_920
timestamp 1604489732
transform 1 0 84678 0 -1 25362
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_932
timestamp 1604489732
transform 1 0 85782 0 -1 25362
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_949
timestamp 1604489732
transform 1 0 87346 0 -1 24274
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_937
timestamp 1604489732
transform 1 0 86242 0 -1 24274
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1555
timestamp 1604489732
transform 1 0 86150 0 -1 24274
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_763
timestamp 1604489732
transform -1 0 87806 0 -1 24274
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_41_950
timestamp 1604489732
transform 1 0 87438 0 1 24274
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_944
timestamp 1604489732
transform 1 0 86886 0 1 24274
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_765
timestamp 1604489732
transform -1 0 87806 0 1 24274
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_949
timestamp 1604489732
transform 1 0 87346 0 -1 25362
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_937
timestamp 1604489732
transform 1 0 86242 0 -1 25362
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1556
timestamp 1604489732
transform 1 0 86150 0 -1 25362
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_767
timestamp 1604489732
transform -1 0 87806 0 -1 25362
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1604489732
transform 1 0 1418 0 -1 26450
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1604489732
transform 1 0 314 0 -1 26450
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1604489732
transform 1 0 1418 0 1 25362
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1604489732
transform 1 0 314 0 1 25362
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1604489732
transform 1 0 38 0 -1 26450
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604489732
transform 1 0 38 0 1 25362
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1604489732
transform 1 0 1418 0 1 26450
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1604489732
transform 1 0 314 0 1 26450
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1604489732
transform 1 0 38 0 1 26450
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1604489732
transform 1 0 1418 0 -1 27538
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1604489732
transform 1 0 314 0 -1 27538
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1604489732
transform 1 0 38 0 -1 27538
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_38
timestamp 1604489732
transform 1 0 3534 0 -1 26450
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_32
timestamp 1604489732
transform 1 0 2982 0 -1 26450
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_27
timestamp 1604489732
transform 1 0 2522 0 -1 26450
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1604489732
transform 1 0 2522 0 1 25362
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1385
timestamp 1604489732
transform 1 0 2890 0 -1 26450
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1604489732
transform 1 0 2522 0 1 26450
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_38
timestamp 1604489732
transform 1 0 3534 0 -1 27538
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_32
timestamp 1604489732
transform 1 0 2982 0 -1 27538
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_27
timestamp 1604489732
transform 1 0 2522 0 -1 27538
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1386
timestamp 1604489732
transform 1 0 2890 0 -1 27538
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604489732
transform -1 0 3902 0 1 25362
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1604489732
transform -1 0 3902 0 -1 26450
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1604489732
transform -1 0 3902 0 1 26450
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1604489732
transform -1 0 3902 0 -1 27538
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_912
timestamp 1604489732
transform 1 0 83942 0 -1 26450
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_908
timestamp 1604489732
transform 1 0 83574 0 -1 26450
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_908
timestamp 1604489732
transform 1 0 83574 0 1 25362
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr1[5]
timestamp 1604489732
transform 1 0 83758 0 -1 26450
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_770
timestamp 1604489732
transform 1 0 83298 0 -1 26450
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_768
timestamp 1604489732
transform 1 0 83298 0 1 25362
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_908
timestamp 1604489732
transform 1 0 83574 0 1 26450
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_772
timestamp 1604489732
transform 1 0 83298 0 1 26450
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_912
timestamp 1604489732
transform 1 0 83942 0 -1 27538
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_908
timestamp 1604489732
transform 1 0 83574 0 -1 27538
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr1[4]
timestamp 1604489732
transform 1 0 83758 0 -1 27538
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_774
timestamp 1604489732
transform 1 0 83298 0 -1 27538
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_920
timestamp 1604489732
transform 1 0 84678 0 1 25362
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_932
timestamp 1604489732
transform 1 0 85782 0 1 25362
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_924
timestamp 1604489732
transform 1 0 85046 0 -1 26450
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_920
timestamp 1604489732
transform 1 0 84678 0 1 26450
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_932
timestamp 1604489732
transform 1 0 85782 0 1 26450
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_924
timestamp 1604489732
transform 1 0 85046 0 -1 27538
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_949
timestamp 1604489732
transform 1 0 87346 0 -1 26450
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_937
timestamp 1604489732
transform 1 0 86242 0 -1 26450
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_950
timestamp 1604489732
transform 1 0 87438 0 1 25362
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_944
timestamp 1604489732
transform 1 0 86886 0 1 25362
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1557
timestamp 1604489732
transform 1 0 86150 0 -1 26450
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_771
timestamp 1604489732
transform -1 0 87806 0 -1 26450
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_769
timestamp 1604489732
transform -1 0 87806 0 1 25362
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_950
timestamp 1604489732
transform 1 0 87438 0 1 26450
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_944
timestamp 1604489732
transform 1 0 86886 0 1 26450
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_773
timestamp 1604489732
transform -1 0 87806 0 1 26450
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_949
timestamp 1604489732
transform 1 0 87346 0 -1 27538
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_937
timestamp 1604489732
transform 1 0 86242 0 -1 27538
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1558
timestamp 1604489732
transform 1 0 86150 0 -1 27538
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_775
timestamp 1604489732
transform -1 0 87806 0 -1 27538
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1604489732
transform 1 0 38 0 1 27538
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1604489732
transform 1 0 38 0 -1 28626
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1604489732
transform 1 0 38 0 1 28626
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1604489732
transform 1 0 314 0 1 27538
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1604489732
transform 1 0 1418 0 1 27538
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1604489732
transform 1 0 314 0 -1 28626
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1604489732
transform 1 0 1418 0 -1 28626
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1604489732
transform 1 0 314 0 1 28626
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1604489732
transform 1 0 1418 0 1 28626
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1387
timestamp 1604489732
transform 1 0 2890 0 -1 28626
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1604489732
transform 1 0 2522 0 1 27538
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_27
timestamp 1604489732
transform 1 0 2522 0 -1 28626
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_32
timestamp 1604489732
transform 1 0 2982 0 -1 28626
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_38
timestamp 1604489732
transform 1 0 3534 0 -1 28626
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1604489732
transform 1 0 2522 0 1 28626
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1604489732
transform -1 0 3902 0 1 27538
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1604489732
transform -1 0 3902 0 -1 28626
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1604489732
transform -1 0 3902 0 1 28626
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_776
timestamp 1604489732
transform 1 0 83298 0 1 27538
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_778
timestamp 1604489732
transform 1 0 83298 0 -1 28626
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_780
timestamp 1604489732
transform 1 0 83298 0 1 28626
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr1[3]
timestamp 1604489732
transform 1 0 83758 0 1 28626
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_908
timestamp 1604489732
transform 1 0 83574 0 1 27538
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_908
timestamp 1604489732
transform 1 0 83574 0 -1 28626
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_908
timestamp 1604489732
transform 1 0 83574 0 1 28626
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_912
timestamp 1604489732
transform 1 0 83942 0 1 28626
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_920
timestamp 1604489732
transform 1 0 84678 0 1 27538
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_932
timestamp 1604489732
transform 1 0 85782 0 1 27538
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_920
timestamp 1604489732
transform 1 0 84678 0 -1 28626
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_932
timestamp 1604489732
transform 1 0 85782 0 -1 28626
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_924
timestamp 1604489732
transform 1 0 85046 0 1 28626
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_950
timestamp 1604489732
transform 1 0 87438 0 1 27538
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_944
timestamp 1604489732
transform 1 0 86886 0 1 27538
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_777
timestamp 1604489732
transform -1 0 87806 0 1 27538
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_949
timestamp 1604489732
transform 1 0 87346 0 -1 28626
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_937
timestamp 1604489732
transform 1 0 86242 0 -1 28626
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1559
timestamp 1604489732
transform 1 0 86150 0 -1 28626
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_779
timestamp 1604489732
transform -1 0 87806 0 -1 28626
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_948
timestamp 1604489732
transform 1 0 87254 0 1 28626
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_936
timestamp 1604489732
transform 1 0 86150 0 1 28626
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_781
timestamp 1604489732
transform -1 0 87806 0 1 28626
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1604489732
transform 1 0 38 0 -1 29714
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1604489732
transform 1 0 38 0 1 29714
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1604489732
transform 1 0 38 0 -1 30802
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1604489732
transform 1 0 314 0 -1 29714
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1604489732
transform 1 0 1418 0 -1 29714
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1604489732
transform 1 0 314 0 1 29714
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1604489732
transform 1 0 1418 0 1 29714
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1604489732
transform 1 0 314 0 -1 30802
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1604489732
transform 1 0 1418 0 -1 30802
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1388
timestamp 1604489732
transform 1 0 2890 0 -1 29714
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1389
timestamp 1604489732
transform 1 0 2890 0 -1 30802
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_27
timestamp 1604489732
transform 1 0 2522 0 -1 29714
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_32
timestamp 1604489732
transform 1 0 2982 0 -1 29714
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_38
timestamp 1604489732
transform 1 0 3534 0 -1 29714
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1604489732
transform 1 0 2522 0 1 29714
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_27
timestamp 1604489732
transform 1 0 2522 0 -1 30802
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_32
timestamp 1604489732
transform 1 0 2982 0 -1 30802
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_38
timestamp 1604489732
transform 1 0 3534 0 -1 30802
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1604489732
transform -1 0 3902 0 -1 29714
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1604489732
transform -1 0 3902 0 1 29714
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1604489732
transform -1 0 3902 0 -1 30802
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_782
timestamp 1604489732
transform 1 0 83298 0 -1 29714
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_784
timestamp 1604489732
transform 1 0 83298 0 1 29714
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_786
timestamp 1604489732
transform 1 0 83298 0 -1 30802
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr1[2]
timestamp 1604489732
transform 1 0 83758 0 1 29714
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_908
timestamp 1604489732
transform 1 0 83574 0 -1 29714
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_908
timestamp 1604489732
transform 1 0 83574 0 1 29714
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_912
timestamp 1604489732
transform 1 0 83942 0 1 29714
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_908
timestamp 1604489732
transform 1 0 83574 0 -1 30802
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_920
timestamp 1604489732
transform 1 0 84678 0 -1 29714
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_932
timestamp 1604489732
transform 1 0 85782 0 -1 29714
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_924
timestamp 1604489732
transform 1 0 85046 0 1 29714
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_920
timestamp 1604489732
transform 1 0 84678 0 -1 30802
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_932
timestamp 1604489732
transform 1 0 85782 0 -1 30802
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_949
timestamp 1604489732
transform 1 0 87346 0 -1 29714
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_937
timestamp 1604489732
transform 1 0 86242 0 -1 29714
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1560
timestamp 1604489732
transform 1 0 86150 0 -1 29714
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_783
timestamp 1604489732
transform -1 0 87806 0 -1 29714
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_948
timestamp 1604489732
transform 1 0 87254 0 1 29714
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_936
timestamp 1604489732
transform 1 0 86150 0 1 29714
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_785
timestamp 1604489732
transform -1 0 87806 0 1 29714
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_949
timestamp 1604489732
transform 1 0 87346 0 -1 30802
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_937
timestamp 1604489732
transform 1 0 86242 0 -1 30802
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1561
timestamp 1604489732
transform 1 0 86150 0 -1 30802
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_787
timestamp 1604489732
transform -1 0 87806 0 -1 30802
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1604489732
transform 1 0 1418 0 1 30802
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1604489732
transform 1 0 314 0 1 30802
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1604489732
transform 1 0 38 0 1 30802
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1604489732
transform 1 0 1418 0 1 31890
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1604489732
transform 1 0 314 0 1 31890
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1604489732
transform 1 0 1418 0 -1 31890
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1604489732
transform 1 0 314 0 -1 31890
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1604489732
transform 1 0 38 0 1 31890
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1604489732
transform 1 0 38 0 -1 31890
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1604489732
transform 1 0 1418 0 -1 32978
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1604489732
transform 1 0 314 0 -1 32978
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1604489732
transform 1 0 38 0 -1 32978
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1604489732
transform 1 0 2522 0 1 30802
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1604489732
transform 1 0 2522 0 1 31890
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_38
timestamp 1604489732
transform 1 0 3534 0 -1 31890
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_32
timestamp 1604489732
transform 1 0 2982 0 -1 31890
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_27
timestamp 1604489732
transform 1 0 2522 0 -1 31890
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1390
timestamp 1604489732
transform 1 0 2890 0 -1 31890
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_38
timestamp 1604489732
transform 1 0 3534 0 -1 32978
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_32
timestamp 1604489732
transform 1 0 2982 0 -1 32978
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_27
timestamp 1604489732
transform 1 0 2522 0 -1 32978
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1391
timestamp 1604489732
transform 1 0 2890 0 -1 32978
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1604489732
transform -1 0 3902 0 1 30802
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1604489732
transform -1 0 3902 0 -1 31890
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1604489732
transform -1 0 3902 0 1 31890
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1604489732
transform -1 0 3902 0 -1 32978
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_908
timestamp 1604489732
transform 1 0 83574 0 1 30802
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_788
timestamp 1604489732
transform 1 0 83298 0 1 30802
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_908
timestamp 1604489732
transform 1 0 83574 0 1 31890
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_912
timestamp 1604489732
transform 1 0 83942 0 -1 31890
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_908
timestamp 1604489732
transform 1 0 83574 0 -1 31890
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr1[1]
timestamp 1604489732
transform 1 0 83758 0 -1 31890
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_792
timestamp 1604489732
transform 1 0 83298 0 1 31890
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_790
timestamp 1604489732
transform 1 0 83298 0 -1 31890
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_908
timestamp 1604489732
transform 1 0 83574 0 -1 32978
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_794
timestamp 1604489732
transform 1 0 83298 0 -1 32978
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_920
timestamp 1604489732
transform 1 0 84678 0 1 30802
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_932
timestamp 1604489732
transform 1 0 85782 0 1 30802
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_924
timestamp 1604489732
transform 1 0 85046 0 -1 31890
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_920
timestamp 1604489732
transform 1 0 84678 0 1 31890
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_932
timestamp 1604489732
transform 1 0 85782 0 1 31890
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_920
timestamp 1604489732
transform 1 0 84678 0 -1 32978
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_932
timestamp 1604489732
transform 1 0 85782 0 -1 32978
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_950
timestamp 1604489732
transform 1 0 87438 0 1 30802
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_944
timestamp 1604489732
transform 1 0 86886 0 1 30802
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_789
timestamp 1604489732
transform -1 0 87806 0 1 30802
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_55_950
timestamp 1604489732
transform 1 0 87438 0 1 31890
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_944
timestamp 1604489732
transform 1 0 86886 0 1 31890
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_949
timestamp 1604489732
transform 1 0 87346 0 -1 31890
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_937
timestamp 1604489732
transform 1 0 86242 0 -1 31890
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1562
timestamp 1604489732
transform 1 0 86150 0 -1 31890
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_793
timestamp 1604489732
transform -1 0 87806 0 1 31890
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_791
timestamp 1604489732
transform -1 0 87806 0 -1 31890
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_949
timestamp 1604489732
transform 1 0 87346 0 -1 32978
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_937
timestamp 1604489732
transform 1 0 86242 0 -1 32978
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1563
timestamp 1604489732
transform 1 0 86150 0 -1 32978
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_795
timestamp 1604489732
transform -1 0 87806 0 -1 32978
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1604489732
transform 1 0 38 0 1 32978
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1604489732
transform 1 0 38 0 -1 34066
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1604489732
transform 1 0 38 0 1 34066
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1604489732
transform 1 0 314 0 1 32978
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1604489732
transform 1 0 1418 0 1 32978
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1604489732
transform 1 0 314 0 -1 34066
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1604489732
transform 1 0 1418 0 -1 34066
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1604489732
transform 1 0 314 0 1 34066
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1604489732
transform 1 0 1418 0 1 34066
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1392
timestamp 1604489732
transform 1 0 2890 0 -1 34066
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1604489732
transform 1 0 2522 0 1 32978
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_27
timestamp 1604489732
transform 1 0 2522 0 -1 34066
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_32
timestamp 1604489732
transform 1 0 2982 0 -1 34066
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_38
timestamp 1604489732
transform 1 0 3534 0 -1 34066
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1604489732
transform 1 0 2522 0 1 34066
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1604489732
transform -1 0 3902 0 1 32978
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1604489732
transform -1 0 3902 0 -1 34066
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1604489732
transform -1 0 3902 0 1 34066
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_796
timestamp 1604489732
transform 1 0 83298 0 1 32978
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_798
timestamp 1604489732
transform 1 0 83298 0 -1 34066
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_800
timestamp 1604489732
transform 1 0 83298 0 1 34066
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_908
timestamp 1604489732
transform 1 0 83574 0 1 32978
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_908
timestamp 1604489732
transform 1 0 83574 0 -1 34066
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_908
timestamp 1604489732
transform 1 0 83574 0 1 34066
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_920
timestamp 1604489732
transform 1 0 84678 0 1 32978
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_932
timestamp 1604489732
transform 1 0 85782 0 1 32978
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_920
timestamp 1604489732
transform 1 0 84678 0 -1 34066
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_932
timestamp 1604489732
transform 1 0 85782 0 -1 34066
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_920
timestamp 1604489732
transform 1 0 84678 0 1 34066
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_932
timestamp 1604489732
transform 1 0 85782 0 1 34066
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_950
timestamp 1604489732
transform 1 0 87438 0 1 32978
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_944
timestamp 1604489732
transform 1 0 86886 0 1 32978
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_797
timestamp 1604489732
transform -1 0 87806 0 1 32978
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_949
timestamp 1604489732
transform 1 0 87346 0 -1 34066
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_937
timestamp 1604489732
transform 1 0 86242 0 -1 34066
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1564
timestamp 1604489732
transform 1 0 86150 0 -1 34066
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_799
timestamp 1604489732
transform -1 0 87806 0 -1 34066
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_59_950
timestamp 1604489732
transform 1 0 87438 0 1 34066
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_944
timestamp 1604489732
transform 1 0 86886 0 1 34066
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_801
timestamp 1604489732
transform -1 0 87806 0 1 34066
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1604489732
transform 1 0 38 0 -1 35154
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1604489732
transform 1 0 38 0 1 35154
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1604489732
transform 1 0 38 0 -1 36242
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1604489732
transform 1 0 314 0 -1 35154
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1604489732
transform 1 0 1418 0 -1 35154
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1604489732
transform 1 0 314 0 1 35154
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1604489732
transform 1 0 1418 0 1 35154
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1604489732
transform 1 0 314 0 -1 36242
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1604489732
transform 1 0 1418 0 -1 36242
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1393
timestamp 1604489732
transform 1 0 2890 0 -1 35154
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1394
timestamp 1604489732
transform 1 0 2890 0 -1 36242
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_27
timestamp 1604489732
transform 1 0 2522 0 -1 35154
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_32
timestamp 1604489732
transform 1 0 2982 0 -1 35154
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_38
timestamp 1604489732
transform 1 0 3534 0 -1 35154
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1604489732
transform 1 0 2522 0 1 35154
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_27
timestamp 1604489732
transform 1 0 2522 0 -1 36242
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_32
timestamp 1604489732
transform 1 0 2982 0 -1 36242
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_38
timestamp 1604489732
transform 1 0 3534 0 -1 36242
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1604489732
transform -1 0 3902 0 -1 35154
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1604489732
transform -1 0 3902 0 1 35154
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1604489732
transform -1 0 3902 0 -1 36242
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_802
timestamp 1604489732
transform 1 0 83298 0 -1 35154
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_804
timestamp 1604489732
transform 1 0 83298 0 1 35154
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_806
timestamp 1604489732
transform 1 0 83298 0 -1 36242
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_908
timestamp 1604489732
transform 1 0 83574 0 -1 35154
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_908
timestamp 1604489732
transform 1 0 83574 0 1 35154
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_908
timestamp 1604489732
transform 1 0 83574 0 -1 36242
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_920
timestamp 1604489732
transform 1 0 84678 0 -1 35154
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_932
timestamp 1604489732
transform 1 0 85782 0 -1 35154
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_920
timestamp 1604489732
transform 1 0 84678 0 1 35154
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_932
timestamp 1604489732
transform 1 0 85782 0 1 35154
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_920
timestamp 1604489732
transform 1 0 84678 0 -1 36242
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_932
timestamp 1604489732
transform 1 0 85782 0 -1 36242
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_949
timestamp 1604489732
transform 1 0 87346 0 -1 35154
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_937
timestamp 1604489732
transform 1 0 86242 0 -1 35154
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1565
timestamp 1604489732
transform 1 0 86150 0 -1 35154
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_803
timestamp 1604489732
transform -1 0 87806 0 -1 35154
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_61_950
timestamp 1604489732
transform 1 0 87438 0 1 35154
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_944
timestamp 1604489732
transform 1 0 86886 0 1 35154
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_805
timestamp 1604489732
transform -1 0 87806 0 1 35154
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_949
timestamp 1604489732
transform 1 0 87346 0 -1 36242
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_937
timestamp 1604489732
transform 1 0 86242 0 -1 36242
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1566
timestamp 1604489732
transform 1 0 86150 0 -1 36242
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_807
timestamp 1604489732
transform -1 0 87806 0 -1 36242
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1604489732
transform 1 0 38 0 1 36242
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1604489732
transform 1 0 38 0 -1 37330
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1604489732
transform 1 0 38 0 1 37330
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1604489732
transform 1 0 314 0 1 36242
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1604489732
transform 1 0 1418 0 1 36242
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1604489732
transform 1 0 314 0 -1 37330
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1604489732
transform 1 0 1418 0 -1 37330
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1604489732
transform 1 0 314 0 1 37330
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1604489732
transform 1 0 1418 0 1 37330
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1395
timestamp 1604489732
transform 1 0 2890 0 -1 37330
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1604489732
transform 1 0 2522 0 1 36242
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_27
timestamp 1604489732
transform 1 0 2522 0 -1 37330
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_32
timestamp 1604489732
transform 1 0 2982 0 -1 37330
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_38
timestamp 1604489732
transform 1 0 3534 0 -1 37330
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1604489732
transform 1 0 2522 0 1 37330
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1604489732
transform -1 0 3902 0 1 36242
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1604489732
transform -1 0 3902 0 -1 37330
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1604489732
transform -1 0 3902 0 1 37330
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_808
timestamp 1604489732
transform 1 0 83298 0 1 36242
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_810
timestamp 1604489732
transform 1 0 83298 0 -1 37330
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_812
timestamp 1604489732
transform 1 0 83298 0 1 37330
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_908
timestamp 1604489732
transform 1 0 83574 0 1 36242
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_908
timestamp 1604489732
transform 1 0 83574 0 -1 37330
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_908
timestamp 1604489732
transform 1 0 83574 0 1 37330
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_920
timestamp 1604489732
transform 1 0 84678 0 1 36242
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_932
timestamp 1604489732
transform 1 0 85782 0 1 36242
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_920
timestamp 1604489732
transform 1 0 84678 0 -1 37330
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_932
timestamp 1604489732
transform 1 0 85782 0 -1 37330
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_920
timestamp 1604489732
transform 1 0 84678 0 1 37330
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_932
timestamp 1604489732
transform 1 0 85782 0 1 37330
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_950
timestamp 1604489732
transform 1 0 87438 0 1 36242
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_944
timestamp 1604489732
transform 1 0 86886 0 1 36242
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_809
timestamp 1604489732
transform -1 0 87806 0 1 36242
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_65_950
timestamp 1604489732
transform 1 0 87438 0 1 37330
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_944
timestamp 1604489732
transform 1 0 86886 0 1 37330
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_949
timestamp 1604489732
transform 1 0 87346 0 -1 37330
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_937
timestamp 1604489732
transform 1 0 86242 0 -1 37330
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1567
timestamp 1604489732
transform 1 0 86150 0 -1 37330
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_813
timestamp 1604489732
transform -1 0 87806 0 1 37330
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_811
timestamp 1604489732
transform -1 0 87806 0 -1 37330
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1604489732
transform 1 0 1418 0 1 38418
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1604489732
transform 1 0 314 0 1 38418
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1604489732
transform 1 0 1418 0 -1 38418
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1604489732
transform 1 0 314 0 -1 38418
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1604489732
transform 1 0 38 0 1 38418
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1604489732
transform 1 0 38 0 -1 38418
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1604489732
transform 1 0 1418 0 -1 39506
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1604489732
transform 1 0 314 0 -1 39506
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1604489732
transform 1 0 38 0 -1 39506
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1604489732
transform 1 0 1418 0 1 39506
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1604489732
transform 1 0 314 0 1 39506
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1604489732
transform 1 0 38 0 1 39506
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1604489732
transform 1 0 2522 0 1 38418
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_38
timestamp 1604489732
transform 1 0 3534 0 -1 38418
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_32
timestamp 1604489732
transform 1 0 2982 0 -1 38418
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_27
timestamp 1604489732
transform 1 0 2522 0 -1 38418
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1396
timestamp 1604489732
transform 1 0 2890 0 -1 38418
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_38
timestamp 1604489732
transform 1 0 3534 0 -1 39506
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_32
timestamp 1604489732
transform 1 0 2982 0 -1 39506
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_27
timestamp 1604489732
transform 1 0 2522 0 -1 39506
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1397
timestamp 1604489732
transform 1 0 2890 0 -1 39506
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1604489732
transform 1 0 2522 0 1 39506
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1604489732
transform -1 0 3902 0 -1 38418
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1604489732
transform -1 0 3902 0 1 38418
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1604489732
transform -1 0 3902 0 -1 39506
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1604489732
transform -1 0 3902 0 1 39506
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_814
timestamp 1604489732
transform 1 0 83298 0 -1 38418
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_816
timestamp 1604489732
transform 1 0 83298 0 1 38418
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_818
timestamp 1604489732
transform 1 0 83298 0 -1 39506
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_820
timestamp 1604489732
transform 1 0 83298 0 1 39506
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_908
timestamp 1604489732
transform 1 0 83574 0 -1 38418
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_908
timestamp 1604489732
transform 1 0 83574 0 1 38418
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_908
timestamp 1604489732
transform 1 0 83574 0 -1 39506
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_908
timestamp 1604489732
transform 1 0 83574 0 1 39506
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_920
timestamp 1604489732
transform 1 0 84678 0 -1 38418
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_932
timestamp 1604489732
transform 1 0 85782 0 -1 38418
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_920
timestamp 1604489732
transform 1 0 84678 0 1 38418
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_932
timestamp 1604489732
transform 1 0 85782 0 1 38418
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_920
timestamp 1604489732
transform 1 0 84678 0 -1 39506
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_932
timestamp 1604489732
transform 1 0 85782 0 -1 39506
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_920
timestamp 1604489732
transform 1 0 84678 0 1 39506
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_932
timestamp 1604489732
transform 1 0 85782 0 1 39506
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_950
timestamp 1604489732
transform 1 0 87438 0 1 38418
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_944
timestamp 1604489732
transform 1 0 86886 0 1 38418
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_949
timestamp 1604489732
transform 1 0 87346 0 -1 38418
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_937
timestamp 1604489732
transform 1 0 86242 0 -1 38418
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1568
timestamp 1604489732
transform 1 0 86150 0 -1 38418
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_817
timestamp 1604489732
transform -1 0 87806 0 1 38418
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_815
timestamp 1604489732
transform -1 0 87806 0 -1 38418
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_68_949
timestamp 1604489732
transform 1 0 87346 0 -1 39506
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_937
timestamp 1604489732
transform 1 0 86242 0 -1 39506
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1569
timestamp 1604489732
transform 1 0 86150 0 -1 39506
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_819
timestamp 1604489732
transform -1 0 87806 0 -1 39506
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_69_950
timestamp 1604489732
transform 1 0 87438 0 1 39506
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_944
timestamp 1604489732
transform 1 0 86886 0 1 39506
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_821
timestamp 1604489732
transform -1 0 87806 0 1 39506
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1604489732
transform 1 0 38 0 -1 40594
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1604489732
transform 1 0 38 0 1 40594
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1604489732
transform 1 0 38 0 -1 41682
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_3
timestamp 1604489732
transform 1 0 314 0 -1 40594
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_15
timestamp 1604489732
transform 1 0 1418 0 -1 40594
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1604489732
transform 1 0 314 0 1 40594
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_15
timestamp 1604489732
transform 1 0 1418 0 1 40594
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1604489732
transform 1 0 314 0 -1 41682
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_15
timestamp 1604489732
transform 1 0 1418 0 -1 41682
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1398
timestamp 1604489732
transform 1 0 2890 0 -1 40594
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1399
timestamp 1604489732
transform 1 0 2890 0 -1 41682
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_27
timestamp 1604489732
transform 1 0 2522 0 -1 40594
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_32
timestamp 1604489732
transform 1 0 2982 0 -1 40594
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_38
timestamp 1604489732
transform 1 0 3534 0 -1 40594
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_27
timestamp 1604489732
transform 1 0 2522 0 1 40594
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_27
timestamp 1604489732
transform 1 0 2522 0 -1 41682
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_32
timestamp 1604489732
transform 1 0 2982 0 -1 41682
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_38
timestamp 1604489732
transform 1 0 3534 0 -1 41682
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1604489732
transform -1 0 3902 0 -1 40594
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1604489732
transform -1 0 3902 0 1 40594
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1604489732
transform -1 0 3902 0 -1 41682
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_822
timestamp 1604489732
transform 1 0 83298 0 -1 40594
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_824
timestamp 1604489732
transform 1 0 83298 0 1 40594
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_826
timestamp 1604489732
transform 1 0 83298 0 -1 41682
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_908
timestamp 1604489732
transform 1 0 83574 0 -1 40594
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_908
timestamp 1604489732
transform 1 0 83574 0 1 40594
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_908
timestamp 1604489732
transform 1 0 83574 0 -1 41682
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_920
timestamp 1604489732
transform 1 0 84678 0 -1 40594
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_932
timestamp 1604489732
transform 1 0 85782 0 -1 40594
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_920
timestamp 1604489732
transform 1 0 84678 0 1 40594
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_932
timestamp 1604489732
transform 1 0 85782 0 1 40594
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_920
timestamp 1604489732
transform 1 0 84678 0 -1 41682
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_932
timestamp 1604489732
transform 1 0 85782 0 -1 41682
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_949
timestamp 1604489732
transform 1 0 87346 0 -1 40594
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_937
timestamp 1604489732
transform 1 0 86242 0 -1 40594
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1570
timestamp 1604489732
transform 1 0 86150 0 -1 40594
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_823
timestamp 1604489732
transform -1 0 87806 0 -1 40594
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_71_950
timestamp 1604489732
transform 1 0 87438 0 1 40594
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_944
timestamp 1604489732
transform 1 0 86886 0 1 40594
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_825
timestamp 1604489732
transform -1 0 87806 0 1 40594
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_72_949
timestamp 1604489732
transform 1 0 87346 0 -1 41682
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_937
timestamp 1604489732
transform 1 0 86242 0 -1 41682
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1571
timestamp 1604489732
transform 1 0 86150 0 -1 41682
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_827
timestamp 1604489732
transform -1 0 87806 0 -1 41682
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1604489732
transform 1 0 38 0 1 41682
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1604489732
transform 1 0 38 0 -1 42770
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1604489732
transform 1 0 38 0 1 42770
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_3
timestamp 1604489732
transform 1 0 314 0 1 41682
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_15
timestamp 1604489732
transform 1 0 1418 0 1 41682
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1604489732
transform 1 0 314 0 -1 42770
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1604489732
transform 1 0 1418 0 -1 42770
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_3
timestamp 1604489732
transform 1 0 314 0 1 42770
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_15
timestamp 1604489732
transform 1 0 1418 0 1 42770
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1400
timestamp 1604489732
transform 1 0 2890 0 -1 42770
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_27
timestamp 1604489732
transform 1 0 2522 0 1 41682
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_27
timestamp 1604489732
transform 1 0 2522 0 -1 42770
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_32
timestamp 1604489732
transform 1 0 2982 0 -1 42770
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_38
timestamp 1604489732
transform 1 0 3534 0 -1 42770
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_27
timestamp 1604489732
transform 1 0 2522 0 1 42770
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1604489732
transform -1 0 3902 0 1 41682
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1604489732
transform -1 0 3902 0 -1 42770
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1604489732
transform -1 0 3902 0 1 42770
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_828
timestamp 1604489732
transform 1 0 83298 0 1 41682
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_830
timestamp 1604489732
transform 1 0 83298 0 -1 42770
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_832
timestamp 1604489732
transform 1 0 83298 0 1 42770
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_908
timestamp 1604489732
transform 1 0 83574 0 1 41682
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_908
timestamp 1604489732
transform 1 0 83574 0 -1 42770
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_908
timestamp 1604489732
transform 1 0 83574 0 1 42770
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_920
timestamp 1604489732
transform 1 0 84678 0 1 41682
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_932
timestamp 1604489732
transform 1 0 85782 0 1 41682
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_920
timestamp 1604489732
transform 1 0 84678 0 -1 42770
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_932
timestamp 1604489732
transform 1 0 85782 0 -1 42770
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_920
timestamp 1604489732
transform 1 0 84678 0 1 42770
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_932
timestamp 1604489732
transform 1 0 85782 0 1 42770
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_950
timestamp 1604489732
transform 1 0 87438 0 1 41682
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_944
timestamp 1604489732
transform 1 0 86886 0 1 41682
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_829
timestamp 1604489732
transform -1 0 87806 0 1 41682
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_74_949
timestamp 1604489732
transform 1 0 87346 0 -1 42770
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_937
timestamp 1604489732
transform 1 0 86242 0 -1 42770
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1572
timestamp 1604489732
transform 1 0 86150 0 -1 42770
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_831
timestamp 1604489732
transform -1 0 87806 0 -1 42770
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_75_950
timestamp 1604489732
transform 1 0 87438 0 1 42770
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_944
timestamp 1604489732
transform 1 0 86886 0 1 42770
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_833
timestamp 1604489732
transform -1 0 87806 0 1 42770
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1604489732
transform 1 0 1418 0 1 43858
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1604489732
transform 1 0 314 0 1 43858
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1604489732
transform 1 0 1418 0 -1 43858
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1604489732
transform 1 0 314 0 -1 43858
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1604489732
transform 1 0 38 0 1 43858
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1604489732
transform 1 0 38 0 -1 43858
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1604489732
transform 1 0 1418 0 -1 44946
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_3
timestamp 1604489732
transform 1 0 314 0 -1 44946
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1604489732
transform 1 0 38 0 -1 44946
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_15
timestamp 1604489732
transform 1 0 1418 0 1 44946
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_3
timestamp 1604489732
transform 1 0 314 0 1 44946
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1604489732
transform 1 0 38 0 1 44946
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1604489732
transform 1 0 2522 0 1 43858
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_38
timestamp 1604489732
transform 1 0 3534 0 -1 43858
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_32
timestamp 1604489732
transform 1 0 2982 0 -1 43858
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_76_27
timestamp 1604489732
transform 1 0 2522 0 -1 43858
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1401
timestamp 1604489732
transform 1 0 2890 0 -1 43858
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_78_38
timestamp 1604489732
transform 1 0 3534 0 -1 44946
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_32
timestamp 1604489732
transform 1 0 2982 0 -1 44946
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_27
timestamp 1604489732
transform 1 0 2522 0 -1 44946
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1402
timestamp 1604489732
transform 1 0 2890 0 -1 44946
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_27
timestamp 1604489732
transform 1 0 2522 0 1 44946
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1604489732
transform -1 0 3902 0 -1 43858
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1604489732
transform -1 0 3902 0 1 43858
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1604489732
transform -1 0 3902 0 -1 44946
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1604489732
transform -1 0 3902 0 1 44946
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_834
timestamp 1604489732
transform 1 0 83298 0 -1 43858
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_836
timestamp 1604489732
transform 1 0 83298 0 1 43858
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_838
timestamp 1604489732
transform 1 0 83298 0 -1 44946
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_840
timestamp 1604489732
transform 1 0 83298 0 1 44946
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_908
timestamp 1604489732
transform 1 0 83574 0 -1 43858
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_908
timestamp 1604489732
transform 1 0 83574 0 1 43858
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_908
timestamp 1604489732
transform 1 0 83574 0 -1 44946
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_908
timestamp 1604489732
transform 1 0 83574 0 1 44946
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_920
timestamp 1604489732
transform 1 0 84678 0 -1 43858
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_932
timestamp 1604489732
transform 1 0 85782 0 -1 43858
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_920
timestamp 1604489732
transform 1 0 84678 0 1 43858
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_932
timestamp 1604489732
transform 1 0 85782 0 1 43858
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_920
timestamp 1604489732
transform 1 0 84678 0 -1 44946
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_932
timestamp 1604489732
transform 1 0 85782 0 -1 44946
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_920
timestamp 1604489732
transform 1 0 84678 0 1 44946
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_932
timestamp 1604489732
transform 1 0 85782 0 1 44946
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_950
timestamp 1604489732
transform 1 0 87438 0 1 43858
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_944
timestamp 1604489732
transform 1 0 86886 0 1 43858
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_76_949
timestamp 1604489732
transform 1 0 87346 0 -1 43858
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_76_937
timestamp 1604489732
transform 1 0 86242 0 -1 43858
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1573
timestamp 1604489732
transform 1 0 86150 0 -1 43858
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_837
timestamp 1604489732
transform -1 0 87806 0 1 43858
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_835
timestamp 1604489732
transform -1 0 87806 0 -1 43858
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_78_949
timestamp 1604489732
transform 1 0 87346 0 -1 44946
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_937
timestamp 1604489732
transform 1 0 86242 0 -1 44946
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1574
timestamp 1604489732
transform 1 0 86150 0 -1 44946
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_839
timestamp 1604489732
transform -1 0 87806 0 -1 44946
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_79_950
timestamp 1604489732
transform 1 0 87438 0 1 44946
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_944
timestamp 1604489732
transform 1 0 86886 0 1 44946
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_841
timestamp 1604489732
transform -1 0 87806 0 1 44946
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1604489732
transform 1 0 38 0 -1 46034
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1604489732
transform 1 0 38 0 1 46034
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1604489732
transform 1 0 38 0 -1 47122
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_3
timestamp 1604489732
transform 1 0 314 0 -1 46034
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_15
timestamp 1604489732
transform 1 0 1418 0 -1 46034
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_3
timestamp 1604489732
transform 1 0 314 0 1 46034
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_15
timestamp 1604489732
transform 1 0 1418 0 1 46034
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_3
timestamp 1604489732
transform 1 0 314 0 -1 47122
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_15
timestamp 1604489732
transform 1 0 1418 0 -1 47122
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1403
timestamp 1604489732
transform 1 0 2890 0 -1 46034
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1404
timestamp 1604489732
transform 1 0 2890 0 -1 47122
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_27
timestamp 1604489732
transform 1 0 2522 0 -1 46034
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_32
timestamp 1604489732
transform 1 0 2982 0 -1 46034
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_38
timestamp 1604489732
transform 1 0 3534 0 -1 46034
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_27
timestamp 1604489732
transform 1 0 2522 0 1 46034
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_27
timestamp 1604489732
transform 1 0 2522 0 -1 47122
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_32
timestamp 1604489732
transform 1 0 2982 0 -1 47122
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_38
timestamp 1604489732
transform 1 0 3534 0 -1 47122
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1604489732
transform -1 0 3902 0 -1 46034
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1604489732
transform -1 0 3902 0 1 46034
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1604489732
transform -1 0 3902 0 -1 47122
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_842
timestamp 1604489732
transform 1 0 83298 0 -1 46034
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_844
timestamp 1604489732
transform 1 0 83298 0 1 46034
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_846
timestamp 1604489732
transform 1 0 83298 0 -1 47122
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_908
timestamp 1604489732
transform 1 0 83574 0 -1 46034
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_908
timestamp 1604489732
transform 1 0 83574 0 1 46034
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_908
timestamp 1604489732
transform 1 0 83574 0 -1 47122
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_920
timestamp 1604489732
transform 1 0 84678 0 -1 46034
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_932
timestamp 1604489732
transform 1 0 85782 0 -1 46034
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_920
timestamp 1604489732
transform 1 0 84678 0 1 46034
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_932
timestamp 1604489732
transform 1 0 85782 0 1 46034
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_920
timestamp 1604489732
transform 1 0 84678 0 -1 47122
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_932
timestamp 1604489732
transform 1 0 85782 0 -1 47122
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_949
timestamp 1604489732
transform 1 0 87346 0 -1 46034
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_937
timestamp 1604489732
transform 1 0 86242 0 -1 46034
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1575
timestamp 1604489732
transform 1 0 86150 0 -1 46034
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_843
timestamp 1604489732
transform -1 0 87806 0 -1 46034
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_81_950
timestamp 1604489732
transform 1 0 87438 0 1 46034
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_944
timestamp 1604489732
transform 1 0 86886 0 1 46034
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_845
timestamp 1604489732
transform -1 0 87806 0 1 46034
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_949
timestamp 1604489732
transform 1 0 87346 0 -1 47122
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_937
timestamp 1604489732
transform 1 0 86242 0 -1 47122
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1576
timestamp 1604489732
transform 1 0 86150 0 -1 47122
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_847
timestamp 1604489732
transform -1 0 87806 0 -1 47122
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1604489732
transform 1 0 38 0 1 47122
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_3
timestamp 1604489732
transform 1 0 314 0 1 47122
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_15
timestamp 1604489732
transform 1 0 1418 0 1 47122
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_27
timestamp 1604489732
transform 1 0 2522 0 1 47122
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1604489732
transform -1 0 3902 0 1 47122
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_848
timestamp 1604489732
transform 1 0 83298 0 1 47122
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_908
timestamp 1604489732
transform 1 0 83574 0 1 47122
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_920
timestamp 1604489732
transform 1 0 84678 0 1 47122
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_932
timestamp 1604489732
transform 1 0 85782 0 1 47122
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_849
timestamp 1604489732
transform -1 0 87806 0 1 47122
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_83_944
timestamp 1604489732
transform 1 0 86886 0 1 47122
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_950
timestamp 1604489732
transform 1 0 87438 0 1 47122
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_15
timestamp 1604489732
transform 1 0 1418 0 1 48210
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_3
timestamp 1604489732
transform 1 0 314 0 1 48210
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_15
timestamp 1604489732
transform 1 0 1418 0 -1 48210
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_3
timestamp 1604489732
transform 1 0 314 0 -1 48210
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1604489732
transform 1 0 38 0 1 48210
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1604489732
transform 1 0 38 0 -1 48210
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_86_15
timestamp 1604489732
transform 1 0 1418 0 -1 49298
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_3
timestamp 1604489732
transform 1 0 314 0 -1 49298
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1604489732
transform 1 0 38 0 -1 49298
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_87_15
timestamp 1604489732
transform 1 0 1418 0 1 49298
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_3
timestamp 1604489732
transform 1 0 314 0 1 49298
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1604489732
transform 1 0 38 0 1 49298
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_85_27
timestamp 1604489732
transform 1 0 2522 0 1 48210
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_38
timestamp 1604489732
transform 1 0 3534 0 -1 48210
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_84_32
timestamp 1604489732
transform 1 0 2982 0 -1 48210
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_84_27
timestamp 1604489732
transform 1 0 2522 0 -1 48210
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1405
timestamp 1604489732
transform 1 0 2890 0 -1 48210
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1604489732
transform -1 0 3902 0 1 48210
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1604489732
transform -1 0 3902 0 -1 48210
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_86_38
timestamp 1604489732
transform 1 0 3534 0 -1 49298
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_86_32
timestamp 1604489732
transform 1 0 2982 0 -1 49298
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_86_27
timestamp 1604489732
transform 1 0 2522 0 -1 49298
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1406
timestamp 1604489732
transform 1 0 2890 0 -1 49298
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1604489732
transform -1 0 3902 0 -1 49298
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_87_27
timestamp 1604489732
transform 1 0 2522 0 1 49298
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1604489732
transform -1 0 3902 0 1 49298
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_850
timestamp 1604489732
transform 1 0 83298 0 -1 48210
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_852
timestamp 1604489732
transform 1 0 83298 0 1 48210
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_854
timestamp 1604489732
transform 1 0 83298 0 -1 49298
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_856
timestamp 1604489732
transform 1 0 83298 0 1 49298
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_908
timestamp 1604489732
transform 1 0 83574 0 -1 48210
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_908
timestamp 1604489732
transform 1 0 83574 0 1 48210
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_908
timestamp 1604489732
transform 1 0 83574 0 -1 49298
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_908
timestamp 1604489732
transform 1 0 83574 0 1 49298
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_932
timestamp 1604489732
transform 1 0 85782 0 1 48210
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_920
timestamp 1604489732
transform 1 0 84678 0 1 48210
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_937
timestamp 1604489732
transform 1 0 86242 0 -1 48210
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_932
timestamp 1604489732
transform 1 0 85782 0 -1 48210
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_920
timestamp 1604489732
transform 1 0 84678 0 -1 48210
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1577
timestamp 1604489732
transform 1 0 86150 0 -1 48210
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_937
timestamp 1604489732
transform 1 0 86242 0 -1 49298
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_932
timestamp 1604489732
transform 1 0 85782 0 -1 49298
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_920
timestamp 1604489732
transform 1 0 84678 0 -1 49298
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1578
timestamp 1604489732
transform 1 0 86150 0 -1 49298
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_932
timestamp 1604489732
transform 1 0 85782 0 1 49298
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_920
timestamp 1604489732
transform 1 0 84678 0 1 49298
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_944
timestamp 1604489732
transform 1 0 86886 0 1 48210
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_950
timestamp 1604489732
transform 1 0 87438 0 1 48210
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_949
timestamp 1604489732
transform 1 0 87346 0 -1 48210
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_853
timestamp 1604489732
transform -1 0 87806 0 1 48210
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_851
timestamp 1604489732
transform -1 0 87806 0 -1 48210
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_86_949
timestamp 1604489732
transform 1 0 87346 0 -1 49298
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_855
timestamp 1604489732
transform -1 0 87806 0 -1 49298
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_87_944
timestamp 1604489732
transform 1 0 86886 0 1 49298
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_950
timestamp 1604489732
transform 1 0 87438 0 1 49298
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_857
timestamp 1604489732
transform -1 0 87806 0 1 49298
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1604489732
transform 1 0 38 0 -1 50386
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1604489732
transform 1 0 38 0 1 50386
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1604489732
transform 1 0 38 0 -1 51474
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_88_3
timestamp 1604489732
transform 1 0 314 0 -1 50386
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_15
timestamp 1604489732
transform 1 0 1418 0 -1 50386
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_3
timestamp 1604489732
transform 1 0 314 0 1 50386
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_15
timestamp 1604489732
transform 1 0 1418 0 1 50386
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_3
timestamp 1604489732
transform 1 0 314 0 -1 51474
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_15
timestamp 1604489732
transform 1 0 1418 0 -1 51474
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_38
timestamp 1604489732
transform 1 0 3534 0 -1 50386
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_88_32
timestamp 1604489732
transform 1 0 2982 0 -1 50386
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_88_27
timestamp 1604489732
transform 1 0 2522 0 -1 50386
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1407
timestamp 1604489732
transform 1 0 2890 0 -1 50386
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1604489732
transform -1 0 3902 0 -1 50386
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_89_27
timestamp 1604489732
transform 1 0 2522 0 1 50386
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1604489732
transform -1 0 3902 0 1 50386
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_90_38
timestamp 1604489732
transform 1 0 3534 0 -1 51474
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_90_32
timestamp 1604489732
transform 1 0 2982 0 -1 51474
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_90_27
timestamp 1604489732
transform 1 0 2522 0 -1 51474
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1408
timestamp 1604489732
transform 1 0 2890 0 -1 51474
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1604489732
transform -1 0 3902 0 -1 51474
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_858
timestamp 1604489732
transform 1 0 83298 0 -1 50386
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_860
timestamp 1604489732
transform 1 0 83298 0 1 50386
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_862
timestamp 1604489732
transform 1 0 83298 0 -1 51474
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_88_908
timestamp 1604489732
transform 1 0 83574 0 -1 50386
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_908
timestamp 1604489732
transform 1 0 83574 0 1 50386
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_908
timestamp 1604489732
transform 1 0 83574 0 -1 51474
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_937
timestamp 1604489732
transform 1 0 86242 0 -1 50386
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_932
timestamp 1604489732
transform 1 0 85782 0 -1 50386
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_88_920
timestamp 1604489732
transform 1 0 84678 0 -1 50386
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1579
timestamp 1604489732
transform 1 0 86150 0 -1 50386
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_932
timestamp 1604489732
transform 1 0 85782 0 1 50386
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_920
timestamp 1604489732
transform 1 0 84678 0 1 50386
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_937
timestamp 1604489732
transform 1 0 86242 0 -1 51474
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_932
timestamp 1604489732
transform 1 0 85782 0 -1 51474
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_90_920
timestamp 1604489732
transform 1 0 84678 0 -1 51474
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1580
timestamp 1604489732
transform 1 0 86150 0 -1 51474
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_859
timestamp 1604489732
transform -1 0 87806 0 -1 50386
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_861
timestamp 1604489732
transform -1 0 87806 0 1 50386
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_863
timestamp 1604489732
transform -1 0 87806 0 -1 51474
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_88_949
timestamp 1604489732
transform 1 0 87346 0 -1 50386
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_89_944
timestamp 1604489732
transform 1 0 86886 0 1 50386
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_950
timestamp 1604489732
transform 1 0 87438 0 1 50386
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_949
timestamp 1604489732
transform 1 0 87346 0 -1 51474
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1604489732
transform 1 0 38 0 1 51474
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1604489732
transform 1 0 38 0 -1 52562
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1604489732
transform 1 0 38 0 1 52562
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_3
timestamp 1604489732
transform 1 0 314 0 1 51474
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_15
timestamp 1604489732
transform 1 0 1418 0 1 51474
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_3
timestamp 1604489732
transform 1 0 314 0 -1 52562
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_15
timestamp 1604489732
transform 1 0 1418 0 -1 52562
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_3
timestamp 1604489732
transform 1 0 314 0 1 52562
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_15
timestamp 1604489732
transform 1 0 1418 0 1 52562
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1604489732
transform -1 0 3902 0 1 51474
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1604489732
transform -1 0 3902 0 -1 52562
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1604489732
transform -1 0 3902 0 1 52562
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1409
timestamp 1604489732
transform 1 0 2890 0 -1 52562
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_27
timestamp 1604489732
transform 1 0 2522 0 1 51474
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_27
timestamp 1604489732
transform 1 0 2522 0 -1 52562
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_92_32
timestamp 1604489732
transform 1 0 2982 0 -1 52562
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_38
timestamp 1604489732
transform 1 0 3534 0 -1 52562
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_27
timestamp 1604489732
transform 1 0 2522 0 1 52562
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_864
timestamp 1604489732
transform 1 0 83298 0 1 51474
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_866
timestamp 1604489732
transform 1 0 83298 0 -1 52562
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_868
timestamp 1604489732
transform 1 0 83298 0 1 52562
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_908
timestamp 1604489732
transform 1 0 83574 0 1 51474
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_908
timestamp 1604489732
transform 1 0 83574 0 -1 52562
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_908
timestamp 1604489732
transform 1 0 83574 0 1 52562
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1581
timestamp 1604489732
transform 1 0 86150 0 -1 52562
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_920
timestamp 1604489732
transform 1 0 84678 0 1 51474
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_932
timestamp 1604489732
transform 1 0 85782 0 1 51474
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_920
timestamp 1604489732
transform 1 0 84678 0 -1 52562
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_932
timestamp 1604489732
transform 1 0 85782 0 -1 52562
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_92_937
timestamp 1604489732
transform 1 0 86242 0 -1 52562
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_920
timestamp 1604489732
transform 1 0 84678 0 1 52562
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_932
timestamp 1604489732
transform 1 0 85782 0 1 52562
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_865
timestamp 1604489732
transform -1 0 87806 0 1 51474
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_867
timestamp 1604489732
transform -1 0 87806 0 -1 52562
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_869
timestamp 1604489732
transform -1 0 87806 0 1 52562
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_91_944
timestamp 1604489732
transform 1 0 86886 0 1 51474
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_950
timestamp 1604489732
transform 1 0 87438 0 1 51474
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_949
timestamp 1604489732
transform 1 0 87346 0 -1 52562
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_93_944
timestamp 1604489732
transform 1 0 86886 0 1 52562
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_950
timestamp 1604489732
transform 1 0 87438 0 1 52562
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_15
timestamp 1604489732
transform 1 0 1418 0 1 53650
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_3
timestamp 1604489732
transform 1 0 314 0 1 53650
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_15
timestamp 1604489732
transform 1 0 1418 0 -1 53650
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_3
timestamp 1604489732
transform 1 0 314 0 -1 53650
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1604489732
transform 1 0 38 0 1 53650
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1604489732
transform 1 0 38 0 -1 53650
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_15
timestamp 1604489732
transform 1 0 1418 0 -1 54738
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_3
timestamp 1604489732
transform 1 0 314 0 -1 54738
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1604489732
transform 1 0 38 0 -1 54738
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_15
timestamp 1604489732
transform 1 0 1418 0 1 54738
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_3
timestamp 1604489732
transform 1 0 314 0 1 54738
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1604489732
transform 1 0 38 0 1 54738
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_95_27
timestamp 1604489732
transform 1 0 2522 0 1 53650
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_38
timestamp 1604489732
transform 1 0 3534 0 -1 53650
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_94_32
timestamp 1604489732
transform 1 0 2982 0 -1 53650
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_94_27
timestamp 1604489732
transform 1 0 2522 0 -1 53650
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1410
timestamp 1604489732
transform 1 0 2890 0 -1 53650
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1604489732
transform -1 0 3902 0 1 53650
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1604489732
transform -1 0 3902 0 -1 53650
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_96_38
timestamp 1604489732
transform 1 0 3534 0 -1 54738
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_96_32
timestamp 1604489732
transform 1 0 2982 0 -1 54738
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_96_27
timestamp 1604489732
transform 1 0 2522 0 -1 54738
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1411
timestamp 1604489732
transform 1 0 2890 0 -1 54738
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1604489732
transform -1 0 3902 0 -1 54738
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_27
timestamp 1604489732
transform 1 0 2522 0 1 54738
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1604489732
transform -1 0 3902 0 1 54738
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_870
timestamp 1604489732
transform 1 0 83298 0 -1 53650
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_872
timestamp 1604489732
transform 1 0 83298 0 1 53650
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_874
timestamp 1604489732
transform 1 0 83298 0 -1 54738
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_876
timestamp 1604489732
transform 1 0 83298 0 1 54738
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_94_908
timestamp 1604489732
transform 1 0 83574 0 -1 53650
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_908
timestamp 1604489732
transform 1 0 83574 0 1 53650
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_908
timestamp 1604489732
transform 1 0 83574 0 -1 54738
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_908
timestamp 1604489732
transform 1 0 83574 0 1 54738
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_932
timestamp 1604489732
transform 1 0 85782 0 1 53650
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_920
timestamp 1604489732
transform 1 0 84678 0 1 53650
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_937
timestamp 1604489732
transform 1 0 86242 0 -1 53650
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_932
timestamp 1604489732
transform 1 0 85782 0 -1 53650
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_94_920
timestamp 1604489732
transform 1 0 84678 0 -1 53650
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1582
timestamp 1604489732
transform 1 0 86150 0 -1 53650
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_937
timestamp 1604489732
transform 1 0 86242 0 -1 54738
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_932
timestamp 1604489732
transform 1 0 85782 0 -1 54738
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_96_920
timestamp 1604489732
transform 1 0 84678 0 -1 54738
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1583
timestamp 1604489732
transform 1 0 86150 0 -1 54738
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_932
timestamp 1604489732
transform 1 0 85782 0 1 54738
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_920
timestamp 1604489732
transform 1 0 84678 0 1 54738
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_944
timestamp 1604489732
transform 1 0 86886 0 1 53650
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_950
timestamp 1604489732
transform 1 0 87438 0 1 53650
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_949
timestamp 1604489732
transform 1 0 87346 0 -1 53650
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_873
timestamp 1604489732
transform -1 0 87806 0 1 53650
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_871
timestamp 1604489732
transform -1 0 87806 0 -1 53650
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_96_949
timestamp 1604489732
transform 1 0 87346 0 -1 54738
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_875
timestamp 1604489732
transform -1 0 87806 0 -1 54738
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_97_944
timestamp 1604489732
transform 1 0 86886 0 1 54738
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_950
timestamp 1604489732
transform 1 0 87438 0 1 54738
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_877
timestamp 1604489732
transform -1 0 87806 0 1 54738
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1604489732
transform 1 0 38 0 -1 55826
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1604489732
transform 1 0 38 0 1 55826
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1604489732
transform 1 0 38 0 -1 56914
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_98_3
timestamp 1604489732
transform 1 0 314 0 -1 55826
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_15
timestamp 1604489732
transform 1 0 1418 0 -1 55826
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_3
timestamp 1604489732
transform 1 0 314 0 1 55826
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_15
timestamp 1604489732
transform 1 0 1418 0 1 55826
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_3
timestamp 1604489732
transform 1 0 314 0 -1 56914
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_15
timestamp 1604489732
transform 1 0 1418 0 -1 56914
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_38
timestamp 1604489732
transform 1 0 3534 0 -1 55826
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_98_32
timestamp 1604489732
transform 1 0 2982 0 -1 55826
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_98_27
timestamp 1604489732
transform 1 0 2522 0 -1 55826
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1412
timestamp 1604489732
transform 1 0 2890 0 -1 55826
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1604489732
transform -1 0 3902 0 -1 55826
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_99_27
timestamp 1604489732
transform 1 0 2522 0 1 55826
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1604489732
transform -1 0 3902 0 1 55826
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_100_38
timestamp 1604489732
transform 1 0 3534 0 -1 56914
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_100_32
timestamp 1604489732
transform 1 0 2982 0 -1 56914
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_100_27
timestamp 1604489732
transform 1 0 2522 0 -1 56914
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1413
timestamp 1604489732
transform 1 0 2890 0 -1 56914
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1604489732
transform -1 0 3902 0 -1 56914
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_878
timestamp 1604489732
transform 1 0 83298 0 -1 55826
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_880
timestamp 1604489732
transform 1 0 83298 0 1 55826
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_882
timestamp 1604489732
transform 1 0 83298 0 -1 56914
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_98_908
timestamp 1604489732
transform 1 0 83574 0 -1 55826
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_908
timestamp 1604489732
transform 1 0 83574 0 1 55826
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_908
timestamp 1604489732
transform 1 0 83574 0 -1 56914
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_937
timestamp 1604489732
transform 1 0 86242 0 -1 55826
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_932
timestamp 1604489732
transform 1 0 85782 0 -1 55826
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_98_920
timestamp 1604489732
transform 1 0 84678 0 -1 55826
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1584
timestamp 1604489732
transform 1 0 86150 0 -1 55826
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_932
timestamp 1604489732
transform 1 0 85782 0 1 55826
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_920
timestamp 1604489732
transform 1 0 84678 0 1 55826
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_937
timestamp 1604489732
transform 1 0 86242 0 -1 56914
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_932
timestamp 1604489732
transform 1 0 85782 0 -1 56914
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_100_920
timestamp 1604489732
transform 1 0 84678 0 -1 56914
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1585
timestamp 1604489732
transform 1 0 86150 0 -1 56914
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_879
timestamp 1604489732
transform -1 0 87806 0 -1 55826
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_881
timestamp 1604489732
transform -1 0 87806 0 1 55826
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_883
timestamp 1604489732
transform -1 0 87806 0 -1 56914
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_98_949
timestamp 1604489732
transform 1 0 87346 0 -1 55826
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_99_944
timestamp 1604489732
transform 1 0 86886 0 1 55826
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_950
timestamp 1604489732
transform 1 0 87438 0 1 55826
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_100_949
timestamp 1604489732
transform 1 0 87346 0 -1 56914
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_101_15
timestamp 1604489732
transform 1 0 1418 0 1 56914
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_3
timestamp 1604489732
transform 1 0 314 0 1 56914
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1604489732
transform 1 0 38 0 1 56914
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_15
timestamp 1604489732
transform 1 0 1418 0 1 58002
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_3
timestamp 1604489732
transform 1 0 314 0 1 58002
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_15
timestamp 1604489732
transform 1 0 1418 0 -1 58002
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_3
timestamp 1604489732
transform 1 0 314 0 -1 58002
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1604489732
transform 1 0 38 0 1 58002
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1604489732
transform 1 0 38 0 -1 58002
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_104_15
timestamp 1604489732
transform 1 0 1418 0 -1 59090
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_3
timestamp 1604489732
transform 1 0 314 0 -1 59090
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1604489732
transform 1 0 38 0 -1 59090
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_27
timestamp 1604489732
transform 1 0 2522 0 1 56914
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1604489732
transform -1 0 3902 0 1 56914
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_27
timestamp 1604489732
transform 1 0 2522 0 1 58002
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_38
timestamp 1604489732
transform 1 0 3534 0 -1 58002
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_102_32
timestamp 1604489732
transform 1 0 2982 0 -1 58002
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_102_27
timestamp 1604489732
transform 1 0 2522 0 -1 58002
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1414
timestamp 1604489732
transform 1 0 2890 0 -1 58002
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1604489732
transform -1 0 3902 0 1 58002
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1604489732
transform -1 0 3902 0 -1 58002
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_104_38
timestamp 1604489732
transform 1 0 3534 0 -1 59090
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_104_32
timestamp 1604489732
transform 1 0 2982 0 -1 59090
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_104_27
timestamp 1604489732
transform 1 0 2522 0 -1 59090
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1415
timestamp 1604489732
transform 1 0 2890 0 -1 59090
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1604489732
transform -1 0 3902 0 -1 59090
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_884
timestamp 1604489732
transform 1 0 83298 0 1 56914
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_886
timestamp 1604489732
transform 1 0 83298 0 -1 58002
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_888
timestamp 1604489732
transform 1 0 83298 0 1 58002
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_890
timestamp 1604489732
transform 1 0 83298 0 -1 59090
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_908
timestamp 1604489732
transform 1 0 83574 0 1 56914
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_908
timestamp 1604489732
transform 1 0 83574 0 -1 58002
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_908
timestamp 1604489732
transform 1 0 83574 0 1 58002
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_908
timestamp 1604489732
transform 1 0 83574 0 -1 59090
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_932
timestamp 1604489732
transform 1 0 85782 0 1 56914
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_920
timestamp 1604489732
transform 1 0 84678 0 1 56914
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_932
timestamp 1604489732
transform 1 0 85782 0 1 58002
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_920
timestamp 1604489732
transform 1 0 84678 0 1 58002
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_937
timestamp 1604489732
transform 1 0 86242 0 -1 58002
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_102_932
timestamp 1604489732
transform 1 0 85782 0 -1 58002
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_102_920
timestamp 1604489732
transform 1 0 84678 0 -1 58002
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1586
timestamp 1604489732
transform 1 0 86150 0 -1 58002
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_937
timestamp 1604489732
transform 1 0 86242 0 -1 59090
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_104_932
timestamp 1604489732
transform 1 0 85782 0 -1 59090
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_104_920
timestamp 1604489732
transform 1 0 84678 0 -1 59090
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1587
timestamp 1604489732
transform 1 0 86150 0 -1 59090
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_944
timestamp 1604489732
transform 1 0 86886 0 1 56914
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_950
timestamp 1604489732
transform 1 0 87438 0 1 56914
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_885
timestamp 1604489732
transform -1 0 87806 0 1 56914
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_103_944
timestamp 1604489732
transform 1 0 86886 0 1 58002
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_950
timestamp 1604489732
transform 1 0 87438 0 1 58002
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_102_949
timestamp 1604489732
transform 1 0 87346 0 -1 58002
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_889
timestamp 1604489732
transform -1 0 87806 0 1 58002
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_887
timestamp 1604489732
transform -1 0 87806 0 -1 58002
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_104_949
timestamp 1604489732
transform 1 0 87346 0 -1 59090
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_891
timestamp 1604489732
transform -1 0 87806 0 -1 59090
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1604489732
transform 1 0 38 0 1 59090
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1604489732
transform 1 0 38 0 -1 60178
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1604489732
transform 1 0 38 0 1 60178
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_105_3
timestamp 1604489732
transform 1 0 314 0 1 59090
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_15
timestamp 1604489732
transform 1 0 1418 0 1 59090
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_3
timestamp 1604489732
transform 1 0 314 0 -1 60178
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_15
timestamp 1604489732
transform 1 0 1418 0 -1 60178
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_3
timestamp 1604489732
transform 1 0 314 0 1 60178
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_15
timestamp 1604489732
transform 1 0 1418 0 1 60178
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1604489732
transform -1 0 3902 0 1 59090
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1604489732
transform -1 0 3902 0 -1 60178
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1604489732
transform -1 0 3902 0 1 60178
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1416
timestamp 1604489732
transform 1 0 2890 0 -1 60178
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_27
timestamp 1604489732
transform 1 0 2522 0 1 59090
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_27
timestamp 1604489732
transform 1 0 2522 0 -1 60178
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_106_32
timestamp 1604489732
transform 1 0 2982 0 -1 60178
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_38
timestamp 1604489732
transform 1 0 3534 0 -1 60178
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_27
timestamp 1604489732
transform 1 0 2522 0 1 60178
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_892
timestamp 1604489732
transform 1 0 83298 0 1 59090
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_894
timestamp 1604489732
transform 1 0 83298 0 -1 60178
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_896
timestamp 1604489732
transform 1 0 83298 0 1 60178
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_105_908
timestamp 1604489732
transform 1 0 83574 0 1 59090
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_908
timestamp 1604489732
transform 1 0 83574 0 -1 60178
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_908
timestamp 1604489732
transform 1 0 83574 0 1 60178
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1588
timestamp 1604489732
transform 1 0 86150 0 -1 60178
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_920
timestamp 1604489732
transform 1 0 84678 0 1 59090
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_932
timestamp 1604489732
transform 1 0 85782 0 1 59090
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_920
timestamp 1604489732
transform 1 0 84678 0 -1 60178
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_932
timestamp 1604489732
transform 1 0 85782 0 -1 60178
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_106_937
timestamp 1604489732
transform 1 0 86242 0 -1 60178
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_920
timestamp 1604489732
transform 1 0 84678 0 1 60178
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_932
timestamp 1604489732
transform 1 0 85782 0 1 60178
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_893
timestamp 1604489732
transform -1 0 87806 0 1 59090
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_895
timestamp 1604489732
transform -1 0 87806 0 -1 60178
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_897
timestamp 1604489732
transform -1 0 87806 0 1 60178
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_105_944
timestamp 1604489732
transform 1 0 86886 0 1 59090
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_950
timestamp 1604489732
transform 1 0 87438 0 1 59090
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_106_949
timestamp 1604489732
transform 1 0 87346 0 -1 60178
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_107_944
timestamp 1604489732
transform 1 0 86886 0 1 60178
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_950
timestamp 1604489732
transform 1 0 87438 0 1 60178
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1604489732
transform 1 0 38 0 -1 61266
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1604489732
transform 1 0 38 0 1 61266
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1604489732
transform 1 0 38 0 -1 62354
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_108_3
timestamp 1604489732
transform 1 0 314 0 -1 61266
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_15
timestamp 1604489732
transform 1 0 1418 0 -1 61266
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_3
timestamp 1604489732
transform 1 0 314 0 1 61266
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_15
timestamp 1604489732
transform 1 0 1418 0 1 61266
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_3
timestamp 1604489732
transform 1 0 314 0 -1 62354
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_15
timestamp 1604489732
transform 1 0 1418 0 -1 62354
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_38
timestamp 1604489732
transform 1 0 3534 0 -1 61266
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_108_32
timestamp 1604489732
transform 1 0 2982 0 -1 61266
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_108_27
timestamp 1604489732
transform 1 0 2522 0 -1 61266
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1417
timestamp 1604489732
transform 1 0 2890 0 -1 61266
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1604489732
transform -1 0 3902 0 -1 61266
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_109_27
timestamp 1604489732
transform 1 0 2522 0 1 61266
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1604489732
transform -1 0 3902 0 1 61266
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_110_38
timestamp 1604489732
transform 1 0 3534 0 -1 62354
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_110_32
timestamp 1604489732
transform 1 0 2982 0 -1 62354
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_110_27
timestamp 1604489732
transform 1 0 2522 0 -1 62354
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1418
timestamp 1604489732
transform 1 0 2890 0 -1 62354
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1604489732
transform -1 0 3902 0 -1 62354
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_898
timestamp 1604489732
transform 1 0 83298 0 -1 61266
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_900
timestamp 1604489732
transform 1 0 83298 0 1 61266
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_902
timestamp 1604489732
transform 1 0 83298 0 -1 62354
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_108_908
timestamp 1604489732
transform 1 0 83574 0 -1 61266
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_908
timestamp 1604489732
transform 1 0 83574 0 1 61266
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_908
timestamp 1604489732
transform 1 0 83574 0 -1 62354
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_937
timestamp 1604489732
transform 1 0 86242 0 -1 61266
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_108_932
timestamp 1604489732
transform 1 0 85782 0 -1 61266
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_108_920
timestamp 1604489732
transform 1 0 84678 0 -1 61266
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1589
timestamp 1604489732
transform 1 0 86150 0 -1 61266
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_932
timestamp 1604489732
transform 1 0 85782 0 1 61266
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_920
timestamp 1604489732
transform 1 0 84678 0 1 61266
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_937
timestamp 1604489732
transform 1 0 86242 0 -1 62354
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_110_932
timestamp 1604489732
transform 1 0 85782 0 -1 62354
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_110_920
timestamp 1604489732
transform 1 0 84678 0 -1 62354
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1590
timestamp 1604489732
transform 1 0 86150 0 -1 62354
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_899
timestamp 1604489732
transform -1 0 87806 0 -1 61266
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_901
timestamp 1604489732
transform -1 0 87806 0 1 61266
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_903
timestamp 1604489732
transform -1 0 87806 0 -1 62354
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_108_949
timestamp 1604489732
transform 1 0 87346 0 -1 61266
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_109_944
timestamp 1604489732
transform 1 0 86886 0 1 61266
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_950
timestamp 1604489732
transform 1 0 87438 0 1 61266
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_110_949
timestamp 1604489732
transform 1 0 87346 0 -1 62354
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_112_15
timestamp 1604489732
transform 1 0 1418 0 -1 63442
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_3
timestamp 1604489732
transform 1 0 314 0 -1 63442
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_15
timestamp 1604489732
transform 1 0 1418 0 1 62354
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_3
timestamp 1604489732
transform 1 0 314 0 1 62354
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1604489732
transform 1 0 38 0 -1 63442
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1604489732
transform 1 0 38 0 1 62354
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_113_15
timestamp 1604489732
transform 1 0 1418 0 1 63442
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_3
timestamp 1604489732
transform 1 0 314 0 1 63442
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1604489732
transform 1 0 38 0 1 63442
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_114_15
timestamp 1604489732
transform 1 0 1418 0 -1 64530
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_3
timestamp 1604489732
transform 1 0 314 0 -1 64530
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1604489732
transform 1 0 38 0 -1 64530
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_112_38
timestamp 1604489732
transform 1 0 3534 0 -1 63442
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_112_32
timestamp 1604489732
transform 1 0 2982 0 -1 63442
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_112_27
timestamp 1604489732
transform 1 0 2522 0 -1 63442
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_111_27
timestamp 1604489732
transform 1 0 2522 0 1 62354
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1419
timestamp 1604489732
transform 1 0 2890 0 -1 63442
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1604489732
transform -1 0 3902 0 -1 63442
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1604489732
transform -1 0 3902 0 1 62354
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_113_27
timestamp 1604489732
transform 1 0 2522 0 1 63442
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1604489732
transform -1 0 3902 0 1 63442
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_114_38
timestamp 1604489732
transform 1 0 3534 0 -1 64530
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_114_32
timestamp 1604489732
transform 1 0 2982 0 -1 64530
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_114_27
timestamp 1604489732
transform 1 0 2522 0 -1 64530
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1420
timestamp 1604489732
transform 1 0 2890 0 -1 64530
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1604489732
transform -1 0 3902 0 -1 64530
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_904
timestamp 1604489732
transform 1 0 83298 0 1 62354
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_906
timestamp 1604489732
transform 1 0 83298 0 -1 63442
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_908
timestamp 1604489732
transform 1 0 83298 0 1 63442
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_910
timestamp 1604489732
transform 1 0 83298 0 -1 64530
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_111_908
timestamp 1604489732
transform 1 0 83574 0 1 62354
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_908
timestamp 1604489732
transform 1 0 83574 0 -1 63442
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_908
timestamp 1604489732
transform 1 0 83574 0 1 63442
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_908
timestamp 1604489732
transform 1 0 83574 0 -1 64530
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_937
timestamp 1604489732
transform 1 0 86242 0 -1 63442
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_112_932
timestamp 1604489732
transform 1 0 85782 0 -1 63442
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_112_920
timestamp 1604489732
transform 1 0 84678 0 -1 63442
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_932
timestamp 1604489732
transform 1 0 85782 0 1 62354
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_920
timestamp 1604489732
transform 1 0 84678 0 1 62354
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1591
timestamp 1604489732
transform 1 0 86150 0 -1 63442
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_932
timestamp 1604489732
transform 1 0 85782 0 1 63442
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_920
timestamp 1604489732
transform 1 0 84678 0 1 63442
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_937
timestamp 1604489732
transform 1 0 86242 0 -1 64530
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_114_932
timestamp 1604489732
transform 1 0 85782 0 -1 64530
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_114_920
timestamp 1604489732
transform 1 0 84678 0 -1 64530
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1592
timestamp 1604489732
transform 1 0 86150 0 -1 64530
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_111_944
timestamp 1604489732
transform 1 0 86886 0 1 62354
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_112_949
timestamp 1604489732
transform 1 0 87346 0 -1 63442
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_111_950
timestamp 1604489732
transform 1 0 87438 0 1 62354
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_907
timestamp 1604489732
transform -1 0 87806 0 -1 63442
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_905
timestamp 1604489732
transform -1 0 87806 0 1 62354
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_113_944
timestamp 1604489732
transform 1 0 86886 0 1 63442
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_950
timestamp 1604489732
transform 1 0 87438 0 1 63442
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_909
timestamp 1604489732
transform -1 0 87806 0 1 63442
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_114_949
timestamp 1604489732
transform 1 0 87346 0 -1 64530
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_911
timestamp 1604489732
transform -1 0 87806 0 -1 64530
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1604489732
transform 1 0 38 0 1 64530
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_230
timestamp 1604489732
transform 1 0 38 0 -1 65618
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_232
timestamp 1604489732
transform 1 0 38 0 1 65618
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_115_3
timestamp 1604489732
transform 1 0 314 0 1 64530
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_15
timestamp 1604489732
transform 1 0 1418 0 1 64530
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_3
timestamp 1604489732
transform 1 0 314 0 -1 65618
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_15
timestamp 1604489732
transform 1 0 1418 0 -1 65618
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_3
timestamp 1604489732
transform 1 0 314 0 1 65618
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_15
timestamp 1604489732
transform 1 0 1418 0 1 65618
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1604489732
transform -1 0 3902 0 1 64530
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_231
timestamp 1604489732
transform -1 0 3902 0 -1 65618
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_233
timestamp 1604489732
transform -1 0 3902 0 1 65618
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1421
timestamp 1604489732
transform 1 0 2890 0 -1 65618
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_27
timestamp 1604489732
transform 1 0 2522 0 1 64530
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_116_27
timestamp 1604489732
transform 1 0 2522 0 -1 65618
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_116_32
timestamp 1604489732
transform 1 0 2982 0 -1 65618
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_38
timestamp 1604489732
transform 1 0 3534 0 -1 65618
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_27
timestamp 1604489732
transform 1 0 2522 0 1 65618
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_912
timestamp 1604489732
transform 1 0 83298 0 1 64530
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_914
timestamp 1604489732
transform 1 0 83298 0 -1 65618
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_916
timestamp 1604489732
transform 1 0 83298 0 1 65618
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_115_908
timestamp 1604489732
transform 1 0 83574 0 1 64530
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_908
timestamp 1604489732
transform 1 0 83574 0 -1 65618
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_908
timestamp 1604489732
transform 1 0 83574 0 1 65618
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1593
timestamp 1604489732
transform 1 0 86150 0 -1 65618
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_920
timestamp 1604489732
transform 1 0 84678 0 1 64530
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_932
timestamp 1604489732
transform 1 0 85782 0 1 64530
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_920
timestamp 1604489732
transform 1 0 84678 0 -1 65618
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_116_932
timestamp 1604489732
transform 1 0 85782 0 -1 65618
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_116_937
timestamp 1604489732
transform 1 0 86242 0 -1 65618
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_920
timestamp 1604489732
transform 1 0 84678 0 1 65618
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_932
timestamp 1604489732
transform 1 0 85782 0 1 65618
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_913
timestamp 1604489732
transform -1 0 87806 0 1 64530
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_915
timestamp 1604489732
transform -1 0 87806 0 -1 65618
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_917
timestamp 1604489732
transform -1 0 87806 0 1 65618
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_115_944
timestamp 1604489732
transform 1 0 86886 0 1 64530
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_950
timestamp 1604489732
transform 1 0 87438 0 1 64530
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_116_949
timestamp 1604489732
transform 1 0 87346 0 -1 65618
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_117_944
timestamp 1604489732
transform 1 0 86886 0 1 65618
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_950
timestamp 1604489732
transform 1 0 87438 0 1 65618
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_234
timestamp 1604489732
transform 1 0 38 0 -1 66706
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_236
timestamp 1604489732
transform 1 0 38 0 1 66706
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_238
timestamp 1604489732
transform 1 0 38 0 -1 67794
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_118_3
timestamp 1604489732
transform 1 0 314 0 -1 66706
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_15
timestamp 1604489732
transform 1 0 1418 0 -1 66706
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_3
timestamp 1604489732
transform 1 0 314 0 1 66706
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_15
timestamp 1604489732
transform 1 0 1418 0 1 66706
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_3
timestamp 1604489732
transform 1 0 314 0 -1 67794
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_15
timestamp 1604489732
transform 1 0 1418 0 -1 67794
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_118_38
timestamp 1604489732
transform 1 0 3534 0 -1 66706
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_118_32
timestamp 1604489732
transform 1 0 2982 0 -1 66706
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_118_27
timestamp 1604489732
transform 1 0 2522 0 -1 66706
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1422
timestamp 1604489732
transform 1 0 2890 0 -1 66706
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_235
timestamp 1604489732
transform -1 0 3902 0 -1 66706
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_119_27
timestamp 1604489732
transform 1 0 2522 0 1 66706
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_237
timestamp 1604489732
transform -1 0 3902 0 1 66706
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_120_38
timestamp 1604489732
transform 1 0 3534 0 -1 67794
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_120_32
timestamp 1604489732
transform 1 0 2982 0 -1 67794
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_120_27
timestamp 1604489732
transform 1 0 2522 0 -1 67794
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1423
timestamp 1604489732
transform 1 0 2890 0 -1 67794
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_239
timestamp 1604489732
transform -1 0 3902 0 -1 67794
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_918
timestamp 1604489732
transform 1 0 83298 0 -1 66706
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_920
timestamp 1604489732
transform 1 0 83298 0 1 66706
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_922
timestamp 1604489732
transform 1 0 83298 0 -1 67794
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_118_908
timestamp 1604489732
transform 1 0 83574 0 -1 66706
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_908
timestamp 1604489732
transform 1 0 83574 0 1 66706
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_908
timestamp 1604489732
transform 1 0 83574 0 -1 67794
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_937
timestamp 1604489732
transform 1 0 86242 0 -1 66706
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_118_932
timestamp 1604489732
transform 1 0 85782 0 -1 66706
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_118_920
timestamp 1604489732
transform 1 0 84678 0 -1 66706
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1594
timestamp 1604489732
transform 1 0 86150 0 -1 66706
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_932
timestamp 1604489732
transform 1 0 85782 0 1 66706
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_920
timestamp 1604489732
transform 1 0 84678 0 1 66706
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_937
timestamp 1604489732
transform 1 0 86242 0 -1 67794
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_120_932
timestamp 1604489732
transform 1 0 85782 0 -1 67794
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_120_920
timestamp 1604489732
transform 1 0 84678 0 -1 67794
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1595
timestamp 1604489732
transform 1 0 86150 0 -1 67794
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_919
timestamp 1604489732
transform -1 0 87806 0 -1 66706
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_921
timestamp 1604489732
transform -1 0 87806 0 1 66706
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_923
timestamp 1604489732
transform -1 0 87806 0 -1 67794
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_118_949
timestamp 1604489732
transform 1 0 87346 0 -1 66706
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_119_944
timestamp 1604489732
transform 1 0 86886 0 1 66706
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_950
timestamp 1604489732
transform 1 0 87438 0 1 66706
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_120_949
timestamp 1604489732
transform 1 0 87346 0 -1 67794
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_122_15
timestamp 1604489732
transform 1 0 1418 0 -1 68882
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_3
timestamp 1604489732
transform 1 0 314 0 -1 68882
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_15
timestamp 1604489732
transform 1 0 1418 0 1 67794
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_3
timestamp 1604489732
transform 1 0 314 0 1 67794
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_242
timestamp 1604489732
transform 1 0 38 0 -1 68882
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_240
timestamp 1604489732
transform 1 0 38 0 1 67794
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_15
timestamp 1604489732
transform 1 0 1418 0 1 68882
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_3
timestamp 1604489732
transform 1 0 314 0 1 68882
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_244
timestamp 1604489732
transform 1 0 38 0 1 68882
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_124_15
timestamp 1604489732
transform 1 0 1418 0 -1 69970
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_3
timestamp 1604489732
transform 1 0 314 0 -1 69970
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_246
timestamp 1604489732
transform 1 0 38 0 -1 69970
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_122_38
timestamp 1604489732
transform 1 0 3534 0 -1 68882
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_122_32
timestamp 1604489732
transform 1 0 2982 0 -1 68882
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_122_27
timestamp 1604489732
transform 1 0 2522 0 -1 68882
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_121_27
timestamp 1604489732
transform 1 0 2522 0 1 67794
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1424
timestamp 1604489732
transform 1 0 2890 0 -1 68882
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_243
timestamp 1604489732
transform -1 0 3902 0 -1 68882
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_241
timestamp 1604489732
transform -1 0 3902 0 1 67794
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_27
timestamp 1604489732
transform 1 0 2522 0 1 68882
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_245
timestamp 1604489732
transform -1 0 3902 0 1 68882
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_124_38
timestamp 1604489732
transform 1 0 3534 0 -1 69970
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_124_32
timestamp 1604489732
transform 1 0 2982 0 -1 69970
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_124_27
timestamp 1604489732
transform 1 0 2522 0 -1 69970
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1425
timestamp 1604489732
transform 1 0 2890 0 -1 69970
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_247
timestamp 1604489732
transform -1 0 3902 0 -1 69970
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_924
timestamp 1604489732
transform 1 0 83298 0 1 67794
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_926
timestamp 1604489732
transform 1 0 83298 0 -1 68882
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_928
timestamp 1604489732
transform 1 0 83298 0 1 68882
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_930
timestamp 1604489732
transform 1 0 83298 0 -1 69970
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_121_908
timestamp 1604489732
transform 1 0 83574 0 1 67794
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_908
timestamp 1604489732
transform 1 0 83574 0 -1 68882
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_908
timestamp 1604489732
transform 1 0 83574 0 1 68882
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_908
timestamp 1604489732
transform 1 0 83574 0 -1 69970
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_937
timestamp 1604489732
transform 1 0 86242 0 -1 68882
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_122_932
timestamp 1604489732
transform 1 0 85782 0 -1 68882
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_122_920
timestamp 1604489732
transform 1 0 84678 0 -1 68882
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_932
timestamp 1604489732
transform 1 0 85782 0 1 67794
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_920
timestamp 1604489732
transform 1 0 84678 0 1 67794
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1596
timestamp 1604489732
transform 1 0 86150 0 -1 68882
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_932
timestamp 1604489732
transform 1 0 85782 0 1 68882
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_920
timestamp 1604489732
transform 1 0 84678 0 1 68882
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_937
timestamp 1604489732
transform 1 0 86242 0 -1 69970
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_124_932
timestamp 1604489732
transform 1 0 85782 0 -1 69970
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_124_920
timestamp 1604489732
transform 1 0 84678 0 -1 69970
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1597
timestamp 1604489732
transform 1 0 86150 0 -1 69970
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_121_944
timestamp 1604489732
transform 1 0 86886 0 1 67794
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_122_949
timestamp 1604489732
transform 1 0 87346 0 -1 68882
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_121_950
timestamp 1604489732
transform 1 0 87438 0 1 67794
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_927
timestamp 1604489732
transform -1 0 87806 0 -1 68882
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_925
timestamp 1604489732
transform -1 0 87806 0 1 67794
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_123_944
timestamp 1604489732
transform 1 0 86886 0 1 68882
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_950
timestamp 1604489732
transform 1 0 87438 0 1 68882
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_929
timestamp 1604489732
transform -1 0 87806 0 1 68882
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_124_949
timestamp 1604489732
transform 1 0 87346 0 -1 69970
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_931
timestamp 1604489732
transform -1 0 87806 0 -1 69970
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_248
timestamp 1604489732
transform 1 0 38 0 1 69970
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_250
timestamp 1604489732
transform 1 0 38 0 -1 71058
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_252
timestamp 1604489732
transform 1 0 38 0 1 71058
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_125_3
timestamp 1604489732
transform 1 0 314 0 1 69970
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_15
timestamp 1604489732
transform 1 0 1418 0 1 69970
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_3
timestamp 1604489732
transform 1 0 314 0 -1 71058
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_15
timestamp 1604489732
transform 1 0 1418 0 -1 71058
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_3
timestamp 1604489732
transform 1 0 314 0 1 71058
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_15
timestamp 1604489732
transform 1 0 1418 0 1 71058
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_249
timestamp 1604489732
transform -1 0 3902 0 1 69970
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_251
timestamp 1604489732
transform -1 0 3902 0 -1 71058
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_253
timestamp 1604489732
transform -1 0 3902 0 1 71058
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1426
timestamp 1604489732
transform 1 0 2890 0 -1 71058
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_27
timestamp 1604489732
transform 1 0 2522 0 1 69970
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_126_27
timestamp 1604489732
transform 1 0 2522 0 -1 71058
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_126_32
timestamp 1604489732
transform 1 0 2982 0 -1 71058
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_38
timestamp 1604489732
transform 1 0 3534 0 -1 71058
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_27
timestamp 1604489732
transform 1 0 2522 0 1 71058
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_932
timestamp 1604489732
transform 1 0 83298 0 1 69970
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_934
timestamp 1604489732
transform 1 0 83298 0 -1 71058
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_936
timestamp 1604489732
transform 1 0 83298 0 1 71058
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_125_908
timestamp 1604489732
transform 1 0 83574 0 1 69970
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_908
timestamp 1604489732
transform 1 0 83574 0 -1 71058
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_908
timestamp 1604489732
transform 1 0 83574 0 1 71058
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1598
timestamp 1604489732
transform 1 0 86150 0 -1 71058
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_920
timestamp 1604489732
transform 1 0 84678 0 1 69970
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_932
timestamp 1604489732
transform 1 0 85782 0 1 69970
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_920
timestamp 1604489732
transform 1 0 84678 0 -1 71058
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_126_932
timestamp 1604489732
transform 1 0 85782 0 -1 71058
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_126_937
timestamp 1604489732
transform 1 0 86242 0 -1 71058
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_920
timestamp 1604489732
transform 1 0 84678 0 1 71058
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_932
timestamp 1604489732
transform 1 0 85782 0 1 71058
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_933
timestamp 1604489732
transform -1 0 87806 0 1 69970
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_935
timestamp 1604489732
transform -1 0 87806 0 -1 71058
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_937
timestamp 1604489732
transform -1 0 87806 0 1 71058
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_125_944
timestamp 1604489732
transform 1 0 86886 0 1 69970
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_950
timestamp 1604489732
transform 1 0 87438 0 1 69970
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_126_949
timestamp 1604489732
transform 1 0 87346 0 -1 71058
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_127_944
timestamp 1604489732
transform 1 0 86886 0 1 71058
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_950
timestamp 1604489732
transform 1 0 87438 0 1 71058
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_15
timestamp 1604489732
transform 1 0 1418 0 -1 72146
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_3
timestamp 1604489732
transform 1 0 314 0 -1 72146
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_254
timestamp 1604489732
transform 1 0 38 0 -1 72146
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_130_15
timestamp 1604489732
transform 1 0 1418 0 -1 73234
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_3
timestamp 1604489732
transform 1 0 314 0 -1 73234
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_15
timestamp 1604489732
transform 1 0 1418 0 1 72146
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_3
timestamp 1604489732
transform 1 0 314 0 1 72146
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_258
timestamp 1604489732
transform 1 0 38 0 -1 73234
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_256
timestamp 1604489732
transform 1 0 38 0 1 72146
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_131_15
timestamp 1604489732
transform 1 0 1418 0 1 73234
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_3
timestamp 1604489732
transform 1 0 314 0 1 73234
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_260
timestamp 1604489732
transform 1 0 38 0 1 73234
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_128_38
timestamp 1604489732
transform 1 0 3534 0 -1 72146
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_128_32
timestamp 1604489732
transform 1 0 2982 0 -1 72146
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_128_27
timestamp 1604489732
transform 1 0 2522 0 -1 72146
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1427
timestamp 1604489732
transform 1 0 2890 0 -1 72146
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_255
timestamp 1604489732
transform -1 0 3902 0 -1 72146
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_130_38
timestamp 1604489732
transform 1 0 3534 0 -1 73234
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_130_32
timestamp 1604489732
transform 1 0 2982 0 -1 73234
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_130_27
timestamp 1604489732
transform 1 0 2522 0 -1 73234
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_129_27
timestamp 1604489732
transform 1 0 2522 0 1 72146
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1428
timestamp 1604489732
transform 1 0 2890 0 -1 73234
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_259
timestamp 1604489732
transform -1 0 3902 0 -1 73234
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_257
timestamp 1604489732
transform -1 0 3902 0 1 72146
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_131_27
timestamp 1604489732
transform 1 0 2522 0 1 73234
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_261
timestamp 1604489732
transform -1 0 3902 0 1 73234
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_938
timestamp 1604489732
transform 1 0 83298 0 -1 72146
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_940
timestamp 1604489732
transform 1 0 83298 0 1 72146
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_942
timestamp 1604489732
transform 1 0 83298 0 -1 73234
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_944
timestamp 1604489732
transform 1 0 83298 0 1 73234
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_128_908
timestamp 1604489732
transform 1 0 83574 0 -1 72146
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_908
timestamp 1604489732
transform 1 0 83574 0 1 72146
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_908
timestamp 1604489732
transform 1 0 83574 0 -1 73234
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_908
timestamp 1604489732
transform 1 0 83574 0 1 73234
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_937
timestamp 1604489732
transform 1 0 86242 0 -1 72146
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_128_932
timestamp 1604489732
transform 1 0 85782 0 -1 72146
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_128_920
timestamp 1604489732
transform 1 0 84678 0 -1 72146
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1599
timestamp 1604489732
transform 1 0 86150 0 -1 72146
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_937
timestamp 1604489732
transform 1 0 86242 0 -1 73234
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_130_932
timestamp 1604489732
transform 1 0 85782 0 -1 73234
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_130_920
timestamp 1604489732
transform 1 0 84678 0 -1 73234
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_932
timestamp 1604489732
transform 1 0 85782 0 1 72146
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_920
timestamp 1604489732
transform 1 0 84678 0 1 72146
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1600
timestamp 1604489732
transform 1 0 86150 0 -1 73234
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_932
timestamp 1604489732
transform 1 0 85782 0 1 73234
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_920
timestamp 1604489732
transform 1 0 84678 0 1 73234
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_128_949
timestamp 1604489732
transform 1 0 87346 0 -1 72146
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_939
timestamp 1604489732
transform -1 0 87806 0 -1 72146
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_129_944
timestamp 1604489732
transform 1 0 86886 0 1 72146
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_130_949
timestamp 1604489732
transform 1 0 87346 0 -1 73234
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_129_950
timestamp 1604489732
transform 1 0 87438 0 1 72146
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_943
timestamp 1604489732
transform -1 0 87806 0 -1 73234
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_941
timestamp 1604489732
transform -1 0 87806 0 1 72146
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_131_944
timestamp 1604489732
transform 1 0 86886 0 1 73234
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_950
timestamp 1604489732
transform 1 0 87438 0 1 73234
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_945
timestamp 1604489732
transform -1 0 87806 0 1 73234
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_262
timestamp 1604489732
transform 1 0 38 0 -1 74322
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_264
timestamp 1604489732
transform 1 0 38 0 1 74322
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_266
timestamp 1604489732
transform 1 0 38 0 -1 75410
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_132_3
timestamp 1604489732
transform 1 0 314 0 -1 74322
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_15
timestamp 1604489732
transform 1 0 1418 0 -1 74322
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_3
timestamp 1604489732
transform 1 0 314 0 1 74322
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_15
timestamp 1604489732
transform 1 0 1418 0 1 74322
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_3
timestamp 1604489732
transform 1 0 314 0 -1 75410
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_15
timestamp 1604489732
transform 1 0 1418 0 -1 75410
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_132_38
timestamp 1604489732
transform 1 0 3534 0 -1 74322
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_132_32
timestamp 1604489732
transform 1 0 2982 0 -1 74322
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_132_27
timestamp 1604489732
transform 1 0 2522 0 -1 74322
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1429
timestamp 1604489732
transform 1 0 2890 0 -1 74322
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_263
timestamp 1604489732
transform -1 0 3902 0 -1 74322
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_133_27
timestamp 1604489732
transform 1 0 2522 0 1 74322
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_265
timestamp 1604489732
transform -1 0 3902 0 1 74322
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_134_38
timestamp 1604489732
transform 1 0 3534 0 -1 75410
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_134_32
timestamp 1604489732
transform 1 0 2982 0 -1 75410
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_134_27
timestamp 1604489732
transform 1 0 2522 0 -1 75410
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1430
timestamp 1604489732
transform 1 0 2890 0 -1 75410
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_267
timestamp 1604489732
transform -1 0 3902 0 -1 75410
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_946
timestamp 1604489732
transform 1 0 83298 0 -1 74322
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_948
timestamp 1604489732
transform 1 0 83298 0 1 74322
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_950
timestamp 1604489732
transform 1 0 83298 0 -1 75410
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_132_908
timestamp 1604489732
transform 1 0 83574 0 -1 74322
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_908
timestamp 1604489732
transform 1 0 83574 0 1 74322
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_908
timestamp 1604489732
transform 1 0 83574 0 -1 75410
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_937
timestamp 1604489732
transform 1 0 86242 0 -1 74322
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_132_932
timestamp 1604489732
transform 1 0 85782 0 -1 74322
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_132_920
timestamp 1604489732
transform 1 0 84678 0 -1 74322
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1601
timestamp 1604489732
transform 1 0 86150 0 -1 74322
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_133_932
timestamp 1604489732
transform 1 0 85782 0 1 74322
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_920
timestamp 1604489732
transform 1 0 84678 0 1 74322
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_937
timestamp 1604489732
transform 1 0 86242 0 -1 75410
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_134_932
timestamp 1604489732
transform 1 0 85782 0 -1 75410
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_134_920
timestamp 1604489732
transform 1 0 84678 0 -1 75410
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1602
timestamp 1604489732
transform 1 0 86150 0 -1 75410
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_947
timestamp 1604489732
transform -1 0 87806 0 -1 74322
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_949
timestamp 1604489732
transform -1 0 87806 0 1 74322
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_951
timestamp 1604489732
transform -1 0 87806 0 -1 75410
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_132_949
timestamp 1604489732
transform 1 0 87346 0 -1 74322
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_133_944
timestamp 1604489732
transform 1 0 86886 0 1 74322
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_950
timestamp 1604489732
transform 1 0 87438 0 1 74322
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_134_949
timestamp 1604489732
transform 1 0 87346 0 -1 75410
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_268
timestamp 1604489732
transform 1 0 38 0 1 75410
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_270
timestamp 1604489732
transform 1 0 38 0 -1 76498
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_272
timestamp 1604489732
transform 1 0 38 0 1 76498
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_135_3
timestamp 1604489732
transform 1 0 314 0 1 75410
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_15
timestamp 1604489732
transform 1 0 1418 0 1 75410
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_3
timestamp 1604489732
transform 1 0 314 0 -1 76498
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_15
timestamp 1604489732
transform 1 0 1418 0 -1 76498
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_3
timestamp 1604489732
transform 1 0 314 0 1 76498
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_15
timestamp 1604489732
transform 1 0 1418 0 1 76498
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_269
timestamp 1604489732
transform -1 0 3902 0 1 75410
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_271
timestamp 1604489732
transform -1 0 3902 0 -1 76498
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_273
timestamp 1604489732
transform -1 0 3902 0 1 76498
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1431
timestamp 1604489732
transform 1 0 2890 0 -1 76498
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_27
timestamp 1604489732
transform 1 0 2522 0 1 75410
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_136_27
timestamp 1604489732
transform 1 0 2522 0 -1 76498
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_136_32
timestamp 1604489732
transform 1 0 2982 0 -1 76498
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_38
timestamp 1604489732
transform 1 0 3534 0 -1 76498
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_27
timestamp 1604489732
transform 1 0 2522 0 1 76498
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_952
timestamp 1604489732
transform 1 0 83298 0 1 75410
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_954
timestamp 1604489732
transform 1 0 83298 0 -1 76498
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_956
timestamp 1604489732
transform 1 0 83298 0 1 76498
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_135_908
timestamp 1604489732
transform 1 0 83574 0 1 75410
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_908
timestamp 1604489732
transform 1 0 83574 0 -1 76498
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_908
timestamp 1604489732
transform 1 0 83574 0 1 76498
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1603
timestamp 1604489732
transform 1 0 86150 0 -1 76498
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_920
timestamp 1604489732
transform 1 0 84678 0 1 75410
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_932
timestamp 1604489732
transform 1 0 85782 0 1 75410
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_920
timestamp 1604489732
transform 1 0 84678 0 -1 76498
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_136_932
timestamp 1604489732
transform 1 0 85782 0 -1 76498
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_136_937
timestamp 1604489732
transform 1 0 86242 0 -1 76498
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_920
timestamp 1604489732
transform 1 0 84678 0 1 76498
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_932
timestamp 1604489732
transform 1 0 85782 0 1 76498
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_953
timestamp 1604489732
transform -1 0 87806 0 1 75410
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_955
timestamp 1604489732
transform -1 0 87806 0 -1 76498
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_957
timestamp 1604489732
transform -1 0 87806 0 1 76498
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_135_944
timestamp 1604489732
transform 1 0 86886 0 1 75410
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_950
timestamp 1604489732
transform 1 0 87438 0 1 75410
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_136_949
timestamp 1604489732
transform 1 0 87346 0 -1 76498
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_137_944
timestamp 1604489732
transform 1 0 86886 0 1 76498
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_950
timestamp 1604489732
transform 1 0 87438 0 1 76498
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_139_15
timestamp 1604489732
transform 1 0 1418 0 1 77586
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_3
timestamp 1604489732
transform 1 0 314 0 1 77586
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_15
timestamp 1604489732
transform 1 0 1418 0 -1 77586
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_3
timestamp 1604489732
transform 1 0 314 0 -1 77586
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_276
timestamp 1604489732
transform 1 0 38 0 1 77586
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_274
timestamp 1604489732
transform 1 0 38 0 -1 77586
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_140_15
timestamp 1604489732
transform 1 0 1418 0 -1 78674
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_3
timestamp 1604489732
transform 1 0 314 0 -1 78674
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_278
timestamp 1604489732
transform 1 0 38 0 -1 78674
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_141_15
timestamp 1604489732
transform 1 0 1418 0 1 78674
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_3
timestamp 1604489732
transform 1 0 314 0 1 78674
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_280
timestamp 1604489732
transform 1 0 38 0 1 78674
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_139_27
timestamp 1604489732
transform 1 0 2522 0 1 77586
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_138_38
timestamp 1604489732
transform 1 0 3534 0 -1 77586
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_138_32
timestamp 1604489732
transform 1 0 2982 0 -1 77586
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_138_27
timestamp 1604489732
transform 1 0 2522 0 -1 77586
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1432
timestamp 1604489732
transform 1 0 2890 0 -1 77586
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_277
timestamp 1604489732
transform -1 0 3902 0 1 77586
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_275
timestamp 1604489732
transform -1 0 3902 0 -1 77586
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_140_38
timestamp 1604489732
transform 1 0 3534 0 -1 78674
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_140_32
timestamp 1604489732
transform 1 0 2982 0 -1 78674
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_140_27
timestamp 1604489732
transform 1 0 2522 0 -1 78674
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1433
timestamp 1604489732
transform 1 0 2890 0 -1 78674
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_279
timestamp 1604489732
transform -1 0 3902 0 -1 78674
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_141_27
timestamp 1604489732
transform 1 0 2522 0 1 78674
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_281
timestamp 1604489732
transform -1 0 3902 0 1 78674
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_958
timestamp 1604489732
transform 1 0 83298 0 -1 77586
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_960
timestamp 1604489732
transform 1 0 83298 0 1 77586
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_962
timestamp 1604489732
transform 1 0 83298 0 -1 78674
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_964
timestamp 1604489732
transform 1 0 83298 0 1 78674
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_138_908
timestamp 1604489732
transform 1 0 83574 0 -1 77586
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_908
timestamp 1604489732
transform 1 0 83574 0 1 77586
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_908
timestamp 1604489732
transform 1 0 83574 0 -1 78674
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_908
timestamp 1604489732
transform 1 0 83574 0 1 78674
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_932
timestamp 1604489732
transform 1 0 85782 0 1 77586
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_920
timestamp 1604489732
transform 1 0 84678 0 1 77586
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_937
timestamp 1604489732
transform 1 0 86242 0 -1 77586
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_138_932
timestamp 1604489732
transform 1 0 85782 0 -1 77586
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_138_920
timestamp 1604489732
transform 1 0 84678 0 -1 77586
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1604
timestamp 1604489732
transform 1 0 86150 0 -1 77586
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_140_937
timestamp 1604489732
transform 1 0 86242 0 -1 78674
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_140_932
timestamp 1604489732
transform 1 0 85782 0 -1 78674
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_140_920
timestamp 1604489732
transform 1 0 84678 0 -1 78674
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1605
timestamp 1604489732
transform 1 0 86150 0 -1 78674
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_141_932
timestamp 1604489732
transform 1 0 85782 0 1 78674
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_920
timestamp 1604489732
transform 1 0 84678 0 1 78674
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_944
timestamp 1604489732
transform 1 0 86886 0 1 77586
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_950
timestamp 1604489732
transform 1 0 87438 0 1 77586
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_138_949
timestamp 1604489732
transform 1 0 87346 0 -1 77586
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_961
timestamp 1604489732
transform -1 0 87806 0 1 77586
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_959
timestamp 1604489732
transform -1 0 87806 0 -1 77586
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_140_949
timestamp 1604489732
transform 1 0 87346 0 -1 78674
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_963
timestamp 1604489732
transform -1 0 87806 0 -1 78674
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_141_944
timestamp 1604489732
transform 1 0 86886 0 1 78674
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_950
timestamp 1604489732
transform 1 0 87438 0 1 78674
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_965
timestamp 1604489732
transform -1 0 87806 0 1 78674
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_282
timestamp 1604489732
transform 1 0 38 0 -1 79762
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_284
timestamp 1604489732
transform 1 0 38 0 1 79762
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_286
timestamp 1604489732
transform 1 0 38 0 -1 80850
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_142_3
timestamp 1604489732
transform 1 0 314 0 -1 79762
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_15
timestamp 1604489732
transform 1 0 1418 0 -1 79762
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_3
timestamp 1604489732
transform 1 0 314 0 1 79762
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_15
timestamp 1604489732
transform 1 0 1418 0 1 79762
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_3
timestamp 1604489732
transform 1 0 314 0 -1 80850
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_15
timestamp 1604489732
transform 1 0 1418 0 -1 80850
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_142_27
timestamp 1604489732
transform 1 0 2522 0 -1 79762
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_142_32
timestamp 1604489732
transform 1 0 2982 0 -1 79762
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1434
timestamp 1604489732
transform 1 0 2890 0 -1 79762
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_142_38
timestamp 1604489732
transform 1 0 3534 0 -1 79762
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_283
timestamp 1604489732
transform -1 0 3902 0 -1 79762
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_143_27
timestamp 1604489732
transform 1 0 2522 0 1 79762
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_143_35
timestamp 1604489732
transform 1 0 3258 0 1 79762
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr0[1]
timestamp 1604489732
transform 1 0 3442 0 1 79762
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_285
timestamp 1604489732
transform -1 0 3902 0 1 79762
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_144_27
timestamp 1604489732
transform 1 0 2522 0 -1 80850
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_144_32
timestamp 1604489732
transform 1 0 2982 0 -1 80850
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1435
timestamp 1604489732
transform 1 0 2890 0 -1 80850
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_144_38
timestamp 1604489732
transform 1 0 3534 0 -1 80850
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_287
timestamp 1604489732
transform -1 0 3902 0 -1 80850
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_966
timestamp 1604489732
transform 1 0 83298 0 -1 79762
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_968
timestamp 1604489732
transform 1 0 83298 0 1 79762
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_970
timestamp 1604489732
transform 1 0 83298 0 -1 80850
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_142_908
timestamp 1604489732
transform 1 0 83574 0 -1 79762
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_908
timestamp 1604489732
transform 1 0 83574 0 1 79762
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_908
timestamp 1604489732
transform 1 0 83574 0 -1 80850
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_937
timestamp 1604489732
transform 1 0 86242 0 -1 79762
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_142_932
timestamp 1604489732
transform 1 0 85782 0 -1 79762
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_142_920
timestamp 1604489732
transform 1 0 84678 0 -1 79762
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1606
timestamp 1604489732
transform 1 0 86150 0 -1 79762
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_143_932
timestamp 1604489732
transform 1 0 85782 0 1 79762
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_920
timestamp 1604489732
transform 1 0 84678 0 1 79762
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_937
timestamp 1604489732
transform 1 0 86242 0 -1 80850
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_144_932
timestamp 1604489732
transform 1 0 85782 0 -1 80850
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_144_920
timestamp 1604489732
transform 1 0 84678 0 -1 80850
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1607
timestamp 1604489732
transform 1 0 86150 0 -1 80850
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_967
timestamp 1604489732
transform -1 0 87806 0 -1 79762
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_969
timestamp 1604489732
transform -1 0 87806 0 1 79762
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_971
timestamp 1604489732
transform -1 0 87806 0 -1 80850
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_142_949
timestamp 1604489732
transform 1 0 87346 0 -1 79762
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_143_944
timestamp 1604489732
transform 1 0 86886 0 1 79762
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_950
timestamp 1604489732
transform 1 0 87438 0 1 79762
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_144_949
timestamp 1604489732
transform 1 0 87346 0 -1 80850
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_288
timestamp 1604489732
transform 1 0 38 0 1 80850
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_290
timestamp 1604489732
transform 1 0 38 0 -1 81938
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_292
timestamp 1604489732
transform 1 0 38 0 1 81938
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_145_3
timestamp 1604489732
transform 1 0 314 0 1 80850
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_15
timestamp 1604489732
transform 1 0 1418 0 1 80850
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_3
timestamp 1604489732
transform 1 0 314 0 -1 81938
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_15
timestamp 1604489732
transform 1 0 1418 0 -1 81938
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_3
timestamp 1604489732
transform 1 0 314 0 1 81938
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_15
timestamp 1604489732
transform 1 0 1418 0 1 81938
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_27
timestamp 1604489732
transform 1 0 2522 0 1 80850
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_289
timestamp 1604489732
transform -1 0 3902 0 1 80850
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_146_38
timestamp 1604489732
transform 1 0 3534 0 -1 81938
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_146_32
timestamp 1604489732
transform 1 0 2982 0 -1 81938
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_146_27
timestamp 1604489732
transform 1 0 2522 0 -1 81938
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1436
timestamp 1604489732
transform 1 0 2890 0 -1 81938
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_291
timestamp 1604489732
transform -1 0 3902 0 -1 81938
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_147_35
timestamp 1604489732
transform 1 0 3258 0 1 81938
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_147_27
timestamp 1604489732
transform 1 0 2522 0 1 81938
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr0[2]
timestamp 1604489732
transform 1 0 3442 0 1 81938
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_293
timestamp 1604489732
transform -1 0 3902 0 1 81938
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_972
timestamp 1604489732
transform 1 0 83298 0 1 80850
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_974
timestamp 1604489732
transform 1 0 83298 0 -1 81938
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_976
timestamp 1604489732
transform 1 0 83298 0 1 81938
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_145_908
timestamp 1604489732
transform 1 0 83574 0 1 80850
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_908
timestamp 1604489732
transform 1 0 83574 0 -1 81938
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_908
timestamp 1604489732
transform 1 0 83574 0 1 81938
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1608
timestamp 1604489732
transform 1 0 86150 0 -1 81938
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_920
timestamp 1604489732
transform 1 0 84678 0 1 80850
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_932
timestamp 1604489732
transform 1 0 85782 0 1 80850
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_920
timestamp 1604489732
transform 1 0 84678 0 -1 81938
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_146_932
timestamp 1604489732
transform 1 0 85782 0 -1 81938
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_146_937
timestamp 1604489732
transform 1 0 86242 0 -1 81938
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_920
timestamp 1604489732
transform 1 0 84678 0 1 81938
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_932
timestamp 1604489732
transform 1 0 85782 0 1 81938
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_973
timestamp 1604489732
transform -1 0 87806 0 1 80850
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_975
timestamp 1604489732
transform -1 0 87806 0 -1 81938
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_977
timestamp 1604489732
transform -1 0 87806 0 1 81938
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_145_944
timestamp 1604489732
transform 1 0 86886 0 1 80850
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_950
timestamp 1604489732
transform 1 0 87438 0 1 80850
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_146_949
timestamp 1604489732
transform 1 0 87346 0 -1 81938
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_147_944
timestamp 1604489732
transform 1 0 86886 0 1 81938
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_950
timestamp 1604489732
transform 1 0 87438 0 1 81938
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_149_15
timestamp 1604489732
transform 1 0 1418 0 1 83026
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_3
timestamp 1604489732
transform 1 0 314 0 1 83026
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_15
timestamp 1604489732
transform 1 0 1418 0 -1 83026
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_3
timestamp 1604489732
transform 1 0 314 0 -1 83026
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_296
timestamp 1604489732
transform 1 0 38 0 1 83026
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_294
timestamp 1604489732
transform 1 0 38 0 -1 83026
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_150_15
timestamp 1604489732
transform 1 0 1418 0 -1 84114
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_3
timestamp 1604489732
transform 1 0 314 0 -1 84114
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_298
timestamp 1604489732
transform 1 0 38 0 -1 84114
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_151_15
timestamp 1604489732
transform 1 0 1418 0 1 84114
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_3
timestamp 1604489732
transform 1 0 314 0 1 84114
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_300
timestamp 1604489732
transform 1 0 38 0 1 84114
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_149_35
timestamp 1604489732
transform 1 0 3258 0 1 83026
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_149_27
timestamp 1604489732
transform 1 0 2522 0 1 83026
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_148_38
timestamp 1604489732
transform 1 0 3534 0 -1 83026
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_148_32
timestamp 1604489732
transform 1 0 2982 0 -1 83026
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_148_27
timestamp 1604489732
transform 1 0 2522 0 -1 83026
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr0[3]
timestamp 1604489732
transform 1 0 3442 0 1 83026
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1437
timestamp 1604489732
transform 1 0 2890 0 -1 83026
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_297
timestamp 1604489732
transform -1 0 3902 0 1 83026
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_295
timestamp 1604489732
transform -1 0 3902 0 -1 83026
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_150_38
timestamp 1604489732
transform 1 0 3534 0 -1 84114
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_150_32
timestamp 1604489732
transform 1 0 2982 0 -1 84114
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_150_27
timestamp 1604489732
transform 1 0 2522 0 -1 84114
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1438
timestamp 1604489732
transform 1 0 2890 0 -1 84114
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_299
timestamp 1604489732
transform -1 0 3902 0 -1 84114
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_151_27
timestamp 1604489732
transform 1 0 2522 0 1 84114
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_301
timestamp 1604489732
transform -1 0 3902 0 1 84114
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_978
timestamp 1604489732
transform 1 0 83298 0 -1 83026
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_980
timestamp 1604489732
transform 1 0 83298 0 1 83026
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_982
timestamp 1604489732
transform 1 0 83298 0 -1 84114
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_984
timestamp 1604489732
transform 1 0 83298 0 1 84114
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_148_908
timestamp 1604489732
transform 1 0 83574 0 -1 83026
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_908
timestamp 1604489732
transform 1 0 83574 0 1 83026
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_908
timestamp 1604489732
transform 1 0 83574 0 -1 84114
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_908
timestamp 1604489732
transform 1 0 83574 0 1 84114
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_932
timestamp 1604489732
transform 1 0 85782 0 1 83026
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_920
timestamp 1604489732
transform 1 0 84678 0 1 83026
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_937
timestamp 1604489732
transform 1 0 86242 0 -1 83026
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_148_932
timestamp 1604489732
transform 1 0 85782 0 -1 83026
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_148_920
timestamp 1604489732
transform 1 0 84678 0 -1 83026
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1609
timestamp 1604489732
transform 1 0 86150 0 -1 83026
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_150_937
timestamp 1604489732
transform 1 0 86242 0 -1 84114
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_150_932
timestamp 1604489732
transform 1 0 85782 0 -1 84114
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_150_920
timestamp 1604489732
transform 1 0 84678 0 -1 84114
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1610
timestamp 1604489732
transform 1 0 86150 0 -1 84114
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_932
timestamp 1604489732
transform 1 0 85782 0 1 84114
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_920
timestamp 1604489732
transform 1 0 84678 0 1 84114
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_944
timestamp 1604489732
transform 1 0 86886 0 1 83026
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_950
timestamp 1604489732
transform 1 0 87438 0 1 83026
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_148_949
timestamp 1604489732
transform 1 0 87346 0 -1 83026
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_981
timestamp 1604489732
transform -1 0 87806 0 1 83026
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_979
timestamp 1604489732
transform -1 0 87806 0 -1 83026
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_150_949
timestamp 1604489732
transform 1 0 87346 0 -1 84114
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_983
timestamp 1604489732
transform -1 0 87806 0 -1 84114
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_151_944
timestamp 1604489732
transform 1 0 86886 0 1 84114
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_950
timestamp 1604489732
transform 1 0 87438 0 1 84114
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_985
timestamp 1604489732
transform -1 0 87806 0 1 84114
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_302
timestamp 1604489732
transform 1 0 38 0 -1 85202
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_304
timestamp 1604489732
transform 1 0 38 0 1 85202
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_306
timestamp 1604489732
transform 1 0 38 0 -1 86290
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_152_3
timestamp 1604489732
transform 1 0 314 0 -1 85202
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_15
timestamp 1604489732
transform 1 0 1418 0 -1 85202
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_3
timestamp 1604489732
transform 1 0 314 0 1 85202
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_15
timestamp 1604489732
transform 1 0 1418 0 1 85202
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_3
timestamp 1604489732
transform 1 0 314 0 -1 86290
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_15
timestamp 1604489732
transform 1 0 1418 0 -1 86290
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_152_36
timestamp 1604489732
transform 1 0 3350 0 -1 85202
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_152_32
timestamp 1604489732
transform 1 0 2982 0 -1 85202
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_152_27
timestamp 1604489732
transform 1 0 2522 0 -1 85202
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr0[4]
timestamp 1604489732
transform 1 0 3442 0 -1 85202
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1439
timestamp 1604489732
transform 1 0 2890 0 -1 85202
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_303
timestamp 1604489732
transform -1 0 3902 0 -1 85202
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_153_27
timestamp 1604489732
transform 1 0 2522 0 1 85202
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_305
timestamp 1604489732
transform -1 0 3902 0 1 85202
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_154_36
timestamp 1604489732
transform 1 0 3350 0 -1 86290
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_154_32
timestamp 1604489732
transform 1 0 2982 0 -1 86290
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_154_27
timestamp 1604489732
transform 1 0 2522 0 -1 86290
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr0[5]
timestamp 1604489732
transform 1 0 3442 0 -1 86290
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1440
timestamp 1604489732
transform 1 0 2890 0 -1 86290
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_307
timestamp 1604489732
transform -1 0 3902 0 -1 86290
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_986
timestamp 1604489732
transform 1 0 83298 0 -1 85202
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_988
timestamp 1604489732
transform 1 0 83298 0 1 85202
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_990
timestamp 1604489732
transform 1 0 83298 0 -1 86290
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_152_908
timestamp 1604489732
transform 1 0 83574 0 -1 85202
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_908
timestamp 1604489732
transform 1 0 83574 0 1 85202
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_908
timestamp 1604489732
transform 1 0 83574 0 -1 86290
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_937
timestamp 1604489732
transform 1 0 86242 0 -1 85202
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_152_932
timestamp 1604489732
transform 1 0 85782 0 -1 85202
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_152_920
timestamp 1604489732
transform 1 0 84678 0 -1 85202
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1611
timestamp 1604489732
transform 1 0 86150 0 -1 85202
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_153_932
timestamp 1604489732
transform 1 0 85782 0 1 85202
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_920
timestamp 1604489732
transform 1 0 84678 0 1 85202
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_937
timestamp 1604489732
transform 1 0 86242 0 -1 86290
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_154_932
timestamp 1604489732
transform 1 0 85782 0 -1 86290
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_154_920
timestamp 1604489732
transform 1 0 84678 0 -1 86290
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1612
timestamp 1604489732
transform 1 0 86150 0 -1 86290
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_987
timestamp 1604489732
transform -1 0 87806 0 -1 85202
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_989
timestamp 1604489732
transform -1 0 87806 0 1 85202
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_991
timestamp 1604489732
transform -1 0 87806 0 -1 86290
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_152_949
timestamp 1604489732
transform 1 0 87346 0 -1 85202
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_153_944
timestamp 1604489732
transform 1 0 86886 0 1 85202
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_950
timestamp 1604489732
transform 1 0 87438 0 1 85202
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_154_949
timestamp 1604489732
transform 1 0 87346 0 -1 86290
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_155_15
timestamp 1604489732
transform 1 0 1418 0 1 86290
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_3
timestamp 1604489732
transform 1 0 314 0 1 86290
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_308
timestamp 1604489732
transform 1 0 38 0 1 86290
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_157_15
timestamp 1604489732
transform 1 0 1418 0 1 87378
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_3
timestamp 1604489732
transform 1 0 314 0 1 87378
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_15
timestamp 1604489732
transform 1 0 1418 0 -1 87378
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_3
timestamp 1604489732
transform 1 0 314 0 -1 87378
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_312
timestamp 1604489732
transform 1 0 38 0 1 87378
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_310
timestamp 1604489732
transform 1 0 38 0 -1 87378
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_158_15
timestamp 1604489732
transform 1 0 1418 0 -1 88466
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_3
timestamp 1604489732
transform 1 0 314 0 -1 88466
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_314
timestamp 1604489732
transform 1 0 38 0 -1 88466
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_155_27
timestamp 1604489732
transform 1 0 2522 0 1 86290
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_309
timestamp 1604489732
transform -1 0 3902 0 1 86290
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_157_35
timestamp 1604489732
transform 1 0 3258 0 1 87378
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_157_27
timestamp 1604489732
transform 1 0 2522 0 1 87378
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_156_38
timestamp 1604489732
transform 1 0 3534 0 -1 87378
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_156_32
timestamp 1604489732
transform 1 0 2982 0 -1 87378
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_156_27
timestamp 1604489732
transform 1 0 2522 0 -1 87378
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr0[6]
timestamp 1604489732
transform 1 0 3442 0 1 87378
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1441
timestamp 1604489732
transform 1 0 2890 0 -1 87378
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_313
timestamp 1604489732
transform -1 0 3902 0 1 87378
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_311
timestamp 1604489732
transform -1 0 3902 0 -1 87378
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_158_38
timestamp 1604489732
transform 1 0 3534 0 -1 88466
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_158_32
timestamp 1604489732
transform 1 0 2982 0 -1 88466
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_158_27
timestamp 1604489732
transform 1 0 2522 0 -1 88466
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1442
timestamp 1604489732
transform 1 0 2890 0 -1 88466
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_315
timestamp 1604489732
transform -1 0 3902 0 -1 88466
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_992
timestamp 1604489732
transform 1 0 83298 0 1 86290
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_994
timestamp 1604489732
transform 1 0 83298 0 -1 87378
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_996
timestamp 1604489732
transform 1 0 83298 0 1 87378
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_998
timestamp 1604489732
transform 1 0 83298 0 -1 88466
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_155_908
timestamp 1604489732
transform 1 0 83574 0 1 86290
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_908
timestamp 1604489732
transform 1 0 83574 0 -1 87378
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_908
timestamp 1604489732
transform 1 0 83574 0 1 87378
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_908
timestamp 1604489732
transform 1 0 83574 0 -1 88466
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_932
timestamp 1604489732
transform 1 0 85782 0 1 86290
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_920
timestamp 1604489732
transform 1 0 84678 0 1 86290
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_932
timestamp 1604489732
transform 1 0 85782 0 1 87378
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_920
timestamp 1604489732
transform 1 0 84678 0 1 87378
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_937
timestamp 1604489732
transform 1 0 86242 0 -1 87378
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_156_932
timestamp 1604489732
transform 1 0 85782 0 -1 87378
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_156_920
timestamp 1604489732
transform 1 0 84678 0 -1 87378
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1613
timestamp 1604489732
transform 1 0 86150 0 -1 87378
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_937
timestamp 1604489732
transform 1 0 86242 0 -1 88466
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_158_932
timestamp 1604489732
transform 1 0 85782 0 -1 88466
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_158_920
timestamp 1604489732
transform 1 0 84678 0 -1 88466
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1614
timestamp 1604489732
transform 1 0 86150 0 -1 88466
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_155_944
timestamp 1604489732
transform 1 0 86886 0 1 86290
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_950
timestamp 1604489732
transform 1 0 87438 0 1 86290
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_993
timestamp 1604489732
transform -1 0 87806 0 1 86290
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_157_944
timestamp 1604489732
transform 1 0 86886 0 1 87378
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_950
timestamp 1604489732
transform 1 0 87438 0 1 87378
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_156_949
timestamp 1604489732
transform 1 0 87346 0 -1 87378
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_997
timestamp 1604489732
transform -1 0 87806 0 1 87378
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_995
timestamp 1604489732
transform -1 0 87806 0 -1 87378
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_158_949
timestamp 1604489732
transform 1 0 87346 0 -1 88466
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_999
timestamp 1604489732
transform -1 0 87806 0 -1 88466
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_316
timestamp 1604489732
transform 1 0 38 0 1 88466
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_318
timestamp 1604489732
transform 1 0 38 0 -1 89554
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_320
timestamp 1604489732
transform 1 0 38 0 1 89554
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_159_3
timestamp 1604489732
transform 1 0 314 0 1 88466
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_15
timestamp 1604489732
transform 1 0 1418 0 1 88466
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_3
timestamp 1604489732
transform 1 0 314 0 -1 89554
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_15
timestamp 1604489732
transform 1 0 1418 0 -1 89554
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_3
timestamp 1604489732
transform 1 0 314 0 1 89554
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_15
timestamp 1604489732
transform 1 0 1418 0 1 89554
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_159_35
timestamp 1604489732
transform 1 0 3258 0 1 88466
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_159_27
timestamp 1604489732
transform 1 0 2522 0 1 88466
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr0[7]
timestamp 1604489732
transform 1 0 3442 0 1 88466
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_317
timestamp 1604489732
transform -1 0 3902 0 1 88466
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_160_38
timestamp 1604489732
transform 1 0 3534 0 -1 89554
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_160_32
timestamp 1604489732
transform 1 0 2982 0 -1 89554
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_160_27
timestamp 1604489732
transform 1 0 2522 0 -1 89554
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1443
timestamp 1604489732
transform 1 0 2890 0 -1 89554
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_319
timestamp 1604489732
transform -1 0 3902 0 -1 89554
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_161_27
timestamp 1604489732
transform 1 0 2522 0 1 89554
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_321
timestamp 1604489732
transform -1 0 3902 0 1 89554
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1000
timestamp 1604489732
transform 1 0 83298 0 1 88466
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1002
timestamp 1604489732
transform 1 0 83298 0 -1 89554
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1004
timestamp 1604489732
transform 1 0 83298 0 1 89554
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_159_908
timestamp 1604489732
transform 1 0 83574 0 1 88466
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_908
timestamp 1604489732
transform 1 0 83574 0 -1 89554
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_908
timestamp 1604489732
transform 1 0 83574 0 1 89554
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1615
timestamp 1604489732
transform 1 0 86150 0 -1 89554
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_159_920
timestamp 1604489732
transform 1 0 84678 0 1 88466
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_932
timestamp 1604489732
transform 1 0 85782 0 1 88466
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_920
timestamp 1604489732
transform 1 0 84678 0 -1 89554
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_160_932
timestamp 1604489732
transform 1 0 85782 0 -1 89554
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_160_937
timestamp 1604489732
transform 1 0 86242 0 -1 89554
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_920
timestamp 1604489732
transform 1 0 84678 0 1 89554
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_932
timestamp 1604489732
transform 1 0 85782 0 1 89554
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1001
timestamp 1604489732
transform -1 0 87806 0 1 88466
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1003
timestamp 1604489732
transform -1 0 87806 0 -1 89554
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1005
timestamp 1604489732
transform -1 0 87806 0 1 89554
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_159_944
timestamp 1604489732
transform 1 0 86886 0 1 88466
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_950
timestamp 1604489732
transform 1 0 87438 0 1 88466
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_160_949
timestamp 1604489732
transform 1 0 87346 0 -1 89554
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_161_944
timestamp 1604489732
transform 1 0 86886 0 1 89554
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_950
timestamp 1604489732
transform 1 0 87438 0 1 89554
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_322
timestamp 1604489732
transform 1 0 38 0 -1 90642
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_324
timestamp 1604489732
transform 1 0 38 0 1 90642
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_326
timestamp 1604489732
transform 1 0 38 0 -1 91730
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_162_3
timestamp 1604489732
transform 1 0 314 0 -1 90642
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_15
timestamp 1604489732
transform 1 0 1418 0 -1 90642
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_3
timestamp 1604489732
transform 1 0 314 0 1 90642
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_15
timestamp 1604489732
transform 1 0 1418 0 1 90642
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_3
timestamp 1604489732
transform 1 0 314 0 -1 91730
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_15
timestamp 1604489732
transform 1 0 1418 0 -1 91730
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_162_38
timestamp 1604489732
transform 1 0 3534 0 -1 90642
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_162_32
timestamp 1604489732
transform 1 0 2982 0 -1 90642
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_162_27
timestamp 1604489732
transform 1 0 2522 0 -1 90642
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1444
timestamp 1604489732
transform 1 0 2890 0 -1 90642
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_323
timestamp 1604489732
transform -1 0 3902 0 -1 90642
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_163_27
timestamp 1604489732
transform 1 0 2522 0 1 90642
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_325
timestamp 1604489732
transform -1 0 3902 0 1 90642
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_164_38
timestamp 1604489732
transform 1 0 3534 0 -1 91730
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_164_32
timestamp 1604489732
transform 1 0 2982 0 -1 91730
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_164_27
timestamp 1604489732
transform 1 0 2522 0 -1 91730
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1445
timestamp 1604489732
transform 1 0 2890 0 -1 91730
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_327
timestamp 1604489732
transform -1 0 3902 0 -1 91730
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1006
timestamp 1604489732
transform 1 0 83298 0 -1 90642
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1008
timestamp 1604489732
transform 1 0 83298 0 1 90642
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1010
timestamp 1604489732
transform 1 0 83298 0 -1 91730
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_162_908
timestamp 1604489732
transform 1 0 83574 0 -1 90642
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_908
timestamp 1604489732
transform 1 0 83574 0 1 90642
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_908
timestamp 1604489732
transform 1 0 83574 0 -1 91730
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_937
timestamp 1604489732
transform 1 0 86242 0 -1 90642
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_162_932
timestamp 1604489732
transform 1 0 85782 0 -1 90642
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_162_920
timestamp 1604489732
transform 1 0 84678 0 -1 90642
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1616
timestamp 1604489732
transform 1 0 86150 0 -1 90642
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_163_932
timestamp 1604489732
transform 1 0 85782 0 1 90642
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_920
timestamp 1604489732
transform 1 0 84678 0 1 90642
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_937
timestamp 1604489732
transform 1 0 86242 0 -1 91730
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_164_932
timestamp 1604489732
transform 1 0 85782 0 -1 91730
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_164_920
timestamp 1604489732
transform 1 0 84678 0 -1 91730
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1617
timestamp 1604489732
transform 1 0 86150 0 -1 91730
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1007
timestamp 1604489732
transform -1 0 87806 0 -1 90642
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1009
timestamp 1604489732
transform -1 0 87806 0 1 90642
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1011
timestamp 1604489732
transform -1 0 87806 0 -1 91730
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_162_949
timestamp 1604489732
transform 1 0 87346 0 -1 90642
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_163_944
timestamp 1604489732
transform 1 0 86886 0 1 90642
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_950
timestamp 1604489732
transform 1 0 87438 0 1 90642
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_164_949
timestamp 1604489732
transform 1 0 87346 0 -1 91730
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_328
timestamp 1604489732
transform 1 0 38 0 1 91730
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_330
timestamp 1604489732
transform 1 0 38 0 -1 92818
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_332
timestamp 1604489732
transform 1 0 38 0 1 92818
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_165_3
timestamp 1604489732
transform 1 0 314 0 1 91730
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_15
timestamp 1604489732
transform 1 0 1418 0 1 91730
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_3
timestamp 1604489732
transform 1 0 314 0 -1 92818
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_15
timestamp 1604489732
transform 1 0 1418 0 -1 92818
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_3
timestamp 1604489732
transform 1 0 314 0 1 92818
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_15
timestamp 1604489732
transform 1 0 1418 0 1 92818
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_329
timestamp 1604489732
transform -1 0 3902 0 1 91730
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_331
timestamp 1604489732
transform -1 0 3902 0 -1 92818
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_333
timestamp 1604489732
transform -1 0 3902 0 1 92818
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1446
timestamp 1604489732
transform 1 0 2890 0 -1 92818
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_27
timestamp 1604489732
transform 1 0 2522 0 1 91730
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_166_27
timestamp 1604489732
transform 1 0 2522 0 -1 92818
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_166_32
timestamp 1604489732
transform 1 0 2982 0 -1 92818
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_38
timestamp 1604489732
transform 1 0 3534 0 -1 92818
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_167_27
timestamp 1604489732
transform 1 0 2522 0 1 92818
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_908
timestamp 1604489732
transform 1 0 83574 0 -1 92818
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_912
timestamp 1604489732
transform 1 0 83942 0 1 91730
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_165_908
timestamp 1604489732
transform 1 0 83574 0 1 91730
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_csb1
timestamp 1604489732
transform 1 0 83758 0 1 91730
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1014
timestamp 1604489732
transform 1 0 83298 0 -1 92818
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1012
timestamp 1604489732
transform 1 0 83298 0 1 91730
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_167_912
timestamp 1604489732
transform 1 0 83942 0 1 92818
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_167_908
timestamp 1604489732
transform 1 0 83574 0 1 92818
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr1[0]
timestamp 1604489732
transform 1 0 83758 0 1 92818
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1016
timestamp 1604489732
transform 1 0 83298 0 1 92818
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1618
timestamp 1604489732
transform 1 0 86150 0 -1 92818
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_924
timestamp 1604489732
transform 1 0 85046 0 1 91730
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_936
timestamp 1604489732
transform 1 0 86150 0 1 91730
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_920
timestamp 1604489732
transform 1 0 84678 0 -1 92818
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_166_932
timestamp 1604489732
transform 1 0 85782 0 -1 92818
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_166_937
timestamp 1604489732
transform 1 0 86242 0 -1 92818
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_924
timestamp 1604489732
transform 1 0 85046 0 1 92818
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_936
timestamp 1604489732
transform 1 0 86150 0 1 92818
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1013
timestamp 1604489732
transform -1 0 87806 0 1 91730
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1015
timestamp 1604489732
transform -1 0 87806 0 -1 92818
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1017
timestamp 1604489732
transform -1 0 87806 0 1 92818
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_165_948
timestamp 1604489732
transform 1 0 87254 0 1 91730
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_166_949
timestamp 1604489732
transform 1 0 87346 0 -1 92818
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_167_948
timestamp 1604489732
transform 1 0 87254 0 1 92818
box -38 -48 314 592
use sram_1rw1r_32_256_8_sky130  SRAM_0
timestamp 1605062100
transform 1 0 4934 0 1 2155
box 0 0 77296 91247
use sky130_fd_sc_hd__decap_12  FILLER_168_15
timestamp 1604489732
transform 1 0 1418 0 -1 93906
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_3
timestamp 1604489732
transform 1 0 314 0 -1 93906
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_334
timestamp 1604489732
transform 1 0 38 0 -1 93906
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_170_15
timestamp 1604489732
transform 1 0 1418 0 -1 94994
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_3
timestamp 1604489732
transform 1 0 314 0 -1 94994
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_15
timestamp 1604489732
transform 1 0 1418 0 1 93906
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_3
timestamp 1604489732
transform 1 0 314 0 1 93906
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_338
timestamp 1604489732
transform 1 0 38 0 -1 94994
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_336
timestamp 1604489732
transform 1 0 38 0 1 93906
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_171_15
timestamp 1604489732
transform 1 0 1418 0 1 94994
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_3
timestamp 1604489732
transform 1 0 314 0 1 94994
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_340
timestamp 1604489732
transform 1 0 38 0 1 94994
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_168_38
timestamp 1604489732
transform 1 0 3534 0 -1 93906
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_168_32
timestamp 1604489732
transform 1 0 2982 0 -1 93906
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_168_27
timestamp 1604489732
transform 1 0 2522 0 -1 93906
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1447
timestamp 1604489732
transform 1 0 2890 0 -1 93906
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_335
timestamp 1604489732
transform -1 0 3902 0 -1 93906
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_170_38
timestamp 1604489732
transform 1 0 3534 0 -1 94994
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_170_32
timestamp 1604489732
transform 1 0 2982 0 -1 94994
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_170_27
timestamp 1604489732
transform 1 0 2522 0 -1 94994
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_169_27
timestamp 1604489732
transform 1 0 2522 0 1 93906
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1448
timestamp 1604489732
transform 1 0 2890 0 -1 94994
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_339
timestamp 1604489732
transform -1 0 3902 0 -1 94994
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_337
timestamp 1604489732
transform -1 0 3902 0 1 93906
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_171_35
timestamp 1604489732
transform 1 0 3258 0 1 94994
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_171_27
timestamp 1604489732
transform 1 0 2522 0 1 94994
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_wmask0[0]
timestamp 1604489732
transform 1 0 3074 0 1 94994
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[2]
timestamp 1604489732
transform 1 0 3442 0 1 94994
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_341
timestamp 1604489732
transform -1 0 3902 0 1 94994
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_168_912
timestamp 1604489732
transform 1 0 83942 0 -1 93906
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_168_908
timestamp 1604489732
transform 1 0 83574 0 -1 93906
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_clk1
timestamp 1604489732
transform 1 0 83758 0 -1 93906
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1018
timestamp 1604489732
transform 1 0 83298 0 -1 93906
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_170_908
timestamp 1604489732
transform 1 0 83574 0 -1 94994
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_908
timestamp 1604489732
transform 1 0 83574 0 1 93906
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1022
timestamp 1604489732
transform 1 0 83298 0 -1 94994
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1020
timestamp 1604489732
transform 1 0 83298 0 1 93906
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_171_908
timestamp 1604489732
transform 1 0 83574 0 1 94994
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1024
timestamp 1604489732
transform 1 0 83298 0 1 94994
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_168_937
timestamp 1604489732
transform 1 0 86242 0 -1 93906
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_924
timestamp 1604489732
transform 1 0 85046 0 -1 93906
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1619
timestamp 1604489732
transform 1 0 86150 0 -1 93906
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_170_937
timestamp 1604489732
transform 1 0 86242 0 -1 94994
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_170_932
timestamp 1604489732
transform 1 0 85782 0 -1 94994
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_170_920
timestamp 1604489732
transform 1 0 84678 0 -1 94994
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_932
timestamp 1604489732
transform 1 0 85782 0 1 93906
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_920
timestamp 1604489732
transform 1 0 84678 0 1 93906
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1620
timestamp 1604489732
transform 1 0 86150 0 -1 94994
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_932
timestamp 1604489732
transform 1 0 85782 0 1 94994
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_920
timestamp 1604489732
transform 1 0 84678 0 1 94994
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_168_949
timestamp 1604489732
transform 1 0 87346 0 -1 93906
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1019
timestamp 1604489732
transform -1 0 87806 0 -1 93906
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_169_944
timestamp 1604489732
transform 1 0 86886 0 1 93906
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_170_949
timestamp 1604489732
transform 1 0 87346 0 -1 94994
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_169_950
timestamp 1604489732
transform 1 0 87438 0 1 93906
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1023
timestamp 1604489732
transform -1 0 87806 0 -1 94994
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1021
timestamp 1604489732
transform -1 0 87806 0 1 93906
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_171_944
timestamp 1604489732
transform 1 0 86886 0 1 94994
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_950
timestamp 1604489732
transform 1 0 87438 0 1 94994
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1025
timestamp 1604489732
transform -1 0 87806 0 1 94994
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_172_15
timestamp 1604489732
transform 1 0 1418 0 -1 96082
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_172_3
timestamp 1604489732
transform 1 0 314 0 -1 96082
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_342
timestamp 1604489732
transform 1 0 38 0 -1 96082
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_173_15
timestamp 1604489732
transform 1 0 1418 0 1 96082
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_173_3
timestamp 1604489732
transform 1 0 314 0 1 96082
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_344
timestamp 1604489732
transform 1 0 38 0 1 96082
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_174_19
timestamp 1604489732
transform 1 0 1786 0 -1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_174_15
timestamp 1604489732
transform 1 0 1418 0 -1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_174_11
timestamp 1604489732
transform 1 0 1050 0 -1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_174_3
timestamp 1604489732
transform 1 0 314 0 -1 97170
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_wmask0[3]
timestamp 1604489732
transform 1 0 866 0 -1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[7]
timestamp 1604489732
transform 1 0 1234 0 -1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[20]
timestamp 1604489732
transform 1 0 1602 0 -1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_346
timestamp 1604489732
transform 1 0 38 0 -1 97170
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_172_23
timestamp 1604489732
transform 1 0 2154 0 -1 96082
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_172_27
timestamp 1604489732
transform 1 0 2522 0 -1 96082
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_wmask0[1]
timestamp 1604489732
transform 1 0 2338 0 -1 96082
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[5]
timestamp 1604489732
transform 1 0 2706 0 -1 96082
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_172_32
timestamp 1604489732
transform 1 0 2982 0 -1 96082
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1449
timestamp 1604489732
transform 1 0 2890 0 -1 96082
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_172_36
timestamp 1604489732
transform 1 0 3350 0 -1 96082
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[16]
timestamp 1604489732
transform 1 0 3442 0 -1 96082
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_343
timestamp 1604489732
transform -1 0 3902 0 -1 96082
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_173_23
timestamp 1604489732
transform 1 0 2154 0 1 96082
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[6]
timestamp 1604489732
transform 1 0 1970 0 1 96082
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_173_27
timestamp 1604489732
transform 1 0 2522 0 1 96082
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[1]
timestamp 1604489732
transform 1 0 2338 0 1 96082
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[18]
timestamp 1604489732
transform 1 0 2706 0 1 96082
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_173_31
timestamp 1604489732
transform 1 0 2890 0 1 96082
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[12]
timestamp 1604489732
transform 1 0 3074 0 1 96082
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_173_35
timestamp 1604489732
transform 1 0 3258 0 1 96082
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[0]
timestamp 1604489732
transform 1 0 3442 0 1 96082
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_345
timestamp 1604489732
transform -1 0 3902 0 1 96082
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_174_23
timestamp 1604489732
transform 1 0 2154 0 -1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[15]
timestamp 1604489732
transform 1 0 1970 0 -1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_174_27
timestamp 1604489732
transform 1 0 2522 0 -1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[14]
timestamp 1604489732
transform 1 0 2338 0 -1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[10]
timestamp 1604489732
transform 1 0 2706 0 -1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_174_32
timestamp 1604489732
transform 1 0 2982 0 -1 97170
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1450
timestamp 1604489732
transform 1 0 2890 0 -1 97170
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_174_36
timestamp 1604489732
transform 1 0 3350 0 -1 97170
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_addr0[0]
timestamp 1604489732
transform 1 0 3442 0 -1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_347
timestamp 1604489732
transform -1 0 3902 0 -1 97170
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_172_912
timestamp 1604489732
transform 1 0 83942 0 -1 96082
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_172_908
timestamp 1604489732
transform 1 0 83574 0 -1 96082
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[31]
timestamp 1604489732
transform 1 0 83758 0 -1 96082
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1026
timestamp 1604489732
transform 1 0 83298 0 -1 96082
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_173_916
timestamp 1604489732
transform 1 0 84310 0 1 96082
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_173_912
timestamp 1604489732
transform 1 0 83942 0 1 96082
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_173_908
timestamp 1604489732
transform 1 0 83574 0 1 96082
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[29]
timestamp 1604489732
transform 1 0 84126 0 1 96082
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[25]
timestamp 1604489732
transform 1 0 83758 0 1 96082
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1028
timestamp 1604489732
transform 1 0 83298 0 1 96082
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_174_916
timestamp 1604489732
transform 1 0 84310 0 -1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_174_912
timestamp 1604489732
transform 1 0 83942 0 -1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_174_908
timestamp 1604489732
transform 1 0 83574 0 -1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[26]
timestamp 1604489732
transform 1 0 84494 0 -1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[23]
timestamp 1604489732
transform 1 0 84126 0 -1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[22]
timestamp 1604489732
transform 1 0 83758 0 -1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1030
timestamp 1604489732
transform 1 0 83298 0 -1 97170
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1621
timestamp 1604489732
transform 1 0 86150 0 -1 96082
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1622
timestamp 1604489732
transform 1 0 86150 0 -1 97170
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[27]
timestamp 1604489732
transform 1 0 84862 0 -1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_172_924
timestamp 1604489732
transform 1 0 85046 0 -1 96082
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_937
timestamp 1604489732
transform 1 0 86242 0 -1 96082
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_928
timestamp 1604489732
transform 1 0 85414 0 1 96082
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_174_920
timestamp 1604489732
transform 1 0 84678 0 -1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_174_924
timestamp 1604489732
transform 1 0 85046 0 -1 97170
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_937
timestamp 1604489732
transform 1 0 86242 0 -1 97170
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1027
timestamp 1604489732
transform -1 0 87806 0 -1 96082
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1029
timestamp 1604489732
transform -1 0 87806 0 1 96082
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1031
timestamp 1604489732
transform -1 0 87806 0 -1 97170
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_172_949
timestamp 1604489732
transform 1 0 87346 0 -1 96082
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_173_940
timestamp 1604489732
transform 1 0 86518 0 1 96082
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_173_948
timestamp 1604489732
transform 1 0 87254 0 1 96082
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_174_949
timestamp 1604489732
transform 1 0 87346 0 -1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_175_19
timestamp 1604489732
transform 1 0 1786 0 1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_175_15
timestamp 1604489732
transform 1 0 1418 0 1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_175_3
timestamp 1604489732
transform 1 0 314 0 1 97170
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_wmask0[2]
timestamp 1604489732
transform 1 0 1602 0 1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_348
timestamp 1604489732
transform 1 0 38 0 1 97170
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_176_15
timestamp 1604489732
transform 1 0 1418 0 -1 98258
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_176_3
timestamp 1604489732
transform 1 0 314 0 -1 98258
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_350
timestamp 1604489732
transform 1 0 38 0 -1 98258
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_177_15
timestamp 1604489732
transform 1 0 1418 0 1 98258
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_3
timestamp 1604489732
transform 1 0 314 0 1 98258
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_352
timestamp 1604489732
transform 1 0 38 0 1 98258
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_175_23
timestamp 1604489732
transform 1 0 2154 0 1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[4]
timestamp 1604489732
transform 1 0 1970 0 1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[19]
timestamp 1604489732
transform 1 0 2338 0 1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_175_31
timestamp 1604489732
transform 1 0 2890 0 1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_175_27
timestamp 1604489732
transform 1 0 2522 0 1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[17]
timestamp 1604489732
transform 1 0 2706 0 1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[11]
timestamp 1604489732
transform 1 0 3074 0 1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_175_35
timestamp 1604489732
transform 1 0 3258 0 1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_clk0
timestamp 1604489732
transform 1 0 3442 0 1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_349
timestamp 1604489732
transform -1 0 3902 0 1 97170
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_176_23
timestamp 1604489732
transform 1 0 2154 0 -1 98258
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[9]
timestamp 1604489732
transform 1 0 2338 0 -1 98258
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_176_32
timestamp 1604489732
transform 1 0 2982 0 -1 98258
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_176_27
timestamp 1604489732
transform 1 0 2522 0 -1 98258
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[3]
timestamp 1604489732
transform 1 0 2706 0 -1 98258
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1451
timestamp 1604489732
transform 1 0 2890 0 -1 98258
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_176_36
timestamp 1604489732
transform 1 0 3350 0 -1 98258
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[13]
timestamp 1604489732
transform 1 0 3442 0 -1 98258
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_351
timestamp 1604489732
transform -1 0 3902 0 -1 98258
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_177_27
timestamp 1604489732
transform 1 0 2522 0 1 98258
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[8]
timestamp 1604489732
transform 1 0 3074 0 1 98258
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_177_35
timestamp 1604489732
transform 1 0 3258 0 1 98258
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[21]
timestamp 1604489732
transform 1 0 3442 0 1 98258
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_353
timestamp 1604489732
transform -1 0 3902 0 1 98258
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_175_916
timestamp 1604489732
transform 1 0 84310 0 1 97170
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_175_912
timestamp 1604489732
transform 1 0 83942 0 1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_175_908
timestamp 1604489732
transform 1 0 83574 0 1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[28]
timestamp 1604489732
transform 1 0 84126 0 1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[24]
timestamp 1604489732
transform 1 0 83758 0 1 97170
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1032
timestamp 1604489732
transform 1 0 83298 0 1 97170
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_176_912
timestamp 1604489732
transform 1 0 83942 0 -1 98258
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_176_908
timestamp 1604489732
transform 1 0 83574 0 -1 98258
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[30]
timestamp 1604489732
transform 1 0 83758 0 -1 98258
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1034
timestamp 1604489732
transform 1 0 83298 0 -1 98258
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_177_908
timestamp 1604489732
transform 1 0 83574 0 1 98258
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1036
timestamp 1604489732
transform 1 0 83298 0 1 98258
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1623
timestamp 1604489732
transform 1 0 86150 0 -1 98258
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_175_928
timestamp 1604489732
transform 1 0 85414 0 1 97170
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_924
timestamp 1604489732
transform 1 0 85046 0 -1 98258
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_937
timestamp 1604489732
transform 1 0 86242 0 -1 98258
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_920
timestamp 1604489732
transform 1 0 84678 0 1 98258
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_932
timestamp 1604489732
transform 1 0 85782 0 1 98258
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1033
timestamp 1604489732
transform -1 0 87806 0 1 97170
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1035
timestamp 1604489732
transform -1 0 87806 0 -1 98258
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1037
timestamp 1604489732
transform -1 0 87806 0 1 98258
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_175_940
timestamp 1604489732
transform 1 0 86518 0 1 97170
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_175_948
timestamp 1604489732
transform 1 0 87254 0 1 97170
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_176_949
timestamp 1604489732
transform 1 0 87346 0 -1 98258
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_177_944
timestamp 1604489732
transform 1 0 86886 0 1 98258
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_950
timestamp 1604489732
transform 1 0 87438 0 1 98258
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_354
timestamp 1604489732
transform 1 0 38 0 -1 99346
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_356
timestamp 1604489732
transform 1 0 38 0 1 99346
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_358
timestamp 1604489732
transform 1 0 38 0 -1 100434
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_178_3
timestamp 1604489732
transform 1 0 314 0 -1 99346
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_15
timestamp 1604489732
transform 1 0 1418 0 -1 99346
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_3
timestamp 1604489732
transform 1 0 314 0 1 99346
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_15
timestamp 1604489732
transform 1 0 1418 0 1 99346
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_3
timestamp 1604489732
transform 1 0 314 0 -1 100434
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_15
timestamp 1604489732
transform 1 0 1418 0 -1 100434
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_178_38
timestamp 1604489732
transform 1 0 3534 0 -1 99346
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_178_32
timestamp 1604489732
transform 1 0 2982 0 -1 99346
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_178_27
timestamp 1604489732
transform 1 0 2522 0 -1 99346
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1452
timestamp 1604489732
transform 1 0 2890 0 -1 99346
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_355
timestamp 1604489732
transform -1 0 3902 0 -1 99346
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_180_38
timestamp 1604489732
transform 1 0 3534 0 -1 100434
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_180_32
timestamp 1604489732
transform 1 0 2982 0 -1 100434
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_180_27
timestamp 1604489732
transform 1 0 2522 0 -1 100434
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_179_27
timestamp 1604489732
transform 1 0 2522 0 1 99346
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1453
timestamp 1604489732
transform 1 0 2890 0 -1 100434
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_359
timestamp 1604489732
transform -1 0 3902 0 -1 100434
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_357
timestamp 1604489732
transform -1 0 3902 0 1 99346
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1038
timestamp 1604489732
transform 1 0 83298 0 -1 99346
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1040
timestamp 1604489732
transform 1 0 83298 0 1 99346
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1042
timestamp 1604489732
transform 1 0 83298 0 -1 100434
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_178_908
timestamp 1604489732
transform 1 0 83574 0 -1 99346
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_908
timestamp 1604489732
transform 1 0 83574 0 1 99346
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_908
timestamp 1604489732
transform 1 0 83574 0 -1 100434
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_937
timestamp 1604489732
transform 1 0 86242 0 -1 99346
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_178_932
timestamp 1604489732
transform 1 0 85782 0 -1 99346
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_178_920
timestamp 1604489732
transform 1 0 84678 0 -1 99346
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1624
timestamp 1604489732
transform 1 0 86150 0 -1 99346
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_180_937
timestamp 1604489732
transform 1 0 86242 0 -1 100434
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_180_932
timestamp 1604489732
transform 1 0 85782 0 -1 100434
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_180_920
timestamp 1604489732
transform 1 0 84678 0 -1 100434
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_932
timestamp 1604489732
transform 1 0 85782 0 1 99346
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_920
timestamp 1604489732
transform 1 0 84678 0 1 99346
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1625
timestamp 1604489732
transform 1 0 86150 0 -1 100434
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1039
timestamp 1604489732
transform -1 0 87806 0 -1 99346
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1041
timestamp 1604489732
transform -1 0 87806 0 1 99346
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1043
timestamp 1604489732
transform -1 0 87806 0 -1 100434
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_178_949
timestamp 1604489732
transform 1 0 87346 0 -1 99346
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_179_944
timestamp 1604489732
transform 1 0 86886 0 1 99346
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_950
timestamp 1604489732
transform 1 0 87438 0 1 99346
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_180_949
timestamp 1604489732
transform 1 0 87346 0 -1 100434
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_182_15
timestamp 1604489732
transform 1 0 1418 0 -1 101522
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_3
timestamp 1604489732
transform 1 0 314 0 -1 101522
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_15
timestamp 1604489732
transform 1 0 1418 0 1 100434
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_3
timestamp 1604489732
transform 1 0 314 0 1 100434
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_362
timestamp 1604489732
transform 1 0 38 0 -1 101522
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_360
timestamp 1604489732
transform 1 0 38 0 1 100434
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_183_15
timestamp 1604489732
transform 1 0 1418 0 1 101522
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_3
timestamp 1604489732
transform 1 0 314 0 1 101522
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_364
timestamp 1604489732
transform 1 0 38 0 1 101522
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_184_15
timestamp 1604489732
transform 1 0 1418 0 -1 102610
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_3
timestamp 1604489732
transform 1 0 314 0 -1 102610
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_366
timestamp 1604489732
transform 1 0 38 0 -1 102610
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_182_38
timestamp 1604489732
transform 1 0 3534 0 -1 101522
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_182_32
timestamp 1604489732
transform 1 0 2982 0 -1 101522
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_182_27
timestamp 1604489732
transform 1 0 2522 0 -1 101522
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_181_27
timestamp 1604489732
transform 1 0 2522 0 1 100434
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1454
timestamp 1604489732
transform 1 0 2890 0 -1 101522
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_363
timestamp 1604489732
transform -1 0 3902 0 -1 101522
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_361
timestamp 1604489732
transform -1 0 3902 0 1 100434
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_183_27
timestamp 1604489732
transform 1 0 2522 0 1 101522
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_365
timestamp 1604489732
transform -1 0 3902 0 1 101522
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_184_38
timestamp 1604489732
transform 1 0 3534 0 -1 102610
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_184_32
timestamp 1604489732
transform 1 0 2982 0 -1 102610
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_184_27
timestamp 1604489732
transform 1 0 2522 0 -1 102610
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1455
timestamp 1604489732
transform 1 0 2890 0 -1 102610
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_367
timestamp 1604489732
transform -1 0 3902 0 -1 102610
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1044
timestamp 1604489732
transform 1 0 83298 0 1 100434
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1046
timestamp 1604489732
transform 1 0 83298 0 -1 101522
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1048
timestamp 1604489732
transform 1 0 83298 0 1 101522
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1050
timestamp 1604489732
transform 1 0 83298 0 -1 102610
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_181_908
timestamp 1604489732
transform 1 0 83574 0 1 100434
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_908
timestamp 1604489732
transform 1 0 83574 0 -1 101522
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_908
timestamp 1604489732
transform 1 0 83574 0 1 101522
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_908
timestamp 1604489732
transform 1 0 83574 0 -1 102610
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_937
timestamp 1604489732
transform 1 0 86242 0 -1 101522
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_182_932
timestamp 1604489732
transform 1 0 85782 0 -1 101522
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_182_920
timestamp 1604489732
transform 1 0 84678 0 -1 101522
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_932
timestamp 1604489732
transform 1 0 85782 0 1 100434
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_920
timestamp 1604489732
transform 1 0 84678 0 1 100434
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1626
timestamp 1604489732
transform 1 0 86150 0 -1 101522
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_183_932
timestamp 1604489732
transform 1 0 85782 0 1 101522
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_920
timestamp 1604489732
transform 1 0 84678 0 1 101522
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_937
timestamp 1604489732
transform 1 0 86242 0 -1 102610
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_184_932
timestamp 1604489732
transform 1 0 85782 0 -1 102610
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_184_920
timestamp 1604489732
transform 1 0 84678 0 -1 102610
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1627
timestamp 1604489732
transform 1 0 86150 0 -1 102610
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_181_944
timestamp 1604489732
transform 1 0 86886 0 1 100434
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_182_949
timestamp 1604489732
transform 1 0 87346 0 -1 101522
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_181_950
timestamp 1604489732
transform 1 0 87438 0 1 100434
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1047
timestamp 1604489732
transform -1 0 87806 0 -1 101522
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1045
timestamp 1604489732
transform -1 0 87806 0 1 100434
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_183_944
timestamp 1604489732
transform 1 0 86886 0 1 101522
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_183_950
timestamp 1604489732
transform 1 0 87438 0 1 101522
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1049
timestamp 1604489732
transform -1 0 87806 0 1 101522
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_184_949
timestamp 1604489732
transform 1 0 87346 0 -1 102610
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1051
timestamp 1604489732
transform -1 0 87806 0 -1 102610
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_368
timestamp 1604489732
transform 1 0 38 0 1 102610
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_370
timestamp 1604489732
transform 1 0 38 0 -1 103698
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_372
timestamp 1604489732
transform 1 0 38 0 1 103698
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_185_3
timestamp 1604489732
transform 1 0 314 0 1 102610
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_15
timestamp 1604489732
transform 1 0 1418 0 1 102610
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_3
timestamp 1604489732
transform 1 0 314 0 -1 103698
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_15
timestamp 1604489732
transform 1 0 1418 0 -1 103698
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_3
timestamp 1604489732
transform 1 0 314 0 1 103698
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_15
timestamp 1604489732
transform 1 0 1418 0 1 103698
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_369
timestamp 1604489732
transform -1 0 3902 0 1 102610
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_371
timestamp 1604489732
transform -1 0 3902 0 -1 103698
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_373
timestamp 1604489732
transform -1 0 3902 0 1 103698
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1456
timestamp 1604489732
transform 1 0 2890 0 -1 103698
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_27
timestamp 1604489732
transform 1 0 2522 0 1 102610
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_186_27
timestamp 1604489732
transform 1 0 2522 0 -1 103698
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_186_32
timestamp 1604489732
transform 1 0 2982 0 -1 103698
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_186_38
timestamp 1604489732
transform 1 0 3534 0 -1 103698
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_187_27
timestamp 1604489732
transform 1 0 2522 0 1 103698
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1052
timestamp 1604489732
transform 1 0 83298 0 1 102610
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1054
timestamp 1604489732
transform 1 0 83298 0 -1 103698
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1056
timestamp 1604489732
transform 1 0 83298 0 1 103698
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_185_908
timestamp 1604489732
transform 1 0 83574 0 1 102610
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_908
timestamp 1604489732
transform 1 0 83574 0 -1 103698
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_908
timestamp 1604489732
transform 1 0 83574 0 1 103698
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1628
timestamp 1604489732
transform 1 0 86150 0 -1 103698
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_920
timestamp 1604489732
transform 1 0 84678 0 1 102610
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_932
timestamp 1604489732
transform 1 0 85782 0 1 102610
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_920
timestamp 1604489732
transform 1 0 84678 0 -1 103698
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_186_932
timestamp 1604489732
transform 1 0 85782 0 -1 103698
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_186_937
timestamp 1604489732
transform 1 0 86242 0 -1 103698
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_920
timestamp 1604489732
transform 1 0 84678 0 1 103698
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_932
timestamp 1604489732
transform 1 0 85782 0 1 103698
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1053
timestamp 1604489732
transform -1 0 87806 0 1 102610
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1055
timestamp 1604489732
transform -1 0 87806 0 -1 103698
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1057
timestamp 1604489732
transform -1 0 87806 0 1 103698
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_185_944
timestamp 1604489732
transform 1 0 86886 0 1 102610
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_185_950
timestamp 1604489732
transform 1 0 87438 0 1 102610
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_186_949
timestamp 1604489732
transform 1 0 87346 0 -1 103698
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_187_944
timestamp 1604489732
transform 1 0 86886 0 1 103698
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_187_950
timestamp 1604489732
transform 1 0 87438 0 1 103698
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_374
timestamp 1604489732
transform 1 0 38 0 -1 104786
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_376
timestamp 1604489732
transform 1 0 38 0 1 104786
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_378
timestamp 1604489732
transform 1 0 38 0 -1 105874
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_188_3
timestamp 1604489732
transform 1 0 314 0 -1 104786
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_15
timestamp 1604489732
transform 1 0 1418 0 -1 104786
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_3
timestamp 1604489732
transform 1 0 314 0 1 104786
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_15
timestamp 1604489732
transform 1 0 1418 0 1 104786
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_3
timestamp 1604489732
transform 1 0 314 0 -1 105874
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_15
timestamp 1604489732
transform 1 0 1418 0 -1 105874
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_188_38
timestamp 1604489732
transform 1 0 3534 0 -1 104786
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_188_32
timestamp 1604489732
transform 1 0 2982 0 -1 104786
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_188_27
timestamp 1604489732
transform 1 0 2522 0 -1 104786
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1457
timestamp 1604489732
transform 1 0 2890 0 -1 104786
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_375
timestamp 1604489732
transform -1 0 3902 0 -1 104786
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_189_27
timestamp 1604489732
transform 1 0 2522 0 1 104786
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_377
timestamp 1604489732
transform -1 0 3902 0 1 104786
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_190_38
timestamp 1604489732
transform 1 0 3534 0 -1 105874
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_190_32
timestamp 1604489732
transform 1 0 2982 0 -1 105874
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_190_27
timestamp 1604489732
transform 1 0 2522 0 -1 105874
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1458
timestamp 1604489732
transform 1 0 2890 0 -1 105874
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_379
timestamp 1604489732
transform -1 0 3902 0 -1 105874
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1058
timestamp 1604489732
transform 1 0 83298 0 -1 104786
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1060
timestamp 1604489732
transform 1 0 83298 0 1 104786
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1062
timestamp 1604489732
transform 1 0 83298 0 -1 105874
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_188_908
timestamp 1604489732
transform 1 0 83574 0 -1 104786
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_908
timestamp 1604489732
transform 1 0 83574 0 1 104786
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_908
timestamp 1604489732
transform 1 0 83574 0 -1 105874
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_937
timestamp 1604489732
transform 1 0 86242 0 -1 104786
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_188_932
timestamp 1604489732
transform 1 0 85782 0 -1 104786
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_188_920
timestamp 1604489732
transform 1 0 84678 0 -1 104786
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1629
timestamp 1604489732
transform 1 0 86150 0 -1 104786
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_189_932
timestamp 1604489732
transform 1 0 85782 0 1 104786
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_920
timestamp 1604489732
transform 1 0 84678 0 1 104786
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_937
timestamp 1604489732
transform 1 0 86242 0 -1 105874
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_190_932
timestamp 1604489732
transform 1 0 85782 0 -1 105874
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_190_920
timestamp 1604489732
transform 1 0 84678 0 -1 105874
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1630
timestamp 1604489732
transform 1 0 86150 0 -1 105874
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1059
timestamp 1604489732
transform -1 0 87806 0 -1 104786
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1061
timestamp 1604489732
transform -1 0 87806 0 1 104786
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1063
timestamp 1604489732
transform -1 0 87806 0 -1 105874
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_188_949
timestamp 1604489732
transform 1 0 87346 0 -1 104786
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_189_944
timestamp 1604489732
transform 1 0 86886 0 1 104786
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_189_950
timestamp 1604489732
transform 1 0 87438 0 1 104786
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_190_949
timestamp 1604489732
transform 1 0 87346 0 -1 105874
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_192_15
timestamp 1604489732
transform 1 0 1418 0 -1 106962
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_3
timestamp 1604489732
transform 1 0 314 0 -1 106962
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_15
timestamp 1604489732
transform 1 0 1418 0 1 105874
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_3
timestamp 1604489732
transform 1 0 314 0 1 105874
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_382
timestamp 1604489732
transform 1 0 38 0 -1 106962
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_380
timestamp 1604489732
transform 1 0 38 0 1 105874
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_193_15
timestamp 1604489732
transform 1 0 1418 0 1 106962
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_3
timestamp 1604489732
transform 1 0 314 0 1 106962
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_384
timestamp 1604489732
transform 1 0 38 0 1 106962
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_194_15
timestamp 1604489732
transform 1 0 1418 0 -1 108050
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_3
timestamp 1604489732
transform 1 0 314 0 -1 108050
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_386
timestamp 1604489732
transform 1 0 38 0 -1 108050
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_192_38
timestamp 1604489732
transform 1 0 3534 0 -1 106962
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_192_32
timestamp 1604489732
transform 1 0 2982 0 -1 106962
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_192_27
timestamp 1604489732
transform 1 0 2522 0 -1 106962
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_191_27
timestamp 1604489732
transform 1 0 2522 0 1 105874
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1459
timestamp 1604489732
transform 1 0 2890 0 -1 106962
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_383
timestamp 1604489732
transform -1 0 3902 0 -1 106962
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_381
timestamp 1604489732
transform -1 0 3902 0 1 105874
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_193_27
timestamp 1604489732
transform 1 0 2522 0 1 106962
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_385
timestamp 1604489732
transform -1 0 3902 0 1 106962
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_194_38
timestamp 1604489732
transform 1 0 3534 0 -1 108050
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_194_32
timestamp 1604489732
transform 1 0 2982 0 -1 108050
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_194_27
timestamp 1604489732
transform 1 0 2522 0 -1 108050
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1460
timestamp 1604489732
transform 1 0 2890 0 -1 108050
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_387
timestamp 1604489732
transform -1 0 3902 0 -1 108050
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1064
timestamp 1604489732
transform 1 0 83298 0 1 105874
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1066
timestamp 1604489732
transform 1 0 83298 0 -1 106962
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1068
timestamp 1604489732
transform 1 0 83298 0 1 106962
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1070
timestamp 1604489732
transform 1 0 83298 0 -1 108050
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_191_908
timestamp 1604489732
transform 1 0 83574 0 1 105874
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_908
timestamp 1604489732
transform 1 0 83574 0 -1 106962
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_908
timestamp 1604489732
transform 1 0 83574 0 1 106962
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_908
timestamp 1604489732
transform 1 0 83574 0 -1 108050
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_937
timestamp 1604489732
transform 1 0 86242 0 -1 106962
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_192_932
timestamp 1604489732
transform 1 0 85782 0 -1 106962
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_192_920
timestamp 1604489732
transform 1 0 84678 0 -1 106962
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_932
timestamp 1604489732
transform 1 0 85782 0 1 105874
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_920
timestamp 1604489732
transform 1 0 84678 0 1 105874
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1631
timestamp 1604489732
transform 1 0 86150 0 -1 106962
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_193_932
timestamp 1604489732
transform 1 0 85782 0 1 106962
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_920
timestamp 1604489732
transform 1 0 84678 0 1 106962
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_937
timestamp 1604489732
transform 1 0 86242 0 -1 108050
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_194_932
timestamp 1604489732
transform 1 0 85782 0 -1 108050
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_194_920
timestamp 1604489732
transform 1 0 84678 0 -1 108050
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1632
timestamp 1604489732
transform 1 0 86150 0 -1 108050
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_191_944
timestamp 1604489732
transform 1 0 86886 0 1 105874
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_192_949
timestamp 1604489732
transform 1 0 87346 0 -1 106962
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_191_950
timestamp 1604489732
transform 1 0 87438 0 1 105874
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1067
timestamp 1604489732
transform -1 0 87806 0 -1 106962
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1065
timestamp 1604489732
transform -1 0 87806 0 1 105874
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_193_944
timestamp 1604489732
transform 1 0 86886 0 1 106962
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_193_950
timestamp 1604489732
transform 1 0 87438 0 1 106962
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1069
timestamp 1604489732
transform -1 0 87806 0 1 106962
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_194_949
timestamp 1604489732
transform 1 0 87346 0 -1 108050
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1071
timestamp 1604489732
transform -1 0 87806 0 -1 108050
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_388
timestamp 1604489732
transform 1 0 38 0 1 108050
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_390
timestamp 1604489732
transform 1 0 38 0 -1 109138
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_392
timestamp 1604489732
transform 1 0 38 0 1 109138
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_195_3
timestamp 1604489732
transform 1 0 314 0 1 108050
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_15
timestamp 1604489732
transform 1 0 1418 0 1 108050
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_3
timestamp 1604489732
transform 1 0 314 0 -1 109138
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_15
timestamp 1604489732
transform 1 0 1418 0 -1 109138
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_3
timestamp 1604489732
transform 1 0 314 0 1 109138
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_15
timestamp 1604489732
transform 1 0 1418 0 1 109138
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_389
timestamp 1604489732
transform -1 0 3902 0 1 108050
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_391
timestamp 1604489732
transform -1 0 3902 0 -1 109138
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_393
timestamp 1604489732
transform -1 0 3902 0 1 109138
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1461
timestamp 1604489732
transform 1 0 2890 0 -1 109138
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_195_27
timestamp 1604489732
transform 1 0 2522 0 1 108050
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_196_27
timestamp 1604489732
transform 1 0 2522 0 -1 109138
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_196_32
timestamp 1604489732
transform 1 0 2982 0 -1 109138
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_196_38
timestamp 1604489732
transform 1 0 3534 0 -1 109138
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_197_27
timestamp 1604489732
transform 1 0 2522 0 1 109138
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1072
timestamp 1604489732
transform 1 0 83298 0 1 108050
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1074
timestamp 1604489732
transform 1 0 83298 0 -1 109138
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1076
timestamp 1604489732
transform 1 0 83298 0 1 109138
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_195_908
timestamp 1604489732
transform 1 0 83574 0 1 108050
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_908
timestamp 1604489732
transform 1 0 83574 0 -1 109138
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_908
timestamp 1604489732
transform 1 0 83574 0 1 109138
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1633
timestamp 1604489732
transform 1 0 86150 0 -1 109138
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_195_920
timestamp 1604489732
transform 1 0 84678 0 1 108050
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_932
timestamp 1604489732
transform 1 0 85782 0 1 108050
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_920
timestamp 1604489732
transform 1 0 84678 0 -1 109138
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_196_932
timestamp 1604489732
transform 1 0 85782 0 -1 109138
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_196_937
timestamp 1604489732
transform 1 0 86242 0 -1 109138
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_920
timestamp 1604489732
transform 1 0 84678 0 1 109138
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_932
timestamp 1604489732
transform 1 0 85782 0 1 109138
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1073
timestamp 1604489732
transform -1 0 87806 0 1 108050
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1075
timestamp 1604489732
transform -1 0 87806 0 -1 109138
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1077
timestamp 1604489732
transform -1 0 87806 0 1 109138
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_195_944
timestamp 1604489732
transform 1 0 86886 0 1 108050
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_195_950
timestamp 1604489732
transform 1 0 87438 0 1 108050
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_196_949
timestamp 1604489732
transform 1 0 87346 0 -1 109138
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_197_944
timestamp 1604489732
transform 1 0 86886 0 1 109138
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_197_950
timestamp 1604489732
transform 1 0 87438 0 1 109138
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_394
timestamp 1604489732
transform 1 0 38 0 -1 110226
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_396
timestamp 1604489732
transform 1 0 38 0 1 110226
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_398
timestamp 1604489732
transform 1 0 38 0 -1 111314
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_198_3
timestamp 1604489732
transform 1 0 314 0 -1 110226
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_15
timestamp 1604489732
transform 1 0 1418 0 -1 110226
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_3
timestamp 1604489732
transform 1 0 314 0 1 110226
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_15
timestamp 1604489732
transform 1 0 1418 0 1 110226
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_3
timestamp 1604489732
transform 1 0 314 0 -1 111314
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_15
timestamp 1604489732
transform 1 0 1418 0 -1 111314
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_198_38
timestamp 1604489732
transform 1 0 3534 0 -1 110226
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_198_32
timestamp 1604489732
transform 1 0 2982 0 -1 110226
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_198_27
timestamp 1604489732
transform 1 0 2522 0 -1 110226
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1462
timestamp 1604489732
transform 1 0 2890 0 -1 110226
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_395
timestamp 1604489732
transform -1 0 3902 0 -1 110226
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_199_27
timestamp 1604489732
transform 1 0 2522 0 1 110226
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_397
timestamp 1604489732
transform -1 0 3902 0 1 110226
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_200_38
timestamp 1604489732
transform 1 0 3534 0 -1 111314
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_200_32
timestamp 1604489732
transform 1 0 2982 0 -1 111314
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_200_27
timestamp 1604489732
transform 1 0 2522 0 -1 111314
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1463
timestamp 1604489732
transform 1 0 2890 0 -1 111314
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_399
timestamp 1604489732
transform -1 0 3902 0 -1 111314
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1078
timestamp 1604489732
transform 1 0 83298 0 -1 110226
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1080
timestamp 1604489732
transform 1 0 83298 0 1 110226
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1082
timestamp 1604489732
transform 1 0 83298 0 -1 111314
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_198_908
timestamp 1604489732
transform 1 0 83574 0 -1 110226
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_908
timestamp 1604489732
transform 1 0 83574 0 1 110226
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_908
timestamp 1604489732
transform 1 0 83574 0 -1 111314
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_937
timestamp 1604489732
transform 1 0 86242 0 -1 110226
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_198_932
timestamp 1604489732
transform 1 0 85782 0 -1 110226
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_198_920
timestamp 1604489732
transform 1 0 84678 0 -1 110226
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1634
timestamp 1604489732
transform 1 0 86150 0 -1 110226
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_199_932
timestamp 1604489732
transform 1 0 85782 0 1 110226
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_920
timestamp 1604489732
transform 1 0 84678 0 1 110226
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_937
timestamp 1604489732
transform 1 0 86242 0 -1 111314
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_200_932
timestamp 1604489732
transform 1 0 85782 0 -1 111314
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_200_920
timestamp 1604489732
transform 1 0 84678 0 -1 111314
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1635
timestamp 1604489732
transform 1 0 86150 0 -1 111314
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1079
timestamp 1604489732
transform -1 0 87806 0 -1 110226
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1081
timestamp 1604489732
transform -1 0 87806 0 1 110226
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1083
timestamp 1604489732
transform -1 0 87806 0 -1 111314
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_198_949
timestamp 1604489732
transform 1 0 87346 0 -1 110226
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_199_944
timestamp 1604489732
transform 1 0 86886 0 1 110226
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_199_950
timestamp 1604489732
transform 1 0 87438 0 1 110226
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_200_949
timestamp 1604489732
transform 1 0 87346 0 -1 111314
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_202_15
timestamp 1604489732
transform 1 0 1418 0 -1 112402
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_3
timestamp 1604489732
transform 1 0 314 0 -1 112402
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_15
timestamp 1604489732
transform 1 0 1418 0 1 111314
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_3
timestamp 1604489732
transform 1 0 314 0 1 111314
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_402
timestamp 1604489732
transform 1 0 38 0 -1 112402
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_400
timestamp 1604489732
transform 1 0 38 0 1 111314
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_203_15
timestamp 1604489732
transform 1 0 1418 0 1 112402
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_3
timestamp 1604489732
transform 1 0 314 0 1 112402
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_404
timestamp 1604489732
transform 1 0 38 0 1 112402
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_204_15
timestamp 1604489732
transform 1 0 1418 0 -1 113490
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_3
timestamp 1604489732
transform 1 0 314 0 -1 113490
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_406
timestamp 1604489732
transform 1 0 38 0 -1 113490
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_202_38
timestamp 1604489732
transform 1 0 3534 0 -1 112402
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_202_32
timestamp 1604489732
transform 1 0 2982 0 -1 112402
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_202_27
timestamp 1604489732
transform 1 0 2522 0 -1 112402
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_201_27
timestamp 1604489732
transform 1 0 2522 0 1 111314
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1464
timestamp 1604489732
transform 1 0 2890 0 -1 112402
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_403
timestamp 1604489732
transform -1 0 3902 0 -1 112402
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_401
timestamp 1604489732
transform -1 0 3902 0 1 111314
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_203_27
timestamp 1604489732
transform 1 0 2522 0 1 112402
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_405
timestamp 1604489732
transform -1 0 3902 0 1 112402
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_204_38
timestamp 1604489732
transform 1 0 3534 0 -1 113490
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_204_32
timestamp 1604489732
transform 1 0 2982 0 -1 113490
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_204_27
timestamp 1604489732
transform 1 0 2522 0 -1 113490
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1465
timestamp 1604489732
transform 1 0 2890 0 -1 113490
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_407
timestamp 1604489732
transform -1 0 3902 0 -1 113490
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1084
timestamp 1604489732
transform 1 0 83298 0 1 111314
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1086
timestamp 1604489732
transform 1 0 83298 0 -1 112402
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1088
timestamp 1604489732
transform 1 0 83298 0 1 112402
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1090
timestamp 1604489732
transform 1 0 83298 0 -1 113490
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_201_908
timestamp 1604489732
transform 1 0 83574 0 1 111314
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_908
timestamp 1604489732
transform 1 0 83574 0 -1 112402
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_908
timestamp 1604489732
transform 1 0 83574 0 1 112402
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_908
timestamp 1604489732
transform 1 0 83574 0 -1 113490
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_937
timestamp 1604489732
transform 1 0 86242 0 -1 112402
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_202_932
timestamp 1604489732
transform 1 0 85782 0 -1 112402
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_202_920
timestamp 1604489732
transform 1 0 84678 0 -1 112402
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_932
timestamp 1604489732
transform 1 0 85782 0 1 111314
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_920
timestamp 1604489732
transform 1 0 84678 0 1 111314
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1636
timestamp 1604489732
transform 1 0 86150 0 -1 112402
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_203_932
timestamp 1604489732
transform 1 0 85782 0 1 112402
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_920
timestamp 1604489732
transform 1 0 84678 0 1 112402
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_937
timestamp 1604489732
transform 1 0 86242 0 -1 113490
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_204_932
timestamp 1604489732
transform 1 0 85782 0 -1 113490
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_204_920
timestamp 1604489732
transform 1 0 84678 0 -1 113490
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1637
timestamp 1604489732
transform 1 0 86150 0 -1 113490
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_201_944
timestamp 1604489732
transform 1 0 86886 0 1 111314
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_202_949
timestamp 1604489732
transform 1 0 87346 0 -1 112402
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_201_950
timestamp 1604489732
transform 1 0 87438 0 1 111314
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1087
timestamp 1604489732
transform -1 0 87806 0 -1 112402
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1085
timestamp 1604489732
transform -1 0 87806 0 1 111314
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_203_944
timestamp 1604489732
transform 1 0 86886 0 1 112402
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_203_950
timestamp 1604489732
transform 1 0 87438 0 1 112402
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1089
timestamp 1604489732
transform -1 0 87806 0 1 112402
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_204_949
timestamp 1604489732
transform 1 0 87346 0 -1 113490
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1091
timestamp 1604489732
transform -1 0 87806 0 -1 113490
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_408
timestamp 1604489732
transform 1 0 38 0 1 113490
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_410
timestamp 1604489732
transform 1 0 38 0 -1 114578
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_412
timestamp 1604489732
transform 1 0 38 0 1 114578
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_205_3
timestamp 1604489732
transform 1 0 314 0 1 113490
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_15
timestamp 1604489732
transform 1 0 1418 0 1 113490
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_3
timestamp 1604489732
transform 1 0 314 0 -1 114578
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_15
timestamp 1604489732
transform 1 0 1418 0 -1 114578
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_3
timestamp 1604489732
transform 1 0 314 0 1 114578
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_15
timestamp 1604489732
transform 1 0 1418 0 1 114578
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_27
timestamp 1604489732
transform 1 0 2522 0 1 113490
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_409
timestamp 1604489732
transform -1 0 3902 0 1 113490
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_206_38
timestamp 1604489732
transform 1 0 3534 0 -1 114578
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_206_32
timestamp 1604489732
transform 1 0 2982 0 -1 114578
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_206_27
timestamp 1604489732
transform 1 0 2522 0 -1 114578
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1466
timestamp 1604489732
transform 1 0 2890 0 -1 114578
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_411
timestamp 1604489732
transform -1 0 3902 0 -1 114578
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_207_35
timestamp 1604489732
transform 1 0 3258 0 1 114578
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_207_27
timestamp 1604489732
transform 1 0 2522 0 1 114578
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_csb0
timestamp 1604489732
transform 1 0 3442 0 1 114578
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_413
timestamp 1604489732
transform -1 0 3902 0 1 114578
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1092
timestamp 1604489732
transform 1 0 83298 0 1 113490
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1094
timestamp 1604489732
transform 1 0 83298 0 -1 114578
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1096
timestamp 1604489732
transform 1 0 83298 0 1 114578
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_205_908
timestamp 1604489732
transform 1 0 83574 0 1 113490
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_908
timestamp 1604489732
transform 1 0 83574 0 -1 114578
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_908
timestamp 1604489732
transform 1 0 83574 0 1 114578
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1638
timestamp 1604489732
transform 1 0 86150 0 -1 114578
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_205_920
timestamp 1604489732
transform 1 0 84678 0 1 113490
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_932
timestamp 1604489732
transform 1 0 85782 0 1 113490
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_920
timestamp 1604489732
transform 1 0 84678 0 -1 114578
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_206_932
timestamp 1604489732
transform 1 0 85782 0 -1 114578
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_206_937
timestamp 1604489732
transform 1 0 86242 0 -1 114578
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_920
timestamp 1604489732
transform 1 0 84678 0 1 114578
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_932
timestamp 1604489732
transform 1 0 85782 0 1 114578
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1093
timestamp 1604489732
transform -1 0 87806 0 1 113490
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1095
timestamp 1604489732
transform -1 0 87806 0 -1 114578
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1097
timestamp 1604489732
transform -1 0 87806 0 1 114578
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_205_944
timestamp 1604489732
transform 1 0 86886 0 1 113490
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_205_950
timestamp 1604489732
transform 1 0 87438 0 1 113490
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_206_949
timestamp 1604489732
transform 1 0 87346 0 -1 114578
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_207_944
timestamp 1604489732
transform 1 0 86886 0 1 114578
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_207_950
timestamp 1604489732
transform 1 0 87438 0 1 114578
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_414
timestamp 1604489732
transform 1 0 38 0 -1 115666
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_416
timestamp 1604489732
transform 1 0 38 0 1 115666
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_418
timestamp 1604489732
transform 1 0 38 0 -1 116754
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_208_3
timestamp 1604489732
transform 1 0 314 0 -1 115666
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_15
timestamp 1604489732
transform 1 0 1418 0 -1 115666
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_3
timestamp 1604489732
transform 1 0 314 0 1 115666
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_15
timestamp 1604489732
transform 1 0 1418 0 1 115666
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_3
timestamp 1604489732
transform 1 0 314 0 -1 116754
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_15
timestamp 1604489732
transform 1 0 1418 0 -1 116754
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_208_38
timestamp 1604489732
transform 1 0 3534 0 -1 115666
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_208_32
timestamp 1604489732
transform 1 0 2982 0 -1 115666
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_208_27
timestamp 1604489732
transform 1 0 2522 0 -1 115666
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1467
timestamp 1604489732
transform 1 0 2890 0 -1 115666
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_415
timestamp 1604489732
transform -1 0 3902 0 -1 115666
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_209_27
timestamp 1604489732
transform 1 0 2522 0 1 115666
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_417
timestamp 1604489732
transform -1 0 3902 0 1 115666
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_210_36
timestamp 1604489732
transform 1 0 3350 0 -1 116754
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_210_32
timestamp 1604489732
transform 1 0 2982 0 -1 116754
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_27
timestamp 1604489732
transform 1 0 2522 0 -1 116754
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_web0
timestamp 1604489732
transform 1 0 3442 0 -1 116754
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1468
timestamp 1604489732
transform 1 0 2890 0 -1 116754
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_419
timestamp 1604489732
transform -1 0 3902 0 -1 116754
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1098
timestamp 1604489732
transform 1 0 83298 0 -1 115666
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1100
timestamp 1604489732
transform 1 0 83298 0 1 115666
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1102
timestamp 1604489732
transform 1 0 83298 0 -1 116754
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_208_908
timestamp 1604489732
transform 1 0 83574 0 -1 115666
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_908
timestamp 1604489732
transform 1 0 83574 0 1 115666
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_908
timestamp 1604489732
transform 1 0 83574 0 -1 116754
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_937
timestamp 1604489732
transform 1 0 86242 0 -1 115666
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_208_932
timestamp 1604489732
transform 1 0 85782 0 -1 115666
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_208_920
timestamp 1604489732
transform 1 0 84678 0 -1 115666
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1639
timestamp 1604489732
transform 1 0 86150 0 -1 115666
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_209_932
timestamp 1604489732
transform 1 0 85782 0 1 115666
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_920
timestamp 1604489732
transform 1 0 84678 0 1 115666
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_937
timestamp 1604489732
transform 1 0 86242 0 -1 116754
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_210_932
timestamp 1604489732
transform 1 0 85782 0 -1 116754
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_210_920
timestamp 1604489732
transform 1 0 84678 0 -1 116754
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1640
timestamp 1604489732
transform 1 0 86150 0 -1 116754
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1099
timestamp 1604489732
transform -1 0 87806 0 -1 115666
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1101
timestamp 1604489732
transform -1 0 87806 0 1 115666
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1103
timestamp 1604489732
transform -1 0 87806 0 -1 116754
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_208_949
timestamp 1604489732
transform 1 0 87346 0 -1 115666
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_209_944
timestamp 1604489732
transform 1 0 86886 0 1 115666
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_209_950
timestamp 1604489732
transform 1 0 87438 0 1 115666
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_210_949
timestamp 1604489732
transform 1 0 87346 0 -1 116754
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_211_15
timestamp 1604489732
transform 1 0 1418 0 1 116754
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_211_3
timestamp 1604489732
transform 1 0 314 0 1 116754
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_420
timestamp 1604489732
transform 1 0 38 0 1 116754
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_213_15
timestamp 1604489732
transform 1 0 1418 0 1 117842
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_213_3
timestamp 1604489732
transform 1 0 314 0 1 117842
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_212_15
timestamp 1604489732
transform 1 0 1418 0 -1 117842
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_212_3
timestamp 1604489732
transform 1 0 314 0 -1 117842
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_424
timestamp 1604489732
transform 1 0 38 0 1 117842
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_422
timestamp 1604489732
transform 1 0 38 0 -1 117842
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_214_15
timestamp 1604489732
transform 1 0 1418 0 -1 118930
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_214_3
timestamp 1604489732
transform 1 0 314 0 -1 118930
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_426
timestamp 1604489732
transform 1 0 38 0 -1 118930
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_211_27
timestamp 1604489732
transform 1 0 2522 0 1 116754
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_421
timestamp 1604489732
transform -1 0 3902 0 1 116754
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_213_27
timestamp 1604489732
transform 1 0 2522 0 1 117842
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_212_38
timestamp 1604489732
transform 1 0 3534 0 -1 117842
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_212_32
timestamp 1604489732
transform 1 0 2982 0 -1 117842
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_212_27
timestamp 1604489732
transform 1 0 2522 0 -1 117842
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1469
timestamp 1604489732
transform 1 0 2890 0 -1 117842
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_425
timestamp 1604489732
transform -1 0 3902 0 1 117842
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_423
timestamp 1604489732
transform -1 0 3902 0 -1 117842
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_214_38
timestamp 1604489732
transform 1 0 3534 0 -1 118930
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_214_32
timestamp 1604489732
transform 1 0 2982 0 -1 118930
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_214_27
timestamp 1604489732
transform 1 0 2522 0 -1 118930
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1470
timestamp 1604489732
transform 1 0 2890 0 -1 118930
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_427
timestamp 1604489732
transform -1 0 3902 0 -1 118930
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1104
timestamp 1604489732
transform 1 0 83298 0 1 116754
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1106
timestamp 1604489732
transform 1 0 83298 0 -1 117842
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1108
timestamp 1604489732
transform 1 0 83298 0 1 117842
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1110
timestamp 1604489732
transform 1 0 83298 0 -1 118930
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_211_908
timestamp 1604489732
transform 1 0 83574 0 1 116754
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_212_908
timestamp 1604489732
transform 1 0 83574 0 -1 117842
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_213_908
timestamp 1604489732
transform 1 0 83574 0 1 117842
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_214_908
timestamp 1604489732
transform 1 0 83574 0 -1 118930
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_211_932
timestamp 1604489732
transform 1 0 85782 0 1 116754
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_211_920
timestamp 1604489732
transform 1 0 84678 0 1 116754
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_213_932
timestamp 1604489732
transform 1 0 85782 0 1 117842
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_213_920
timestamp 1604489732
transform 1 0 84678 0 1 117842
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_212_937
timestamp 1604489732
transform 1 0 86242 0 -1 117842
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_212_932
timestamp 1604489732
transform 1 0 85782 0 -1 117842
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_212_920
timestamp 1604489732
transform 1 0 84678 0 -1 117842
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1641
timestamp 1604489732
transform 1 0 86150 0 -1 117842
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_214_937
timestamp 1604489732
transform 1 0 86242 0 -1 118930
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_214_932
timestamp 1604489732
transform 1 0 85782 0 -1 118930
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_214_920
timestamp 1604489732
transform 1 0 84678 0 -1 118930
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1642
timestamp 1604489732
transform 1 0 86150 0 -1 118930
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_211_944
timestamp 1604489732
transform 1 0 86886 0 1 116754
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_211_950
timestamp 1604489732
transform 1 0 87438 0 1 116754
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1105
timestamp 1604489732
transform -1 0 87806 0 1 116754
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_213_944
timestamp 1604489732
transform 1 0 86886 0 1 117842
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_213_950
timestamp 1604489732
transform 1 0 87438 0 1 117842
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_212_949
timestamp 1604489732
transform 1 0 87346 0 -1 117842
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1109
timestamp 1604489732
transform -1 0 87806 0 1 117842
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1107
timestamp 1604489732
transform -1 0 87806 0 -1 117842
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_214_949
timestamp 1604489732
transform 1 0 87346 0 -1 118930
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1111
timestamp 1604489732
transform -1 0 87806 0 -1 118930
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_428
timestamp 1604489732
transform 1 0 38 0 1 118930
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_430
timestamp 1604489732
transform 1 0 38 0 -1 120018
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_432
timestamp 1604489732
transform 1 0 38 0 1 120018
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_215_3
timestamp 1604489732
transform 1 0 314 0 1 118930
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_215_15
timestamp 1604489732
transform 1 0 1418 0 1 118930
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_216_3
timestamp 1604489732
transform 1 0 314 0 -1 120018
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_216_15
timestamp 1604489732
transform 1 0 1418 0 -1 120018
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_217_3
timestamp 1604489732
transform 1 0 314 0 1 120018
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_217_15
timestamp 1604489732
transform 1 0 1418 0 1 120018
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_429
timestamp 1604489732
transform -1 0 3902 0 1 118930
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_431
timestamp 1604489732
transform -1 0 3902 0 -1 120018
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_433
timestamp 1604489732
transform -1 0 3902 0 1 120018
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1471
timestamp 1604489732
transform 1 0 2890 0 -1 120018
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_215_27
timestamp 1604489732
transform 1 0 2522 0 1 118930
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_216_27
timestamp 1604489732
transform 1 0 2522 0 -1 120018
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_216_32
timestamp 1604489732
transform 1 0 2982 0 -1 120018
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_216_38
timestamp 1604489732
transform 1 0 3534 0 -1 120018
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_217_27
timestamp 1604489732
transform 1 0 2522 0 1 120018
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1112
timestamp 1604489732
transform 1 0 83298 0 1 118930
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1114
timestamp 1604489732
transform 1 0 83298 0 -1 120018
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1116
timestamp 1604489732
transform 1 0 83298 0 1 120018
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_215_908
timestamp 1604489732
transform 1 0 83574 0 1 118930
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_216_908
timestamp 1604489732
transform 1 0 83574 0 -1 120018
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_217_908
timestamp 1604489732
transform 1 0 83574 0 1 120018
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1643
timestamp 1604489732
transform 1 0 86150 0 -1 120018
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_215_920
timestamp 1604489732
transform 1 0 84678 0 1 118930
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_215_932
timestamp 1604489732
transform 1 0 85782 0 1 118930
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_216_920
timestamp 1604489732
transform 1 0 84678 0 -1 120018
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_216_932
timestamp 1604489732
transform 1 0 85782 0 -1 120018
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_216_937
timestamp 1604489732
transform 1 0 86242 0 -1 120018
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_217_920
timestamp 1604489732
transform 1 0 84678 0 1 120018
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_217_932
timestamp 1604489732
transform 1 0 85782 0 1 120018
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1113
timestamp 1604489732
transform -1 0 87806 0 1 118930
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1115
timestamp 1604489732
transform -1 0 87806 0 -1 120018
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1117
timestamp 1604489732
transform -1 0 87806 0 1 120018
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_215_944
timestamp 1604489732
transform 1 0 86886 0 1 118930
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_215_950
timestamp 1604489732
transform 1 0 87438 0 1 118930
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_216_949
timestamp 1604489732
transform 1 0 87346 0 -1 120018
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_217_944
timestamp 1604489732
transform 1 0 86886 0 1 120018
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_217_950
timestamp 1604489732
transform 1 0 87438 0 1 120018
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_434
timestamp 1604489732
transform 1 0 38 0 -1 121106
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_436
timestamp 1604489732
transform 1 0 38 0 1 121106
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_438
timestamp 1604489732
transform 1 0 38 0 -1 122194
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_218_3
timestamp 1604489732
transform 1 0 314 0 -1 121106
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_218_15
timestamp 1604489732
transform 1 0 1418 0 -1 121106
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_219_3
timestamp 1604489732
transform 1 0 314 0 1 121106
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_219_15
timestamp 1604489732
transform 1 0 1418 0 1 121106
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_220_3
timestamp 1604489732
transform 1 0 314 0 -1 122194
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_220_15
timestamp 1604489732
transform 1 0 1418 0 -1 122194
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_218_38
timestamp 1604489732
transform 1 0 3534 0 -1 121106
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_218_32
timestamp 1604489732
transform 1 0 2982 0 -1 121106
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_218_27
timestamp 1604489732
transform 1 0 2522 0 -1 121106
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1472
timestamp 1604489732
transform 1 0 2890 0 -1 121106
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_435
timestamp 1604489732
transform -1 0 3902 0 -1 121106
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_219_27
timestamp 1604489732
transform 1 0 2522 0 1 121106
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_437
timestamp 1604489732
transform -1 0 3902 0 1 121106
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_220_38
timestamp 1604489732
transform 1 0 3534 0 -1 122194
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_220_32
timestamp 1604489732
transform 1 0 2982 0 -1 122194
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_220_27
timestamp 1604489732
transform 1 0 2522 0 -1 122194
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1473
timestamp 1604489732
transform 1 0 2890 0 -1 122194
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_439
timestamp 1604489732
transform -1 0 3902 0 -1 122194
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1118
timestamp 1604489732
transform 1 0 83298 0 -1 121106
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1120
timestamp 1604489732
transform 1 0 83298 0 1 121106
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1122
timestamp 1604489732
transform 1 0 83298 0 -1 122194
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_218_908
timestamp 1604489732
transform 1 0 83574 0 -1 121106
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_219_908
timestamp 1604489732
transform 1 0 83574 0 1 121106
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_220_908
timestamp 1604489732
transform 1 0 83574 0 -1 122194
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_218_937
timestamp 1604489732
transform 1 0 86242 0 -1 121106
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_218_932
timestamp 1604489732
transform 1 0 85782 0 -1 121106
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_218_920
timestamp 1604489732
transform 1 0 84678 0 -1 121106
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1644
timestamp 1604489732
transform 1 0 86150 0 -1 121106
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_219_932
timestamp 1604489732
transform 1 0 85782 0 1 121106
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_219_920
timestamp 1604489732
transform 1 0 84678 0 1 121106
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_220_937
timestamp 1604489732
transform 1 0 86242 0 -1 122194
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_220_932
timestamp 1604489732
transform 1 0 85782 0 -1 122194
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_220_920
timestamp 1604489732
transform 1 0 84678 0 -1 122194
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1645
timestamp 1604489732
transform 1 0 86150 0 -1 122194
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1119
timestamp 1604489732
transform -1 0 87806 0 -1 121106
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1121
timestamp 1604489732
transform -1 0 87806 0 1 121106
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1123
timestamp 1604489732
transform -1 0 87806 0 -1 122194
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_218_949
timestamp 1604489732
transform 1 0 87346 0 -1 121106
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_219_944
timestamp 1604489732
transform 1 0 86886 0 1 121106
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_219_950
timestamp 1604489732
transform 1 0 87438 0 1 121106
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_220_949
timestamp 1604489732
transform 1 0 87346 0 -1 122194
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_440
timestamp 1604489732
transform 1 0 38 0 1 122194
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_442
timestamp 1604489732
transform 1 0 38 0 -1 123282
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_444
timestamp 1604489732
transform 1 0 38 0 1 123282
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_221_3
timestamp 1604489732
transform 1 0 314 0 1 122194
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_221_15
timestamp 1604489732
transform 1 0 1418 0 1 122194
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_222_3
timestamp 1604489732
transform 1 0 314 0 -1 123282
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_222_15
timestamp 1604489732
transform 1 0 1418 0 -1 123282
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_223_3
timestamp 1604489732
transform 1 0 314 0 1 123282
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_223_15
timestamp 1604489732
transform 1 0 1418 0 1 123282
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_441
timestamp 1604489732
transform -1 0 3902 0 1 122194
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_443
timestamp 1604489732
transform -1 0 3902 0 -1 123282
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_445
timestamp 1604489732
transform -1 0 3902 0 1 123282
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1474
timestamp 1604489732
transform 1 0 2890 0 -1 123282
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_221_27
timestamp 1604489732
transform 1 0 2522 0 1 122194
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_222_27
timestamp 1604489732
transform 1 0 2522 0 -1 123282
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_222_32
timestamp 1604489732
transform 1 0 2982 0 -1 123282
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_222_38
timestamp 1604489732
transform 1 0 3534 0 -1 123282
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_223_27
timestamp 1604489732
transform 1 0 2522 0 1 123282
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1124
timestamp 1604489732
transform 1 0 83298 0 1 122194
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1126
timestamp 1604489732
transform 1 0 83298 0 -1 123282
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1128
timestamp 1604489732
transform 1 0 83298 0 1 123282
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_221_908
timestamp 1604489732
transform 1 0 83574 0 1 122194
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_222_908
timestamp 1604489732
transform 1 0 83574 0 -1 123282
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_223_908
timestamp 1604489732
transform 1 0 83574 0 1 123282
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1646
timestamp 1604489732
transform 1 0 86150 0 -1 123282
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_221_920
timestamp 1604489732
transform 1 0 84678 0 1 122194
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_221_932
timestamp 1604489732
transform 1 0 85782 0 1 122194
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_222_920
timestamp 1604489732
transform 1 0 84678 0 -1 123282
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_222_932
timestamp 1604489732
transform 1 0 85782 0 -1 123282
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_222_937
timestamp 1604489732
transform 1 0 86242 0 -1 123282
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_223_920
timestamp 1604489732
transform 1 0 84678 0 1 123282
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_223_932
timestamp 1604489732
transform 1 0 85782 0 1 123282
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1125
timestamp 1604489732
transform -1 0 87806 0 1 122194
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1127
timestamp 1604489732
transform -1 0 87806 0 -1 123282
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1129
timestamp 1604489732
transform -1 0 87806 0 1 123282
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_221_944
timestamp 1604489732
transform 1 0 86886 0 1 122194
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_221_950
timestamp 1604489732
transform 1 0 87438 0 1 122194
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_222_949
timestamp 1604489732
transform 1 0 87346 0 -1 123282
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_223_944
timestamp 1604489732
transform 1 0 86886 0 1 123282
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_223_950
timestamp 1604489732
transform 1 0 87438 0 1 123282
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_225_15
timestamp 1604489732
transform 1 0 1418 0 1 124370
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_225_3
timestamp 1604489732
transform 1 0 314 0 1 124370
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_224_15
timestamp 1604489732
transform 1 0 1418 0 -1 124370
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_224_3
timestamp 1604489732
transform 1 0 314 0 -1 124370
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_448
timestamp 1604489732
transform 1 0 38 0 1 124370
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_446
timestamp 1604489732
transform 1 0 38 0 -1 124370
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_226_15
timestamp 1604489732
transform 1 0 1418 0 -1 125458
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_226_3
timestamp 1604489732
transform 1 0 314 0 -1 125458
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_450
timestamp 1604489732
transform 1 0 38 0 -1 125458
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_227_15
timestamp 1604489732
transform 1 0 1418 0 1 125458
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_227_3
timestamp 1604489732
transform 1 0 314 0 1 125458
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_452
timestamp 1604489732
transform 1 0 38 0 1 125458
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_225_27
timestamp 1604489732
transform 1 0 2522 0 1 124370
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_224_38
timestamp 1604489732
transform 1 0 3534 0 -1 124370
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_224_32
timestamp 1604489732
transform 1 0 2982 0 -1 124370
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_224_27
timestamp 1604489732
transform 1 0 2522 0 -1 124370
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1475
timestamp 1604489732
transform 1 0 2890 0 -1 124370
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_449
timestamp 1604489732
transform -1 0 3902 0 1 124370
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_447
timestamp 1604489732
transform -1 0 3902 0 -1 124370
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_226_38
timestamp 1604489732
transform 1 0 3534 0 -1 125458
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_226_32
timestamp 1604489732
transform 1 0 2982 0 -1 125458
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_226_27
timestamp 1604489732
transform 1 0 2522 0 -1 125458
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1476
timestamp 1604489732
transform 1 0 2890 0 -1 125458
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_451
timestamp 1604489732
transform -1 0 3902 0 -1 125458
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_227_27
timestamp 1604489732
transform 1 0 2522 0 1 125458
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_453
timestamp 1604489732
transform -1 0 3902 0 1 125458
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1130
timestamp 1604489732
transform 1 0 83298 0 -1 124370
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1132
timestamp 1604489732
transform 1 0 83298 0 1 124370
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1134
timestamp 1604489732
transform 1 0 83298 0 -1 125458
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1136
timestamp 1604489732
transform 1 0 83298 0 1 125458
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_224_908
timestamp 1604489732
transform 1 0 83574 0 -1 124370
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_225_908
timestamp 1604489732
transform 1 0 83574 0 1 124370
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_226_908
timestamp 1604489732
transform 1 0 83574 0 -1 125458
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_227_908
timestamp 1604489732
transform 1 0 83574 0 1 125458
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_225_932
timestamp 1604489732
transform 1 0 85782 0 1 124370
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_225_920
timestamp 1604489732
transform 1 0 84678 0 1 124370
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_224_937
timestamp 1604489732
transform 1 0 86242 0 -1 124370
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_224_932
timestamp 1604489732
transform 1 0 85782 0 -1 124370
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_224_920
timestamp 1604489732
transform 1 0 84678 0 -1 124370
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1647
timestamp 1604489732
transform 1 0 86150 0 -1 124370
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_226_937
timestamp 1604489732
transform 1 0 86242 0 -1 125458
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_226_932
timestamp 1604489732
transform 1 0 85782 0 -1 125458
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_226_920
timestamp 1604489732
transform 1 0 84678 0 -1 125458
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1648
timestamp 1604489732
transform 1 0 86150 0 -1 125458
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_227_932
timestamp 1604489732
transform 1 0 85782 0 1 125458
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_227_920
timestamp 1604489732
transform 1 0 84678 0 1 125458
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_225_944
timestamp 1604489732
transform 1 0 86886 0 1 124370
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_225_950
timestamp 1604489732
transform 1 0 87438 0 1 124370
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_224_949
timestamp 1604489732
transform 1 0 87346 0 -1 124370
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1133
timestamp 1604489732
transform -1 0 87806 0 1 124370
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1131
timestamp 1604489732
transform -1 0 87806 0 -1 124370
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_226_949
timestamp 1604489732
transform 1 0 87346 0 -1 125458
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1135
timestamp 1604489732
transform -1 0 87806 0 -1 125458
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_227_944
timestamp 1604489732
transform 1 0 86886 0 1 125458
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_227_950
timestamp 1604489732
transform 1 0 87438 0 1 125458
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1137
timestamp 1604489732
transform -1 0 87806 0 1 125458
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_454
timestamp 1604489732
transform 1 0 38 0 -1 126546
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_456
timestamp 1604489732
transform 1 0 38 0 1 126546
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_458
timestamp 1604489732
transform 1 0 38 0 -1 127634
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_228_3
timestamp 1604489732
transform 1 0 314 0 -1 126546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_228_15
timestamp 1604489732
transform 1 0 1418 0 -1 126546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_229_3
timestamp 1604489732
transform 1 0 314 0 1 126546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_229_15
timestamp 1604489732
transform 1 0 1418 0 1 126546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_230_3
timestamp 1604489732
transform 1 0 314 0 -1 127634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_230_15
timestamp 1604489732
transform 1 0 1418 0 -1 127634
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_228_38
timestamp 1604489732
transform 1 0 3534 0 -1 126546
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_228_32
timestamp 1604489732
transform 1 0 2982 0 -1 126546
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_228_27
timestamp 1604489732
transform 1 0 2522 0 -1 126546
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1477
timestamp 1604489732
transform 1 0 2890 0 -1 126546
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_455
timestamp 1604489732
transform -1 0 3902 0 -1 126546
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_229_27
timestamp 1604489732
transform 1 0 2522 0 1 126546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_457
timestamp 1604489732
transform -1 0 3902 0 1 126546
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_230_38
timestamp 1604489732
transform 1 0 3534 0 -1 127634
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_230_32
timestamp 1604489732
transform 1 0 2982 0 -1 127634
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_230_27
timestamp 1604489732
transform 1 0 2522 0 -1 127634
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1478
timestamp 1604489732
transform 1 0 2890 0 -1 127634
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_459
timestamp 1604489732
transform -1 0 3902 0 -1 127634
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1138
timestamp 1604489732
transform 1 0 83298 0 -1 126546
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1140
timestamp 1604489732
transform 1 0 83298 0 1 126546
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1142
timestamp 1604489732
transform 1 0 83298 0 -1 127634
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_228_908
timestamp 1604489732
transform 1 0 83574 0 -1 126546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_229_908
timestamp 1604489732
transform 1 0 83574 0 1 126546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_230_908
timestamp 1604489732
transform 1 0 83574 0 -1 127634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_228_937
timestamp 1604489732
transform 1 0 86242 0 -1 126546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_228_932
timestamp 1604489732
transform 1 0 85782 0 -1 126546
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_228_920
timestamp 1604489732
transform 1 0 84678 0 -1 126546
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1649
timestamp 1604489732
transform 1 0 86150 0 -1 126546
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_229_932
timestamp 1604489732
transform 1 0 85782 0 1 126546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_229_920
timestamp 1604489732
transform 1 0 84678 0 1 126546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_230_937
timestamp 1604489732
transform 1 0 86242 0 -1 127634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_230_932
timestamp 1604489732
transform 1 0 85782 0 -1 127634
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_230_920
timestamp 1604489732
transform 1 0 84678 0 -1 127634
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1650
timestamp 1604489732
transform 1 0 86150 0 -1 127634
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1139
timestamp 1604489732
transform -1 0 87806 0 -1 126546
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1141
timestamp 1604489732
transform -1 0 87806 0 1 126546
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1143
timestamp 1604489732
transform -1 0 87806 0 -1 127634
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_228_949
timestamp 1604489732
transform 1 0 87346 0 -1 126546
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_229_944
timestamp 1604489732
transform 1 0 86886 0 1 126546
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_229_950
timestamp 1604489732
transform 1 0 87438 0 1 126546
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_230_949
timestamp 1604489732
transform 1 0 87346 0 -1 127634
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_460
timestamp 1604489732
transform 1 0 38 0 1 127634
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_462
timestamp 1604489732
transform 1 0 38 0 -1 128722
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_464
timestamp 1604489732
transform 1 0 38 0 1 128722
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_231_3
timestamp 1604489732
transform 1 0 314 0 1 127634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_231_15
timestamp 1604489732
transform 1 0 1418 0 1 127634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_232_3
timestamp 1604489732
transform 1 0 314 0 -1 128722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_232_15
timestamp 1604489732
transform 1 0 1418 0 -1 128722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_233_3
timestamp 1604489732
transform 1 0 314 0 1 128722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_233_15
timestamp 1604489732
transform 1 0 1418 0 1 128722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_461
timestamp 1604489732
transform -1 0 3902 0 1 127634
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_463
timestamp 1604489732
transform -1 0 3902 0 -1 128722
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_465
timestamp 1604489732
transform -1 0 3902 0 1 128722
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1479
timestamp 1604489732
transform 1 0 2890 0 -1 128722
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_231_27
timestamp 1604489732
transform 1 0 2522 0 1 127634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_232_27
timestamp 1604489732
transform 1 0 2522 0 -1 128722
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_232_32
timestamp 1604489732
transform 1 0 2982 0 -1 128722
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_232_38
timestamp 1604489732
transform 1 0 3534 0 -1 128722
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_233_27
timestamp 1604489732
transform 1 0 2522 0 1 128722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1144
timestamp 1604489732
transform 1 0 83298 0 1 127634
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1146
timestamp 1604489732
transform 1 0 83298 0 -1 128722
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1148
timestamp 1604489732
transform 1 0 83298 0 1 128722
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_231_908
timestamp 1604489732
transform 1 0 83574 0 1 127634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_232_908
timestamp 1604489732
transform 1 0 83574 0 -1 128722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_233_908
timestamp 1604489732
transform 1 0 83574 0 1 128722
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1651
timestamp 1604489732
transform 1 0 86150 0 -1 128722
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_231_920
timestamp 1604489732
transform 1 0 84678 0 1 127634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_231_932
timestamp 1604489732
transform 1 0 85782 0 1 127634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_232_920
timestamp 1604489732
transform 1 0 84678 0 -1 128722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_232_932
timestamp 1604489732
transform 1 0 85782 0 -1 128722
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_232_937
timestamp 1604489732
transform 1 0 86242 0 -1 128722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_233_920
timestamp 1604489732
transform 1 0 84678 0 1 128722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_233_932
timestamp 1604489732
transform 1 0 85782 0 1 128722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1145
timestamp 1604489732
transform -1 0 87806 0 1 127634
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1147
timestamp 1604489732
transform -1 0 87806 0 -1 128722
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1149
timestamp 1604489732
transform -1 0 87806 0 1 128722
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_231_944
timestamp 1604489732
transform 1 0 86886 0 1 127634
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_231_950
timestamp 1604489732
transform 1 0 87438 0 1 127634
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_232_949
timestamp 1604489732
transform 1 0 87346 0 -1 128722
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_233_944
timestamp 1604489732
transform 1 0 86886 0 1 128722
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_233_950
timestamp 1604489732
transform 1 0 87438 0 1 128722
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_235_15
timestamp 1604489732
transform 1 0 1418 0 1 129810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_235_3
timestamp 1604489732
transform 1 0 314 0 1 129810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_234_15
timestamp 1604489732
transform 1 0 1418 0 -1 129810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_234_3
timestamp 1604489732
transform 1 0 314 0 -1 129810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_468
timestamp 1604489732
transform 1 0 38 0 1 129810
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_466
timestamp 1604489732
transform 1 0 38 0 -1 129810
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_236_15
timestamp 1604489732
transform 1 0 1418 0 -1 130898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_236_3
timestamp 1604489732
transform 1 0 314 0 -1 130898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_470
timestamp 1604489732
transform 1 0 38 0 -1 130898
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_237_15
timestamp 1604489732
transform 1 0 1418 0 1 130898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_237_3
timestamp 1604489732
transform 1 0 314 0 1 130898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_472
timestamp 1604489732
transform 1 0 38 0 1 130898
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_235_27
timestamp 1604489732
transform 1 0 2522 0 1 129810
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_234_38
timestamp 1604489732
transform 1 0 3534 0 -1 129810
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_234_32
timestamp 1604489732
transform 1 0 2982 0 -1 129810
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_234_27
timestamp 1604489732
transform 1 0 2522 0 -1 129810
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1480
timestamp 1604489732
transform 1 0 2890 0 -1 129810
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_469
timestamp 1604489732
transform -1 0 3902 0 1 129810
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_467
timestamp 1604489732
transform -1 0 3902 0 -1 129810
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_236_38
timestamp 1604489732
transform 1 0 3534 0 -1 130898
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_236_32
timestamp 1604489732
transform 1 0 2982 0 -1 130898
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_236_27
timestamp 1604489732
transform 1 0 2522 0 -1 130898
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1481
timestamp 1604489732
transform 1 0 2890 0 -1 130898
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_471
timestamp 1604489732
transform -1 0 3902 0 -1 130898
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_237_27
timestamp 1604489732
transform 1 0 2522 0 1 130898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_473
timestamp 1604489732
transform -1 0 3902 0 1 130898
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1150
timestamp 1604489732
transform 1 0 83298 0 -1 129810
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1152
timestamp 1604489732
transform 1 0 83298 0 1 129810
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1154
timestamp 1604489732
transform 1 0 83298 0 -1 130898
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1156
timestamp 1604489732
transform 1 0 83298 0 1 130898
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_234_908
timestamp 1604489732
transform 1 0 83574 0 -1 129810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_235_908
timestamp 1604489732
transform 1 0 83574 0 1 129810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_236_908
timestamp 1604489732
transform 1 0 83574 0 -1 130898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_237_908
timestamp 1604489732
transform 1 0 83574 0 1 130898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_235_932
timestamp 1604489732
transform 1 0 85782 0 1 129810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_235_920
timestamp 1604489732
transform 1 0 84678 0 1 129810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_234_937
timestamp 1604489732
transform 1 0 86242 0 -1 129810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_234_932
timestamp 1604489732
transform 1 0 85782 0 -1 129810
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_234_920
timestamp 1604489732
transform 1 0 84678 0 -1 129810
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1652
timestamp 1604489732
transform 1 0 86150 0 -1 129810
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_236_937
timestamp 1604489732
transform 1 0 86242 0 -1 130898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_236_932
timestamp 1604489732
transform 1 0 85782 0 -1 130898
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_236_920
timestamp 1604489732
transform 1 0 84678 0 -1 130898
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1653
timestamp 1604489732
transform 1 0 86150 0 -1 130898
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_237_932
timestamp 1604489732
transform 1 0 85782 0 1 130898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_237_920
timestamp 1604489732
transform 1 0 84678 0 1 130898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_235_944
timestamp 1604489732
transform 1 0 86886 0 1 129810
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_235_950
timestamp 1604489732
transform 1 0 87438 0 1 129810
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_234_949
timestamp 1604489732
transform 1 0 87346 0 -1 129810
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1153
timestamp 1604489732
transform -1 0 87806 0 1 129810
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1151
timestamp 1604489732
transform -1 0 87806 0 -1 129810
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_236_949
timestamp 1604489732
transform 1 0 87346 0 -1 130898
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1155
timestamp 1604489732
transform -1 0 87806 0 -1 130898
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_237_944
timestamp 1604489732
transform 1 0 86886 0 1 130898
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_237_950
timestamp 1604489732
transform 1 0 87438 0 1 130898
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1157
timestamp 1604489732
transform -1 0 87806 0 1 130898
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_474
timestamp 1604489732
transform 1 0 38 0 -1 131986
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_476
timestamp 1604489732
transform 1 0 38 0 1 131986
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_478
timestamp 1604489732
transform 1 0 38 0 -1 133074
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_238_3
timestamp 1604489732
transform 1 0 314 0 -1 131986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_238_15
timestamp 1604489732
transform 1 0 1418 0 -1 131986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_239_3
timestamp 1604489732
transform 1 0 314 0 1 131986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_239_15
timestamp 1604489732
transform 1 0 1418 0 1 131986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_240_3
timestamp 1604489732
transform 1 0 314 0 -1 133074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_240_15
timestamp 1604489732
transform 1 0 1418 0 -1 133074
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_238_38
timestamp 1604489732
transform 1 0 3534 0 -1 131986
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_238_32
timestamp 1604489732
transform 1 0 2982 0 -1 131986
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_238_27
timestamp 1604489732
transform 1 0 2522 0 -1 131986
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1482
timestamp 1604489732
transform 1 0 2890 0 -1 131986
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_475
timestamp 1604489732
transform -1 0 3902 0 -1 131986
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_239_27
timestamp 1604489732
transform 1 0 2522 0 1 131986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_477
timestamp 1604489732
transform -1 0 3902 0 1 131986
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_240_38
timestamp 1604489732
transform 1 0 3534 0 -1 133074
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_240_32
timestamp 1604489732
transform 1 0 2982 0 -1 133074
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_240_27
timestamp 1604489732
transform 1 0 2522 0 -1 133074
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1483
timestamp 1604489732
transform 1 0 2890 0 -1 133074
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_479
timestamp 1604489732
transform -1 0 3902 0 -1 133074
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1158
timestamp 1604489732
transform 1 0 83298 0 -1 131986
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1160
timestamp 1604489732
transform 1 0 83298 0 1 131986
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1162
timestamp 1604489732
transform 1 0 83298 0 -1 133074
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_238_908
timestamp 1604489732
transform 1 0 83574 0 -1 131986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_239_908
timestamp 1604489732
transform 1 0 83574 0 1 131986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_240_908
timestamp 1604489732
transform 1 0 83574 0 -1 133074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_238_937
timestamp 1604489732
transform 1 0 86242 0 -1 131986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_238_932
timestamp 1604489732
transform 1 0 85782 0 -1 131986
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_238_920
timestamp 1604489732
transform 1 0 84678 0 -1 131986
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1654
timestamp 1604489732
transform 1 0 86150 0 -1 131986
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_239_932
timestamp 1604489732
transform 1 0 85782 0 1 131986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_239_920
timestamp 1604489732
transform 1 0 84678 0 1 131986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_240_937
timestamp 1604489732
transform 1 0 86242 0 -1 133074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_240_932
timestamp 1604489732
transform 1 0 85782 0 -1 133074
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_240_920
timestamp 1604489732
transform 1 0 84678 0 -1 133074
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1655
timestamp 1604489732
transform 1 0 86150 0 -1 133074
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1159
timestamp 1604489732
transform -1 0 87806 0 -1 131986
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1161
timestamp 1604489732
transform -1 0 87806 0 1 131986
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1163
timestamp 1604489732
transform -1 0 87806 0 -1 133074
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_238_949
timestamp 1604489732
transform 1 0 87346 0 -1 131986
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_239_944
timestamp 1604489732
transform 1 0 86886 0 1 131986
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_239_950
timestamp 1604489732
transform 1 0 87438 0 1 131986
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_240_949
timestamp 1604489732
transform 1 0 87346 0 -1 133074
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_480
timestamp 1604489732
transform 1 0 38 0 1 133074
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_482
timestamp 1604489732
transform 1 0 38 0 -1 134162
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_484
timestamp 1604489732
transform 1 0 38 0 1 134162
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_241_3
timestamp 1604489732
transform 1 0 314 0 1 133074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_241_15
timestamp 1604489732
transform 1 0 1418 0 1 133074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_242_3
timestamp 1604489732
transform 1 0 314 0 -1 134162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_242_15
timestamp 1604489732
transform 1 0 1418 0 -1 134162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_243_3
timestamp 1604489732
transform 1 0 314 0 1 134162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_243_15
timestamp 1604489732
transform 1 0 1418 0 1 134162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_481
timestamp 1604489732
transform -1 0 3902 0 1 133074
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_483
timestamp 1604489732
transform -1 0 3902 0 -1 134162
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_485
timestamp 1604489732
transform -1 0 3902 0 1 134162
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1484
timestamp 1604489732
transform 1 0 2890 0 -1 134162
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_241_27
timestamp 1604489732
transform 1 0 2522 0 1 133074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_242_27
timestamp 1604489732
transform 1 0 2522 0 -1 134162
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_242_32
timestamp 1604489732
transform 1 0 2982 0 -1 134162
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_242_38
timestamp 1604489732
transform 1 0 3534 0 -1 134162
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_243_27
timestamp 1604489732
transform 1 0 2522 0 1 134162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1164
timestamp 1604489732
transform 1 0 83298 0 1 133074
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1166
timestamp 1604489732
transform 1 0 83298 0 -1 134162
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1168
timestamp 1604489732
transform 1 0 83298 0 1 134162
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_241_908
timestamp 1604489732
transform 1 0 83574 0 1 133074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_242_908
timestamp 1604489732
transform 1 0 83574 0 -1 134162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_243_908
timestamp 1604489732
transform 1 0 83574 0 1 134162
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1656
timestamp 1604489732
transform 1 0 86150 0 -1 134162
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_241_920
timestamp 1604489732
transform 1 0 84678 0 1 133074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_241_932
timestamp 1604489732
transform 1 0 85782 0 1 133074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_242_920
timestamp 1604489732
transform 1 0 84678 0 -1 134162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_242_932
timestamp 1604489732
transform 1 0 85782 0 -1 134162
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_242_937
timestamp 1604489732
transform 1 0 86242 0 -1 134162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_243_920
timestamp 1604489732
transform 1 0 84678 0 1 134162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_243_932
timestamp 1604489732
transform 1 0 85782 0 1 134162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1165
timestamp 1604489732
transform -1 0 87806 0 1 133074
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1167
timestamp 1604489732
transform -1 0 87806 0 -1 134162
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1169
timestamp 1604489732
transform -1 0 87806 0 1 134162
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_241_944
timestamp 1604489732
transform 1 0 86886 0 1 133074
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_241_950
timestamp 1604489732
transform 1 0 87438 0 1 133074
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_242_949
timestamp 1604489732
transform 1 0 87346 0 -1 134162
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_243_944
timestamp 1604489732
transform 1 0 86886 0 1 134162
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_243_950
timestamp 1604489732
transform 1 0 87438 0 1 134162
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_245_15
timestamp 1604489732
transform 1 0 1418 0 1 135250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_245_3
timestamp 1604489732
transform 1 0 314 0 1 135250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_244_15
timestamp 1604489732
transform 1 0 1418 0 -1 135250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_244_3
timestamp 1604489732
transform 1 0 314 0 -1 135250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_488
timestamp 1604489732
transform 1 0 38 0 1 135250
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_486
timestamp 1604489732
transform 1 0 38 0 -1 135250
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_246_15
timestamp 1604489732
transform 1 0 1418 0 -1 136338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_246_3
timestamp 1604489732
transform 1 0 314 0 -1 136338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_490
timestamp 1604489732
transform 1 0 38 0 -1 136338
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_247_15
timestamp 1604489732
transform 1 0 1418 0 1 136338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_247_3
timestamp 1604489732
transform 1 0 314 0 1 136338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_492
timestamp 1604489732
transform 1 0 38 0 1 136338
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_245_27
timestamp 1604489732
transform 1 0 2522 0 1 135250
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_244_38
timestamp 1604489732
transform 1 0 3534 0 -1 135250
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_244_32
timestamp 1604489732
transform 1 0 2982 0 -1 135250
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_244_27
timestamp 1604489732
transform 1 0 2522 0 -1 135250
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1485
timestamp 1604489732
transform 1 0 2890 0 -1 135250
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_489
timestamp 1604489732
transform -1 0 3902 0 1 135250
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_487
timestamp 1604489732
transform -1 0 3902 0 -1 135250
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_246_38
timestamp 1604489732
transform 1 0 3534 0 -1 136338
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_246_32
timestamp 1604489732
transform 1 0 2982 0 -1 136338
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_246_27
timestamp 1604489732
transform 1 0 2522 0 -1 136338
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1486
timestamp 1604489732
transform 1 0 2890 0 -1 136338
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_491
timestamp 1604489732
transform -1 0 3902 0 -1 136338
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_247_27
timestamp 1604489732
transform 1 0 2522 0 1 136338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_493
timestamp 1604489732
transform -1 0 3902 0 1 136338
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1170
timestamp 1604489732
transform 1 0 83298 0 -1 135250
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1172
timestamp 1604489732
transform 1 0 83298 0 1 135250
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1174
timestamp 1604489732
transform 1 0 83298 0 -1 136338
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1176
timestamp 1604489732
transform 1 0 83298 0 1 136338
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_244_908
timestamp 1604489732
transform 1 0 83574 0 -1 135250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_245_908
timestamp 1604489732
transform 1 0 83574 0 1 135250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_246_908
timestamp 1604489732
transform 1 0 83574 0 -1 136338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_247_908
timestamp 1604489732
transform 1 0 83574 0 1 136338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_245_932
timestamp 1604489732
transform 1 0 85782 0 1 135250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_245_920
timestamp 1604489732
transform 1 0 84678 0 1 135250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_244_937
timestamp 1604489732
transform 1 0 86242 0 -1 135250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_244_932
timestamp 1604489732
transform 1 0 85782 0 -1 135250
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_244_920
timestamp 1604489732
transform 1 0 84678 0 -1 135250
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1657
timestamp 1604489732
transform 1 0 86150 0 -1 135250
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_246_937
timestamp 1604489732
transform 1 0 86242 0 -1 136338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_246_932
timestamp 1604489732
transform 1 0 85782 0 -1 136338
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_246_920
timestamp 1604489732
transform 1 0 84678 0 -1 136338
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1658
timestamp 1604489732
transform 1 0 86150 0 -1 136338
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_247_932
timestamp 1604489732
transform 1 0 85782 0 1 136338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_247_920
timestamp 1604489732
transform 1 0 84678 0 1 136338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_245_944
timestamp 1604489732
transform 1 0 86886 0 1 135250
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_245_950
timestamp 1604489732
transform 1 0 87438 0 1 135250
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_244_949
timestamp 1604489732
transform 1 0 87346 0 -1 135250
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1173
timestamp 1604489732
transform -1 0 87806 0 1 135250
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1171
timestamp 1604489732
transform -1 0 87806 0 -1 135250
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_246_949
timestamp 1604489732
transform 1 0 87346 0 -1 136338
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1175
timestamp 1604489732
transform -1 0 87806 0 -1 136338
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_247_944
timestamp 1604489732
transform 1 0 86886 0 1 136338
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_950
timestamp 1604489732
transform 1 0 87438 0 1 136338
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1177
timestamp 1604489732
transform -1 0 87806 0 1 136338
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_494
timestamp 1604489732
transform 1 0 38 0 -1 137426
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_496
timestamp 1604489732
transform 1 0 38 0 1 137426
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_498
timestamp 1604489732
transform 1 0 38 0 -1 138514
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_248_3
timestamp 1604489732
transform 1 0 314 0 -1 137426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_248_15
timestamp 1604489732
transform 1 0 1418 0 -1 137426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_249_3
timestamp 1604489732
transform 1 0 314 0 1 137426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_249_15
timestamp 1604489732
transform 1 0 1418 0 1 137426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_250_3
timestamp 1604489732
transform 1 0 314 0 -1 138514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_250_15
timestamp 1604489732
transform 1 0 1418 0 -1 138514
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_248_38
timestamp 1604489732
transform 1 0 3534 0 -1 137426
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_248_32
timestamp 1604489732
transform 1 0 2982 0 -1 137426
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_248_27
timestamp 1604489732
transform 1 0 2522 0 -1 137426
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1487
timestamp 1604489732
transform 1 0 2890 0 -1 137426
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_495
timestamp 1604489732
transform -1 0 3902 0 -1 137426
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_249_27
timestamp 1604489732
transform 1 0 2522 0 1 137426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_497
timestamp 1604489732
transform -1 0 3902 0 1 137426
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_250_38
timestamp 1604489732
transform 1 0 3534 0 -1 138514
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_250_32
timestamp 1604489732
transform 1 0 2982 0 -1 138514
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_250_27
timestamp 1604489732
transform 1 0 2522 0 -1 138514
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1488
timestamp 1604489732
transform 1 0 2890 0 -1 138514
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_499
timestamp 1604489732
transform -1 0 3902 0 -1 138514
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1178
timestamp 1604489732
transform 1 0 83298 0 -1 137426
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1180
timestamp 1604489732
transform 1 0 83298 0 1 137426
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1182
timestamp 1604489732
transform 1 0 83298 0 -1 138514
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_248_908
timestamp 1604489732
transform 1 0 83574 0 -1 137426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_249_908
timestamp 1604489732
transform 1 0 83574 0 1 137426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_250_908
timestamp 1604489732
transform 1 0 83574 0 -1 138514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_248_937
timestamp 1604489732
transform 1 0 86242 0 -1 137426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_248_932
timestamp 1604489732
transform 1 0 85782 0 -1 137426
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_248_920
timestamp 1604489732
transform 1 0 84678 0 -1 137426
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1659
timestamp 1604489732
transform 1 0 86150 0 -1 137426
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_249_932
timestamp 1604489732
transform 1 0 85782 0 1 137426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_249_920
timestamp 1604489732
transform 1 0 84678 0 1 137426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_250_937
timestamp 1604489732
transform 1 0 86242 0 -1 138514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_250_932
timestamp 1604489732
transform 1 0 85782 0 -1 138514
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_250_920
timestamp 1604489732
transform 1 0 84678 0 -1 138514
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1660
timestamp 1604489732
transform 1 0 86150 0 -1 138514
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1179
timestamp 1604489732
transform -1 0 87806 0 -1 137426
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1181
timestamp 1604489732
transform -1 0 87806 0 1 137426
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1183
timestamp 1604489732
transform -1 0 87806 0 -1 138514
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_248_949
timestamp 1604489732
transform 1 0 87346 0 -1 137426
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_249_944
timestamp 1604489732
transform 1 0 86886 0 1 137426
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_950
timestamp 1604489732
transform 1 0 87438 0 1 137426
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_250_949
timestamp 1604489732
transform 1 0 87346 0 -1 138514
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_500
timestamp 1604489732
transform 1 0 38 0 1 138514
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_251_3
timestamp 1604489732
transform 1 0 314 0 1 138514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_251_15
timestamp 1604489732
transform 1 0 1418 0 1 138514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_501
timestamp 1604489732
transform -1 0 3902 0 1 138514
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_251_27
timestamp 1604489732
transform 1 0 2522 0 1 138514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1184
timestamp 1604489732
transform 1 0 83298 0 1 138514
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_251_908
timestamp 1604489732
transform 1 0 83574 0 1 138514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_251_920
timestamp 1604489732
transform 1 0 84678 0 1 138514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_251_932
timestamp 1604489732
transform 1 0 85782 0 1 138514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1185
timestamp 1604489732
transform -1 0 87806 0 1 138514
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_251_944
timestamp 1604489732
transform 1 0 86886 0 1 138514
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_950
timestamp 1604489732
transform 1 0 87438 0 1 138514
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_502
timestamp 1604489732
transform 1 0 38 0 -1 139602
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_504
timestamp 1604489732
transform 1 0 38 0 1 139602
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_506
timestamp 1604489732
transform 1 0 38 0 -1 140690
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_252_3
timestamp 1604489732
transform 1 0 314 0 -1 139602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_252_15
timestamp 1604489732
transform 1 0 1418 0 -1 139602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_253_3
timestamp 1604489732
transform 1 0 314 0 1 139602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_253_15
timestamp 1604489732
transform 1 0 1418 0 1 139602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_254_3
timestamp 1604489732
transform 1 0 314 0 -1 140690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_254_15
timestamp 1604489732
transform 1 0 1418 0 -1 140690
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_252_38
timestamp 1604489732
transform 1 0 3534 0 -1 139602
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_252_32
timestamp 1604489732
transform 1 0 2982 0 -1 139602
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_252_27
timestamp 1604489732
transform 1 0 2522 0 -1 139602
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1489
timestamp 1604489732
transform 1 0 2890 0 -1 139602
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_503
timestamp 1604489732
transform -1 0 3902 0 -1 139602
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_253_27
timestamp 1604489732
transform 1 0 2522 0 1 139602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_505
timestamp 1604489732
transform -1 0 3902 0 1 139602
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_254_38
timestamp 1604489732
transform 1 0 3534 0 -1 140690
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_254_32
timestamp 1604489732
transform 1 0 2982 0 -1 140690
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_254_27
timestamp 1604489732
transform 1 0 2522 0 -1 140690
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1490
timestamp 1604489732
transform 1 0 2890 0 -1 140690
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_507
timestamp 1604489732
transform -1 0 3902 0 -1 140690
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1186
timestamp 1604489732
transform 1 0 83298 0 -1 139602
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1188
timestamp 1604489732
transform 1 0 83298 0 1 139602
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1190
timestamp 1604489732
transform 1 0 83298 0 -1 140690
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_252_908
timestamp 1604489732
transform 1 0 83574 0 -1 139602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_253_908
timestamp 1604489732
transform 1 0 83574 0 1 139602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_254_908
timestamp 1604489732
transform 1 0 83574 0 -1 140690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_252_937
timestamp 1604489732
transform 1 0 86242 0 -1 139602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_252_932
timestamp 1604489732
transform 1 0 85782 0 -1 139602
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_252_920
timestamp 1604489732
transform 1 0 84678 0 -1 139602
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1661
timestamp 1604489732
transform 1 0 86150 0 -1 139602
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_253_932
timestamp 1604489732
transform 1 0 85782 0 1 139602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_253_920
timestamp 1604489732
transform 1 0 84678 0 1 139602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_254_937
timestamp 1604489732
transform 1 0 86242 0 -1 140690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_254_932
timestamp 1604489732
transform 1 0 85782 0 -1 140690
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_254_920
timestamp 1604489732
transform 1 0 84678 0 -1 140690
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1662
timestamp 1604489732
transform 1 0 86150 0 -1 140690
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1187
timestamp 1604489732
transform -1 0 87806 0 -1 139602
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1189
timestamp 1604489732
transform -1 0 87806 0 1 139602
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1191
timestamp 1604489732
transform -1 0 87806 0 -1 140690
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_252_949
timestamp 1604489732
transform 1 0 87346 0 -1 139602
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_253_944
timestamp 1604489732
transform 1 0 86886 0 1 139602
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_950
timestamp 1604489732
transform 1 0 87438 0 1 139602
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_254_949
timestamp 1604489732
transform 1 0 87346 0 -1 140690
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_256_15
timestamp 1604489732
transform 1 0 1418 0 -1 141778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_256_3
timestamp 1604489732
transform 1 0 314 0 -1 141778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_255_15
timestamp 1604489732
transform 1 0 1418 0 1 140690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_255_3
timestamp 1604489732
transform 1 0 314 0 1 140690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_510
timestamp 1604489732
transform 1 0 38 0 -1 141778
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_508
timestamp 1604489732
transform 1 0 38 0 1 140690
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_257_15
timestamp 1604489732
transform 1 0 1418 0 1 141778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_257_3
timestamp 1604489732
transform 1 0 314 0 1 141778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_512
timestamp 1604489732
transform 1 0 38 0 1 141778
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_258_15
timestamp 1604489732
transform 1 0 1418 0 -1 142866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_258_3
timestamp 1604489732
transform 1 0 314 0 -1 142866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_514
timestamp 1604489732
transform 1 0 38 0 -1 142866
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_256_38
timestamp 1604489732
transform 1 0 3534 0 -1 141778
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_256_32
timestamp 1604489732
transform 1 0 2982 0 -1 141778
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_256_27
timestamp 1604489732
transform 1 0 2522 0 -1 141778
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_255_27
timestamp 1604489732
transform 1 0 2522 0 1 140690
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1491
timestamp 1604489732
transform 1 0 2890 0 -1 141778
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_511
timestamp 1604489732
transform -1 0 3902 0 -1 141778
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_509
timestamp 1604489732
transform -1 0 3902 0 1 140690
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_257_27
timestamp 1604489732
transform 1 0 2522 0 1 141778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_513
timestamp 1604489732
transform -1 0 3902 0 1 141778
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_258_38
timestamp 1604489732
transform 1 0 3534 0 -1 142866
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_258_32
timestamp 1604489732
transform 1 0 2982 0 -1 142866
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_258_27
timestamp 1604489732
transform 1 0 2522 0 -1 142866
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1492
timestamp 1604489732
transform 1 0 2890 0 -1 142866
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_515
timestamp 1604489732
transform -1 0 3902 0 -1 142866
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1192
timestamp 1604489732
transform 1 0 83298 0 1 140690
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1194
timestamp 1604489732
transform 1 0 83298 0 -1 141778
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1196
timestamp 1604489732
transform 1 0 83298 0 1 141778
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1198
timestamp 1604489732
transform 1 0 83298 0 -1 142866
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_255_908
timestamp 1604489732
transform 1 0 83574 0 1 140690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_256_908
timestamp 1604489732
transform 1 0 83574 0 -1 141778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_257_908
timestamp 1604489732
transform 1 0 83574 0 1 141778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_258_908
timestamp 1604489732
transform 1 0 83574 0 -1 142866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_256_937
timestamp 1604489732
transform 1 0 86242 0 -1 141778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_256_932
timestamp 1604489732
transform 1 0 85782 0 -1 141778
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_256_920
timestamp 1604489732
transform 1 0 84678 0 -1 141778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_255_932
timestamp 1604489732
transform 1 0 85782 0 1 140690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_255_920
timestamp 1604489732
transform 1 0 84678 0 1 140690
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1663
timestamp 1604489732
transform 1 0 86150 0 -1 141778
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_257_932
timestamp 1604489732
transform 1 0 85782 0 1 141778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_257_920
timestamp 1604489732
transform 1 0 84678 0 1 141778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_258_937
timestamp 1604489732
transform 1 0 86242 0 -1 142866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_258_932
timestamp 1604489732
transform 1 0 85782 0 -1 142866
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_258_920
timestamp 1604489732
transform 1 0 84678 0 -1 142866
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1664
timestamp 1604489732
transform 1 0 86150 0 -1 142866
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_255_944
timestamp 1604489732
transform 1 0 86886 0 1 140690
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_256_949
timestamp 1604489732
transform 1 0 87346 0 -1 141778
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_255_950
timestamp 1604489732
transform 1 0 87438 0 1 140690
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1195
timestamp 1604489732
transform -1 0 87806 0 -1 141778
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1193
timestamp 1604489732
transform -1 0 87806 0 1 140690
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_257_944
timestamp 1604489732
transform 1 0 86886 0 1 141778
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_950
timestamp 1604489732
transform 1 0 87438 0 1 141778
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1197
timestamp 1604489732
transform -1 0 87806 0 1 141778
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_258_949
timestamp 1604489732
transform 1 0 87346 0 -1 142866
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1199
timestamp 1604489732
transform -1 0 87806 0 -1 142866
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_516
timestamp 1604489732
transform 1 0 38 0 1 142866
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_518
timestamp 1604489732
transform 1 0 38 0 -1 143954
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_520
timestamp 1604489732
transform 1 0 38 0 1 143954
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_259_3
timestamp 1604489732
transform 1 0 314 0 1 142866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_259_15
timestamp 1604489732
transform 1 0 1418 0 1 142866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_260_3
timestamp 1604489732
transform 1 0 314 0 -1 143954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_260_15
timestamp 1604489732
transform 1 0 1418 0 -1 143954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_261_3
timestamp 1604489732
transform 1 0 314 0 1 143954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_261_15
timestamp 1604489732
transform 1 0 1418 0 1 143954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_517
timestamp 1604489732
transform -1 0 3902 0 1 142866
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_519
timestamp 1604489732
transform -1 0 3902 0 -1 143954
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_521
timestamp 1604489732
transform -1 0 3902 0 1 143954
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1493
timestamp 1604489732
transform 1 0 2890 0 -1 143954
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_259_27
timestamp 1604489732
transform 1 0 2522 0 1 142866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_260_27
timestamp 1604489732
transform 1 0 2522 0 -1 143954
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_260_32
timestamp 1604489732
transform 1 0 2982 0 -1 143954
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_38
timestamp 1604489732
transform 1 0 3534 0 -1 143954
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_261_27
timestamp 1604489732
transform 1 0 2522 0 1 143954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1200
timestamp 1604489732
transform 1 0 83298 0 1 142866
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1202
timestamp 1604489732
transform 1 0 83298 0 -1 143954
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1204
timestamp 1604489732
transform 1 0 83298 0 1 143954
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_259_908
timestamp 1604489732
transform 1 0 83574 0 1 142866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_260_908
timestamp 1604489732
transform 1 0 83574 0 -1 143954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_261_908
timestamp 1604489732
transform 1 0 83574 0 1 143954
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1665
timestamp 1604489732
transform 1 0 86150 0 -1 143954
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_259_920
timestamp 1604489732
transform 1 0 84678 0 1 142866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_259_932
timestamp 1604489732
transform 1 0 85782 0 1 142866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_260_920
timestamp 1604489732
transform 1 0 84678 0 -1 143954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_260_932
timestamp 1604489732
transform 1 0 85782 0 -1 143954
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_260_937
timestamp 1604489732
transform 1 0 86242 0 -1 143954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_261_920
timestamp 1604489732
transform 1 0 84678 0 1 143954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_261_932
timestamp 1604489732
transform 1 0 85782 0 1 143954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1201
timestamp 1604489732
transform -1 0 87806 0 1 142866
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1203
timestamp 1604489732
transform -1 0 87806 0 -1 143954
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1205
timestamp 1604489732
transform -1 0 87806 0 1 143954
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_259_944
timestamp 1604489732
transform 1 0 86886 0 1 142866
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_950
timestamp 1604489732
transform 1 0 87438 0 1 142866
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_260_949
timestamp 1604489732
transform 1 0 87346 0 -1 143954
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_261_944
timestamp 1604489732
transform 1 0 86886 0 1 143954
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_950
timestamp 1604489732
transform 1 0 87438 0 1 143954
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_262_15
timestamp 1604489732
transform 1 0 1418 0 -1 145042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_262_3
timestamp 1604489732
transform 1 0 314 0 -1 145042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_522
timestamp 1604489732
transform 1 0 38 0 -1 145042
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_264_15
timestamp 1604489732
transform 1 0 1418 0 -1 146130
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_264_3
timestamp 1604489732
transform 1 0 314 0 -1 146130
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_263_15
timestamp 1604489732
transform 1 0 1418 0 1 145042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_263_3
timestamp 1604489732
transform 1 0 314 0 1 145042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_526
timestamp 1604489732
transform 1 0 38 0 -1 146130
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_524
timestamp 1604489732
transform 1 0 38 0 1 145042
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_265_15
timestamp 1604489732
transform 1 0 1418 0 1 146130
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_265_3
timestamp 1604489732
transform 1 0 314 0 1 146130
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_528
timestamp 1604489732
transform 1 0 38 0 1 146130
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_262_38
timestamp 1604489732
transform 1 0 3534 0 -1 145042
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_262_32
timestamp 1604489732
transform 1 0 2982 0 -1 145042
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_262_27
timestamp 1604489732
transform 1 0 2522 0 -1 145042
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1494
timestamp 1604489732
transform 1 0 2890 0 -1 145042
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_523
timestamp 1604489732
transform -1 0 3902 0 -1 145042
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_264_38
timestamp 1604489732
transform 1 0 3534 0 -1 146130
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_264_32
timestamp 1604489732
transform 1 0 2982 0 -1 146130
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_264_27
timestamp 1604489732
transform 1 0 2522 0 -1 146130
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_263_27
timestamp 1604489732
transform 1 0 2522 0 1 145042
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1495
timestamp 1604489732
transform 1 0 2890 0 -1 146130
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_527
timestamp 1604489732
transform -1 0 3902 0 -1 146130
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_525
timestamp 1604489732
transform -1 0 3902 0 1 145042
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_265_27
timestamp 1604489732
transform 1 0 2522 0 1 146130
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_529
timestamp 1604489732
transform -1 0 3902 0 1 146130
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1206
timestamp 1604489732
transform 1 0 83298 0 -1 145042
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1208
timestamp 1604489732
transform 1 0 83298 0 1 145042
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1210
timestamp 1604489732
transform 1 0 83298 0 -1 146130
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1212
timestamp 1604489732
transform 1 0 83298 0 1 146130
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_262_908
timestamp 1604489732
transform 1 0 83574 0 -1 145042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_263_908
timestamp 1604489732
transform 1 0 83574 0 1 145042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_264_908
timestamp 1604489732
transform 1 0 83574 0 -1 146130
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_265_908
timestamp 1604489732
transform 1 0 83574 0 1 146130
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_262_937
timestamp 1604489732
transform 1 0 86242 0 -1 145042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_262_932
timestamp 1604489732
transform 1 0 85782 0 -1 145042
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_262_920
timestamp 1604489732
transform 1 0 84678 0 -1 145042
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1666
timestamp 1604489732
transform 1 0 86150 0 -1 145042
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_264_937
timestamp 1604489732
transform 1 0 86242 0 -1 146130
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_264_932
timestamp 1604489732
transform 1 0 85782 0 -1 146130
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_264_920
timestamp 1604489732
transform 1 0 84678 0 -1 146130
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_263_932
timestamp 1604489732
transform 1 0 85782 0 1 145042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_263_920
timestamp 1604489732
transform 1 0 84678 0 1 145042
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1667
timestamp 1604489732
transform 1 0 86150 0 -1 146130
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_265_932
timestamp 1604489732
transform 1 0 85782 0 1 146130
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_265_920
timestamp 1604489732
transform 1 0 84678 0 1 146130
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_262_949
timestamp 1604489732
transform 1 0 87346 0 -1 145042
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1207
timestamp 1604489732
transform -1 0 87806 0 -1 145042
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_263_944
timestamp 1604489732
transform 1 0 86886 0 1 145042
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_264_949
timestamp 1604489732
transform 1 0 87346 0 -1 146130
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_263_950
timestamp 1604489732
transform 1 0 87438 0 1 145042
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1211
timestamp 1604489732
transform -1 0 87806 0 -1 146130
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1209
timestamp 1604489732
transform -1 0 87806 0 1 145042
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_265_944
timestamp 1604489732
transform 1 0 86886 0 1 146130
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_950
timestamp 1604489732
transform 1 0 87438 0 1 146130
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1213
timestamp 1604489732
transform -1 0 87806 0 1 146130
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_530
timestamp 1604489732
transform 1 0 38 0 -1 147218
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_532
timestamp 1604489732
transform 1 0 38 0 1 147218
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_534
timestamp 1604489732
transform 1 0 38 0 -1 148306
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_266_3
timestamp 1604489732
transform 1 0 314 0 -1 147218
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_266_15
timestamp 1604489732
transform 1 0 1418 0 -1 147218
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_267_3
timestamp 1604489732
transform 1 0 314 0 1 147218
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_267_15
timestamp 1604489732
transform 1 0 1418 0 1 147218
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_268_3
timestamp 1604489732
transform 1 0 314 0 -1 148306
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_268_15
timestamp 1604489732
transform 1 0 1418 0 -1 148306
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_266_38
timestamp 1604489732
transform 1 0 3534 0 -1 147218
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_266_32
timestamp 1604489732
transform 1 0 2982 0 -1 147218
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_266_27
timestamp 1604489732
transform 1 0 2522 0 -1 147218
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1496
timestamp 1604489732
transform 1 0 2890 0 -1 147218
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_531
timestamp 1604489732
transform -1 0 3902 0 -1 147218
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_267_27
timestamp 1604489732
transform 1 0 2522 0 1 147218
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_533
timestamp 1604489732
transform -1 0 3902 0 1 147218
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_268_38
timestamp 1604489732
transform 1 0 3534 0 -1 148306
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_268_32
timestamp 1604489732
transform 1 0 2982 0 -1 148306
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_268_27
timestamp 1604489732
transform 1 0 2522 0 -1 148306
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1497
timestamp 1604489732
transform 1 0 2890 0 -1 148306
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_535
timestamp 1604489732
transform -1 0 3902 0 -1 148306
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1214
timestamp 1604489732
transform 1 0 83298 0 -1 147218
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1216
timestamp 1604489732
transform 1 0 83298 0 1 147218
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1218
timestamp 1604489732
transform 1 0 83298 0 -1 148306
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_266_908
timestamp 1604489732
transform 1 0 83574 0 -1 147218
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_267_908
timestamp 1604489732
transform 1 0 83574 0 1 147218
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_268_908
timestamp 1604489732
transform 1 0 83574 0 -1 148306
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_266_937
timestamp 1604489732
transform 1 0 86242 0 -1 147218
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_266_932
timestamp 1604489732
transform 1 0 85782 0 -1 147218
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_266_920
timestamp 1604489732
transform 1 0 84678 0 -1 147218
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1668
timestamp 1604489732
transform 1 0 86150 0 -1 147218
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_267_932
timestamp 1604489732
transform 1 0 85782 0 1 147218
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_267_920
timestamp 1604489732
transform 1 0 84678 0 1 147218
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_268_937
timestamp 1604489732
transform 1 0 86242 0 -1 148306
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_268_932
timestamp 1604489732
transform 1 0 85782 0 -1 148306
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_268_920
timestamp 1604489732
transform 1 0 84678 0 -1 148306
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1669
timestamp 1604489732
transform 1 0 86150 0 -1 148306
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1215
timestamp 1604489732
transform -1 0 87806 0 -1 147218
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1217
timestamp 1604489732
transform -1 0 87806 0 1 147218
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1219
timestamp 1604489732
transform -1 0 87806 0 -1 148306
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_266_949
timestamp 1604489732
transform 1 0 87346 0 -1 147218
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_267_944
timestamp 1604489732
transform 1 0 86886 0 1 147218
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_267_950
timestamp 1604489732
transform 1 0 87438 0 1 147218
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_268_949
timestamp 1604489732
transform 1 0 87346 0 -1 148306
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_536
timestamp 1604489732
transform 1 0 38 0 1 148306
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_538
timestamp 1604489732
transform 1 0 38 0 -1 149394
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_540
timestamp 1604489732
transform 1 0 38 0 1 149394
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_269_3
timestamp 1604489732
transform 1 0 314 0 1 148306
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_269_15
timestamp 1604489732
transform 1 0 1418 0 1 148306
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_270_3
timestamp 1604489732
transform 1 0 314 0 -1 149394
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_270_15
timestamp 1604489732
transform 1 0 1418 0 -1 149394
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_271_3
timestamp 1604489732
transform 1 0 314 0 1 149394
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_271_15
timestamp 1604489732
transform 1 0 1418 0 1 149394
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_537
timestamp 1604489732
transform -1 0 3902 0 1 148306
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_539
timestamp 1604489732
transform -1 0 3902 0 -1 149394
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_541
timestamp 1604489732
transform -1 0 3902 0 1 149394
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1498
timestamp 1604489732
transform 1 0 2890 0 -1 149394
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_269_27
timestamp 1604489732
transform 1 0 2522 0 1 148306
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_270_27
timestamp 1604489732
transform 1 0 2522 0 -1 149394
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_270_32
timestamp 1604489732
transform 1 0 2982 0 -1 149394
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_270_38
timestamp 1604489732
transform 1 0 3534 0 -1 149394
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_271_27
timestamp 1604489732
transform 1 0 2522 0 1 149394
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1220
timestamp 1604489732
transform 1 0 83298 0 1 148306
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1222
timestamp 1604489732
transform 1 0 83298 0 -1 149394
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1224
timestamp 1604489732
transform 1 0 83298 0 1 149394
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_269_908
timestamp 1604489732
transform 1 0 83574 0 1 148306
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_270_908
timestamp 1604489732
transform 1 0 83574 0 -1 149394
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_271_908
timestamp 1604489732
transform 1 0 83574 0 1 149394
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1670
timestamp 1604489732
transform 1 0 86150 0 -1 149394
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_269_920
timestamp 1604489732
transform 1 0 84678 0 1 148306
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_269_932
timestamp 1604489732
transform 1 0 85782 0 1 148306
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_270_920
timestamp 1604489732
transform 1 0 84678 0 -1 149394
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_270_932
timestamp 1604489732
transform 1 0 85782 0 -1 149394
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_270_937
timestamp 1604489732
transform 1 0 86242 0 -1 149394
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_271_920
timestamp 1604489732
transform 1 0 84678 0 1 149394
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_271_932
timestamp 1604489732
transform 1 0 85782 0 1 149394
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1221
timestamp 1604489732
transform -1 0 87806 0 1 148306
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1223
timestamp 1604489732
transform -1 0 87806 0 -1 149394
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1225
timestamp 1604489732
transform -1 0 87806 0 1 149394
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_269_944
timestamp 1604489732
transform 1 0 86886 0 1 148306
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_269_950
timestamp 1604489732
transform 1 0 87438 0 1 148306
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_270_949
timestamp 1604489732
transform 1 0 87346 0 -1 149394
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_271_944
timestamp 1604489732
transform 1 0 86886 0 1 149394
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_271_950
timestamp 1604489732
transform 1 0 87438 0 1 149394
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_273_15
timestamp 1604489732
transform 1 0 1418 0 1 150482
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_273_3
timestamp 1604489732
transform 1 0 314 0 1 150482
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_272_15
timestamp 1604489732
transform 1 0 1418 0 -1 150482
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_272_3
timestamp 1604489732
transform 1 0 314 0 -1 150482
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_544
timestamp 1604489732
transform 1 0 38 0 1 150482
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_542
timestamp 1604489732
transform 1 0 38 0 -1 150482
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_274_15
timestamp 1604489732
transform 1 0 1418 0 -1 151570
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_274_3
timestamp 1604489732
transform 1 0 314 0 -1 151570
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_546
timestamp 1604489732
transform 1 0 38 0 -1 151570
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_275_15
timestamp 1604489732
transform 1 0 1418 0 1 151570
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_275_3
timestamp 1604489732
transform 1 0 314 0 1 151570
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_548
timestamp 1604489732
transform 1 0 38 0 1 151570
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_273_27
timestamp 1604489732
transform 1 0 2522 0 1 150482
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_272_38
timestamp 1604489732
transform 1 0 3534 0 -1 150482
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_272_32
timestamp 1604489732
transform 1 0 2982 0 -1 150482
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_272_27
timestamp 1604489732
transform 1 0 2522 0 -1 150482
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1499
timestamp 1604489732
transform 1 0 2890 0 -1 150482
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_545
timestamp 1604489732
transform -1 0 3902 0 1 150482
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_543
timestamp 1604489732
transform -1 0 3902 0 -1 150482
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_274_38
timestamp 1604489732
transform 1 0 3534 0 -1 151570
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_274_32
timestamp 1604489732
transform 1 0 2982 0 -1 151570
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_274_27
timestamp 1604489732
transform 1 0 2522 0 -1 151570
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1500
timestamp 1604489732
transform 1 0 2890 0 -1 151570
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_547
timestamp 1604489732
transform -1 0 3902 0 -1 151570
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_275_27
timestamp 1604489732
transform 1 0 2522 0 1 151570
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_549
timestamp 1604489732
transform -1 0 3902 0 1 151570
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1226
timestamp 1604489732
transform 1 0 83298 0 -1 150482
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1228
timestamp 1604489732
transform 1 0 83298 0 1 150482
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1230
timestamp 1604489732
transform 1 0 83298 0 -1 151570
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1232
timestamp 1604489732
transform 1 0 83298 0 1 151570
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_272_908
timestamp 1604489732
transform 1 0 83574 0 -1 150482
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_273_908
timestamp 1604489732
transform 1 0 83574 0 1 150482
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_274_908
timestamp 1604489732
transform 1 0 83574 0 -1 151570
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_275_908
timestamp 1604489732
transform 1 0 83574 0 1 151570
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_273_932
timestamp 1604489732
transform 1 0 85782 0 1 150482
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_273_920
timestamp 1604489732
transform 1 0 84678 0 1 150482
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_272_937
timestamp 1604489732
transform 1 0 86242 0 -1 150482
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_272_932
timestamp 1604489732
transform 1 0 85782 0 -1 150482
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_272_920
timestamp 1604489732
transform 1 0 84678 0 -1 150482
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1671
timestamp 1604489732
transform 1 0 86150 0 -1 150482
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_274_937
timestamp 1604489732
transform 1 0 86242 0 -1 151570
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_274_932
timestamp 1604489732
transform 1 0 85782 0 -1 151570
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_274_920
timestamp 1604489732
transform 1 0 84678 0 -1 151570
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1672
timestamp 1604489732
transform 1 0 86150 0 -1 151570
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_275_932
timestamp 1604489732
transform 1 0 85782 0 1 151570
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_275_920
timestamp 1604489732
transform 1 0 84678 0 1 151570
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_273_944
timestamp 1604489732
transform 1 0 86886 0 1 150482
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_273_950
timestamp 1604489732
transform 1 0 87438 0 1 150482
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_272_949
timestamp 1604489732
transform 1 0 87346 0 -1 150482
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1229
timestamp 1604489732
transform -1 0 87806 0 1 150482
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1227
timestamp 1604489732
transform -1 0 87806 0 -1 150482
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_274_949
timestamp 1604489732
transform 1 0 87346 0 -1 151570
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1231
timestamp 1604489732
transform -1 0 87806 0 -1 151570
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_275_944
timestamp 1604489732
transform 1 0 86886 0 1 151570
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_275_950
timestamp 1604489732
transform 1 0 87438 0 1 151570
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1233
timestamp 1604489732
transform -1 0 87806 0 1 151570
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_550
timestamp 1604489732
transform 1 0 38 0 -1 152658
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_552
timestamp 1604489732
transform 1 0 38 0 1 152658
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_554
timestamp 1604489732
transform 1 0 38 0 -1 153746
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_276_3
timestamp 1604489732
transform 1 0 314 0 -1 152658
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_276_15
timestamp 1604489732
transform 1 0 1418 0 -1 152658
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_277_3
timestamp 1604489732
transform 1 0 314 0 1 152658
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_277_15
timestamp 1604489732
transform 1 0 1418 0 1 152658
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_278_3
timestamp 1604489732
transform 1 0 314 0 -1 153746
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_278_15
timestamp 1604489732
transform 1 0 1418 0 -1 153746
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_276_38
timestamp 1604489732
transform 1 0 3534 0 -1 152658
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_276_32
timestamp 1604489732
transform 1 0 2982 0 -1 152658
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_276_27
timestamp 1604489732
transform 1 0 2522 0 -1 152658
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1501
timestamp 1604489732
transform 1 0 2890 0 -1 152658
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_551
timestamp 1604489732
transform -1 0 3902 0 -1 152658
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_277_27
timestamp 1604489732
transform 1 0 2522 0 1 152658
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_553
timestamp 1604489732
transform -1 0 3902 0 1 152658
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_278_38
timestamp 1604489732
transform 1 0 3534 0 -1 153746
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_278_32
timestamp 1604489732
transform 1 0 2982 0 -1 153746
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_278_27
timestamp 1604489732
transform 1 0 2522 0 -1 153746
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1502
timestamp 1604489732
transform 1 0 2890 0 -1 153746
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_555
timestamp 1604489732
transform -1 0 3902 0 -1 153746
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1234
timestamp 1604489732
transform 1 0 83298 0 -1 152658
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1236
timestamp 1604489732
transform 1 0 83298 0 1 152658
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1238
timestamp 1604489732
transform 1 0 83298 0 -1 153746
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_276_908
timestamp 1604489732
transform 1 0 83574 0 -1 152658
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_277_908
timestamp 1604489732
transform 1 0 83574 0 1 152658
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_278_908
timestamp 1604489732
transform 1 0 83574 0 -1 153746
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_276_937
timestamp 1604489732
transform 1 0 86242 0 -1 152658
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_276_932
timestamp 1604489732
transform 1 0 85782 0 -1 152658
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_276_920
timestamp 1604489732
transform 1 0 84678 0 -1 152658
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1673
timestamp 1604489732
transform 1 0 86150 0 -1 152658
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_277_932
timestamp 1604489732
transform 1 0 85782 0 1 152658
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_277_920
timestamp 1604489732
transform 1 0 84678 0 1 152658
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_278_937
timestamp 1604489732
transform 1 0 86242 0 -1 153746
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_278_932
timestamp 1604489732
transform 1 0 85782 0 -1 153746
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_278_920
timestamp 1604489732
transform 1 0 84678 0 -1 153746
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1674
timestamp 1604489732
transform 1 0 86150 0 -1 153746
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1235
timestamp 1604489732
transform -1 0 87806 0 -1 152658
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1237
timestamp 1604489732
transform -1 0 87806 0 1 152658
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1239
timestamp 1604489732
transform -1 0 87806 0 -1 153746
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_276_949
timestamp 1604489732
transform 1 0 87346 0 -1 152658
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_277_944
timestamp 1604489732
transform 1 0 86886 0 1 152658
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_277_950
timestamp 1604489732
transform 1 0 87438 0 1 152658
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_278_949
timestamp 1604489732
transform 1 0 87346 0 -1 153746
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_556
timestamp 1604489732
transform 1 0 38 0 1 153746
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_558
timestamp 1604489732
transform 1 0 38 0 -1 154834
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_560
timestamp 1604489732
transform 1 0 38 0 1 154834
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_279_3
timestamp 1604489732
transform 1 0 314 0 1 153746
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_279_15
timestamp 1604489732
transform 1 0 1418 0 1 153746
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_280_3
timestamp 1604489732
transform 1 0 314 0 -1 154834
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_280_15
timestamp 1604489732
transform 1 0 1418 0 -1 154834
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_281_3
timestamp 1604489732
transform 1 0 314 0 1 154834
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_281_15
timestamp 1604489732
transform 1 0 1418 0 1 154834
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_557
timestamp 1604489732
transform -1 0 3902 0 1 153746
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_559
timestamp 1604489732
transform -1 0 3902 0 -1 154834
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_561
timestamp 1604489732
transform -1 0 3902 0 1 154834
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1503
timestamp 1604489732
transform 1 0 2890 0 -1 154834
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_279_27
timestamp 1604489732
transform 1 0 2522 0 1 153746
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_280_27
timestamp 1604489732
transform 1 0 2522 0 -1 154834
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_280_32
timestamp 1604489732
transform 1 0 2982 0 -1 154834
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_280_38
timestamp 1604489732
transform 1 0 3534 0 -1 154834
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_281_27
timestamp 1604489732
transform 1 0 2522 0 1 154834
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1240
timestamp 1604489732
transform 1 0 83298 0 1 153746
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1242
timestamp 1604489732
transform 1 0 83298 0 -1 154834
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1244
timestamp 1604489732
transform 1 0 83298 0 1 154834
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_279_908
timestamp 1604489732
transform 1 0 83574 0 1 153746
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_280_908
timestamp 1604489732
transform 1 0 83574 0 -1 154834
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_281_908
timestamp 1604489732
transform 1 0 83574 0 1 154834
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1675
timestamp 1604489732
transform 1 0 86150 0 -1 154834
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_279_920
timestamp 1604489732
transform 1 0 84678 0 1 153746
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_279_932
timestamp 1604489732
transform 1 0 85782 0 1 153746
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_280_920
timestamp 1604489732
transform 1 0 84678 0 -1 154834
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_280_932
timestamp 1604489732
transform 1 0 85782 0 -1 154834
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_280_937
timestamp 1604489732
transform 1 0 86242 0 -1 154834
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_281_920
timestamp 1604489732
transform 1 0 84678 0 1 154834
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_281_932
timestamp 1604489732
transform 1 0 85782 0 1 154834
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1241
timestamp 1604489732
transform -1 0 87806 0 1 153746
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1243
timestamp 1604489732
transform -1 0 87806 0 -1 154834
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1245
timestamp 1604489732
transform -1 0 87806 0 1 154834
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_279_944
timestamp 1604489732
transform 1 0 86886 0 1 153746
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_279_950
timestamp 1604489732
transform 1 0 87438 0 1 153746
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_280_949
timestamp 1604489732
transform 1 0 87346 0 -1 154834
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_281_944
timestamp 1604489732
transform 1 0 86886 0 1 154834
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_281_950
timestamp 1604489732
transform 1 0 87438 0 1 154834
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_283_15
timestamp 1604489732
transform 1 0 1418 0 1 155922
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_283_3
timestamp 1604489732
transform 1 0 314 0 1 155922
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_282_15
timestamp 1604489732
transform 1 0 1418 0 -1 155922
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_282_3
timestamp 1604489732
transform 1 0 314 0 -1 155922
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_564
timestamp 1604489732
transform 1 0 38 0 1 155922
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_562
timestamp 1604489732
transform 1 0 38 0 -1 155922
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_284_15
timestamp 1604489732
transform 1 0 1418 0 -1 157010
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_284_3
timestamp 1604489732
transform 1 0 314 0 -1 157010
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_566
timestamp 1604489732
transform 1 0 38 0 -1 157010
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_285_15
timestamp 1604489732
transform 1 0 1418 0 1 157010
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_285_3
timestamp 1604489732
transform 1 0 314 0 1 157010
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_568
timestamp 1604489732
transform 1 0 38 0 1 157010
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_283_27
timestamp 1604489732
transform 1 0 2522 0 1 155922
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_282_38
timestamp 1604489732
transform 1 0 3534 0 -1 155922
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_282_32
timestamp 1604489732
transform 1 0 2982 0 -1 155922
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_282_27
timestamp 1604489732
transform 1 0 2522 0 -1 155922
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1504
timestamp 1604489732
transform 1 0 2890 0 -1 155922
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_565
timestamp 1604489732
transform -1 0 3902 0 1 155922
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_563
timestamp 1604489732
transform -1 0 3902 0 -1 155922
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_284_38
timestamp 1604489732
transform 1 0 3534 0 -1 157010
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_284_32
timestamp 1604489732
transform 1 0 2982 0 -1 157010
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_284_27
timestamp 1604489732
transform 1 0 2522 0 -1 157010
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1505
timestamp 1604489732
transform 1 0 2890 0 -1 157010
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_567
timestamp 1604489732
transform -1 0 3902 0 -1 157010
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_285_27
timestamp 1604489732
transform 1 0 2522 0 1 157010
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_569
timestamp 1604489732
transform -1 0 3902 0 1 157010
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1246
timestamp 1604489732
transform 1 0 83298 0 -1 155922
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1248
timestamp 1604489732
transform 1 0 83298 0 1 155922
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1250
timestamp 1604489732
transform 1 0 83298 0 -1 157010
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1252
timestamp 1604489732
transform 1 0 83298 0 1 157010
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_282_908
timestamp 1604489732
transform 1 0 83574 0 -1 155922
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_283_908
timestamp 1604489732
transform 1 0 83574 0 1 155922
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_284_908
timestamp 1604489732
transform 1 0 83574 0 -1 157010
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_285_908
timestamp 1604489732
transform 1 0 83574 0 1 157010
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_283_932
timestamp 1604489732
transform 1 0 85782 0 1 155922
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_283_920
timestamp 1604489732
transform 1 0 84678 0 1 155922
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_282_937
timestamp 1604489732
transform 1 0 86242 0 -1 155922
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_282_932
timestamp 1604489732
transform 1 0 85782 0 -1 155922
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_282_920
timestamp 1604489732
transform 1 0 84678 0 -1 155922
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1676
timestamp 1604489732
transform 1 0 86150 0 -1 155922
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_284_937
timestamp 1604489732
transform 1 0 86242 0 -1 157010
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_284_932
timestamp 1604489732
transform 1 0 85782 0 -1 157010
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_284_920
timestamp 1604489732
transform 1 0 84678 0 -1 157010
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1677
timestamp 1604489732
transform 1 0 86150 0 -1 157010
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_285_932
timestamp 1604489732
transform 1 0 85782 0 1 157010
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_285_920
timestamp 1604489732
transform 1 0 84678 0 1 157010
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_283_944
timestamp 1604489732
transform 1 0 86886 0 1 155922
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_283_950
timestamp 1604489732
transform 1 0 87438 0 1 155922
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_282_949
timestamp 1604489732
transform 1 0 87346 0 -1 155922
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1249
timestamp 1604489732
transform -1 0 87806 0 1 155922
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1247
timestamp 1604489732
transform -1 0 87806 0 -1 155922
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_284_949
timestamp 1604489732
transform 1 0 87346 0 -1 157010
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1251
timestamp 1604489732
transform -1 0 87806 0 -1 157010
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_285_944
timestamp 1604489732
transform 1 0 86886 0 1 157010
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_285_950
timestamp 1604489732
transform 1 0 87438 0 1 157010
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1253
timestamp 1604489732
transform -1 0 87806 0 1 157010
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_570
timestamp 1604489732
transform 1 0 38 0 -1 158098
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_572
timestamp 1604489732
transform 1 0 38 0 1 158098
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_574
timestamp 1604489732
transform 1 0 38 0 -1 159186
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_286_3
timestamp 1604489732
transform 1 0 314 0 -1 158098
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_286_15
timestamp 1604489732
transform 1 0 1418 0 -1 158098
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_287_3
timestamp 1604489732
transform 1 0 314 0 1 158098
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_287_15
timestamp 1604489732
transform 1 0 1418 0 1 158098
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_288_3
timestamp 1604489732
transform 1 0 314 0 -1 159186
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_288_15
timestamp 1604489732
transform 1 0 1418 0 -1 159186
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_286_38
timestamp 1604489732
transform 1 0 3534 0 -1 158098
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_286_32
timestamp 1604489732
transform 1 0 2982 0 -1 158098
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_286_27
timestamp 1604489732
transform 1 0 2522 0 -1 158098
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1506
timestamp 1604489732
transform 1 0 2890 0 -1 158098
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_571
timestamp 1604489732
transform -1 0 3902 0 -1 158098
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_287_27
timestamp 1604489732
transform 1 0 2522 0 1 158098
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_573
timestamp 1604489732
transform -1 0 3902 0 1 158098
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_288_38
timestamp 1604489732
transform 1 0 3534 0 -1 159186
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_288_32
timestamp 1604489732
transform 1 0 2982 0 -1 159186
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_288_27
timestamp 1604489732
transform 1 0 2522 0 -1 159186
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1507
timestamp 1604489732
transform 1 0 2890 0 -1 159186
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_575
timestamp 1604489732
transform -1 0 3902 0 -1 159186
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1254
timestamp 1604489732
transform 1 0 83298 0 -1 158098
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1256
timestamp 1604489732
transform 1 0 83298 0 1 158098
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1258
timestamp 1604489732
transform 1 0 83298 0 -1 159186
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_286_908
timestamp 1604489732
transform 1 0 83574 0 -1 158098
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_287_908
timestamp 1604489732
transform 1 0 83574 0 1 158098
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_288_908
timestamp 1604489732
transform 1 0 83574 0 -1 159186
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_286_937
timestamp 1604489732
transform 1 0 86242 0 -1 158098
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_286_932
timestamp 1604489732
transform 1 0 85782 0 -1 158098
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_286_920
timestamp 1604489732
transform 1 0 84678 0 -1 158098
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1678
timestamp 1604489732
transform 1 0 86150 0 -1 158098
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_287_932
timestamp 1604489732
transform 1 0 85782 0 1 158098
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_287_920
timestamp 1604489732
transform 1 0 84678 0 1 158098
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_288_937
timestamp 1604489732
transform 1 0 86242 0 -1 159186
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_288_932
timestamp 1604489732
transform 1 0 85782 0 -1 159186
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_288_920
timestamp 1604489732
transform 1 0 84678 0 -1 159186
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1679
timestamp 1604489732
transform 1 0 86150 0 -1 159186
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1255
timestamp 1604489732
transform -1 0 87806 0 -1 158098
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1257
timestamp 1604489732
transform -1 0 87806 0 1 158098
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1259
timestamp 1604489732
transform -1 0 87806 0 -1 159186
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_286_949
timestamp 1604489732
transform 1 0 87346 0 -1 158098
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_287_944
timestamp 1604489732
transform 1 0 86886 0 1 158098
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_287_950
timestamp 1604489732
transform 1 0 87438 0 1 158098
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_288_949
timestamp 1604489732
transform 1 0 87346 0 -1 159186
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_289_15
timestamp 1604489732
transform 1 0 1418 0 1 159186
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_289_3
timestamp 1604489732
transform 1 0 314 0 1 159186
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_576
timestamp 1604489732
transform 1 0 38 0 1 159186
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_291_15
timestamp 1604489732
transform 1 0 1418 0 1 160274
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_291_3
timestamp 1604489732
transform 1 0 314 0 1 160274
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_290_15
timestamp 1604489732
transform 1 0 1418 0 -1 160274
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_290_3
timestamp 1604489732
transform 1 0 314 0 -1 160274
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_580
timestamp 1604489732
transform 1 0 38 0 1 160274
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_578
timestamp 1604489732
transform 1 0 38 0 -1 160274
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_292_15
timestamp 1604489732
transform 1 0 1418 0 -1 161362
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_292_3
timestamp 1604489732
transform 1 0 314 0 -1 161362
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_582
timestamp 1604489732
transform 1 0 38 0 -1 161362
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_289_27
timestamp 1604489732
transform 1 0 2522 0 1 159186
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_577
timestamp 1604489732
transform -1 0 3902 0 1 159186
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_291_27
timestamp 1604489732
transform 1 0 2522 0 1 160274
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_290_38
timestamp 1604489732
transform 1 0 3534 0 -1 160274
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_290_32
timestamp 1604489732
transform 1 0 2982 0 -1 160274
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_290_27
timestamp 1604489732
transform 1 0 2522 0 -1 160274
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1508
timestamp 1604489732
transform 1 0 2890 0 -1 160274
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_581
timestamp 1604489732
transform -1 0 3902 0 1 160274
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_579
timestamp 1604489732
transform -1 0 3902 0 -1 160274
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_292_38
timestamp 1604489732
transform 1 0 3534 0 -1 161362
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_292_32
timestamp 1604489732
transform 1 0 2982 0 -1 161362
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_292_27
timestamp 1604489732
transform 1 0 2522 0 -1 161362
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1509
timestamp 1604489732
transform 1 0 2890 0 -1 161362
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_583
timestamp 1604489732
transform -1 0 3902 0 -1 161362
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1260
timestamp 1604489732
transform 1 0 83298 0 1 159186
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1262
timestamp 1604489732
transform 1 0 83298 0 -1 160274
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1264
timestamp 1604489732
transform 1 0 83298 0 1 160274
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1266
timestamp 1604489732
transform 1 0 83298 0 -1 161362
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_289_908
timestamp 1604489732
transform 1 0 83574 0 1 159186
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_290_908
timestamp 1604489732
transform 1 0 83574 0 -1 160274
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_291_908
timestamp 1604489732
transform 1 0 83574 0 1 160274
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_292_908
timestamp 1604489732
transform 1 0 83574 0 -1 161362
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_289_932
timestamp 1604489732
transform 1 0 85782 0 1 159186
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_289_920
timestamp 1604489732
transform 1 0 84678 0 1 159186
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_291_932
timestamp 1604489732
transform 1 0 85782 0 1 160274
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_291_920
timestamp 1604489732
transform 1 0 84678 0 1 160274
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_290_937
timestamp 1604489732
transform 1 0 86242 0 -1 160274
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_290_932
timestamp 1604489732
transform 1 0 85782 0 -1 160274
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_290_920
timestamp 1604489732
transform 1 0 84678 0 -1 160274
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1680
timestamp 1604489732
transform 1 0 86150 0 -1 160274
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_292_937
timestamp 1604489732
transform 1 0 86242 0 -1 161362
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_292_932
timestamp 1604489732
transform 1 0 85782 0 -1 161362
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_292_920
timestamp 1604489732
transform 1 0 84678 0 -1 161362
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1681
timestamp 1604489732
transform 1 0 86150 0 -1 161362
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_289_944
timestamp 1604489732
transform 1 0 86886 0 1 159186
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_289_950
timestamp 1604489732
transform 1 0 87438 0 1 159186
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1261
timestamp 1604489732
transform -1 0 87806 0 1 159186
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_291_944
timestamp 1604489732
transform 1 0 86886 0 1 160274
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_291_950
timestamp 1604489732
transform 1 0 87438 0 1 160274
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_290_949
timestamp 1604489732
transform 1 0 87346 0 -1 160274
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1265
timestamp 1604489732
transform -1 0 87806 0 1 160274
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1263
timestamp 1604489732
transform -1 0 87806 0 -1 160274
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_292_949
timestamp 1604489732
transform 1 0 87346 0 -1 161362
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1267
timestamp 1604489732
transform -1 0 87806 0 -1 161362
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_584
timestamp 1604489732
transform 1 0 38 0 1 161362
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_586
timestamp 1604489732
transform 1 0 38 0 -1 162450
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_588
timestamp 1604489732
transform 1 0 38 0 1 162450
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_293_3
timestamp 1604489732
transform 1 0 314 0 1 161362
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_293_15
timestamp 1604489732
transform 1 0 1418 0 1 161362
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_294_3
timestamp 1604489732
transform 1 0 314 0 -1 162450
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_294_15
timestamp 1604489732
transform 1 0 1418 0 -1 162450
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_295_3
timestamp 1604489732
transform 1 0 314 0 1 162450
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_295_15
timestamp 1604489732
transform 1 0 1418 0 1 162450
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_585
timestamp 1604489732
transform -1 0 3902 0 1 161362
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_587
timestamp 1604489732
transform -1 0 3902 0 -1 162450
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_589
timestamp 1604489732
transform -1 0 3902 0 1 162450
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1510
timestamp 1604489732
transform 1 0 2890 0 -1 162450
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_293_27
timestamp 1604489732
transform 1 0 2522 0 1 161362
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_294_27
timestamp 1604489732
transform 1 0 2522 0 -1 162450
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_294_32
timestamp 1604489732
transform 1 0 2982 0 -1 162450
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_294_38
timestamp 1604489732
transform 1 0 3534 0 -1 162450
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_295_27
timestamp 1604489732
transform 1 0 2522 0 1 162450
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1268
timestamp 1604489732
transform 1 0 83298 0 1 161362
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1270
timestamp 1604489732
transform 1 0 83298 0 -1 162450
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1272
timestamp 1604489732
transform 1 0 83298 0 1 162450
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_293_908
timestamp 1604489732
transform 1 0 83574 0 1 161362
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_294_908
timestamp 1604489732
transform 1 0 83574 0 -1 162450
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_295_908
timestamp 1604489732
transform 1 0 83574 0 1 162450
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1682
timestamp 1604489732
transform 1 0 86150 0 -1 162450
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_293_920
timestamp 1604489732
transform 1 0 84678 0 1 161362
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_293_932
timestamp 1604489732
transform 1 0 85782 0 1 161362
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_294_920
timestamp 1604489732
transform 1 0 84678 0 -1 162450
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_294_932
timestamp 1604489732
transform 1 0 85782 0 -1 162450
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_294_937
timestamp 1604489732
transform 1 0 86242 0 -1 162450
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_295_920
timestamp 1604489732
transform 1 0 84678 0 1 162450
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_295_932
timestamp 1604489732
transform 1 0 85782 0 1 162450
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1269
timestamp 1604489732
transform -1 0 87806 0 1 161362
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1271
timestamp 1604489732
transform -1 0 87806 0 -1 162450
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1273
timestamp 1604489732
transform -1 0 87806 0 1 162450
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_293_944
timestamp 1604489732
transform 1 0 86886 0 1 161362
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_293_950
timestamp 1604489732
transform 1 0 87438 0 1 161362
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_294_949
timestamp 1604489732
transform 1 0 87346 0 -1 162450
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_295_944
timestamp 1604489732
transform 1 0 86886 0 1 162450
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_295_950
timestamp 1604489732
transform 1 0 87438 0 1 162450
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_590
timestamp 1604489732
transform 1 0 38 0 -1 163538
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_592
timestamp 1604489732
transform 1 0 38 0 1 163538
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_594
timestamp 1604489732
transform 1 0 38 0 -1 164626
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_296_3
timestamp 1604489732
transform 1 0 314 0 -1 163538
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_296_15
timestamp 1604489732
transform 1 0 1418 0 -1 163538
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_297_3
timestamp 1604489732
transform 1 0 314 0 1 163538
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_297_15
timestamp 1604489732
transform 1 0 1418 0 1 163538
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_298_3
timestamp 1604489732
transform 1 0 314 0 -1 164626
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_298_15
timestamp 1604489732
transform 1 0 1418 0 -1 164626
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_296_38
timestamp 1604489732
transform 1 0 3534 0 -1 163538
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_296_32
timestamp 1604489732
transform 1 0 2982 0 -1 163538
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_296_27
timestamp 1604489732
transform 1 0 2522 0 -1 163538
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1511
timestamp 1604489732
transform 1 0 2890 0 -1 163538
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_591
timestamp 1604489732
transform -1 0 3902 0 -1 163538
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_297_27
timestamp 1604489732
transform 1 0 2522 0 1 163538
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_593
timestamp 1604489732
transform -1 0 3902 0 1 163538
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_298_38
timestamp 1604489732
transform 1 0 3534 0 -1 164626
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_298_32
timestamp 1604489732
transform 1 0 2982 0 -1 164626
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_298_27
timestamp 1604489732
transform 1 0 2522 0 -1 164626
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1512
timestamp 1604489732
transform 1 0 2890 0 -1 164626
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_595
timestamp 1604489732
transform -1 0 3902 0 -1 164626
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1274
timestamp 1604489732
transform 1 0 83298 0 -1 163538
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1276
timestamp 1604489732
transform 1 0 83298 0 1 163538
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1278
timestamp 1604489732
transform 1 0 83298 0 -1 164626
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_296_908
timestamp 1604489732
transform 1 0 83574 0 -1 163538
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_297_908
timestamp 1604489732
transform 1 0 83574 0 1 163538
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_298_908
timestamp 1604489732
transform 1 0 83574 0 -1 164626
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_296_937
timestamp 1604489732
transform 1 0 86242 0 -1 163538
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_296_932
timestamp 1604489732
transform 1 0 85782 0 -1 163538
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_296_920
timestamp 1604489732
transform 1 0 84678 0 -1 163538
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1683
timestamp 1604489732
transform 1 0 86150 0 -1 163538
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_297_932
timestamp 1604489732
transform 1 0 85782 0 1 163538
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_297_920
timestamp 1604489732
transform 1 0 84678 0 1 163538
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_298_937
timestamp 1604489732
transform 1 0 86242 0 -1 164626
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_298_932
timestamp 1604489732
transform 1 0 85782 0 -1 164626
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_298_920
timestamp 1604489732
transform 1 0 84678 0 -1 164626
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1684
timestamp 1604489732
transform 1 0 86150 0 -1 164626
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1275
timestamp 1604489732
transform -1 0 87806 0 -1 163538
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1277
timestamp 1604489732
transform -1 0 87806 0 1 163538
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1279
timestamp 1604489732
transform -1 0 87806 0 -1 164626
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_296_949
timestamp 1604489732
transform 1 0 87346 0 -1 163538
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_297_944
timestamp 1604489732
transform 1 0 86886 0 1 163538
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_297_950
timestamp 1604489732
transform 1 0 87438 0 1 163538
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_298_949
timestamp 1604489732
transform 1 0 87346 0 -1 164626
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_300_15
timestamp 1604489732
transform 1 0 1418 0 -1 165714
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_300_3
timestamp 1604489732
transform 1 0 314 0 -1 165714
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_299_15
timestamp 1604489732
transform 1 0 1418 0 1 164626
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_299_3
timestamp 1604489732
transform 1 0 314 0 1 164626
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_598
timestamp 1604489732
transform 1 0 38 0 -1 165714
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_596
timestamp 1604489732
transform 1 0 38 0 1 164626
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_301_15
timestamp 1604489732
transform 1 0 1418 0 1 165714
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_301_3
timestamp 1604489732
transform 1 0 314 0 1 165714
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_600
timestamp 1604489732
transform 1 0 38 0 1 165714
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_302_15
timestamp 1604489732
transform 1 0 1418 0 -1 166802
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_302_3
timestamp 1604489732
transform 1 0 314 0 -1 166802
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_602
timestamp 1604489732
transform 1 0 38 0 -1 166802
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_300_38
timestamp 1604489732
transform 1 0 3534 0 -1 165714
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_300_32
timestamp 1604489732
transform 1 0 2982 0 -1 165714
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_300_27
timestamp 1604489732
transform 1 0 2522 0 -1 165714
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_299_27
timestamp 1604489732
transform 1 0 2522 0 1 164626
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1513
timestamp 1604489732
transform 1 0 2890 0 -1 165714
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_599
timestamp 1604489732
transform -1 0 3902 0 -1 165714
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_597
timestamp 1604489732
transform -1 0 3902 0 1 164626
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_301_27
timestamp 1604489732
transform 1 0 2522 0 1 165714
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_601
timestamp 1604489732
transform -1 0 3902 0 1 165714
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_302_38
timestamp 1604489732
transform 1 0 3534 0 -1 166802
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_302_32
timestamp 1604489732
transform 1 0 2982 0 -1 166802
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_302_27
timestamp 1604489732
transform 1 0 2522 0 -1 166802
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1514
timestamp 1604489732
transform 1 0 2890 0 -1 166802
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_603
timestamp 1604489732
transform -1 0 3902 0 -1 166802
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1280
timestamp 1604489732
transform 1 0 83298 0 1 164626
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1282
timestamp 1604489732
transform 1 0 83298 0 -1 165714
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1284
timestamp 1604489732
transform 1 0 83298 0 1 165714
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1286
timestamp 1604489732
transform 1 0 83298 0 -1 166802
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_299_908
timestamp 1604489732
transform 1 0 83574 0 1 164626
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_300_908
timestamp 1604489732
transform 1 0 83574 0 -1 165714
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_301_908
timestamp 1604489732
transform 1 0 83574 0 1 165714
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_302_908
timestamp 1604489732
transform 1 0 83574 0 -1 166802
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_300_937
timestamp 1604489732
transform 1 0 86242 0 -1 165714
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_300_932
timestamp 1604489732
transform 1 0 85782 0 -1 165714
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_300_920
timestamp 1604489732
transform 1 0 84678 0 -1 165714
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_299_932
timestamp 1604489732
transform 1 0 85782 0 1 164626
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_299_920
timestamp 1604489732
transform 1 0 84678 0 1 164626
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1685
timestamp 1604489732
transform 1 0 86150 0 -1 165714
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_301_932
timestamp 1604489732
transform 1 0 85782 0 1 165714
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_301_920
timestamp 1604489732
transform 1 0 84678 0 1 165714
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_302_937
timestamp 1604489732
transform 1 0 86242 0 -1 166802
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_302_932
timestamp 1604489732
transform 1 0 85782 0 -1 166802
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_302_920
timestamp 1604489732
transform 1 0 84678 0 -1 166802
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1686
timestamp 1604489732
transform 1 0 86150 0 -1 166802
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_299_944
timestamp 1604489732
transform 1 0 86886 0 1 164626
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_300_949
timestamp 1604489732
transform 1 0 87346 0 -1 165714
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_299_950
timestamp 1604489732
transform 1 0 87438 0 1 164626
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1283
timestamp 1604489732
transform -1 0 87806 0 -1 165714
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1281
timestamp 1604489732
transform -1 0 87806 0 1 164626
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_301_944
timestamp 1604489732
transform 1 0 86886 0 1 165714
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_301_950
timestamp 1604489732
transform 1 0 87438 0 1 165714
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1285
timestamp 1604489732
transform -1 0 87806 0 1 165714
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_302_949
timestamp 1604489732
transform 1 0 87346 0 -1 166802
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1287
timestamp 1604489732
transform -1 0 87806 0 -1 166802
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_604
timestamp 1604489732
transform 1 0 38 0 1 166802
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_606
timestamp 1604489732
transform 1 0 38 0 -1 167890
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_608
timestamp 1604489732
transform 1 0 38 0 1 167890
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_303_3
timestamp 1604489732
transform 1 0 314 0 1 166802
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_303_15
timestamp 1604489732
transform 1 0 1418 0 1 166802
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_304_3
timestamp 1604489732
transform 1 0 314 0 -1 167890
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_304_15
timestamp 1604489732
transform 1 0 1418 0 -1 167890
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_305_3
timestamp 1604489732
transform 1 0 314 0 1 167890
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_305_15
timestamp 1604489732
transform 1 0 1418 0 1 167890
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_605
timestamp 1604489732
transform -1 0 3902 0 1 166802
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_607
timestamp 1604489732
transform -1 0 3902 0 -1 167890
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_609
timestamp 1604489732
transform -1 0 3902 0 1 167890
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1515
timestamp 1604489732
transform 1 0 2890 0 -1 167890
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_303_27
timestamp 1604489732
transform 1 0 2522 0 1 166802
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_304_27
timestamp 1604489732
transform 1 0 2522 0 -1 167890
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_304_32
timestamp 1604489732
transform 1 0 2982 0 -1 167890
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_304_38
timestamp 1604489732
transform 1 0 3534 0 -1 167890
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_305_27
timestamp 1604489732
transform 1 0 2522 0 1 167890
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1288
timestamp 1604489732
transform 1 0 83298 0 1 166802
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1290
timestamp 1604489732
transform 1 0 83298 0 -1 167890
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1292
timestamp 1604489732
transform 1 0 83298 0 1 167890
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_303_908
timestamp 1604489732
transform 1 0 83574 0 1 166802
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_304_908
timestamp 1604489732
transform 1 0 83574 0 -1 167890
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_305_908
timestamp 1604489732
transform 1 0 83574 0 1 167890
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1687
timestamp 1604489732
transform 1 0 86150 0 -1 167890
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_303_920
timestamp 1604489732
transform 1 0 84678 0 1 166802
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_303_932
timestamp 1604489732
transform 1 0 85782 0 1 166802
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_304_920
timestamp 1604489732
transform 1 0 84678 0 -1 167890
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_304_932
timestamp 1604489732
transform 1 0 85782 0 -1 167890
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_304_937
timestamp 1604489732
transform 1 0 86242 0 -1 167890
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_305_920
timestamp 1604489732
transform 1 0 84678 0 1 167890
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_305_932
timestamp 1604489732
transform 1 0 85782 0 1 167890
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1289
timestamp 1604489732
transform -1 0 87806 0 1 166802
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1291
timestamp 1604489732
transform -1 0 87806 0 -1 167890
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1293
timestamp 1604489732
transform -1 0 87806 0 1 167890
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_303_944
timestamp 1604489732
transform 1 0 86886 0 1 166802
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_303_950
timestamp 1604489732
transform 1 0 87438 0 1 166802
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_304_949
timestamp 1604489732
transform 1 0 87346 0 -1 167890
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_305_944
timestamp 1604489732
transform 1 0 86886 0 1 167890
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_305_950
timestamp 1604489732
transform 1 0 87438 0 1 167890
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_306_15
timestamp 1604489732
transform 1 0 1418 0 -1 168978
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_306_3
timestamp 1604489732
transform 1 0 314 0 -1 168978
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_610
timestamp 1604489732
transform 1 0 38 0 -1 168978
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_307_15
timestamp 1604489732
transform 1 0 1418 0 1 168978
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_307_3
timestamp 1604489732
transform 1 0 314 0 1 168978
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_612
timestamp 1604489732
transform 1 0 38 0 1 168978
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_309_15
timestamp 1604489732
transform 1 0 1418 0 1 170066
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_309_3
timestamp 1604489732
transform 1 0 314 0 1 170066
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_308_15
timestamp 1604489732
transform 1 0 1418 0 -1 170066
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_308_3
timestamp 1604489732
transform 1 0 314 0 -1 170066
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_616
timestamp 1604489732
transform 1 0 38 0 1 170066
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_614
timestamp 1604489732
transform 1 0 38 0 -1 170066
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_306_38
timestamp 1604489732
transform 1 0 3534 0 -1 168978
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_306_32
timestamp 1604489732
transform 1 0 2982 0 -1 168978
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_306_27
timestamp 1604489732
transform 1 0 2522 0 -1 168978
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1516
timestamp 1604489732
transform 1 0 2890 0 -1 168978
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_611
timestamp 1604489732
transform -1 0 3902 0 -1 168978
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_307_27
timestamp 1604489732
transform 1 0 2522 0 1 168978
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_613
timestamp 1604489732
transform -1 0 3902 0 1 168978
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_309_27
timestamp 1604489732
transform 1 0 2522 0 1 170066
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_308_38
timestamp 1604489732
transform 1 0 3534 0 -1 170066
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_308_32
timestamp 1604489732
transform 1 0 2982 0 -1 170066
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_308_27
timestamp 1604489732
transform 1 0 2522 0 -1 170066
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1517
timestamp 1604489732
transform 1 0 2890 0 -1 170066
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_617
timestamp 1604489732
transform -1 0 3902 0 1 170066
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_615
timestamp 1604489732
transform -1 0 3902 0 -1 170066
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1294
timestamp 1604489732
transform 1 0 83298 0 -1 168978
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1296
timestamp 1604489732
transform 1 0 83298 0 1 168978
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1298
timestamp 1604489732
transform 1 0 83298 0 -1 170066
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1300
timestamp 1604489732
transform 1 0 83298 0 1 170066
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_306_908
timestamp 1604489732
transform 1 0 83574 0 -1 168978
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_307_908
timestamp 1604489732
transform 1 0 83574 0 1 168978
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_308_908
timestamp 1604489732
transform 1 0 83574 0 -1 170066
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_309_908
timestamp 1604489732
transform 1 0 83574 0 1 170066
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_306_937
timestamp 1604489732
transform 1 0 86242 0 -1 168978
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_306_932
timestamp 1604489732
transform 1 0 85782 0 -1 168978
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_306_920
timestamp 1604489732
transform 1 0 84678 0 -1 168978
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1688
timestamp 1604489732
transform 1 0 86150 0 -1 168978
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_307_932
timestamp 1604489732
transform 1 0 85782 0 1 168978
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_307_920
timestamp 1604489732
transform 1 0 84678 0 1 168978
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_309_932
timestamp 1604489732
transform 1 0 85782 0 1 170066
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_309_920
timestamp 1604489732
transform 1 0 84678 0 1 170066
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_308_937
timestamp 1604489732
transform 1 0 86242 0 -1 170066
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_308_932
timestamp 1604489732
transform 1 0 85782 0 -1 170066
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_308_920
timestamp 1604489732
transform 1 0 84678 0 -1 170066
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1689
timestamp 1604489732
transform 1 0 86150 0 -1 170066
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_306_949
timestamp 1604489732
transform 1 0 87346 0 -1 168978
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1295
timestamp 1604489732
transform -1 0 87806 0 -1 168978
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_307_944
timestamp 1604489732
transform 1 0 86886 0 1 168978
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_307_950
timestamp 1604489732
transform 1 0 87438 0 1 168978
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1297
timestamp 1604489732
transform -1 0 87806 0 1 168978
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_309_944
timestamp 1604489732
transform 1 0 86886 0 1 170066
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_309_950
timestamp 1604489732
transform 1 0 87438 0 1 170066
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_308_949
timestamp 1604489732
transform 1 0 87346 0 -1 170066
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1301
timestamp 1604489732
transform -1 0 87806 0 1 170066
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1299
timestamp 1604489732
transform -1 0 87806 0 -1 170066
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_618
timestamp 1604489732
transform 1 0 38 0 -1 171154
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_620
timestamp 1604489732
transform 1 0 38 0 1 171154
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_622
timestamp 1604489732
transform 1 0 38 0 -1 172242
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_310_3
timestamp 1604489732
transform 1 0 314 0 -1 171154
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_310_15
timestamp 1604489732
transform 1 0 1418 0 -1 171154
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_311_3
timestamp 1604489732
transform 1 0 314 0 1 171154
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_311_15
timestamp 1604489732
transform 1 0 1418 0 1 171154
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_312_3
timestamp 1604489732
transform 1 0 314 0 -1 172242
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_312_15
timestamp 1604489732
transform 1 0 1418 0 -1 172242
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_310_38
timestamp 1604489732
transform 1 0 3534 0 -1 171154
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_310_32
timestamp 1604489732
transform 1 0 2982 0 -1 171154
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_310_27
timestamp 1604489732
transform 1 0 2522 0 -1 171154
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1518
timestamp 1604489732
transform 1 0 2890 0 -1 171154
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_619
timestamp 1604489732
transform -1 0 3902 0 -1 171154
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_311_27
timestamp 1604489732
transform 1 0 2522 0 1 171154
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_621
timestamp 1604489732
transform -1 0 3902 0 1 171154
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_312_38
timestamp 1604489732
transform 1 0 3534 0 -1 172242
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_312_32
timestamp 1604489732
transform 1 0 2982 0 -1 172242
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_312_27
timestamp 1604489732
transform 1 0 2522 0 -1 172242
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1519
timestamp 1604489732
transform 1 0 2890 0 -1 172242
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_623
timestamp 1604489732
transform -1 0 3902 0 -1 172242
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1302
timestamp 1604489732
transform 1 0 83298 0 -1 171154
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1304
timestamp 1604489732
transform 1 0 83298 0 1 171154
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1306
timestamp 1604489732
transform 1 0 83298 0 -1 172242
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_310_908
timestamp 1604489732
transform 1 0 83574 0 -1 171154
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_311_908
timestamp 1604489732
transform 1 0 83574 0 1 171154
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_312_908
timestamp 1604489732
transform 1 0 83574 0 -1 172242
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_310_937
timestamp 1604489732
transform 1 0 86242 0 -1 171154
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_310_932
timestamp 1604489732
transform 1 0 85782 0 -1 171154
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_310_920
timestamp 1604489732
transform 1 0 84678 0 -1 171154
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1690
timestamp 1604489732
transform 1 0 86150 0 -1 171154
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_311_932
timestamp 1604489732
transform 1 0 85782 0 1 171154
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_311_920
timestamp 1604489732
transform 1 0 84678 0 1 171154
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_312_937
timestamp 1604489732
transform 1 0 86242 0 -1 172242
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_312_932
timestamp 1604489732
transform 1 0 85782 0 -1 172242
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_312_920
timestamp 1604489732
transform 1 0 84678 0 -1 172242
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1691
timestamp 1604489732
transform 1 0 86150 0 -1 172242
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1303
timestamp 1604489732
transform -1 0 87806 0 -1 171154
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1305
timestamp 1604489732
transform -1 0 87806 0 1 171154
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1307
timestamp 1604489732
transform -1 0 87806 0 -1 172242
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_310_949
timestamp 1604489732
transform 1 0 87346 0 -1 171154
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_311_944
timestamp 1604489732
transform 1 0 86886 0 1 171154
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_311_950
timestamp 1604489732
transform 1 0 87438 0 1 171154
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_312_949
timestamp 1604489732
transform 1 0 87346 0 -1 172242
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_624
timestamp 1604489732
transform 1 0 38 0 1 172242
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_626
timestamp 1604489732
transform 1 0 38 0 -1 173330
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_628
timestamp 1604489732
transform 1 0 38 0 1 173330
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_313_3
timestamp 1604489732
transform 1 0 314 0 1 172242
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_313_15
timestamp 1604489732
transform 1 0 1418 0 1 172242
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_314_3
timestamp 1604489732
transform 1 0 314 0 -1 173330
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_314_15
timestamp 1604489732
transform 1 0 1418 0 -1 173330
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_315_3
timestamp 1604489732
transform 1 0 314 0 1 173330
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_315_15
timestamp 1604489732
transform 1 0 1418 0 1 173330
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_625
timestamp 1604489732
transform -1 0 3902 0 1 172242
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_627
timestamp 1604489732
transform -1 0 3902 0 -1 173330
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_629
timestamp 1604489732
transform -1 0 3902 0 1 173330
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1520
timestamp 1604489732
transform 1 0 2890 0 -1 173330
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_313_27
timestamp 1604489732
transform 1 0 2522 0 1 172242
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_314_27
timestamp 1604489732
transform 1 0 2522 0 -1 173330
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_314_32
timestamp 1604489732
transform 1 0 2982 0 -1 173330
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_314_38
timestamp 1604489732
transform 1 0 3534 0 -1 173330
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_315_27
timestamp 1604489732
transform 1 0 2522 0 1 173330
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1308
timestamp 1604489732
transform 1 0 83298 0 1 172242
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1310
timestamp 1604489732
transform 1 0 83298 0 -1 173330
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1312
timestamp 1604489732
transform 1 0 83298 0 1 173330
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_313_908
timestamp 1604489732
transform 1 0 83574 0 1 172242
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_314_908
timestamp 1604489732
transform 1 0 83574 0 -1 173330
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_315_908
timestamp 1604489732
transform 1 0 83574 0 1 173330
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1692
timestamp 1604489732
transform 1 0 86150 0 -1 173330
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_313_920
timestamp 1604489732
transform 1 0 84678 0 1 172242
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_313_932
timestamp 1604489732
transform 1 0 85782 0 1 172242
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_314_920
timestamp 1604489732
transform 1 0 84678 0 -1 173330
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_314_932
timestamp 1604489732
transform 1 0 85782 0 -1 173330
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_314_937
timestamp 1604489732
transform 1 0 86242 0 -1 173330
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_315_920
timestamp 1604489732
transform 1 0 84678 0 1 173330
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_315_932
timestamp 1604489732
transform 1 0 85782 0 1 173330
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1309
timestamp 1604489732
transform -1 0 87806 0 1 172242
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1311
timestamp 1604489732
transform -1 0 87806 0 -1 173330
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1313
timestamp 1604489732
transform -1 0 87806 0 1 173330
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_313_944
timestamp 1604489732
transform 1 0 86886 0 1 172242
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_313_950
timestamp 1604489732
transform 1 0 87438 0 1 172242
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_314_949
timestamp 1604489732
transform 1 0 87346 0 -1 173330
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_315_944
timestamp 1604489732
transform 1 0 86886 0 1 173330
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_315_950
timestamp 1604489732
transform 1 0 87438 0 1 173330
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_316_15
timestamp 1604489732
transform 1 0 1418 0 -1 174418
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_316_3
timestamp 1604489732
transform 1 0 314 0 -1 174418
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_630
timestamp 1604489732
transform 1 0 38 0 -1 174418
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_318_15
timestamp 1604489732
transform 1 0 1418 0 -1 175506
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_318_3
timestamp 1604489732
transform 1 0 314 0 -1 175506
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_317_15
timestamp 1604489732
transform 1 0 1418 0 1 174418
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_317_3
timestamp 1604489732
transform 1 0 314 0 1 174418
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_634
timestamp 1604489732
transform 1 0 38 0 -1 175506
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_632
timestamp 1604489732
transform 1 0 38 0 1 174418
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_319_15
timestamp 1604489732
transform 1 0 1418 0 1 175506
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_319_3
timestamp 1604489732
transform 1 0 314 0 1 175506
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_636
timestamp 1604489732
transform 1 0 38 0 1 175506
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_316_36
timestamp 1604489732
transform 1 0 3350 0 -1 174418
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_316_32
timestamp 1604489732
transform 1 0 2982 0 -1 174418
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_316_27
timestamp 1604489732
transform 1 0 2522 0 -1 174418
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_addr0[1]
timestamp 1604489732
transform 1 0 3442 0 -1 174418
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1521
timestamp 1604489732
transform 1 0 2890 0 -1 174418
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_631
timestamp 1604489732
transform -1 0 3902 0 -1 174418
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_318_38
timestamp 1604489732
transform 1 0 3534 0 -1 175506
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_318_32
timestamp 1604489732
transform 1 0 2982 0 -1 175506
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_318_27
timestamp 1604489732
transform 1 0 2522 0 -1 175506
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_317_27
timestamp 1604489732
transform 1 0 2522 0 1 174418
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1522
timestamp 1604489732
transform 1 0 2890 0 -1 175506
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_635
timestamp 1604489732
transform -1 0 3902 0 -1 175506
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_633
timestamp 1604489732
transform -1 0 3902 0 1 174418
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_319_35
timestamp 1604489732
transform 1 0 3258 0 1 175506
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_319_27
timestamp 1604489732
transform 1 0 2522 0 1 175506
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_addr0[2]
timestamp 1604489732
transform 1 0 3442 0 1 175506
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_637
timestamp 1604489732
transform -1 0 3902 0 1 175506
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1314
timestamp 1604489732
transform 1 0 83298 0 -1 174418
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1316
timestamp 1604489732
transform 1 0 83298 0 1 174418
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1318
timestamp 1604489732
transform 1 0 83298 0 -1 175506
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1320
timestamp 1604489732
transform 1 0 83298 0 1 175506
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_316_908
timestamp 1604489732
transform 1 0 83574 0 -1 174418
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_317_908
timestamp 1604489732
transform 1 0 83574 0 1 174418
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_318_908
timestamp 1604489732
transform 1 0 83574 0 -1 175506
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_319_908
timestamp 1604489732
transform 1 0 83574 0 1 175506
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_316_937
timestamp 1604489732
transform 1 0 86242 0 -1 174418
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_316_932
timestamp 1604489732
transform 1 0 85782 0 -1 174418
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_316_920
timestamp 1604489732
transform 1 0 84678 0 -1 174418
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1693
timestamp 1604489732
transform 1 0 86150 0 -1 174418
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_318_937
timestamp 1604489732
transform 1 0 86242 0 -1 175506
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_318_932
timestamp 1604489732
transform 1 0 85782 0 -1 175506
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_318_920
timestamp 1604489732
transform 1 0 84678 0 -1 175506
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_317_932
timestamp 1604489732
transform 1 0 85782 0 1 174418
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_317_920
timestamp 1604489732
transform 1 0 84678 0 1 174418
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1694
timestamp 1604489732
transform 1 0 86150 0 -1 175506
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_319_932
timestamp 1604489732
transform 1 0 85782 0 1 175506
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_319_920
timestamp 1604489732
transform 1 0 84678 0 1 175506
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_316_949
timestamp 1604489732
transform 1 0 87346 0 -1 174418
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1315
timestamp 1604489732
transform -1 0 87806 0 -1 174418
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_317_944
timestamp 1604489732
transform 1 0 86886 0 1 174418
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_318_949
timestamp 1604489732
transform 1 0 87346 0 -1 175506
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_317_950
timestamp 1604489732
transform 1 0 87438 0 1 174418
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1319
timestamp 1604489732
transform -1 0 87806 0 -1 175506
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1317
timestamp 1604489732
transform -1 0 87806 0 1 174418
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_319_944
timestamp 1604489732
transform 1 0 86886 0 1 175506
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_319_950
timestamp 1604489732
transform 1 0 87438 0 1 175506
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1321
timestamp 1604489732
transform -1 0 87806 0 1 175506
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_638
timestamp 1604489732
transform 1 0 38 0 -1 176594
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_640
timestamp 1604489732
transform 1 0 38 0 1 176594
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_642
timestamp 1604489732
transform 1 0 38 0 -1 177682
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_320_3
timestamp 1604489732
transform 1 0 314 0 -1 176594
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_320_15
timestamp 1604489732
transform 1 0 1418 0 -1 176594
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_321_3
timestamp 1604489732
transform 1 0 314 0 1 176594
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_321_15
timestamp 1604489732
transform 1 0 1418 0 1 176594
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_322_3
timestamp 1604489732
transform 1 0 314 0 -1 177682
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_322_15
timestamp 1604489732
transform 1 0 1418 0 -1 177682
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_320_27
timestamp 1604489732
transform 1 0 2522 0 -1 176594
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_320_32
timestamp 1604489732
transform 1 0 2982 0 -1 176594
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1523
timestamp 1604489732
transform 1 0 2890 0 -1 176594
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_320_38
timestamp 1604489732
transform 1 0 3534 0 -1 176594
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_639
timestamp 1604489732
transform -1 0 3902 0 -1 176594
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_321_27
timestamp 1604489732
transform 1 0 2522 0 1 176594
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_321_35
timestamp 1604489732
transform 1 0 3258 0 1 176594
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_addr0[3]
timestamp 1604489732
transform 1 0 3442 0 1 176594
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_641
timestamp 1604489732
transform -1 0 3902 0 1 176594
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_322_27
timestamp 1604489732
transform 1 0 2522 0 -1 177682
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_322_32
timestamp 1604489732
transform 1 0 2982 0 -1 177682
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1524
timestamp 1604489732
transform 1 0 2890 0 -1 177682
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_322_38
timestamp 1604489732
transform 1 0 3534 0 -1 177682
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_643
timestamp 1604489732
transform -1 0 3902 0 -1 177682
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1322
timestamp 1604489732
transform 1 0 83298 0 -1 176594
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1324
timestamp 1604489732
transform 1 0 83298 0 1 176594
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1326
timestamp 1604489732
transform 1 0 83298 0 -1 177682
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_320_908
timestamp 1604489732
transform 1 0 83574 0 -1 176594
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_321_908
timestamp 1604489732
transform 1 0 83574 0 1 176594
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_322_908
timestamp 1604489732
transform 1 0 83574 0 -1 177682
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_320_937
timestamp 1604489732
transform 1 0 86242 0 -1 176594
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_320_932
timestamp 1604489732
transform 1 0 85782 0 -1 176594
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_320_920
timestamp 1604489732
transform 1 0 84678 0 -1 176594
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1695
timestamp 1604489732
transform 1 0 86150 0 -1 176594
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_321_932
timestamp 1604489732
transform 1 0 85782 0 1 176594
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_321_920
timestamp 1604489732
transform 1 0 84678 0 1 176594
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_322_937
timestamp 1604489732
transform 1 0 86242 0 -1 177682
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_322_932
timestamp 1604489732
transform 1 0 85782 0 -1 177682
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_322_920
timestamp 1604489732
transform 1 0 84678 0 -1 177682
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1696
timestamp 1604489732
transform 1 0 86150 0 -1 177682
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1323
timestamp 1604489732
transform -1 0 87806 0 -1 176594
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1325
timestamp 1604489732
transform -1 0 87806 0 1 176594
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1327
timestamp 1604489732
transform -1 0 87806 0 -1 177682
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_320_949
timestamp 1604489732
transform 1 0 87346 0 -1 176594
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_321_944
timestamp 1604489732
transform 1 0 86886 0 1 176594
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_321_950
timestamp 1604489732
transform 1 0 87438 0 1 176594
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_322_949
timestamp 1604489732
transform 1 0 87346 0 -1 177682
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_644
timestamp 1604489732
transform 1 0 38 0 1 177682
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_646
timestamp 1604489732
transform 1 0 38 0 -1 178770
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_648
timestamp 1604489732
transform 1 0 38 0 1 178770
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_323_3
timestamp 1604489732
transform 1 0 314 0 1 177682
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_323_15
timestamp 1604489732
transform 1 0 1418 0 1 177682
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_324_3
timestamp 1604489732
transform 1 0 314 0 -1 178770
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_324_15
timestamp 1604489732
transform 1 0 1418 0 -1 178770
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_325_3
timestamp 1604489732
transform 1 0 314 0 1 178770
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_325_15
timestamp 1604489732
transform 1 0 1418 0 1 178770
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_323_27
timestamp 1604489732
transform 1 0 2522 0 1 177682
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_645
timestamp 1604489732
transform -1 0 3902 0 1 177682
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_324_38
timestamp 1604489732
transform 1 0 3534 0 -1 178770
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_324_32
timestamp 1604489732
transform 1 0 2982 0 -1 178770
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_324_27
timestamp 1604489732
transform 1 0 2522 0 -1 178770
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1525
timestamp 1604489732
transform 1 0 2890 0 -1 178770
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_647
timestamp 1604489732
transform -1 0 3902 0 -1 178770
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_325_35
timestamp 1604489732
transform 1 0 3258 0 1 178770
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_325_27
timestamp 1604489732
transform 1 0 2522 0 1 178770
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_addr0[4]
timestamp 1604489732
transform 1 0 3442 0 1 178770
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_649
timestamp 1604489732
transform -1 0 3902 0 1 178770
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1328
timestamp 1604489732
transform 1 0 83298 0 1 177682
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1330
timestamp 1604489732
transform 1 0 83298 0 -1 178770
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1332
timestamp 1604489732
transform 1 0 83298 0 1 178770
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_323_908
timestamp 1604489732
transform 1 0 83574 0 1 177682
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_324_908
timestamp 1604489732
transform 1 0 83574 0 -1 178770
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_325_908
timestamp 1604489732
transform 1 0 83574 0 1 178770
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1697
timestamp 1604489732
transform 1 0 86150 0 -1 178770
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_323_920
timestamp 1604489732
transform 1 0 84678 0 1 177682
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_323_932
timestamp 1604489732
transform 1 0 85782 0 1 177682
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_324_920
timestamp 1604489732
transform 1 0 84678 0 -1 178770
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_324_932
timestamp 1604489732
transform 1 0 85782 0 -1 178770
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_324_937
timestamp 1604489732
transform 1 0 86242 0 -1 178770
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_325_920
timestamp 1604489732
transform 1 0 84678 0 1 178770
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_325_932
timestamp 1604489732
transform 1 0 85782 0 1 178770
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1329
timestamp 1604489732
transform -1 0 87806 0 1 177682
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1331
timestamp 1604489732
transform -1 0 87806 0 -1 178770
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1333
timestamp 1604489732
transform -1 0 87806 0 1 178770
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_323_944
timestamp 1604489732
transform 1 0 86886 0 1 177682
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_323_950
timestamp 1604489732
transform 1 0 87438 0 1 177682
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_324_949
timestamp 1604489732
transform 1 0 87346 0 -1 178770
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_325_944
timestamp 1604489732
transform 1 0 86886 0 1 178770
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_325_950
timestamp 1604489732
transform 1 0 87438 0 1 178770
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_327_15
timestamp 1604489732
transform 1 0 1418 0 1 179858
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_327_3
timestamp 1604489732
transform 1 0 314 0 1 179858
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_326_15
timestamp 1604489732
transform 1 0 1418 0 -1 179858
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_326_3
timestamp 1604489732
transform 1 0 314 0 -1 179858
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_652
timestamp 1604489732
transform 1 0 38 0 1 179858
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_650
timestamp 1604489732
transform 1 0 38 0 -1 179858
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_328_15
timestamp 1604489732
transform 1 0 1418 0 -1 180946
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_328_3
timestamp 1604489732
transform 1 0 314 0 -1 180946
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_654
timestamp 1604489732
transform 1 0 38 0 -1 180946
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_329_15
timestamp 1604489732
transform 1 0 1418 0 1 180946
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_329_3
timestamp 1604489732
transform 1 0 314 0 1 180946
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_656
timestamp 1604489732
transform 1 0 38 0 1 180946
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_327_35
timestamp 1604489732
transform 1 0 3258 0 1 179858
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_327_27
timestamp 1604489732
transform 1 0 2522 0 1 179858
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_326_38
timestamp 1604489732
transform 1 0 3534 0 -1 179858
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_326_32
timestamp 1604489732
transform 1 0 2982 0 -1 179858
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_326_27
timestamp 1604489732
transform 1 0 2522 0 -1 179858
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_addr0[5]
timestamp 1604489732
transform 1 0 3442 0 1 179858
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1526
timestamp 1604489732
transform 1 0 2890 0 -1 179858
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_653
timestamp 1604489732
transform -1 0 3902 0 1 179858
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_651
timestamp 1604489732
transform -1 0 3902 0 -1 179858
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_328_38
timestamp 1604489732
transform 1 0 3534 0 -1 180946
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_328_32
timestamp 1604489732
transform 1 0 2982 0 -1 180946
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_328_27
timestamp 1604489732
transform 1 0 2522 0 -1 180946
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1527
timestamp 1604489732
transform 1 0 2890 0 -1 180946
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_655
timestamp 1604489732
transform -1 0 3902 0 -1 180946
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_329_27
timestamp 1604489732
transform 1 0 2522 0 1 180946
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_657
timestamp 1604489732
transform -1 0 3902 0 1 180946
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1334
timestamp 1604489732
transform 1 0 83298 0 -1 179858
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1336
timestamp 1604489732
transform 1 0 83298 0 1 179858
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1338
timestamp 1604489732
transform 1 0 83298 0 -1 180946
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1340
timestamp 1604489732
transform 1 0 83298 0 1 180946
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_326_908
timestamp 1604489732
transform 1 0 83574 0 -1 179858
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_327_908
timestamp 1604489732
transform 1 0 83574 0 1 179858
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_328_908
timestamp 1604489732
transform 1 0 83574 0 -1 180946
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_329_908
timestamp 1604489732
transform 1 0 83574 0 1 180946
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_327_932
timestamp 1604489732
transform 1 0 85782 0 1 179858
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_327_920
timestamp 1604489732
transform 1 0 84678 0 1 179858
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_326_937
timestamp 1604489732
transform 1 0 86242 0 -1 179858
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_326_932
timestamp 1604489732
transform 1 0 85782 0 -1 179858
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_326_920
timestamp 1604489732
transform 1 0 84678 0 -1 179858
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1698
timestamp 1604489732
transform 1 0 86150 0 -1 179858
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_328_937
timestamp 1604489732
transform 1 0 86242 0 -1 180946
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_328_932
timestamp 1604489732
transform 1 0 85782 0 -1 180946
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_328_920
timestamp 1604489732
transform 1 0 84678 0 -1 180946
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1699
timestamp 1604489732
transform 1 0 86150 0 -1 180946
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_329_932
timestamp 1604489732
transform 1 0 85782 0 1 180946
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_329_920
timestamp 1604489732
transform 1 0 84678 0 1 180946
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_327_944
timestamp 1604489732
transform 1 0 86886 0 1 179858
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_327_950
timestamp 1604489732
transform 1 0 87438 0 1 179858
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_326_949
timestamp 1604489732
transform 1 0 87346 0 -1 179858
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1337
timestamp 1604489732
transform -1 0 87806 0 1 179858
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1335
timestamp 1604489732
transform -1 0 87806 0 -1 179858
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_328_949
timestamp 1604489732
transform 1 0 87346 0 -1 180946
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1339
timestamp 1604489732
transform -1 0 87806 0 -1 180946
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_329_944
timestamp 1604489732
transform 1 0 86886 0 1 180946
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_329_950
timestamp 1604489732
transform 1 0 87438 0 1 180946
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1341
timestamp 1604489732
transform -1 0 87806 0 1 180946
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_658
timestamp 1604489732
transform 1 0 38 0 -1 182034
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_660
timestamp 1604489732
transform 1 0 38 0 1 182034
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_662
timestamp 1604489732
transform 1 0 38 0 -1 183122
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_330_3
timestamp 1604489732
transform 1 0 314 0 -1 182034
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_330_15
timestamp 1604489732
transform 1 0 1418 0 -1 182034
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_331_3
timestamp 1604489732
transform 1 0 314 0 1 182034
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_331_15
timestamp 1604489732
transform 1 0 1418 0 1 182034
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_332_3
timestamp 1604489732
transform 1 0 314 0 -1 183122
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_332_15
timestamp 1604489732
transform 1 0 1418 0 -1 183122
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_330_36
timestamp 1604489732
transform 1 0 3350 0 -1 182034
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_330_32
timestamp 1604489732
transform 1 0 2982 0 -1 182034
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_330_27
timestamp 1604489732
transform 1 0 2522 0 -1 182034
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_addr0[6]
timestamp 1604489732
transform 1 0 3442 0 -1 182034
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1528
timestamp 1604489732
transform 1 0 2890 0 -1 182034
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_659
timestamp 1604489732
transform -1 0 3902 0 -1 182034
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_331_27
timestamp 1604489732
transform 1 0 2522 0 1 182034
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_661
timestamp 1604489732
transform -1 0 3902 0 1 182034
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_332_36
timestamp 1604489732
transform 1 0 3350 0 -1 183122
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_332_32
timestamp 1604489732
transform 1 0 2982 0 -1 183122
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_332_27
timestamp 1604489732
transform 1 0 2522 0 -1 183122
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_addr0[7]
timestamp 1604489732
transform 1 0 3442 0 -1 183122
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1529
timestamp 1604489732
transform 1 0 2890 0 -1 183122
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_663
timestamp 1604489732
transform -1 0 3902 0 -1 183122
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1342
timestamp 1604489732
transform 1 0 83298 0 -1 182034
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1344
timestamp 1604489732
transform 1 0 83298 0 1 182034
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1346
timestamp 1604489732
transform 1 0 83298 0 -1 183122
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_330_908
timestamp 1604489732
transform 1 0 83574 0 -1 182034
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_331_908
timestamp 1604489732
transform 1 0 83574 0 1 182034
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_332_908
timestamp 1604489732
transform 1 0 83574 0 -1 183122
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_330_937
timestamp 1604489732
transform 1 0 86242 0 -1 182034
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_330_932
timestamp 1604489732
transform 1 0 85782 0 -1 182034
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_330_920
timestamp 1604489732
transform 1 0 84678 0 -1 182034
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1700
timestamp 1604489732
transform 1 0 86150 0 -1 182034
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_331_932
timestamp 1604489732
transform 1 0 85782 0 1 182034
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_331_920
timestamp 1604489732
transform 1 0 84678 0 1 182034
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_332_937
timestamp 1604489732
transform 1 0 86242 0 -1 183122
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_332_932
timestamp 1604489732
transform 1 0 85782 0 -1 183122
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_332_920
timestamp 1604489732
transform 1 0 84678 0 -1 183122
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1701
timestamp 1604489732
transform 1 0 86150 0 -1 183122
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1343
timestamp 1604489732
transform -1 0 87806 0 -1 182034
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1345
timestamp 1604489732
transform -1 0 87806 0 1 182034
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1347
timestamp 1604489732
transform -1 0 87806 0 -1 183122
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_330_949
timestamp 1604489732
transform 1 0 87346 0 -1 182034
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_331_944
timestamp 1604489732
transform 1 0 86886 0 1 182034
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_331_950
timestamp 1604489732
transform 1 0 87438 0 1 182034
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_332_949
timestamp 1604489732
transform 1 0 87346 0 -1 183122
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_664
timestamp 1604489732
transform 1 0 38 0 1 183122
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_666
timestamp 1604489732
transform 1 0 38 0 -1 184210
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_668
timestamp 1604489732
transform 1 0 38 0 1 184210
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_333_3
timestamp 1604489732
transform 1 0 314 0 1 183122
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_333_15
timestamp 1604489732
transform 1 0 1418 0 1 183122
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_334_3
timestamp 1604489732
transform 1 0 314 0 -1 184210
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_334_15
timestamp 1604489732
transform 1 0 1418 0 -1 184210
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_335_3
timestamp 1604489732
transform 1 0 314 0 1 184210
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_335_15
timestamp 1604489732
transform 1 0 1418 0 1 184210
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_665
timestamp 1604489732
transform -1 0 3902 0 1 183122
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_667
timestamp 1604489732
transform -1 0 3902 0 -1 184210
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_669
timestamp 1604489732
transform -1 0 3902 0 1 184210
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1530
timestamp 1604489732
transform 1 0 2890 0 -1 184210
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_333_27
timestamp 1604489732
transform 1 0 2522 0 1 183122
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_334_27
timestamp 1604489732
transform 1 0 2522 0 -1 184210
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_334_32
timestamp 1604489732
transform 1 0 2982 0 -1 184210
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_334_38
timestamp 1604489732
transform 1 0 3534 0 -1 184210
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_335_27
timestamp 1604489732
transform 1 0 2522 0 1 184210
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1348
timestamp 1604489732
transform 1 0 83298 0 1 183122
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1350
timestamp 1604489732
transform 1 0 83298 0 -1 184210
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1352
timestamp 1604489732
transform 1 0 83298 0 1 184210
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_333_908
timestamp 1604489732
transform 1 0 83574 0 1 183122
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_334_908
timestamp 1604489732
transform 1 0 83574 0 -1 184210
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_335_908
timestamp 1604489732
transform 1 0 83574 0 1 184210
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1702
timestamp 1604489732
transform 1 0 86150 0 -1 184210
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_333_920
timestamp 1604489732
transform 1 0 84678 0 1 183122
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_333_932
timestamp 1604489732
transform 1 0 85782 0 1 183122
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_334_920
timestamp 1604489732
transform 1 0 84678 0 -1 184210
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_334_932
timestamp 1604489732
transform 1 0 85782 0 -1 184210
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_334_937
timestamp 1604489732
transform 1 0 86242 0 -1 184210
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_335_920
timestamp 1604489732
transform 1 0 84678 0 1 184210
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_335_932
timestamp 1604489732
transform 1 0 85782 0 1 184210
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1349
timestamp 1604489732
transform -1 0 87806 0 1 183122
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1351
timestamp 1604489732
transform -1 0 87806 0 -1 184210
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1353
timestamp 1604489732
transform -1 0 87806 0 1 184210
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_333_944
timestamp 1604489732
transform 1 0 86886 0 1 183122
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_333_950
timestamp 1604489732
transform 1 0 87438 0 1 183122
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_334_949
timestamp 1604489732
transform 1 0 87346 0 -1 184210
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_335_944
timestamp 1604489732
transform 1 0 86886 0 1 184210
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_335_950
timestamp 1604489732
transform 1 0 87438 0 1 184210
box -38 -48 130 592
use sram_1rw1r_32_256_8_sky130  SRAM_1
timestamp 1605062100
transform 1 0 4934 0 1 96202
box 0 0 77296 91247
use sky130_fd_sc_hd__decap_3  PHY_670
timestamp 1604489732
transform 1 0 38 0 -1 185298
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_672
timestamp 1604489732
transform 1 0 38 0 1 185298
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_674
timestamp 1604489732
transform 1 0 38 0 -1 186386
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_336_3
timestamp 1604489732
transform 1 0 314 0 -1 185298
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_336_15
timestamp 1604489732
transform 1 0 1418 0 -1 185298
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_337_3
timestamp 1604489732
transform 1 0 314 0 1 185298
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_337_15
timestamp 1604489732
transform 1 0 1418 0 1 185298
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_338_3
timestamp 1604489732
transform 1 0 314 0 -1 186386
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_338_15
timestamp 1604489732
transform 1 0 1418 0 -1 186386
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_336_38
timestamp 1604489732
transform 1 0 3534 0 -1 185298
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_336_32
timestamp 1604489732
transform 1 0 2982 0 -1 185298
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_336_27
timestamp 1604489732
transform 1 0 2522 0 -1 185298
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1531
timestamp 1604489732
transform 1 0 2890 0 -1 185298
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_671
timestamp 1604489732
transform -1 0 3902 0 -1 185298
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_337_27
timestamp 1604489732
transform 1 0 2522 0 1 185298
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_673
timestamp 1604489732
transform -1 0 3902 0 1 185298
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_338_38
timestamp 1604489732
transform 1 0 3534 0 -1 186386
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_338_32
timestamp 1604489732
transform 1 0 2982 0 -1 186386
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_338_27
timestamp 1604489732
transform 1 0 2522 0 -1 186386
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1532
timestamp 1604489732
transform 1 0 2890 0 -1 186386
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_675
timestamp 1604489732
transform -1 0 3902 0 -1 186386
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_676
timestamp 1604489732
transform 1 0 38 0 1 186386
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_678
timestamp 1604489732
transform 1 0 38 0 -1 187474
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_339_3
timestamp 1604489732
transform 1 0 314 0 1 186386
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_339_15
timestamp 1604489732
transform 1 0 1418 0 1 186386
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_340_3
timestamp 1604489732
transform 1 0 314 0 -1 187474
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_340_15
timestamp 1604489732
transform 1 0 1418 0 -1 187474
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_677
timestamp 1604489732
transform -1 0 3902 0 1 186386
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_679
timestamp 1604489732
transform -1 0 3902 0 -1 187474
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1533
timestamp 1604489732
transform 1 0 2890 0 -1 187474
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_339_27
timestamp 1604489732
transform 1 0 2522 0 1 186386
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_340_27
timestamp 1604489732
transform 1 0 2522 0 -1 187474
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_340_32
timestamp 1604489732
transform 1 0 2982 0 -1 187474
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_340_38
timestamp 1604489732
transform 1 0 3534 0 -1 187474
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_337_908
timestamp 1604489732
transform 1 0 83574 0 1 185298
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_336_908
timestamp 1604489732
transform 1 0 83574 0 -1 185298
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1356
timestamp 1604489732
transform 1 0 83298 0 1 185298
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1354
timestamp 1604489732
transform 1 0 83298 0 -1 185298
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_339_908
timestamp 1604489732
transform 1 0 83574 0 1 186386
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_338_908
timestamp 1604489732
transform 1 0 83574 0 -1 186386
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1360
timestamp 1604489732
transform 1 0 83298 0 1 186386
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1358
timestamp 1604489732
transform 1 0 83298 0 -1 186386
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_340_908
timestamp 1604489732
transform 1 0 83574 0 -1 187474
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1362
timestamp 1604489732
transform 1 0 83298 0 -1 187474
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_336_937
timestamp 1604489732
transform 1 0 86242 0 -1 185298
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_336_932
timestamp 1604489732
transform 1 0 85782 0 -1 185298
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_336_920
timestamp 1604489732
transform 1 0 84678 0 -1 185298
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1703
timestamp 1604489732
transform 1 0 86150 0 -1 185298
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_337_932
timestamp 1604489732
transform 1 0 85782 0 1 185298
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_337_920
timestamp 1604489732
transform 1 0 84678 0 1 185298
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_339_932
timestamp 1604489732
transform 1 0 85782 0 1 186386
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_339_920
timestamp 1604489732
transform 1 0 84678 0 1 186386
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_338_937
timestamp 1604489732
transform 1 0 86242 0 -1 186386
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_338_932
timestamp 1604489732
transform 1 0 85782 0 -1 186386
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_338_920
timestamp 1604489732
transform 1 0 84678 0 -1 186386
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1704
timestamp 1604489732
transform 1 0 86150 0 -1 186386
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_336_949
timestamp 1604489732
transform 1 0 87346 0 -1 185298
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1355
timestamp 1604489732
transform -1 0 87806 0 -1 185298
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_337_944
timestamp 1604489732
transform 1 0 86886 0 1 185298
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_337_950
timestamp 1604489732
transform 1 0 87438 0 1 185298
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1357
timestamp 1604489732
transform -1 0 87806 0 1 185298
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_339_944
timestamp 1604489732
transform 1 0 86886 0 1 186386
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_338_949
timestamp 1604489732
transform 1 0 87346 0 -1 186386
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_339_950
timestamp 1604489732
transform 1 0 87438 0 1 186386
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1361
timestamp 1604489732
transform -1 0 87806 0 1 186386
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1359
timestamp 1604489732
transform -1 0 87806 0 -1 186386
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1705
timestamp 1604489732
transform 1 0 86150 0 -1 187474
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_340_920
timestamp 1604489732
transform 1 0 84678 0 -1 187474
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_340_932
timestamp 1604489732
transform 1 0 85782 0 -1 187474
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_340_937
timestamp 1604489732
transform 1 0 86242 0 -1 187474
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1363
timestamp 1604489732
transform -1 0 87806 0 -1 187474
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_340_949
timestamp 1604489732
transform 1 0 87346 0 -1 187474
box -38 -48 222 592
<< labels >>
rlabel metal3 s 88454 346 88934 466 6 mgmt_addr[0]
port 0 nsew default input
rlabel metal3 s 88454 1434 88934 1554 6 mgmt_addr[1]
port 1 nsew default input
rlabel metal3 s 88454 2658 88934 2778 6 mgmt_addr[2]
port 2 nsew default input
rlabel metal3 s 88454 3882 88934 4002 6 mgmt_addr[3]
port 3 nsew default input
rlabel metal3 s 88454 5106 88934 5226 6 mgmt_addr[4]
port 4 nsew default input
rlabel metal3 s 88454 6330 88934 6450 6 mgmt_addr[5]
port 5 nsew default input
rlabel metal3 s 88454 7554 88934 7674 6 mgmt_addr[6]
port 6 nsew default input
rlabel metal3 s 88454 8642 88934 8762 6 mgmt_addr[7]
port 7 nsew default input
rlabel metal3 s 88454 9866 88934 9986 6 mgmt_addr_ro[0]
port 8 nsew default input
rlabel metal3 s 88454 11090 88934 11210 6 mgmt_addr_ro[1]
port 9 nsew default input
rlabel metal3 s 88454 12314 88934 12434 6 mgmt_addr_ro[2]
port 10 nsew default input
rlabel metal3 s 88454 13538 88934 13658 6 mgmt_addr_ro[3]
port 11 nsew default input
rlabel metal3 s 88454 14762 88934 14882 6 mgmt_addr_ro[4]
port 12 nsew default input
rlabel metal3 s 88454 15850 88934 15970 6 mgmt_addr_ro[5]
port 13 nsew default input
rlabel metal3 s 88454 17074 88934 17194 6 mgmt_addr_ro[6]
port 14 nsew default input
rlabel metal3 s 88454 18298 88934 18418 6 mgmt_addr_ro[7]
port 15 nsew default input
rlabel metal3 s 88454 19522 88934 19642 6 mgmt_clk
port 16 nsew default input
rlabel metal3 s 88454 20746 88934 20866 6 mgmt_ena[0]
port 17 nsew default input
rlabel metal3 s 88454 21970 88934 22090 6 mgmt_ena[1]
port 18 nsew default input
rlabel metal3 s 88454 23058 88934 23178 6 mgmt_ena_ro
port 19 nsew default input
rlabel metal3 s 88454 24282 88934 24402 6 mgmt_rdata[0]
port 20 nsew default tristate
rlabel metal3 s 88454 36386 88934 36506 6 mgmt_rdata[10]
port 21 nsew default tristate
rlabel metal3 s 88454 37610 88934 37730 6 mgmt_rdata[11]
port 22 nsew default tristate
rlabel metal3 s 88454 38698 88934 38818 6 mgmt_rdata[12]
port 23 nsew default tristate
rlabel metal3 s 88454 39922 88934 40042 6 mgmt_rdata[13]
port 24 nsew default tristate
rlabel metal3 s 88454 41146 88934 41266 6 mgmt_rdata[14]
port 25 nsew default tristate
rlabel metal3 s 88454 42370 88934 42490 6 mgmt_rdata[15]
port 26 nsew default tristate
rlabel metal3 s 88454 43594 88934 43714 6 mgmt_rdata[16]
port 27 nsew default tristate
rlabel metal3 s 88454 44818 88934 44938 6 mgmt_rdata[17]
port 28 nsew default tristate
rlabel metal3 s 88454 45906 88934 46026 6 mgmt_rdata[18]
port 29 nsew default tristate
rlabel metal3 s 88454 47130 88934 47250 6 mgmt_rdata[19]
port 30 nsew default tristate
rlabel metal3 s 88454 25506 88934 25626 6 mgmt_rdata[1]
port 31 nsew default tristate
rlabel metal3 s 88454 48354 88934 48474 6 mgmt_rdata[20]
port 32 nsew default tristate
rlabel metal3 s 88454 49578 88934 49698 6 mgmt_rdata[21]
port 33 nsew default tristate
rlabel metal3 s 88454 50802 88934 50922 6 mgmt_rdata[22]
port 34 nsew default tristate
rlabel metal3 s 88454 52026 88934 52146 6 mgmt_rdata[23]
port 35 nsew default tristate
rlabel metal3 s 88454 53250 88934 53370 6 mgmt_rdata[24]
port 36 nsew default tristate
rlabel metal3 s 88454 54338 88934 54458 6 mgmt_rdata[25]
port 37 nsew default tristate
rlabel metal3 s 88454 55562 88934 55682 6 mgmt_rdata[26]
port 38 nsew default tristate
rlabel metal3 s 88454 56786 88934 56906 6 mgmt_rdata[27]
port 39 nsew default tristate
rlabel metal3 s 88454 58010 88934 58130 6 mgmt_rdata[28]
port 40 nsew default tristate
rlabel metal3 s 88454 59234 88934 59354 6 mgmt_rdata[29]
port 41 nsew default tristate
rlabel metal3 s 88454 26730 88934 26850 6 mgmt_rdata[2]
port 42 nsew default tristate
rlabel metal3 s 88454 60458 88934 60578 6 mgmt_rdata[30]
port 43 nsew default tristate
rlabel metal3 s 88454 61546 88934 61666 6 mgmt_rdata[31]
port 44 nsew default tristate
rlabel metal3 s 88454 62770 88934 62890 6 mgmt_rdata[32]
port 45 nsew default tristate
rlabel metal3 s 88454 63994 88934 64114 6 mgmt_rdata[33]
port 46 nsew default tristate
rlabel metal3 s 88454 65218 88934 65338 6 mgmt_rdata[34]
port 47 nsew default tristate
rlabel metal3 s 88454 66442 88934 66562 6 mgmt_rdata[35]
port 48 nsew default tristate
rlabel metal3 s 88454 67666 88934 67786 6 mgmt_rdata[36]
port 49 nsew default tristate
rlabel metal3 s 88454 68754 88934 68874 6 mgmt_rdata[37]
port 50 nsew default tristate
rlabel metal3 s 88454 69978 88934 70098 6 mgmt_rdata[38]
port 51 nsew default tristate
rlabel metal3 s 88454 71202 88934 71322 6 mgmt_rdata[39]
port 52 nsew default tristate
rlabel metal3 s 88454 27954 88934 28074 6 mgmt_rdata[3]
port 53 nsew default tristate
rlabel metal3 s 88454 72426 88934 72546 6 mgmt_rdata[40]
port 54 nsew default tristate
rlabel metal3 s 88454 73650 88934 73770 6 mgmt_rdata[41]
port 55 nsew default tristate
rlabel metal3 s 88454 74874 88934 74994 6 mgmt_rdata[42]
port 56 nsew default tristate
rlabel metal3 s 88454 76098 88934 76218 6 mgmt_rdata[43]
port 57 nsew default tristate
rlabel metal3 s 88454 77186 88934 77306 6 mgmt_rdata[44]
port 58 nsew default tristate
rlabel metal3 s 88454 78410 88934 78530 6 mgmt_rdata[45]
port 59 nsew default tristate
rlabel metal3 s 88454 79634 88934 79754 6 mgmt_rdata[46]
port 60 nsew default tristate
rlabel metal3 s 88454 80858 88934 80978 6 mgmt_rdata[47]
port 61 nsew default tristate
rlabel metal3 s 88454 82082 88934 82202 6 mgmt_rdata[48]
port 62 nsew default tristate
rlabel metal3 s 88454 83306 88934 83426 6 mgmt_rdata[49]
port 63 nsew default tristate
rlabel metal3 s 88454 29178 88934 29298 6 mgmt_rdata[4]
port 64 nsew default tristate
rlabel metal3 s 88454 84394 88934 84514 6 mgmt_rdata[50]
port 65 nsew default tristate
rlabel metal3 s 88454 85618 88934 85738 6 mgmt_rdata[51]
port 66 nsew default tristate
rlabel metal3 s 88454 86842 88934 86962 6 mgmt_rdata[52]
port 67 nsew default tristate
rlabel metal3 s 88454 88066 88934 88186 6 mgmt_rdata[53]
port 68 nsew default tristate
rlabel metal3 s 88454 89290 88934 89410 6 mgmt_rdata[54]
port 69 nsew default tristate
rlabel metal3 s 88454 90514 88934 90634 6 mgmt_rdata[55]
port 70 nsew default tristate
rlabel metal3 s 88454 91602 88934 91722 6 mgmt_rdata[56]
port 71 nsew default tristate
rlabel metal3 s 88454 92826 88934 92946 6 mgmt_rdata[57]
port 72 nsew default tristate
rlabel metal3 s 88454 94050 88934 94170 6 mgmt_rdata[58]
port 73 nsew default tristate
rlabel metal3 s 88454 95274 88934 95394 6 mgmt_rdata[59]
port 74 nsew default tristate
rlabel metal3 s 88454 30402 88934 30522 6 mgmt_rdata[5]
port 75 nsew default tristate
rlabel metal3 s 88454 96498 88934 96618 6 mgmt_rdata[60]
port 76 nsew default tristate
rlabel metal3 s 88454 97722 88934 97842 6 mgmt_rdata[61]
port 77 nsew default tristate
rlabel metal3 s 88454 98946 88934 99066 6 mgmt_rdata[62]
port 78 nsew default tristate
rlabel metal3 s 88454 100034 88934 100154 6 mgmt_rdata[63]
port 79 nsew default tristate
rlabel metal3 s 88454 31490 88934 31610 6 mgmt_rdata[6]
port 80 nsew default tristate
rlabel metal3 s 88454 32714 88934 32834 6 mgmt_rdata[7]
port 81 nsew default tristate
rlabel metal3 s 88454 33938 88934 34058 6 mgmt_rdata[8]
port 82 nsew default tristate
rlabel metal3 s 88454 35162 88934 35282 6 mgmt_rdata[9]
port 83 nsew default tristate
rlabel metal3 s 88454 101258 88934 101378 6 mgmt_rdata_ro[0]
port 84 nsew default tristate
rlabel metal3 s 88454 113362 88934 113482 6 mgmt_rdata_ro[10]
port 85 nsew default tristate
rlabel metal3 s 88454 114450 88934 114570 6 mgmt_rdata_ro[11]
port 86 nsew default tristate
rlabel metal3 s 88454 115674 88934 115794 6 mgmt_rdata_ro[12]
port 87 nsew default tristate
rlabel metal3 s 88454 116898 88934 117018 6 mgmt_rdata_ro[13]
port 88 nsew default tristate
rlabel metal3 s 88454 118122 88934 118242 6 mgmt_rdata_ro[14]
port 89 nsew default tristate
rlabel metal3 s 88454 119346 88934 119466 6 mgmt_rdata_ro[15]
port 90 nsew default tristate
rlabel metal3 s 88454 120570 88934 120690 6 mgmt_rdata_ro[16]
port 91 nsew default tristate
rlabel metal3 s 88454 121794 88934 121914 6 mgmt_rdata_ro[17]
port 92 nsew default tristate
rlabel metal3 s 88454 122882 88934 123002 6 mgmt_rdata_ro[18]
port 93 nsew default tristate
rlabel metal3 s 88454 124106 88934 124226 6 mgmt_rdata_ro[19]
port 94 nsew default tristate
rlabel metal3 s 88454 102482 88934 102602 6 mgmt_rdata_ro[1]
port 95 nsew default tristate
rlabel metal3 s 88454 125330 88934 125450 6 mgmt_rdata_ro[20]
port 96 nsew default tristate
rlabel metal3 s 88454 126554 88934 126674 6 mgmt_rdata_ro[21]
port 97 nsew default tristate
rlabel metal3 s 88454 127778 88934 127898 6 mgmt_rdata_ro[22]
port 98 nsew default tristate
rlabel metal3 s 88454 129002 88934 129122 6 mgmt_rdata_ro[23]
port 99 nsew default tristate
rlabel metal3 s 88454 130090 88934 130210 6 mgmt_rdata_ro[24]
port 100 nsew default tristate
rlabel metal3 s 88454 131314 88934 131434 6 mgmt_rdata_ro[25]
port 101 nsew default tristate
rlabel metal3 s 88454 132538 88934 132658 6 mgmt_rdata_ro[26]
port 102 nsew default tristate
rlabel metal3 s 88454 133762 88934 133882 6 mgmt_rdata_ro[27]
port 103 nsew default tristate
rlabel metal3 s 88454 134986 88934 135106 6 mgmt_rdata_ro[28]
port 104 nsew default tristate
rlabel metal3 s 88454 136210 88934 136330 6 mgmt_rdata_ro[29]
port 105 nsew default tristate
rlabel metal3 s 88454 103706 88934 103826 6 mgmt_rdata_ro[2]
port 106 nsew default tristate
rlabel metal3 s 88454 137298 88934 137418 6 mgmt_rdata_ro[30]
port 107 nsew default tristate
rlabel metal3 s 88454 138522 88934 138642 6 mgmt_rdata_ro[31]
port 108 nsew default tristate
rlabel metal3 s 88454 104930 88934 105050 6 mgmt_rdata_ro[3]
port 109 nsew default tristate
rlabel metal3 s 88454 106154 88934 106274 6 mgmt_rdata_ro[4]
port 110 nsew default tristate
rlabel metal3 s 88454 107242 88934 107362 6 mgmt_rdata_ro[5]
port 111 nsew default tristate
rlabel metal3 s 88454 108466 88934 108586 6 mgmt_rdata_ro[6]
port 112 nsew default tristate
rlabel metal3 s 88454 109690 88934 109810 6 mgmt_rdata_ro[7]
port 113 nsew default tristate
rlabel metal3 s 88454 110914 88934 111034 6 mgmt_rdata_ro[8]
port 114 nsew default tristate
rlabel metal3 s 88454 112138 88934 112258 6 mgmt_rdata_ro[9]
port 115 nsew default tristate
rlabel metal3 s 88454 139746 88934 139866 6 mgmt_wdata[0]
port 116 nsew default input
rlabel metal3 s 88454 151850 88934 151970 6 mgmt_wdata[10]
port 117 nsew default input
rlabel metal3 s 88454 152938 88934 153058 6 mgmt_wdata[11]
port 118 nsew default input
rlabel metal3 s 88454 154162 88934 154282 6 mgmt_wdata[12]
port 119 nsew default input
rlabel metal3 s 88454 155386 88934 155506 6 mgmt_wdata[13]
port 120 nsew default input
rlabel metal3 s 88454 156610 88934 156730 6 mgmt_wdata[14]
port 121 nsew default input
rlabel metal3 s 88454 157834 88934 157954 6 mgmt_wdata[15]
port 122 nsew default input
rlabel metal3 s 88454 159058 88934 159178 6 mgmt_wdata[16]
port 123 nsew default input
rlabel metal3 s 88454 160146 88934 160266 6 mgmt_wdata[17]
port 124 nsew default input
rlabel metal3 s 88454 161370 88934 161490 6 mgmt_wdata[18]
port 125 nsew default input
rlabel metal3 s 88454 162594 88934 162714 6 mgmt_wdata[19]
port 126 nsew default input
rlabel metal3 s 88454 140970 88934 141090 6 mgmt_wdata[1]
port 127 nsew default input
rlabel metal3 s 88454 163818 88934 163938 6 mgmt_wdata[20]
port 128 nsew default input
rlabel metal3 s 88454 165042 88934 165162 6 mgmt_wdata[21]
port 129 nsew default input
rlabel metal3 s 88454 166266 88934 166386 6 mgmt_wdata[22]
port 130 nsew default input
rlabel metal3 s 88454 167490 88934 167610 6 mgmt_wdata[23]
port 131 nsew default input
rlabel metal3 s 88454 168578 88934 168698 6 mgmt_wdata[24]
port 132 nsew default input
rlabel metal3 s 88454 169802 88934 169922 6 mgmt_wdata[25]
port 133 nsew default input
rlabel metal3 s 88454 171026 88934 171146 6 mgmt_wdata[26]
port 134 nsew default input
rlabel metal3 s 88454 172250 88934 172370 6 mgmt_wdata[27]
port 135 nsew default input
rlabel metal3 s 88454 173474 88934 173594 6 mgmt_wdata[28]
port 136 nsew default input
rlabel metal3 s 88454 174698 88934 174818 6 mgmt_wdata[29]
port 137 nsew default input
rlabel metal3 s 88454 142194 88934 142314 6 mgmt_wdata[2]
port 138 nsew default input
rlabel metal3 s 88454 175786 88934 175906 6 mgmt_wdata[30]
port 139 nsew default input
rlabel metal3 s 88454 177010 88934 177130 6 mgmt_wdata[31]
port 140 nsew default input
rlabel metal3 s 88454 143418 88934 143538 6 mgmt_wdata[3]
port 141 nsew default input
rlabel metal3 s 88454 144642 88934 144762 6 mgmt_wdata[4]
port 142 nsew default input
rlabel metal3 s 88454 145730 88934 145850 6 mgmt_wdata[5]
port 143 nsew default input
rlabel metal3 s 88454 146954 88934 147074 6 mgmt_wdata[6]
port 144 nsew default input
rlabel metal3 s 88454 148178 88934 148298 6 mgmt_wdata[7]
port 145 nsew default input
rlabel metal3 s 88454 149402 88934 149522 6 mgmt_wdata[8]
port 146 nsew default input
rlabel metal3 s 88454 150626 88934 150746 6 mgmt_wdata[9]
port 147 nsew default input
rlabel metal3 s 88454 178234 88934 178354 6 mgmt_wen[0]
port 148 nsew default input
rlabel metal3 s 88454 179458 88934 179578 6 mgmt_wen[1]
port 149 nsew default input
rlabel metal3 s 88454 180682 88934 180802 6 mgmt_wen_mask[0]
port 150 nsew default input
rlabel metal3 s 88454 181906 88934 182026 6 mgmt_wen_mask[1]
port 151 nsew default input
rlabel metal3 s 88454 182994 88934 183114 6 mgmt_wen_mask[2]
port 152 nsew default input
rlabel metal3 s 88454 184218 88934 184338 6 mgmt_wen_mask[3]
port 153 nsew default input
rlabel metal3 s 88454 185442 88934 185562 6 mgmt_wen_mask[4]
port 154 nsew default input
rlabel metal3 s 88454 186666 88934 186786 6 mgmt_wen_mask[5]
port 155 nsew default input
rlabel metal3 s 88454 187890 88934 188010 6 mgmt_wen_mask[6]
port 156 nsew default input
rlabel metal3 s 88454 189114 88934 189234 6 mgmt_wen_mask[7]
port 157 nsew default input
rlabel metal5 s 38 5092 87806 5412 6 VPWR
port 158 nsew default input
rlabel metal5 s 38 10092 87806 10412 6 VGND
port 159 nsew default input
<< properties >>
string FIXED_BBOX 0 0 88934 189234
<< end >>
