caravel.cdl.NG.unfolded.no.empty