magic
tech sky130A
magscale 1 2
timestamp 1606421840
<< error_p >>
rect -3510 799 -3452 805
rect -3392 799 -3334 805
rect -3274 799 -3216 805
rect -3156 799 -3098 805
rect -3038 799 -2980 805
rect -2920 799 -2862 805
rect -2802 799 -2744 805
rect -2684 799 -2626 805
rect -2566 799 -2508 805
rect -2448 799 -2390 805
rect -2330 799 -2272 805
rect -2212 799 -2154 805
rect -2094 799 -2036 805
rect -1976 799 -1918 805
rect -1858 799 -1800 805
rect -1740 799 -1682 805
rect -1622 799 -1564 805
rect -1504 799 -1446 805
rect -1386 799 -1328 805
rect -1268 799 -1210 805
rect -1150 799 -1092 805
rect -1032 799 -974 805
rect -914 799 -856 805
rect -796 799 -738 805
rect -678 799 -620 805
rect -560 799 -502 805
rect -442 799 -384 805
rect -324 799 -266 805
rect -206 799 -148 805
rect -88 799 -30 805
rect 30 799 88 805
rect 148 799 206 805
rect 266 799 324 805
rect 384 799 442 805
rect 502 799 560 805
rect 620 799 678 805
rect 738 799 796 805
rect 856 799 914 805
rect 974 799 1032 805
rect 1092 799 1150 805
rect 1210 799 1268 805
rect 1328 799 1386 805
rect 1446 799 1504 805
rect 1564 799 1622 805
rect 1682 799 1740 805
rect 1800 799 1858 805
rect 1918 799 1976 805
rect 2036 799 2094 805
rect 2154 799 2212 805
rect 2272 799 2330 805
rect 2390 799 2448 805
rect 2508 799 2566 805
rect 2626 799 2684 805
rect 2744 799 2802 805
rect 2862 799 2920 805
rect 2980 799 3038 805
rect 3098 799 3156 805
rect 3216 799 3274 805
rect 3334 799 3392 805
rect 3452 799 3510 805
rect -3510 765 -3498 799
rect -3392 765 -3380 799
rect -3274 765 -3262 799
rect -3156 765 -3144 799
rect -3038 765 -3026 799
rect -2920 765 -2908 799
rect -2802 765 -2790 799
rect -2684 765 -2672 799
rect -2566 765 -2554 799
rect -2448 765 -2436 799
rect -2330 765 -2318 799
rect -2212 765 -2200 799
rect -2094 765 -2082 799
rect -1976 765 -1964 799
rect -1858 765 -1846 799
rect -1740 765 -1728 799
rect -1622 765 -1610 799
rect -1504 765 -1492 799
rect -1386 765 -1374 799
rect -1268 765 -1256 799
rect -1150 765 -1138 799
rect -1032 765 -1020 799
rect -914 765 -902 799
rect -796 765 -784 799
rect -678 765 -666 799
rect -560 765 -548 799
rect -442 765 -430 799
rect -324 765 -312 799
rect -206 765 -194 799
rect -88 765 -76 799
rect 30 765 42 799
rect 148 765 160 799
rect 266 765 278 799
rect 384 765 396 799
rect 502 765 514 799
rect 620 765 632 799
rect 738 765 750 799
rect 856 765 868 799
rect 974 765 986 799
rect 1092 765 1104 799
rect 1210 765 1222 799
rect 1328 765 1340 799
rect 1446 765 1458 799
rect 1564 765 1576 799
rect 1682 765 1694 799
rect 1800 765 1812 799
rect 1918 765 1930 799
rect 2036 765 2048 799
rect 2154 765 2166 799
rect 2272 765 2284 799
rect 2390 765 2402 799
rect 2508 765 2520 799
rect 2626 765 2638 799
rect 2744 765 2756 799
rect 2862 765 2874 799
rect 2980 765 2992 799
rect 3098 765 3110 799
rect 3216 765 3228 799
rect 3334 765 3346 799
rect 3452 765 3464 799
rect -3510 759 -3452 765
rect -3392 759 -3334 765
rect -3274 759 -3216 765
rect -3156 759 -3098 765
rect -3038 759 -2980 765
rect -2920 759 -2862 765
rect -2802 759 -2744 765
rect -2684 759 -2626 765
rect -2566 759 -2508 765
rect -2448 759 -2390 765
rect -2330 759 -2272 765
rect -2212 759 -2154 765
rect -2094 759 -2036 765
rect -1976 759 -1918 765
rect -1858 759 -1800 765
rect -1740 759 -1682 765
rect -1622 759 -1564 765
rect -1504 759 -1446 765
rect -1386 759 -1328 765
rect -1268 759 -1210 765
rect -1150 759 -1092 765
rect -1032 759 -974 765
rect -914 759 -856 765
rect -796 759 -738 765
rect -678 759 -620 765
rect -560 759 -502 765
rect -442 759 -384 765
rect -324 759 -266 765
rect -206 759 -148 765
rect -88 759 -30 765
rect 30 759 88 765
rect 148 759 206 765
rect 266 759 324 765
rect 384 759 442 765
rect 502 759 560 765
rect 620 759 678 765
rect 738 759 796 765
rect 856 759 914 765
rect 974 759 1032 765
rect 1092 759 1150 765
rect 1210 759 1268 765
rect 1328 759 1386 765
rect 1446 759 1504 765
rect 1564 759 1622 765
rect 1682 759 1740 765
rect 1800 759 1858 765
rect 1918 759 1976 765
rect 2036 759 2094 765
rect 2154 759 2212 765
rect 2272 759 2330 765
rect 2390 759 2448 765
rect 2508 759 2566 765
rect 2626 759 2684 765
rect 2744 759 2802 765
rect 2862 759 2920 765
rect 2980 759 3038 765
rect 3098 759 3156 765
rect 3216 759 3274 765
rect 3334 759 3392 765
rect 3452 759 3510 765
rect -3510 71 -3452 77
rect -3392 71 -3334 77
rect -3274 71 -3216 77
rect -3156 71 -3098 77
rect -3038 71 -2980 77
rect -2920 71 -2862 77
rect -2802 71 -2744 77
rect -2684 71 -2626 77
rect -2566 71 -2508 77
rect -2448 71 -2390 77
rect -2330 71 -2272 77
rect -2212 71 -2154 77
rect -2094 71 -2036 77
rect -1976 71 -1918 77
rect -1858 71 -1800 77
rect -1740 71 -1682 77
rect -1622 71 -1564 77
rect -1504 71 -1446 77
rect -1386 71 -1328 77
rect -1268 71 -1210 77
rect -1150 71 -1092 77
rect -1032 71 -974 77
rect -914 71 -856 77
rect -796 71 -738 77
rect -678 71 -620 77
rect -560 71 -502 77
rect -442 71 -384 77
rect -324 71 -266 77
rect -206 71 -148 77
rect -88 71 -30 77
rect 30 71 88 77
rect 148 71 206 77
rect 266 71 324 77
rect 384 71 442 77
rect 502 71 560 77
rect 620 71 678 77
rect 738 71 796 77
rect 856 71 914 77
rect 974 71 1032 77
rect 1092 71 1150 77
rect 1210 71 1268 77
rect 1328 71 1386 77
rect 1446 71 1504 77
rect 1564 71 1622 77
rect 1682 71 1740 77
rect 1800 71 1858 77
rect 1918 71 1976 77
rect 2036 71 2094 77
rect 2154 71 2212 77
rect 2272 71 2330 77
rect 2390 71 2448 77
rect 2508 71 2566 77
rect 2626 71 2684 77
rect 2744 71 2802 77
rect 2862 71 2920 77
rect 2980 71 3038 77
rect 3098 71 3156 77
rect 3216 71 3274 77
rect 3334 71 3392 77
rect 3452 71 3510 77
rect -3510 37 -3498 71
rect -3392 37 -3380 71
rect -3274 37 -3262 71
rect -3156 37 -3144 71
rect -3038 37 -3026 71
rect -2920 37 -2908 71
rect -2802 37 -2790 71
rect -2684 37 -2672 71
rect -2566 37 -2554 71
rect -2448 37 -2436 71
rect -2330 37 -2318 71
rect -2212 37 -2200 71
rect -2094 37 -2082 71
rect -1976 37 -1964 71
rect -1858 37 -1846 71
rect -1740 37 -1728 71
rect -1622 37 -1610 71
rect -1504 37 -1492 71
rect -1386 37 -1374 71
rect -1268 37 -1256 71
rect -1150 37 -1138 71
rect -1032 37 -1020 71
rect -914 37 -902 71
rect -796 37 -784 71
rect -678 37 -666 71
rect -560 37 -548 71
rect -442 37 -430 71
rect -324 37 -312 71
rect -206 37 -194 71
rect -88 37 -76 71
rect 30 37 42 71
rect 148 37 160 71
rect 266 37 278 71
rect 384 37 396 71
rect 502 37 514 71
rect 620 37 632 71
rect 738 37 750 71
rect 856 37 868 71
rect 974 37 986 71
rect 1092 37 1104 71
rect 1210 37 1222 71
rect 1328 37 1340 71
rect 1446 37 1458 71
rect 1564 37 1576 71
rect 1682 37 1694 71
rect 1800 37 1812 71
rect 1918 37 1930 71
rect 2036 37 2048 71
rect 2154 37 2166 71
rect 2272 37 2284 71
rect 2390 37 2402 71
rect 2508 37 2520 71
rect 2626 37 2638 71
rect 2744 37 2756 71
rect 2862 37 2874 71
rect 2980 37 2992 71
rect 3098 37 3110 71
rect 3216 37 3228 71
rect 3334 37 3346 71
rect 3452 37 3464 71
rect -3510 31 -3452 37
rect -3392 31 -3334 37
rect -3274 31 -3216 37
rect -3156 31 -3098 37
rect -3038 31 -2980 37
rect -2920 31 -2862 37
rect -2802 31 -2744 37
rect -2684 31 -2626 37
rect -2566 31 -2508 37
rect -2448 31 -2390 37
rect -2330 31 -2272 37
rect -2212 31 -2154 37
rect -2094 31 -2036 37
rect -1976 31 -1918 37
rect -1858 31 -1800 37
rect -1740 31 -1682 37
rect -1622 31 -1564 37
rect -1504 31 -1446 37
rect -1386 31 -1328 37
rect -1268 31 -1210 37
rect -1150 31 -1092 37
rect -1032 31 -974 37
rect -914 31 -856 37
rect -796 31 -738 37
rect -678 31 -620 37
rect -560 31 -502 37
rect -442 31 -384 37
rect -324 31 -266 37
rect -206 31 -148 37
rect -88 31 -30 37
rect 30 31 88 37
rect 148 31 206 37
rect 266 31 324 37
rect 384 31 442 37
rect 502 31 560 37
rect 620 31 678 37
rect 738 31 796 37
rect 856 31 914 37
rect 974 31 1032 37
rect 1092 31 1150 37
rect 1210 31 1268 37
rect 1328 31 1386 37
rect 1446 31 1504 37
rect 1564 31 1622 37
rect 1682 31 1740 37
rect 1800 31 1858 37
rect 1918 31 1976 37
rect 2036 31 2094 37
rect 2154 31 2212 37
rect 2272 31 2330 37
rect 2390 31 2448 37
rect 2508 31 2566 37
rect 2626 31 2684 37
rect 2744 31 2802 37
rect 2862 31 2920 37
rect 2980 31 3038 37
rect 3098 31 3156 37
rect 3216 31 3274 37
rect 3334 31 3392 37
rect 3452 31 3510 37
rect -3510 -37 -3452 -31
rect -3392 -37 -3334 -31
rect -3274 -37 -3216 -31
rect -3156 -37 -3098 -31
rect -3038 -37 -2980 -31
rect -2920 -37 -2862 -31
rect -2802 -37 -2744 -31
rect -2684 -37 -2626 -31
rect -2566 -37 -2508 -31
rect -2448 -37 -2390 -31
rect -2330 -37 -2272 -31
rect -2212 -37 -2154 -31
rect -2094 -37 -2036 -31
rect -1976 -37 -1918 -31
rect -1858 -37 -1800 -31
rect -1740 -37 -1682 -31
rect -1622 -37 -1564 -31
rect -1504 -37 -1446 -31
rect -1386 -37 -1328 -31
rect -1268 -37 -1210 -31
rect -1150 -37 -1092 -31
rect -1032 -37 -974 -31
rect -914 -37 -856 -31
rect -796 -37 -738 -31
rect -678 -37 -620 -31
rect -560 -37 -502 -31
rect -442 -37 -384 -31
rect -324 -37 -266 -31
rect -206 -37 -148 -31
rect -88 -37 -30 -31
rect 30 -37 88 -31
rect 148 -37 206 -31
rect 266 -37 324 -31
rect 384 -37 442 -31
rect 502 -37 560 -31
rect 620 -37 678 -31
rect 738 -37 796 -31
rect 856 -37 914 -31
rect 974 -37 1032 -31
rect 1092 -37 1150 -31
rect 1210 -37 1268 -31
rect 1328 -37 1386 -31
rect 1446 -37 1504 -31
rect 1564 -37 1622 -31
rect 1682 -37 1740 -31
rect 1800 -37 1858 -31
rect 1918 -37 1976 -31
rect 2036 -37 2094 -31
rect 2154 -37 2212 -31
rect 2272 -37 2330 -31
rect 2390 -37 2448 -31
rect 2508 -37 2566 -31
rect 2626 -37 2684 -31
rect 2744 -37 2802 -31
rect 2862 -37 2920 -31
rect 2980 -37 3038 -31
rect 3098 -37 3156 -31
rect 3216 -37 3274 -31
rect 3334 -37 3392 -31
rect 3452 -37 3510 -31
rect -3510 -71 -3498 -37
rect -3392 -71 -3380 -37
rect -3274 -71 -3262 -37
rect -3156 -71 -3144 -37
rect -3038 -71 -3026 -37
rect -2920 -71 -2908 -37
rect -2802 -71 -2790 -37
rect -2684 -71 -2672 -37
rect -2566 -71 -2554 -37
rect -2448 -71 -2436 -37
rect -2330 -71 -2318 -37
rect -2212 -71 -2200 -37
rect -2094 -71 -2082 -37
rect -1976 -71 -1964 -37
rect -1858 -71 -1846 -37
rect -1740 -71 -1728 -37
rect -1622 -71 -1610 -37
rect -1504 -71 -1492 -37
rect -1386 -71 -1374 -37
rect -1268 -71 -1256 -37
rect -1150 -71 -1138 -37
rect -1032 -71 -1020 -37
rect -914 -71 -902 -37
rect -796 -71 -784 -37
rect -678 -71 -666 -37
rect -560 -71 -548 -37
rect -442 -71 -430 -37
rect -324 -71 -312 -37
rect -206 -71 -194 -37
rect -88 -71 -76 -37
rect 30 -71 42 -37
rect 148 -71 160 -37
rect 266 -71 278 -37
rect 384 -71 396 -37
rect 502 -71 514 -37
rect 620 -71 632 -37
rect 738 -71 750 -37
rect 856 -71 868 -37
rect 974 -71 986 -37
rect 1092 -71 1104 -37
rect 1210 -71 1222 -37
rect 1328 -71 1340 -37
rect 1446 -71 1458 -37
rect 1564 -71 1576 -37
rect 1682 -71 1694 -37
rect 1800 -71 1812 -37
rect 1918 -71 1930 -37
rect 2036 -71 2048 -37
rect 2154 -71 2166 -37
rect 2272 -71 2284 -37
rect 2390 -71 2402 -37
rect 2508 -71 2520 -37
rect 2626 -71 2638 -37
rect 2744 -71 2756 -37
rect 2862 -71 2874 -37
rect 2980 -71 2992 -37
rect 3098 -71 3110 -37
rect 3216 -71 3228 -37
rect 3334 -71 3346 -37
rect 3452 -71 3464 -37
rect -3510 -77 -3452 -71
rect -3392 -77 -3334 -71
rect -3274 -77 -3216 -71
rect -3156 -77 -3098 -71
rect -3038 -77 -2980 -71
rect -2920 -77 -2862 -71
rect -2802 -77 -2744 -71
rect -2684 -77 -2626 -71
rect -2566 -77 -2508 -71
rect -2448 -77 -2390 -71
rect -2330 -77 -2272 -71
rect -2212 -77 -2154 -71
rect -2094 -77 -2036 -71
rect -1976 -77 -1918 -71
rect -1858 -77 -1800 -71
rect -1740 -77 -1682 -71
rect -1622 -77 -1564 -71
rect -1504 -77 -1446 -71
rect -1386 -77 -1328 -71
rect -1268 -77 -1210 -71
rect -1150 -77 -1092 -71
rect -1032 -77 -974 -71
rect -914 -77 -856 -71
rect -796 -77 -738 -71
rect -678 -77 -620 -71
rect -560 -77 -502 -71
rect -442 -77 -384 -71
rect -324 -77 -266 -71
rect -206 -77 -148 -71
rect -88 -77 -30 -71
rect 30 -77 88 -71
rect 148 -77 206 -71
rect 266 -77 324 -71
rect 384 -77 442 -71
rect 502 -77 560 -71
rect 620 -77 678 -71
rect 738 -77 796 -71
rect 856 -77 914 -71
rect 974 -77 1032 -71
rect 1092 -77 1150 -71
rect 1210 -77 1268 -71
rect 1328 -77 1386 -71
rect 1446 -77 1504 -71
rect 1564 -77 1622 -71
rect 1682 -77 1740 -71
rect 1800 -77 1858 -71
rect 1918 -77 1976 -71
rect 2036 -77 2094 -71
rect 2154 -77 2212 -71
rect 2272 -77 2330 -71
rect 2390 -77 2448 -71
rect 2508 -77 2566 -71
rect 2626 -77 2684 -71
rect 2744 -77 2802 -71
rect 2862 -77 2920 -71
rect 2980 -77 3038 -71
rect 3098 -77 3156 -71
rect 3216 -77 3274 -71
rect 3334 -77 3392 -71
rect 3452 -77 3510 -71
rect -3510 -765 -3452 -759
rect -3392 -765 -3334 -759
rect -3274 -765 -3216 -759
rect -3156 -765 -3098 -759
rect -3038 -765 -2980 -759
rect -2920 -765 -2862 -759
rect -2802 -765 -2744 -759
rect -2684 -765 -2626 -759
rect -2566 -765 -2508 -759
rect -2448 -765 -2390 -759
rect -2330 -765 -2272 -759
rect -2212 -765 -2154 -759
rect -2094 -765 -2036 -759
rect -1976 -765 -1918 -759
rect -1858 -765 -1800 -759
rect -1740 -765 -1682 -759
rect -1622 -765 -1564 -759
rect -1504 -765 -1446 -759
rect -1386 -765 -1328 -759
rect -1268 -765 -1210 -759
rect -1150 -765 -1092 -759
rect -1032 -765 -974 -759
rect -914 -765 -856 -759
rect -796 -765 -738 -759
rect -678 -765 -620 -759
rect -560 -765 -502 -759
rect -442 -765 -384 -759
rect -324 -765 -266 -759
rect -206 -765 -148 -759
rect -88 -765 -30 -759
rect 30 -765 88 -759
rect 148 -765 206 -759
rect 266 -765 324 -759
rect 384 -765 442 -759
rect 502 -765 560 -759
rect 620 -765 678 -759
rect 738 -765 796 -759
rect 856 -765 914 -759
rect 974 -765 1032 -759
rect 1092 -765 1150 -759
rect 1210 -765 1268 -759
rect 1328 -765 1386 -759
rect 1446 -765 1504 -759
rect 1564 -765 1622 -759
rect 1682 -765 1740 -759
rect 1800 -765 1858 -759
rect 1918 -765 1976 -759
rect 2036 -765 2094 -759
rect 2154 -765 2212 -759
rect 2272 -765 2330 -759
rect 2390 -765 2448 -759
rect 2508 -765 2566 -759
rect 2626 -765 2684 -759
rect 2744 -765 2802 -759
rect 2862 -765 2920 -759
rect 2980 -765 3038 -759
rect 3098 -765 3156 -759
rect 3216 -765 3274 -759
rect 3334 -765 3392 -759
rect 3452 -765 3510 -759
rect -3510 -799 -3498 -765
rect -3392 -799 -3380 -765
rect -3274 -799 -3262 -765
rect -3156 -799 -3144 -765
rect -3038 -799 -3026 -765
rect -2920 -799 -2908 -765
rect -2802 -799 -2790 -765
rect -2684 -799 -2672 -765
rect -2566 -799 -2554 -765
rect -2448 -799 -2436 -765
rect -2330 -799 -2318 -765
rect -2212 -799 -2200 -765
rect -2094 -799 -2082 -765
rect -1976 -799 -1964 -765
rect -1858 -799 -1846 -765
rect -1740 -799 -1728 -765
rect -1622 -799 -1610 -765
rect -1504 -799 -1492 -765
rect -1386 -799 -1374 -765
rect -1268 -799 -1256 -765
rect -1150 -799 -1138 -765
rect -1032 -799 -1020 -765
rect -914 -799 -902 -765
rect -796 -799 -784 -765
rect -678 -799 -666 -765
rect -560 -799 -548 -765
rect -442 -799 -430 -765
rect -324 -799 -312 -765
rect -206 -799 -194 -765
rect -88 -799 -76 -765
rect 30 -799 42 -765
rect 148 -799 160 -765
rect 266 -799 278 -765
rect 384 -799 396 -765
rect 502 -799 514 -765
rect 620 -799 632 -765
rect 738 -799 750 -765
rect 856 -799 868 -765
rect 974 -799 986 -765
rect 1092 -799 1104 -765
rect 1210 -799 1222 -765
rect 1328 -799 1340 -765
rect 1446 -799 1458 -765
rect 1564 -799 1576 -765
rect 1682 -799 1694 -765
rect 1800 -799 1812 -765
rect 1918 -799 1930 -765
rect 2036 -799 2048 -765
rect 2154 -799 2166 -765
rect 2272 -799 2284 -765
rect 2390 -799 2402 -765
rect 2508 -799 2520 -765
rect 2626 -799 2638 -765
rect 2744 -799 2756 -765
rect 2862 -799 2874 -765
rect 2980 -799 2992 -765
rect 3098 -799 3110 -765
rect 3216 -799 3228 -765
rect 3334 -799 3346 -765
rect 3452 -799 3464 -765
rect -3510 -805 -3452 -799
rect -3392 -805 -3334 -799
rect -3274 -805 -3216 -799
rect -3156 -805 -3098 -799
rect -3038 -805 -2980 -799
rect -2920 -805 -2862 -799
rect -2802 -805 -2744 -799
rect -2684 -805 -2626 -799
rect -2566 -805 -2508 -799
rect -2448 -805 -2390 -799
rect -2330 -805 -2272 -799
rect -2212 -805 -2154 -799
rect -2094 -805 -2036 -799
rect -1976 -805 -1918 -799
rect -1858 -805 -1800 -799
rect -1740 -805 -1682 -799
rect -1622 -805 -1564 -799
rect -1504 -805 -1446 -799
rect -1386 -805 -1328 -799
rect -1268 -805 -1210 -799
rect -1150 -805 -1092 -799
rect -1032 -805 -974 -799
rect -914 -805 -856 -799
rect -796 -805 -738 -799
rect -678 -805 -620 -799
rect -560 -805 -502 -799
rect -442 -805 -384 -799
rect -324 -805 -266 -799
rect -206 -805 -148 -799
rect -88 -805 -30 -799
rect 30 -805 88 -799
rect 148 -805 206 -799
rect 266 -805 324 -799
rect 384 -805 442 -799
rect 502 -805 560 -799
rect 620 -805 678 -799
rect 738 -805 796 -799
rect 856 -805 914 -799
rect 974 -805 1032 -799
rect 1092 -805 1150 -799
rect 1210 -805 1268 -799
rect 1328 -805 1386 -799
rect 1446 -805 1504 -799
rect 1564 -805 1622 -799
rect 1682 -805 1740 -799
rect 1800 -805 1858 -799
rect 1918 -805 1976 -799
rect 2036 -805 2094 -799
rect 2154 -805 2212 -799
rect 2272 -805 2330 -799
rect 2390 -805 2448 -799
rect 2508 -805 2566 -799
rect 2626 -805 2684 -799
rect 2744 -805 2802 -799
rect 2862 -805 2920 -799
rect 2980 -805 3038 -799
rect 3098 -805 3156 -799
rect 3216 -805 3274 -799
rect 3334 -805 3392 -799
rect 3452 -805 3510 -799
<< nwell >>
rect -3707 -937 3707 937
<< pmos >>
rect -3511 118 -3451 718
rect -3393 118 -3333 718
rect -3275 118 -3215 718
rect -3157 118 -3097 718
rect -3039 118 -2979 718
rect -2921 118 -2861 718
rect -2803 118 -2743 718
rect -2685 118 -2625 718
rect -2567 118 -2507 718
rect -2449 118 -2389 718
rect -2331 118 -2271 718
rect -2213 118 -2153 718
rect -2095 118 -2035 718
rect -1977 118 -1917 718
rect -1859 118 -1799 718
rect -1741 118 -1681 718
rect -1623 118 -1563 718
rect -1505 118 -1445 718
rect -1387 118 -1327 718
rect -1269 118 -1209 718
rect -1151 118 -1091 718
rect -1033 118 -973 718
rect -915 118 -855 718
rect -797 118 -737 718
rect -679 118 -619 718
rect -561 118 -501 718
rect -443 118 -383 718
rect -325 118 -265 718
rect -207 118 -147 718
rect -89 118 -29 718
rect 29 118 89 718
rect 147 118 207 718
rect 265 118 325 718
rect 383 118 443 718
rect 501 118 561 718
rect 619 118 679 718
rect 737 118 797 718
rect 855 118 915 718
rect 973 118 1033 718
rect 1091 118 1151 718
rect 1209 118 1269 718
rect 1327 118 1387 718
rect 1445 118 1505 718
rect 1563 118 1623 718
rect 1681 118 1741 718
rect 1799 118 1859 718
rect 1917 118 1977 718
rect 2035 118 2095 718
rect 2153 118 2213 718
rect 2271 118 2331 718
rect 2389 118 2449 718
rect 2507 118 2567 718
rect 2625 118 2685 718
rect 2743 118 2803 718
rect 2861 118 2921 718
rect 2979 118 3039 718
rect 3097 118 3157 718
rect 3215 118 3275 718
rect 3333 118 3393 718
rect 3451 118 3511 718
rect -3511 -718 -3451 -118
rect -3393 -718 -3333 -118
rect -3275 -718 -3215 -118
rect -3157 -718 -3097 -118
rect -3039 -718 -2979 -118
rect -2921 -718 -2861 -118
rect -2803 -718 -2743 -118
rect -2685 -718 -2625 -118
rect -2567 -718 -2507 -118
rect -2449 -718 -2389 -118
rect -2331 -718 -2271 -118
rect -2213 -718 -2153 -118
rect -2095 -718 -2035 -118
rect -1977 -718 -1917 -118
rect -1859 -718 -1799 -118
rect -1741 -718 -1681 -118
rect -1623 -718 -1563 -118
rect -1505 -718 -1445 -118
rect -1387 -718 -1327 -118
rect -1269 -718 -1209 -118
rect -1151 -718 -1091 -118
rect -1033 -718 -973 -118
rect -915 -718 -855 -118
rect -797 -718 -737 -118
rect -679 -718 -619 -118
rect -561 -718 -501 -118
rect -443 -718 -383 -118
rect -325 -718 -265 -118
rect -207 -718 -147 -118
rect -89 -718 -29 -118
rect 29 -718 89 -118
rect 147 -718 207 -118
rect 265 -718 325 -118
rect 383 -718 443 -118
rect 501 -718 561 -118
rect 619 -718 679 -118
rect 737 -718 797 -118
rect 855 -718 915 -118
rect 973 -718 1033 -118
rect 1091 -718 1151 -118
rect 1209 -718 1269 -118
rect 1327 -718 1387 -118
rect 1445 -718 1505 -118
rect 1563 -718 1623 -118
rect 1681 -718 1741 -118
rect 1799 -718 1859 -118
rect 1917 -718 1977 -118
rect 2035 -718 2095 -118
rect 2153 -718 2213 -118
rect 2271 -718 2331 -118
rect 2389 -718 2449 -118
rect 2507 -718 2567 -118
rect 2625 -718 2685 -118
rect 2743 -718 2803 -118
rect 2861 -718 2921 -118
rect 2979 -718 3039 -118
rect 3097 -718 3157 -118
rect 3215 -718 3275 -118
rect 3333 -718 3393 -118
rect 3451 -718 3511 -118
<< pdiff >>
rect -3569 706 -3511 718
rect -3569 130 -3557 706
rect -3523 130 -3511 706
rect -3569 118 -3511 130
rect -3451 706 -3393 718
rect -3451 130 -3439 706
rect -3405 130 -3393 706
rect -3451 118 -3393 130
rect -3333 706 -3275 718
rect -3333 130 -3321 706
rect -3287 130 -3275 706
rect -3333 118 -3275 130
rect -3215 706 -3157 718
rect -3215 130 -3203 706
rect -3169 130 -3157 706
rect -3215 118 -3157 130
rect -3097 706 -3039 718
rect -3097 130 -3085 706
rect -3051 130 -3039 706
rect -3097 118 -3039 130
rect -2979 706 -2921 718
rect -2979 130 -2967 706
rect -2933 130 -2921 706
rect -2979 118 -2921 130
rect -2861 706 -2803 718
rect -2861 130 -2849 706
rect -2815 130 -2803 706
rect -2861 118 -2803 130
rect -2743 706 -2685 718
rect -2743 130 -2731 706
rect -2697 130 -2685 706
rect -2743 118 -2685 130
rect -2625 706 -2567 718
rect -2625 130 -2613 706
rect -2579 130 -2567 706
rect -2625 118 -2567 130
rect -2507 706 -2449 718
rect -2507 130 -2495 706
rect -2461 130 -2449 706
rect -2507 118 -2449 130
rect -2389 706 -2331 718
rect -2389 130 -2377 706
rect -2343 130 -2331 706
rect -2389 118 -2331 130
rect -2271 706 -2213 718
rect -2271 130 -2259 706
rect -2225 130 -2213 706
rect -2271 118 -2213 130
rect -2153 706 -2095 718
rect -2153 130 -2141 706
rect -2107 130 -2095 706
rect -2153 118 -2095 130
rect -2035 706 -1977 718
rect -2035 130 -2023 706
rect -1989 130 -1977 706
rect -2035 118 -1977 130
rect -1917 706 -1859 718
rect -1917 130 -1905 706
rect -1871 130 -1859 706
rect -1917 118 -1859 130
rect -1799 706 -1741 718
rect -1799 130 -1787 706
rect -1753 130 -1741 706
rect -1799 118 -1741 130
rect -1681 706 -1623 718
rect -1681 130 -1669 706
rect -1635 130 -1623 706
rect -1681 118 -1623 130
rect -1563 706 -1505 718
rect -1563 130 -1551 706
rect -1517 130 -1505 706
rect -1563 118 -1505 130
rect -1445 706 -1387 718
rect -1445 130 -1433 706
rect -1399 130 -1387 706
rect -1445 118 -1387 130
rect -1327 706 -1269 718
rect -1327 130 -1315 706
rect -1281 130 -1269 706
rect -1327 118 -1269 130
rect -1209 706 -1151 718
rect -1209 130 -1197 706
rect -1163 130 -1151 706
rect -1209 118 -1151 130
rect -1091 706 -1033 718
rect -1091 130 -1079 706
rect -1045 130 -1033 706
rect -1091 118 -1033 130
rect -973 706 -915 718
rect -973 130 -961 706
rect -927 130 -915 706
rect -973 118 -915 130
rect -855 706 -797 718
rect -855 130 -843 706
rect -809 130 -797 706
rect -855 118 -797 130
rect -737 706 -679 718
rect -737 130 -725 706
rect -691 130 -679 706
rect -737 118 -679 130
rect -619 706 -561 718
rect -619 130 -607 706
rect -573 130 -561 706
rect -619 118 -561 130
rect -501 706 -443 718
rect -501 130 -489 706
rect -455 130 -443 706
rect -501 118 -443 130
rect -383 706 -325 718
rect -383 130 -371 706
rect -337 130 -325 706
rect -383 118 -325 130
rect -265 706 -207 718
rect -265 130 -253 706
rect -219 130 -207 706
rect -265 118 -207 130
rect -147 706 -89 718
rect -147 130 -135 706
rect -101 130 -89 706
rect -147 118 -89 130
rect -29 706 29 718
rect -29 130 -17 706
rect 17 130 29 706
rect -29 118 29 130
rect 89 706 147 718
rect 89 130 101 706
rect 135 130 147 706
rect 89 118 147 130
rect 207 706 265 718
rect 207 130 219 706
rect 253 130 265 706
rect 207 118 265 130
rect 325 706 383 718
rect 325 130 337 706
rect 371 130 383 706
rect 325 118 383 130
rect 443 706 501 718
rect 443 130 455 706
rect 489 130 501 706
rect 443 118 501 130
rect 561 706 619 718
rect 561 130 573 706
rect 607 130 619 706
rect 561 118 619 130
rect 679 706 737 718
rect 679 130 691 706
rect 725 130 737 706
rect 679 118 737 130
rect 797 706 855 718
rect 797 130 809 706
rect 843 130 855 706
rect 797 118 855 130
rect 915 706 973 718
rect 915 130 927 706
rect 961 130 973 706
rect 915 118 973 130
rect 1033 706 1091 718
rect 1033 130 1045 706
rect 1079 130 1091 706
rect 1033 118 1091 130
rect 1151 706 1209 718
rect 1151 130 1163 706
rect 1197 130 1209 706
rect 1151 118 1209 130
rect 1269 706 1327 718
rect 1269 130 1281 706
rect 1315 130 1327 706
rect 1269 118 1327 130
rect 1387 706 1445 718
rect 1387 130 1399 706
rect 1433 130 1445 706
rect 1387 118 1445 130
rect 1505 706 1563 718
rect 1505 130 1517 706
rect 1551 130 1563 706
rect 1505 118 1563 130
rect 1623 706 1681 718
rect 1623 130 1635 706
rect 1669 130 1681 706
rect 1623 118 1681 130
rect 1741 706 1799 718
rect 1741 130 1753 706
rect 1787 130 1799 706
rect 1741 118 1799 130
rect 1859 706 1917 718
rect 1859 130 1871 706
rect 1905 130 1917 706
rect 1859 118 1917 130
rect 1977 706 2035 718
rect 1977 130 1989 706
rect 2023 130 2035 706
rect 1977 118 2035 130
rect 2095 706 2153 718
rect 2095 130 2107 706
rect 2141 130 2153 706
rect 2095 118 2153 130
rect 2213 706 2271 718
rect 2213 130 2225 706
rect 2259 130 2271 706
rect 2213 118 2271 130
rect 2331 706 2389 718
rect 2331 130 2343 706
rect 2377 130 2389 706
rect 2331 118 2389 130
rect 2449 706 2507 718
rect 2449 130 2461 706
rect 2495 130 2507 706
rect 2449 118 2507 130
rect 2567 706 2625 718
rect 2567 130 2579 706
rect 2613 130 2625 706
rect 2567 118 2625 130
rect 2685 706 2743 718
rect 2685 130 2697 706
rect 2731 130 2743 706
rect 2685 118 2743 130
rect 2803 706 2861 718
rect 2803 130 2815 706
rect 2849 130 2861 706
rect 2803 118 2861 130
rect 2921 706 2979 718
rect 2921 130 2933 706
rect 2967 130 2979 706
rect 2921 118 2979 130
rect 3039 706 3097 718
rect 3039 130 3051 706
rect 3085 130 3097 706
rect 3039 118 3097 130
rect 3157 706 3215 718
rect 3157 130 3169 706
rect 3203 130 3215 706
rect 3157 118 3215 130
rect 3275 706 3333 718
rect 3275 130 3287 706
rect 3321 130 3333 706
rect 3275 118 3333 130
rect 3393 706 3451 718
rect 3393 130 3405 706
rect 3439 130 3451 706
rect 3393 118 3451 130
rect 3511 706 3569 718
rect 3511 130 3523 706
rect 3557 130 3569 706
rect 3511 118 3569 130
rect -3569 -130 -3511 -118
rect -3569 -706 -3557 -130
rect -3523 -706 -3511 -130
rect -3569 -718 -3511 -706
rect -3451 -130 -3393 -118
rect -3451 -706 -3439 -130
rect -3405 -706 -3393 -130
rect -3451 -718 -3393 -706
rect -3333 -130 -3275 -118
rect -3333 -706 -3321 -130
rect -3287 -706 -3275 -130
rect -3333 -718 -3275 -706
rect -3215 -130 -3157 -118
rect -3215 -706 -3203 -130
rect -3169 -706 -3157 -130
rect -3215 -718 -3157 -706
rect -3097 -130 -3039 -118
rect -3097 -706 -3085 -130
rect -3051 -706 -3039 -130
rect -3097 -718 -3039 -706
rect -2979 -130 -2921 -118
rect -2979 -706 -2967 -130
rect -2933 -706 -2921 -130
rect -2979 -718 -2921 -706
rect -2861 -130 -2803 -118
rect -2861 -706 -2849 -130
rect -2815 -706 -2803 -130
rect -2861 -718 -2803 -706
rect -2743 -130 -2685 -118
rect -2743 -706 -2731 -130
rect -2697 -706 -2685 -130
rect -2743 -718 -2685 -706
rect -2625 -130 -2567 -118
rect -2625 -706 -2613 -130
rect -2579 -706 -2567 -130
rect -2625 -718 -2567 -706
rect -2507 -130 -2449 -118
rect -2507 -706 -2495 -130
rect -2461 -706 -2449 -130
rect -2507 -718 -2449 -706
rect -2389 -130 -2331 -118
rect -2389 -706 -2377 -130
rect -2343 -706 -2331 -130
rect -2389 -718 -2331 -706
rect -2271 -130 -2213 -118
rect -2271 -706 -2259 -130
rect -2225 -706 -2213 -130
rect -2271 -718 -2213 -706
rect -2153 -130 -2095 -118
rect -2153 -706 -2141 -130
rect -2107 -706 -2095 -130
rect -2153 -718 -2095 -706
rect -2035 -130 -1977 -118
rect -2035 -706 -2023 -130
rect -1989 -706 -1977 -130
rect -2035 -718 -1977 -706
rect -1917 -130 -1859 -118
rect -1917 -706 -1905 -130
rect -1871 -706 -1859 -130
rect -1917 -718 -1859 -706
rect -1799 -130 -1741 -118
rect -1799 -706 -1787 -130
rect -1753 -706 -1741 -130
rect -1799 -718 -1741 -706
rect -1681 -130 -1623 -118
rect -1681 -706 -1669 -130
rect -1635 -706 -1623 -130
rect -1681 -718 -1623 -706
rect -1563 -130 -1505 -118
rect -1563 -706 -1551 -130
rect -1517 -706 -1505 -130
rect -1563 -718 -1505 -706
rect -1445 -130 -1387 -118
rect -1445 -706 -1433 -130
rect -1399 -706 -1387 -130
rect -1445 -718 -1387 -706
rect -1327 -130 -1269 -118
rect -1327 -706 -1315 -130
rect -1281 -706 -1269 -130
rect -1327 -718 -1269 -706
rect -1209 -130 -1151 -118
rect -1209 -706 -1197 -130
rect -1163 -706 -1151 -130
rect -1209 -718 -1151 -706
rect -1091 -130 -1033 -118
rect -1091 -706 -1079 -130
rect -1045 -706 -1033 -130
rect -1091 -718 -1033 -706
rect -973 -130 -915 -118
rect -973 -706 -961 -130
rect -927 -706 -915 -130
rect -973 -718 -915 -706
rect -855 -130 -797 -118
rect -855 -706 -843 -130
rect -809 -706 -797 -130
rect -855 -718 -797 -706
rect -737 -130 -679 -118
rect -737 -706 -725 -130
rect -691 -706 -679 -130
rect -737 -718 -679 -706
rect -619 -130 -561 -118
rect -619 -706 -607 -130
rect -573 -706 -561 -130
rect -619 -718 -561 -706
rect -501 -130 -443 -118
rect -501 -706 -489 -130
rect -455 -706 -443 -130
rect -501 -718 -443 -706
rect -383 -130 -325 -118
rect -383 -706 -371 -130
rect -337 -706 -325 -130
rect -383 -718 -325 -706
rect -265 -130 -207 -118
rect -265 -706 -253 -130
rect -219 -706 -207 -130
rect -265 -718 -207 -706
rect -147 -130 -89 -118
rect -147 -706 -135 -130
rect -101 -706 -89 -130
rect -147 -718 -89 -706
rect -29 -130 29 -118
rect -29 -706 -17 -130
rect 17 -706 29 -130
rect -29 -718 29 -706
rect 89 -130 147 -118
rect 89 -706 101 -130
rect 135 -706 147 -130
rect 89 -718 147 -706
rect 207 -130 265 -118
rect 207 -706 219 -130
rect 253 -706 265 -130
rect 207 -718 265 -706
rect 325 -130 383 -118
rect 325 -706 337 -130
rect 371 -706 383 -130
rect 325 -718 383 -706
rect 443 -130 501 -118
rect 443 -706 455 -130
rect 489 -706 501 -130
rect 443 -718 501 -706
rect 561 -130 619 -118
rect 561 -706 573 -130
rect 607 -706 619 -130
rect 561 -718 619 -706
rect 679 -130 737 -118
rect 679 -706 691 -130
rect 725 -706 737 -130
rect 679 -718 737 -706
rect 797 -130 855 -118
rect 797 -706 809 -130
rect 843 -706 855 -130
rect 797 -718 855 -706
rect 915 -130 973 -118
rect 915 -706 927 -130
rect 961 -706 973 -130
rect 915 -718 973 -706
rect 1033 -130 1091 -118
rect 1033 -706 1045 -130
rect 1079 -706 1091 -130
rect 1033 -718 1091 -706
rect 1151 -130 1209 -118
rect 1151 -706 1163 -130
rect 1197 -706 1209 -130
rect 1151 -718 1209 -706
rect 1269 -130 1327 -118
rect 1269 -706 1281 -130
rect 1315 -706 1327 -130
rect 1269 -718 1327 -706
rect 1387 -130 1445 -118
rect 1387 -706 1399 -130
rect 1433 -706 1445 -130
rect 1387 -718 1445 -706
rect 1505 -130 1563 -118
rect 1505 -706 1517 -130
rect 1551 -706 1563 -130
rect 1505 -718 1563 -706
rect 1623 -130 1681 -118
rect 1623 -706 1635 -130
rect 1669 -706 1681 -130
rect 1623 -718 1681 -706
rect 1741 -130 1799 -118
rect 1741 -706 1753 -130
rect 1787 -706 1799 -130
rect 1741 -718 1799 -706
rect 1859 -130 1917 -118
rect 1859 -706 1871 -130
rect 1905 -706 1917 -130
rect 1859 -718 1917 -706
rect 1977 -130 2035 -118
rect 1977 -706 1989 -130
rect 2023 -706 2035 -130
rect 1977 -718 2035 -706
rect 2095 -130 2153 -118
rect 2095 -706 2107 -130
rect 2141 -706 2153 -130
rect 2095 -718 2153 -706
rect 2213 -130 2271 -118
rect 2213 -706 2225 -130
rect 2259 -706 2271 -130
rect 2213 -718 2271 -706
rect 2331 -130 2389 -118
rect 2331 -706 2343 -130
rect 2377 -706 2389 -130
rect 2331 -718 2389 -706
rect 2449 -130 2507 -118
rect 2449 -706 2461 -130
rect 2495 -706 2507 -130
rect 2449 -718 2507 -706
rect 2567 -130 2625 -118
rect 2567 -706 2579 -130
rect 2613 -706 2625 -130
rect 2567 -718 2625 -706
rect 2685 -130 2743 -118
rect 2685 -706 2697 -130
rect 2731 -706 2743 -130
rect 2685 -718 2743 -706
rect 2803 -130 2861 -118
rect 2803 -706 2815 -130
rect 2849 -706 2861 -130
rect 2803 -718 2861 -706
rect 2921 -130 2979 -118
rect 2921 -706 2933 -130
rect 2967 -706 2979 -130
rect 2921 -718 2979 -706
rect 3039 -130 3097 -118
rect 3039 -706 3051 -130
rect 3085 -706 3097 -130
rect 3039 -718 3097 -706
rect 3157 -130 3215 -118
rect 3157 -706 3169 -130
rect 3203 -706 3215 -130
rect 3157 -718 3215 -706
rect 3275 -130 3333 -118
rect 3275 -706 3287 -130
rect 3321 -706 3333 -130
rect 3275 -718 3333 -706
rect 3393 -130 3451 -118
rect 3393 -706 3405 -130
rect 3439 -706 3451 -130
rect 3393 -718 3451 -706
rect 3511 -130 3569 -118
rect 3511 -706 3523 -130
rect 3557 -706 3569 -130
rect 3511 -718 3569 -706
<< pdiffc >>
rect -3557 130 -3523 706
rect -3439 130 -3405 706
rect -3321 130 -3287 706
rect -3203 130 -3169 706
rect -3085 130 -3051 706
rect -2967 130 -2933 706
rect -2849 130 -2815 706
rect -2731 130 -2697 706
rect -2613 130 -2579 706
rect -2495 130 -2461 706
rect -2377 130 -2343 706
rect -2259 130 -2225 706
rect -2141 130 -2107 706
rect -2023 130 -1989 706
rect -1905 130 -1871 706
rect -1787 130 -1753 706
rect -1669 130 -1635 706
rect -1551 130 -1517 706
rect -1433 130 -1399 706
rect -1315 130 -1281 706
rect -1197 130 -1163 706
rect -1079 130 -1045 706
rect -961 130 -927 706
rect -843 130 -809 706
rect -725 130 -691 706
rect -607 130 -573 706
rect -489 130 -455 706
rect -371 130 -337 706
rect -253 130 -219 706
rect -135 130 -101 706
rect -17 130 17 706
rect 101 130 135 706
rect 219 130 253 706
rect 337 130 371 706
rect 455 130 489 706
rect 573 130 607 706
rect 691 130 725 706
rect 809 130 843 706
rect 927 130 961 706
rect 1045 130 1079 706
rect 1163 130 1197 706
rect 1281 130 1315 706
rect 1399 130 1433 706
rect 1517 130 1551 706
rect 1635 130 1669 706
rect 1753 130 1787 706
rect 1871 130 1905 706
rect 1989 130 2023 706
rect 2107 130 2141 706
rect 2225 130 2259 706
rect 2343 130 2377 706
rect 2461 130 2495 706
rect 2579 130 2613 706
rect 2697 130 2731 706
rect 2815 130 2849 706
rect 2933 130 2967 706
rect 3051 130 3085 706
rect 3169 130 3203 706
rect 3287 130 3321 706
rect 3405 130 3439 706
rect 3523 130 3557 706
rect -3557 -706 -3523 -130
rect -3439 -706 -3405 -130
rect -3321 -706 -3287 -130
rect -3203 -706 -3169 -130
rect -3085 -706 -3051 -130
rect -2967 -706 -2933 -130
rect -2849 -706 -2815 -130
rect -2731 -706 -2697 -130
rect -2613 -706 -2579 -130
rect -2495 -706 -2461 -130
rect -2377 -706 -2343 -130
rect -2259 -706 -2225 -130
rect -2141 -706 -2107 -130
rect -2023 -706 -1989 -130
rect -1905 -706 -1871 -130
rect -1787 -706 -1753 -130
rect -1669 -706 -1635 -130
rect -1551 -706 -1517 -130
rect -1433 -706 -1399 -130
rect -1315 -706 -1281 -130
rect -1197 -706 -1163 -130
rect -1079 -706 -1045 -130
rect -961 -706 -927 -130
rect -843 -706 -809 -130
rect -725 -706 -691 -130
rect -607 -706 -573 -130
rect -489 -706 -455 -130
rect -371 -706 -337 -130
rect -253 -706 -219 -130
rect -135 -706 -101 -130
rect -17 -706 17 -130
rect 101 -706 135 -130
rect 219 -706 253 -130
rect 337 -706 371 -130
rect 455 -706 489 -130
rect 573 -706 607 -130
rect 691 -706 725 -130
rect 809 -706 843 -130
rect 927 -706 961 -130
rect 1045 -706 1079 -130
rect 1163 -706 1197 -130
rect 1281 -706 1315 -130
rect 1399 -706 1433 -130
rect 1517 -706 1551 -130
rect 1635 -706 1669 -130
rect 1753 -706 1787 -130
rect 1871 -706 1905 -130
rect 1989 -706 2023 -130
rect 2107 -706 2141 -130
rect 2225 -706 2259 -130
rect 2343 -706 2377 -130
rect 2461 -706 2495 -130
rect 2579 -706 2613 -130
rect 2697 -706 2731 -130
rect 2815 -706 2849 -130
rect 2933 -706 2967 -130
rect 3051 -706 3085 -130
rect 3169 -706 3203 -130
rect 3287 -706 3321 -130
rect 3405 -706 3439 -130
rect 3523 -706 3557 -130
<< nsubdiff >>
rect -3671 867 -3575 901
rect 3575 867 3671 901
rect -3671 805 -3637 867
rect 3637 805 3671 867
rect -3671 -867 -3637 -805
rect 3637 -867 3671 -805
rect -3671 -901 -3575 -867
rect 3575 -901 3671 -867
<< nsubdiffcont >>
rect -3575 867 3575 901
rect -3671 -805 -3637 805
rect 3637 -805 3671 805
rect -3575 -901 3575 -867
<< poly >>
rect -3514 799 -3448 815
rect -3514 765 -3498 799
rect -3464 765 -3448 799
rect -3514 749 -3448 765
rect -3396 799 -3330 815
rect -3396 765 -3380 799
rect -3346 765 -3330 799
rect -3396 749 -3330 765
rect -3278 799 -3212 815
rect -3278 765 -3262 799
rect -3228 765 -3212 799
rect -3278 749 -3212 765
rect -3160 799 -3094 815
rect -3160 765 -3144 799
rect -3110 765 -3094 799
rect -3160 749 -3094 765
rect -3042 799 -2976 815
rect -3042 765 -3026 799
rect -2992 765 -2976 799
rect -3042 749 -2976 765
rect -2924 799 -2858 815
rect -2924 765 -2908 799
rect -2874 765 -2858 799
rect -2924 749 -2858 765
rect -2806 799 -2740 815
rect -2806 765 -2790 799
rect -2756 765 -2740 799
rect -2806 749 -2740 765
rect -2688 799 -2622 815
rect -2688 765 -2672 799
rect -2638 765 -2622 799
rect -2688 749 -2622 765
rect -2570 799 -2504 815
rect -2570 765 -2554 799
rect -2520 765 -2504 799
rect -2570 749 -2504 765
rect -2452 799 -2386 815
rect -2452 765 -2436 799
rect -2402 765 -2386 799
rect -2452 749 -2386 765
rect -2334 799 -2268 815
rect -2334 765 -2318 799
rect -2284 765 -2268 799
rect -2334 749 -2268 765
rect -2216 799 -2150 815
rect -2216 765 -2200 799
rect -2166 765 -2150 799
rect -2216 749 -2150 765
rect -2098 799 -2032 815
rect -2098 765 -2082 799
rect -2048 765 -2032 799
rect -2098 749 -2032 765
rect -1980 799 -1914 815
rect -1980 765 -1964 799
rect -1930 765 -1914 799
rect -1980 749 -1914 765
rect -1862 799 -1796 815
rect -1862 765 -1846 799
rect -1812 765 -1796 799
rect -1862 749 -1796 765
rect -1744 799 -1678 815
rect -1744 765 -1728 799
rect -1694 765 -1678 799
rect -1744 749 -1678 765
rect -1626 799 -1560 815
rect -1626 765 -1610 799
rect -1576 765 -1560 799
rect -1626 749 -1560 765
rect -1508 799 -1442 815
rect -1508 765 -1492 799
rect -1458 765 -1442 799
rect -1508 749 -1442 765
rect -1390 799 -1324 815
rect -1390 765 -1374 799
rect -1340 765 -1324 799
rect -1390 749 -1324 765
rect -1272 799 -1206 815
rect -1272 765 -1256 799
rect -1222 765 -1206 799
rect -1272 749 -1206 765
rect -1154 799 -1088 815
rect -1154 765 -1138 799
rect -1104 765 -1088 799
rect -1154 749 -1088 765
rect -1036 799 -970 815
rect -1036 765 -1020 799
rect -986 765 -970 799
rect -1036 749 -970 765
rect -918 799 -852 815
rect -918 765 -902 799
rect -868 765 -852 799
rect -918 749 -852 765
rect -800 799 -734 815
rect -800 765 -784 799
rect -750 765 -734 799
rect -800 749 -734 765
rect -682 799 -616 815
rect -682 765 -666 799
rect -632 765 -616 799
rect -682 749 -616 765
rect -564 799 -498 815
rect -564 765 -548 799
rect -514 765 -498 799
rect -564 749 -498 765
rect -446 799 -380 815
rect -446 765 -430 799
rect -396 765 -380 799
rect -446 749 -380 765
rect -328 799 -262 815
rect -328 765 -312 799
rect -278 765 -262 799
rect -328 749 -262 765
rect -210 799 -144 815
rect -210 765 -194 799
rect -160 765 -144 799
rect -210 749 -144 765
rect -92 799 -26 815
rect -92 765 -76 799
rect -42 765 -26 799
rect -92 749 -26 765
rect 26 799 92 815
rect 26 765 42 799
rect 76 765 92 799
rect 26 749 92 765
rect 144 799 210 815
rect 144 765 160 799
rect 194 765 210 799
rect 144 749 210 765
rect 262 799 328 815
rect 262 765 278 799
rect 312 765 328 799
rect 262 749 328 765
rect 380 799 446 815
rect 380 765 396 799
rect 430 765 446 799
rect 380 749 446 765
rect 498 799 564 815
rect 498 765 514 799
rect 548 765 564 799
rect 498 749 564 765
rect 616 799 682 815
rect 616 765 632 799
rect 666 765 682 799
rect 616 749 682 765
rect 734 799 800 815
rect 734 765 750 799
rect 784 765 800 799
rect 734 749 800 765
rect 852 799 918 815
rect 852 765 868 799
rect 902 765 918 799
rect 852 749 918 765
rect 970 799 1036 815
rect 970 765 986 799
rect 1020 765 1036 799
rect 970 749 1036 765
rect 1088 799 1154 815
rect 1088 765 1104 799
rect 1138 765 1154 799
rect 1088 749 1154 765
rect 1206 799 1272 815
rect 1206 765 1222 799
rect 1256 765 1272 799
rect 1206 749 1272 765
rect 1324 799 1390 815
rect 1324 765 1340 799
rect 1374 765 1390 799
rect 1324 749 1390 765
rect 1442 799 1508 815
rect 1442 765 1458 799
rect 1492 765 1508 799
rect 1442 749 1508 765
rect 1560 799 1626 815
rect 1560 765 1576 799
rect 1610 765 1626 799
rect 1560 749 1626 765
rect 1678 799 1744 815
rect 1678 765 1694 799
rect 1728 765 1744 799
rect 1678 749 1744 765
rect 1796 799 1862 815
rect 1796 765 1812 799
rect 1846 765 1862 799
rect 1796 749 1862 765
rect 1914 799 1980 815
rect 1914 765 1930 799
rect 1964 765 1980 799
rect 1914 749 1980 765
rect 2032 799 2098 815
rect 2032 765 2048 799
rect 2082 765 2098 799
rect 2032 749 2098 765
rect 2150 799 2216 815
rect 2150 765 2166 799
rect 2200 765 2216 799
rect 2150 749 2216 765
rect 2268 799 2334 815
rect 2268 765 2284 799
rect 2318 765 2334 799
rect 2268 749 2334 765
rect 2386 799 2452 815
rect 2386 765 2402 799
rect 2436 765 2452 799
rect 2386 749 2452 765
rect 2504 799 2570 815
rect 2504 765 2520 799
rect 2554 765 2570 799
rect 2504 749 2570 765
rect 2622 799 2688 815
rect 2622 765 2638 799
rect 2672 765 2688 799
rect 2622 749 2688 765
rect 2740 799 2806 815
rect 2740 765 2756 799
rect 2790 765 2806 799
rect 2740 749 2806 765
rect 2858 799 2924 815
rect 2858 765 2874 799
rect 2908 765 2924 799
rect 2858 749 2924 765
rect 2976 799 3042 815
rect 2976 765 2992 799
rect 3026 765 3042 799
rect 2976 749 3042 765
rect 3094 799 3160 815
rect 3094 765 3110 799
rect 3144 765 3160 799
rect 3094 749 3160 765
rect 3212 799 3278 815
rect 3212 765 3228 799
rect 3262 765 3278 799
rect 3212 749 3278 765
rect 3330 799 3396 815
rect 3330 765 3346 799
rect 3380 765 3396 799
rect 3330 749 3396 765
rect 3448 799 3514 815
rect 3448 765 3464 799
rect 3498 765 3514 799
rect 3448 749 3514 765
rect -3511 718 -3451 749
rect -3393 718 -3333 749
rect -3275 718 -3215 749
rect -3157 718 -3097 749
rect -3039 718 -2979 749
rect -2921 718 -2861 749
rect -2803 718 -2743 749
rect -2685 718 -2625 749
rect -2567 718 -2507 749
rect -2449 718 -2389 749
rect -2331 718 -2271 749
rect -2213 718 -2153 749
rect -2095 718 -2035 749
rect -1977 718 -1917 749
rect -1859 718 -1799 749
rect -1741 718 -1681 749
rect -1623 718 -1563 749
rect -1505 718 -1445 749
rect -1387 718 -1327 749
rect -1269 718 -1209 749
rect -1151 718 -1091 749
rect -1033 718 -973 749
rect -915 718 -855 749
rect -797 718 -737 749
rect -679 718 -619 749
rect -561 718 -501 749
rect -443 718 -383 749
rect -325 718 -265 749
rect -207 718 -147 749
rect -89 718 -29 749
rect 29 718 89 749
rect 147 718 207 749
rect 265 718 325 749
rect 383 718 443 749
rect 501 718 561 749
rect 619 718 679 749
rect 737 718 797 749
rect 855 718 915 749
rect 973 718 1033 749
rect 1091 718 1151 749
rect 1209 718 1269 749
rect 1327 718 1387 749
rect 1445 718 1505 749
rect 1563 718 1623 749
rect 1681 718 1741 749
rect 1799 718 1859 749
rect 1917 718 1977 749
rect 2035 718 2095 749
rect 2153 718 2213 749
rect 2271 718 2331 749
rect 2389 718 2449 749
rect 2507 718 2567 749
rect 2625 718 2685 749
rect 2743 718 2803 749
rect 2861 718 2921 749
rect 2979 718 3039 749
rect 3097 718 3157 749
rect 3215 718 3275 749
rect 3333 718 3393 749
rect 3451 718 3511 749
rect -3511 87 -3451 118
rect -3393 87 -3333 118
rect -3275 87 -3215 118
rect -3157 87 -3097 118
rect -3039 87 -2979 118
rect -2921 87 -2861 118
rect -2803 87 -2743 118
rect -2685 87 -2625 118
rect -2567 87 -2507 118
rect -2449 87 -2389 118
rect -2331 87 -2271 118
rect -2213 87 -2153 118
rect -2095 87 -2035 118
rect -1977 87 -1917 118
rect -1859 87 -1799 118
rect -1741 87 -1681 118
rect -1623 87 -1563 118
rect -1505 87 -1445 118
rect -1387 87 -1327 118
rect -1269 87 -1209 118
rect -1151 87 -1091 118
rect -1033 87 -973 118
rect -915 87 -855 118
rect -797 87 -737 118
rect -679 87 -619 118
rect -561 87 -501 118
rect -443 87 -383 118
rect -325 87 -265 118
rect -207 87 -147 118
rect -89 87 -29 118
rect 29 87 89 118
rect 147 87 207 118
rect 265 87 325 118
rect 383 87 443 118
rect 501 87 561 118
rect 619 87 679 118
rect 737 87 797 118
rect 855 87 915 118
rect 973 87 1033 118
rect 1091 87 1151 118
rect 1209 87 1269 118
rect 1327 87 1387 118
rect 1445 87 1505 118
rect 1563 87 1623 118
rect 1681 87 1741 118
rect 1799 87 1859 118
rect 1917 87 1977 118
rect 2035 87 2095 118
rect 2153 87 2213 118
rect 2271 87 2331 118
rect 2389 87 2449 118
rect 2507 87 2567 118
rect 2625 87 2685 118
rect 2743 87 2803 118
rect 2861 87 2921 118
rect 2979 87 3039 118
rect 3097 87 3157 118
rect 3215 87 3275 118
rect 3333 87 3393 118
rect 3451 87 3511 118
rect -3514 71 -3448 87
rect -3514 37 -3498 71
rect -3464 37 -3448 71
rect -3514 21 -3448 37
rect -3396 71 -3330 87
rect -3396 37 -3380 71
rect -3346 37 -3330 71
rect -3396 21 -3330 37
rect -3278 71 -3212 87
rect -3278 37 -3262 71
rect -3228 37 -3212 71
rect -3278 21 -3212 37
rect -3160 71 -3094 87
rect -3160 37 -3144 71
rect -3110 37 -3094 71
rect -3160 21 -3094 37
rect -3042 71 -2976 87
rect -3042 37 -3026 71
rect -2992 37 -2976 71
rect -3042 21 -2976 37
rect -2924 71 -2858 87
rect -2924 37 -2908 71
rect -2874 37 -2858 71
rect -2924 21 -2858 37
rect -2806 71 -2740 87
rect -2806 37 -2790 71
rect -2756 37 -2740 71
rect -2806 21 -2740 37
rect -2688 71 -2622 87
rect -2688 37 -2672 71
rect -2638 37 -2622 71
rect -2688 21 -2622 37
rect -2570 71 -2504 87
rect -2570 37 -2554 71
rect -2520 37 -2504 71
rect -2570 21 -2504 37
rect -2452 71 -2386 87
rect -2452 37 -2436 71
rect -2402 37 -2386 71
rect -2452 21 -2386 37
rect -2334 71 -2268 87
rect -2334 37 -2318 71
rect -2284 37 -2268 71
rect -2334 21 -2268 37
rect -2216 71 -2150 87
rect -2216 37 -2200 71
rect -2166 37 -2150 71
rect -2216 21 -2150 37
rect -2098 71 -2032 87
rect -2098 37 -2082 71
rect -2048 37 -2032 71
rect -2098 21 -2032 37
rect -1980 71 -1914 87
rect -1980 37 -1964 71
rect -1930 37 -1914 71
rect -1980 21 -1914 37
rect -1862 71 -1796 87
rect -1862 37 -1846 71
rect -1812 37 -1796 71
rect -1862 21 -1796 37
rect -1744 71 -1678 87
rect -1744 37 -1728 71
rect -1694 37 -1678 71
rect -1744 21 -1678 37
rect -1626 71 -1560 87
rect -1626 37 -1610 71
rect -1576 37 -1560 71
rect -1626 21 -1560 37
rect -1508 71 -1442 87
rect -1508 37 -1492 71
rect -1458 37 -1442 71
rect -1508 21 -1442 37
rect -1390 71 -1324 87
rect -1390 37 -1374 71
rect -1340 37 -1324 71
rect -1390 21 -1324 37
rect -1272 71 -1206 87
rect -1272 37 -1256 71
rect -1222 37 -1206 71
rect -1272 21 -1206 37
rect -1154 71 -1088 87
rect -1154 37 -1138 71
rect -1104 37 -1088 71
rect -1154 21 -1088 37
rect -1036 71 -970 87
rect -1036 37 -1020 71
rect -986 37 -970 71
rect -1036 21 -970 37
rect -918 71 -852 87
rect -918 37 -902 71
rect -868 37 -852 71
rect -918 21 -852 37
rect -800 71 -734 87
rect -800 37 -784 71
rect -750 37 -734 71
rect -800 21 -734 37
rect -682 71 -616 87
rect -682 37 -666 71
rect -632 37 -616 71
rect -682 21 -616 37
rect -564 71 -498 87
rect -564 37 -548 71
rect -514 37 -498 71
rect -564 21 -498 37
rect -446 71 -380 87
rect -446 37 -430 71
rect -396 37 -380 71
rect -446 21 -380 37
rect -328 71 -262 87
rect -328 37 -312 71
rect -278 37 -262 71
rect -328 21 -262 37
rect -210 71 -144 87
rect -210 37 -194 71
rect -160 37 -144 71
rect -210 21 -144 37
rect -92 71 -26 87
rect -92 37 -76 71
rect -42 37 -26 71
rect -92 21 -26 37
rect 26 71 92 87
rect 26 37 42 71
rect 76 37 92 71
rect 26 21 92 37
rect 144 71 210 87
rect 144 37 160 71
rect 194 37 210 71
rect 144 21 210 37
rect 262 71 328 87
rect 262 37 278 71
rect 312 37 328 71
rect 262 21 328 37
rect 380 71 446 87
rect 380 37 396 71
rect 430 37 446 71
rect 380 21 446 37
rect 498 71 564 87
rect 498 37 514 71
rect 548 37 564 71
rect 498 21 564 37
rect 616 71 682 87
rect 616 37 632 71
rect 666 37 682 71
rect 616 21 682 37
rect 734 71 800 87
rect 734 37 750 71
rect 784 37 800 71
rect 734 21 800 37
rect 852 71 918 87
rect 852 37 868 71
rect 902 37 918 71
rect 852 21 918 37
rect 970 71 1036 87
rect 970 37 986 71
rect 1020 37 1036 71
rect 970 21 1036 37
rect 1088 71 1154 87
rect 1088 37 1104 71
rect 1138 37 1154 71
rect 1088 21 1154 37
rect 1206 71 1272 87
rect 1206 37 1222 71
rect 1256 37 1272 71
rect 1206 21 1272 37
rect 1324 71 1390 87
rect 1324 37 1340 71
rect 1374 37 1390 71
rect 1324 21 1390 37
rect 1442 71 1508 87
rect 1442 37 1458 71
rect 1492 37 1508 71
rect 1442 21 1508 37
rect 1560 71 1626 87
rect 1560 37 1576 71
rect 1610 37 1626 71
rect 1560 21 1626 37
rect 1678 71 1744 87
rect 1678 37 1694 71
rect 1728 37 1744 71
rect 1678 21 1744 37
rect 1796 71 1862 87
rect 1796 37 1812 71
rect 1846 37 1862 71
rect 1796 21 1862 37
rect 1914 71 1980 87
rect 1914 37 1930 71
rect 1964 37 1980 71
rect 1914 21 1980 37
rect 2032 71 2098 87
rect 2032 37 2048 71
rect 2082 37 2098 71
rect 2032 21 2098 37
rect 2150 71 2216 87
rect 2150 37 2166 71
rect 2200 37 2216 71
rect 2150 21 2216 37
rect 2268 71 2334 87
rect 2268 37 2284 71
rect 2318 37 2334 71
rect 2268 21 2334 37
rect 2386 71 2452 87
rect 2386 37 2402 71
rect 2436 37 2452 71
rect 2386 21 2452 37
rect 2504 71 2570 87
rect 2504 37 2520 71
rect 2554 37 2570 71
rect 2504 21 2570 37
rect 2622 71 2688 87
rect 2622 37 2638 71
rect 2672 37 2688 71
rect 2622 21 2688 37
rect 2740 71 2806 87
rect 2740 37 2756 71
rect 2790 37 2806 71
rect 2740 21 2806 37
rect 2858 71 2924 87
rect 2858 37 2874 71
rect 2908 37 2924 71
rect 2858 21 2924 37
rect 2976 71 3042 87
rect 2976 37 2992 71
rect 3026 37 3042 71
rect 2976 21 3042 37
rect 3094 71 3160 87
rect 3094 37 3110 71
rect 3144 37 3160 71
rect 3094 21 3160 37
rect 3212 71 3278 87
rect 3212 37 3228 71
rect 3262 37 3278 71
rect 3212 21 3278 37
rect 3330 71 3396 87
rect 3330 37 3346 71
rect 3380 37 3396 71
rect 3330 21 3396 37
rect 3448 71 3514 87
rect 3448 37 3464 71
rect 3498 37 3514 71
rect 3448 21 3514 37
rect -3514 -37 -3448 -21
rect -3514 -71 -3498 -37
rect -3464 -71 -3448 -37
rect -3514 -87 -3448 -71
rect -3396 -37 -3330 -21
rect -3396 -71 -3380 -37
rect -3346 -71 -3330 -37
rect -3396 -87 -3330 -71
rect -3278 -37 -3212 -21
rect -3278 -71 -3262 -37
rect -3228 -71 -3212 -37
rect -3278 -87 -3212 -71
rect -3160 -37 -3094 -21
rect -3160 -71 -3144 -37
rect -3110 -71 -3094 -37
rect -3160 -87 -3094 -71
rect -3042 -37 -2976 -21
rect -3042 -71 -3026 -37
rect -2992 -71 -2976 -37
rect -3042 -87 -2976 -71
rect -2924 -37 -2858 -21
rect -2924 -71 -2908 -37
rect -2874 -71 -2858 -37
rect -2924 -87 -2858 -71
rect -2806 -37 -2740 -21
rect -2806 -71 -2790 -37
rect -2756 -71 -2740 -37
rect -2806 -87 -2740 -71
rect -2688 -37 -2622 -21
rect -2688 -71 -2672 -37
rect -2638 -71 -2622 -37
rect -2688 -87 -2622 -71
rect -2570 -37 -2504 -21
rect -2570 -71 -2554 -37
rect -2520 -71 -2504 -37
rect -2570 -87 -2504 -71
rect -2452 -37 -2386 -21
rect -2452 -71 -2436 -37
rect -2402 -71 -2386 -37
rect -2452 -87 -2386 -71
rect -2334 -37 -2268 -21
rect -2334 -71 -2318 -37
rect -2284 -71 -2268 -37
rect -2334 -87 -2268 -71
rect -2216 -37 -2150 -21
rect -2216 -71 -2200 -37
rect -2166 -71 -2150 -37
rect -2216 -87 -2150 -71
rect -2098 -37 -2032 -21
rect -2098 -71 -2082 -37
rect -2048 -71 -2032 -37
rect -2098 -87 -2032 -71
rect -1980 -37 -1914 -21
rect -1980 -71 -1964 -37
rect -1930 -71 -1914 -37
rect -1980 -87 -1914 -71
rect -1862 -37 -1796 -21
rect -1862 -71 -1846 -37
rect -1812 -71 -1796 -37
rect -1862 -87 -1796 -71
rect -1744 -37 -1678 -21
rect -1744 -71 -1728 -37
rect -1694 -71 -1678 -37
rect -1744 -87 -1678 -71
rect -1626 -37 -1560 -21
rect -1626 -71 -1610 -37
rect -1576 -71 -1560 -37
rect -1626 -87 -1560 -71
rect -1508 -37 -1442 -21
rect -1508 -71 -1492 -37
rect -1458 -71 -1442 -37
rect -1508 -87 -1442 -71
rect -1390 -37 -1324 -21
rect -1390 -71 -1374 -37
rect -1340 -71 -1324 -37
rect -1390 -87 -1324 -71
rect -1272 -37 -1206 -21
rect -1272 -71 -1256 -37
rect -1222 -71 -1206 -37
rect -1272 -87 -1206 -71
rect -1154 -37 -1088 -21
rect -1154 -71 -1138 -37
rect -1104 -71 -1088 -37
rect -1154 -87 -1088 -71
rect -1036 -37 -970 -21
rect -1036 -71 -1020 -37
rect -986 -71 -970 -37
rect -1036 -87 -970 -71
rect -918 -37 -852 -21
rect -918 -71 -902 -37
rect -868 -71 -852 -37
rect -918 -87 -852 -71
rect -800 -37 -734 -21
rect -800 -71 -784 -37
rect -750 -71 -734 -37
rect -800 -87 -734 -71
rect -682 -37 -616 -21
rect -682 -71 -666 -37
rect -632 -71 -616 -37
rect -682 -87 -616 -71
rect -564 -37 -498 -21
rect -564 -71 -548 -37
rect -514 -71 -498 -37
rect -564 -87 -498 -71
rect -446 -37 -380 -21
rect -446 -71 -430 -37
rect -396 -71 -380 -37
rect -446 -87 -380 -71
rect -328 -37 -262 -21
rect -328 -71 -312 -37
rect -278 -71 -262 -37
rect -328 -87 -262 -71
rect -210 -37 -144 -21
rect -210 -71 -194 -37
rect -160 -71 -144 -37
rect -210 -87 -144 -71
rect -92 -37 -26 -21
rect -92 -71 -76 -37
rect -42 -71 -26 -37
rect -92 -87 -26 -71
rect 26 -37 92 -21
rect 26 -71 42 -37
rect 76 -71 92 -37
rect 26 -87 92 -71
rect 144 -37 210 -21
rect 144 -71 160 -37
rect 194 -71 210 -37
rect 144 -87 210 -71
rect 262 -37 328 -21
rect 262 -71 278 -37
rect 312 -71 328 -37
rect 262 -87 328 -71
rect 380 -37 446 -21
rect 380 -71 396 -37
rect 430 -71 446 -37
rect 380 -87 446 -71
rect 498 -37 564 -21
rect 498 -71 514 -37
rect 548 -71 564 -37
rect 498 -87 564 -71
rect 616 -37 682 -21
rect 616 -71 632 -37
rect 666 -71 682 -37
rect 616 -87 682 -71
rect 734 -37 800 -21
rect 734 -71 750 -37
rect 784 -71 800 -37
rect 734 -87 800 -71
rect 852 -37 918 -21
rect 852 -71 868 -37
rect 902 -71 918 -37
rect 852 -87 918 -71
rect 970 -37 1036 -21
rect 970 -71 986 -37
rect 1020 -71 1036 -37
rect 970 -87 1036 -71
rect 1088 -37 1154 -21
rect 1088 -71 1104 -37
rect 1138 -71 1154 -37
rect 1088 -87 1154 -71
rect 1206 -37 1272 -21
rect 1206 -71 1222 -37
rect 1256 -71 1272 -37
rect 1206 -87 1272 -71
rect 1324 -37 1390 -21
rect 1324 -71 1340 -37
rect 1374 -71 1390 -37
rect 1324 -87 1390 -71
rect 1442 -37 1508 -21
rect 1442 -71 1458 -37
rect 1492 -71 1508 -37
rect 1442 -87 1508 -71
rect 1560 -37 1626 -21
rect 1560 -71 1576 -37
rect 1610 -71 1626 -37
rect 1560 -87 1626 -71
rect 1678 -37 1744 -21
rect 1678 -71 1694 -37
rect 1728 -71 1744 -37
rect 1678 -87 1744 -71
rect 1796 -37 1862 -21
rect 1796 -71 1812 -37
rect 1846 -71 1862 -37
rect 1796 -87 1862 -71
rect 1914 -37 1980 -21
rect 1914 -71 1930 -37
rect 1964 -71 1980 -37
rect 1914 -87 1980 -71
rect 2032 -37 2098 -21
rect 2032 -71 2048 -37
rect 2082 -71 2098 -37
rect 2032 -87 2098 -71
rect 2150 -37 2216 -21
rect 2150 -71 2166 -37
rect 2200 -71 2216 -37
rect 2150 -87 2216 -71
rect 2268 -37 2334 -21
rect 2268 -71 2284 -37
rect 2318 -71 2334 -37
rect 2268 -87 2334 -71
rect 2386 -37 2452 -21
rect 2386 -71 2402 -37
rect 2436 -71 2452 -37
rect 2386 -87 2452 -71
rect 2504 -37 2570 -21
rect 2504 -71 2520 -37
rect 2554 -71 2570 -37
rect 2504 -87 2570 -71
rect 2622 -37 2688 -21
rect 2622 -71 2638 -37
rect 2672 -71 2688 -37
rect 2622 -87 2688 -71
rect 2740 -37 2806 -21
rect 2740 -71 2756 -37
rect 2790 -71 2806 -37
rect 2740 -87 2806 -71
rect 2858 -37 2924 -21
rect 2858 -71 2874 -37
rect 2908 -71 2924 -37
rect 2858 -87 2924 -71
rect 2976 -37 3042 -21
rect 2976 -71 2992 -37
rect 3026 -71 3042 -37
rect 2976 -87 3042 -71
rect 3094 -37 3160 -21
rect 3094 -71 3110 -37
rect 3144 -71 3160 -37
rect 3094 -87 3160 -71
rect 3212 -37 3278 -21
rect 3212 -71 3228 -37
rect 3262 -71 3278 -37
rect 3212 -87 3278 -71
rect 3330 -37 3396 -21
rect 3330 -71 3346 -37
rect 3380 -71 3396 -37
rect 3330 -87 3396 -71
rect 3448 -37 3514 -21
rect 3448 -71 3464 -37
rect 3498 -71 3514 -37
rect 3448 -87 3514 -71
rect -3511 -118 -3451 -87
rect -3393 -118 -3333 -87
rect -3275 -118 -3215 -87
rect -3157 -118 -3097 -87
rect -3039 -118 -2979 -87
rect -2921 -118 -2861 -87
rect -2803 -118 -2743 -87
rect -2685 -118 -2625 -87
rect -2567 -118 -2507 -87
rect -2449 -118 -2389 -87
rect -2331 -118 -2271 -87
rect -2213 -118 -2153 -87
rect -2095 -118 -2035 -87
rect -1977 -118 -1917 -87
rect -1859 -118 -1799 -87
rect -1741 -118 -1681 -87
rect -1623 -118 -1563 -87
rect -1505 -118 -1445 -87
rect -1387 -118 -1327 -87
rect -1269 -118 -1209 -87
rect -1151 -118 -1091 -87
rect -1033 -118 -973 -87
rect -915 -118 -855 -87
rect -797 -118 -737 -87
rect -679 -118 -619 -87
rect -561 -118 -501 -87
rect -443 -118 -383 -87
rect -325 -118 -265 -87
rect -207 -118 -147 -87
rect -89 -118 -29 -87
rect 29 -118 89 -87
rect 147 -118 207 -87
rect 265 -118 325 -87
rect 383 -118 443 -87
rect 501 -118 561 -87
rect 619 -118 679 -87
rect 737 -118 797 -87
rect 855 -118 915 -87
rect 973 -118 1033 -87
rect 1091 -118 1151 -87
rect 1209 -118 1269 -87
rect 1327 -118 1387 -87
rect 1445 -118 1505 -87
rect 1563 -118 1623 -87
rect 1681 -118 1741 -87
rect 1799 -118 1859 -87
rect 1917 -118 1977 -87
rect 2035 -118 2095 -87
rect 2153 -118 2213 -87
rect 2271 -118 2331 -87
rect 2389 -118 2449 -87
rect 2507 -118 2567 -87
rect 2625 -118 2685 -87
rect 2743 -118 2803 -87
rect 2861 -118 2921 -87
rect 2979 -118 3039 -87
rect 3097 -118 3157 -87
rect 3215 -118 3275 -87
rect 3333 -118 3393 -87
rect 3451 -118 3511 -87
rect -3511 -749 -3451 -718
rect -3393 -749 -3333 -718
rect -3275 -749 -3215 -718
rect -3157 -749 -3097 -718
rect -3039 -749 -2979 -718
rect -2921 -749 -2861 -718
rect -2803 -749 -2743 -718
rect -2685 -749 -2625 -718
rect -2567 -749 -2507 -718
rect -2449 -749 -2389 -718
rect -2331 -749 -2271 -718
rect -2213 -749 -2153 -718
rect -2095 -749 -2035 -718
rect -1977 -749 -1917 -718
rect -1859 -749 -1799 -718
rect -1741 -749 -1681 -718
rect -1623 -749 -1563 -718
rect -1505 -749 -1445 -718
rect -1387 -749 -1327 -718
rect -1269 -749 -1209 -718
rect -1151 -749 -1091 -718
rect -1033 -749 -973 -718
rect -915 -749 -855 -718
rect -797 -749 -737 -718
rect -679 -749 -619 -718
rect -561 -749 -501 -718
rect -443 -749 -383 -718
rect -325 -749 -265 -718
rect -207 -749 -147 -718
rect -89 -749 -29 -718
rect 29 -749 89 -718
rect 147 -749 207 -718
rect 265 -749 325 -718
rect 383 -749 443 -718
rect 501 -749 561 -718
rect 619 -749 679 -718
rect 737 -749 797 -718
rect 855 -749 915 -718
rect 973 -749 1033 -718
rect 1091 -749 1151 -718
rect 1209 -749 1269 -718
rect 1327 -749 1387 -718
rect 1445 -749 1505 -718
rect 1563 -749 1623 -718
rect 1681 -749 1741 -718
rect 1799 -749 1859 -718
rect 1917 -749 1977 -718
rect 2035 -749 2095 -718
rect 2153 -749 2213 -718
rect 2271 -749 2331 -718
rect 2389 -749 2449 -718
rect 2507 -749 2567 -718
rect 2625 -749 2685 -718
rect 2743 -749 2803 -718
rect 2861 -749 2921 -718
rect 2979 -749 3039 -718
rect 3097 -749 3157 -718
rect 3215 -749 3275 -718
rect 3333 -749 3393 -718
rect 3451 -749 3511 -718
rect -3514 -765 -3448 -749
rect -3514 -799 -3498 -765
rect -3464 -799 -3448 -765
rect -3514 -815 -3448 -799
rect -3396 -765 -3330 -749
rect -3396 -799 -3380 -765
rect -3346 -799 -3330 -765
rect -3396 -815 -3330 -799
rect -3278 -765 -3212 -749
rect -3278 -799 -3262 -765
rect -3228 -799 -3212 -765
rect -3278 -815 -3212 -799
rect -3160 -765 -3094 -749
rect -3160 -799 -3144 -765
rect -3110 -799 -3094 -765
rect -3160 -815 -3094 -799
rect -3042 -765 -2976 -749
rect -3042 -799 -3026 -765
rect -2992 -799 -2976 -765
rect -3042 -815 -2976 -799
rect -2924 -765 -2858 -749
rect -2924 -799 -2908 -765
rect -2874 -799 -2858 -765
rect -2924 -815 -2858 -799
rect -2806 -765 -2740 -749
rect -2806 -799 -2790 -765
rect -2756 -799 -2740 -765
rect -2806 -815 -2740 -799
rect -2688 -765 -2622 -749
rect -2688 -799 -2672 -765
rect -2638 -799 -2622 -765
rect -2688 -815 -2622 -799
rect -2570 -765 -2504 -749
rect -2570 -799 -2554 -765
rect -2520 -799 -2504 -765
rect -2570 -815 -2504 -799
rect -2452 -765 -2386 -749
rect -2452 -799 -2436 -765
rect -2402 -799 -2386 -765
rect -2452 -815 -2386 -799
rect -2334 -765 -2268 -749
rect -2334 -799 -2318 -765
rect -2284 -799 -2268 -765
rect -2334 -815 -2268 -799
rect -2216 -765 -2150 -749
rect -2216 -799 -2200 -765
rect -2166 -799 -2150 -765
rect -2216 -815 -2150 -799
rect -2098 -765 -2032 -749
rect -2098 -799 -2082 -765
rect -2048 -799 -2032 -765
rect -2098 -815 -2032 -799
rect -1980 -765 -1914 -749
rect -1980 -799 -1964 -765
rect -1930 -799 -1914 -765
rect -1980 -815 -1914 -799
rect -1862 -765 -1796 -749
rect -1862 -799 -1846 -765
rect -1812 -799 -1796 -765
rect -1862 -815 -1796 -799
rect -1744 -765 -1678 -749
rect -1744 -799 -1728 -765
rect -1694 -799 -1678 -765
rect -1744 -815 -1678 -799
rect -1626 -765 -1560 -749
rect -1626 -799 -1610 -765
rect -1576 -799 -1560 -765
rect -1626 -815 -1560 -799
rect -1508 -765 -1442 -749
rect -1508 -799 -1492 -765
rect -1458 -799 -1442 -765
rect -1508 -815 -1442 -799
rect -1390 -765 -1324 -749
rect -1390 -799 -1374 -765
rect -1340 -799 -1324 -765
rect -1390 -815 -1324 -799
rect -1272 -765 -1206 -749
rect -1272 -799 -1256 -765
rect -1222 -799 -1206 -765
rect -1272 -815 -1206 -799
rect -1154 -765 -1088 -749
rect -1154 -799 -1138 -765
rect -1104 -799 -1088 -765
rect -1154 -815 -1088 -799
rect -1036 -765 -970 -749
rect -1036 -799 -1020 -765
rect -986 -799 -970 -765
rect -1036 -815 -970 -799
rect -918 -765 -852 -749
rect -918 -799 -902 -765
rect -868 -799 -852 -765
rect -918 -815 -852 -799
rect -800 -765 -734 -749
rect -800 -799 -784 -765
rect -750 -799 -734 -765
rect -800 -815 -734 -799
rect -682 -765 -616 -749
rect -682 -799 -666 -765
rect -632 -799 -616 -765
rect -682 -815 -616 -799
rect -564 -765 -498 -749
rect -564 -799 -548 -765
rect -514 -799 -498 -765
rect -564 -815 -498 -799
rect -446 -765 -380 -749
rect -446 -799 -430 -765
rect -396 -799 -380 -765
rect -446 -815 -380 -799
rect -328 -765 -262 -749
rect -328 -799 -312 -765
rect -278 -799 -262 -765
rect -328 -815 -262 -799
rect -210 -765 -144 -749
rect -210 -799 -194 -765
rect -160 -799 -144 -765
rect -210 -815 -144 -799
rect -92 -765 -26 -749
rect -92 -799 -76 -765
rect -42 -799 -26 -765
rect -92 -815 -26 -799
rect 26 -765 92 -749
rect 26 -799 42 -765
rect 76 -799 92 -765
rect 26 -815 92 -799
rect 144 -765 210 -749
rect 144 -799 160 -765
rect 194 -799 210 -765
rect 144 -815 210 -799
rect 262 -765 328 -749
rect 262 -799 278 -765
rect 312 -799 328 -765
rect 262 -815 328 -799
rect 380 -765 446 -749
rect 380 -799 396 -765
rect 430 -799 446 -765
rect 380 -815 446 -799
rect 498 -765 564 -749
rect 498 -799 514 -765
rect 548 -799 564 -765
rect 498 -815 564 -799
rect 616 -765 682 -749
rect 616 -799 632 -765
rect 666 -799 682 -765
rect 616 -815 682 -799
rect 734 -765 800 -749
rect 734 -799 750 -765
rect 784 -799 800 -765
rect 734 -815 800 -799
rect 852 -765 918 -749
rect 852 -799 868 -765
rect 902 -799 918 -765
rect 852 -815 918 -799
rect 970 -765 1036 -749
rect 970 -799 986 -765
rect 1020 -799 1036 -765
rect 970 -815 1036 -799
rect 1088 -765 1154 -749
rect 1088 -799 1104 -765
rect 1138 -799 1154 -765
rect 1088 -815 1154 -799
rect 1206 -765 1272 -749
rect 1206 -799 1222 -765
rect 1256 -799 1272 -765
rect 1206 -815 1272 -799
rect 1324 -765 1390 -749
rect 1324 -799 1340 -765
rect 1374 -799 1390 -765
rect 1324 -815 1390 -799
rect 1442 -765 1508 -749
rect 1442 -799 1458 -765
rect 1492 -799 1508 -765
rect 1442 -815 1508 -799
rect 1560 -765 1626 -749
rect 1560 -799 1576 -765
rect 1610 -799 1626 -765
rect 1560 -815 1626 -799
rect 1678 -765 1744 -749
rect 1678 -799 1694 -765
rect 1728 -799 1744 -765
rect 1678 -815 1744 -799
rect 1796 -765 1862 -749
rect 1796 -799 1812 -765
rect 1846 -799 1862 -765
rect 1796 -815 1862 -799
rect 1914 -765 1980 -749
rect 1914 -799 1930 -765
rect 1964 -799 1980 -765
rect 1914 -815 1980 -799
rect 2032 -765 2098 -749
rect 2032 -799 2048 -765
rect 2082 -799 2098 -765
rect 2032 -815 2098 -799
rect 2150 -765 2216 -749
rect 2150 -799 2166 -765
rect 2200 -799 2216 -765
rect 2150 -815 2216 -799
rect 2268 -765 2334 -749
rect 2268 -799 2284 -765
rect 2318 -799 2334 -765
rect 2268 -815 2334 -799
rect 2386 -765 2452 -749
rect 2386 -799 2402 -765
rect 2436 -799 2452 -765
rect 2386 -815 2452 -799
rect 2504 -765 2570 -749
rect 2504 -799 2520 -765
rect 2554 -799 2570 -765
rect 2504 -815 2570 -799
rect 2622 -765 2688 -749
rect 2622 -799 2638 -765
rect 2672 -799 2688 -765
rect 2622 -815 2688 -799
rect 2740 -765 2806 -749
rect 2740 -799 2756 -765
rect 2790 -799 2806 -765
rect 2740 -815 2806 -799
rect 2858 -765 2924 -749
rect 2858 -799 2874 -765
rect 2908 -799 2924 -765
rect 2858 -815 2924 -799
rect 2976 -765 3042 -749
rect 2976 -799 2992 -765
rect 3026 -799 3042 -765
rect 2976 -815 3042 -799
rect 3094 -765 3160 -749
rect 3094 -799 3110 -765
rect 3144 -799 3160 -765
rect 3094 -815 3160 -799
rect 3212 -765 3278 -749
rect 3212 -799 3228 -765
rect 3262 -799 3278 -765
rect 3212 -815 3278 -799
rect 3330 -765 3396 -749
rect 3330 -799 3346 -765
rect 3380 -799 3396 -765
rect 3330 -815 3396 -799
rect 3448 -765 3514 -749
rect 3448 -799 3464 -765
rect 3498 -799 3514 -765
rect 3448 -815 3514 -799
<< polycont >>
rect -3498 765 -3464 799
rect -3380 765 -3346 799
rect -3262 765 -3228 799
rect -3144 765 -3110 799
rect -3026 765 -2992 799
rect -2908 765 -2874 799
rect -2790 765 -2756 799
rect -2672 765 -2638 799
rect -2554 765 -2520 799
rect -2436 765 -2402 799
rect -2318 765 -2284 799
rect -2200 765 -2166 799
rect -2082 765 -2048 799
rect -1964 765 -1930 799
rect -1846 765 -1812 799
rect -1728 765 -1694 799
rect -1610 765 -1576 799
rect -1492 765 -1458 799
rect -1374 765 -1340 799
rect -1256 765 -1222 799
rect -1138 765 -1104 799
rect -1020 765 -986 799
rect -902 765 -868 799
rect -784 765 -750 799
rect -666 765 -632 799
rect -548 765 -514 799
rect -430 765 -396 799
rect -312 765 -278 799
rect -194 765 -160 799
rect -76 765 -42 799
rect 42 765 76 799
rect 160 765 194 799
rect 278 765 312 799
rect 396 765 430 799
rect 514 765 548 799
rect 632 765 666 799
rect 750 765 784 799
rect 868 765 902 799
rect 986 765 1020 799
rect 1104 765 1138 799
rect 1222 765 1256 799
rect 1340 765 1374 799
rect 1458 765 1492 799
rect 1576 765 1610 799
rect 1694 765 1728 799
rect 1812 765 1846 799
rect 1930 765 1964 799
rect 2048 765 2082 799
rect 2166 765 2200 799
rect 2284 765 2318 799
rect 2402 765 2436 799
rect 2520 765 2554 799
rect 2638 765 2672 799
rect 2756 765 2790 799
rect 2874 765 2908 799
rect 2992 765 3026 799
rect 3110 765 3144 799
rect 3228 765 3262 799
rect 3346 765 3380 799
rect 3464 765 3498 799
rect -3498 37 -3464 71
rect -3380 37 -3346 71
rect -3262 37 -3228 71
rect -3144 37 -3110 71
rect -3026 37 -2992 71
rect -2908 37 -2874 71
rect -2790 37 -2756 71
rect -2672 37 -2638 71
rect -2554 37 -2520 71
rect -2436 37 -2402 71
rect -2318 37 -2284 71
rect -2200 37 -2166 71
rect -2082 37 -2048 71
rect -1964 37 -1930 71
rect -1846 37 -1812 71
rect -1728 37 -1694 71
rect -1610 37 -1576 71
rect -1492 37 -1458 71
rect -1374 37 -1340 71
rect -1256 37 -1222 71
rect -1138 37 -1104 71
rect -1020 37 -986 71
rect -902 37 -868 71
rect -784 37 -750 71
rect -666 37 -632 71
rect -548 37 -514 71
rect -430 37 -396 71
rect -312 37 -278 71
rect -194 37 -160 71
rect -76 37 -42 71
rect 42 37 76 71
rect 160 37 194 71
rect 278 37 312 71
rect 396 37 430 71
rect 514 37 548 71
rect 632 37 666 71
rect 750 37 784 71
rect 868 37 902 71
rect 986 37 1020 71
rect 1104 37 1138 71
rect 1222 37 1256 71
rect 1340 37 1374 71
rect 1458 37 1492 71
rect 1576 37 1610 71
rect 1694 37 1728 71
rect 1812 37 1846 71
rect 1930 37 1964 71
rect 2048 37 2082 71
rect 2166 37 2200 71
rect 2284 37 2318 71
rect 2402 37 2436 71
rect 2520 37 2554 71
rect 2638 37 2672 71
rect 2756 37 2790 71
rect 2874 37 2908 71
rect 2992 37 3026 71
rect 3110 37 3144 71
rect 3228 37 3262 71
rect 3346 37 3380 71
rect 3464 37 3498 71
rect -3498 -71 -3464 -37
rect -3380 -71 -3346 -37
rect -3262 -71 -3228 -37
rect -3144 -71 -3110 -37
rect -3026 -71 -2992 -37
rect -2908 -71 -2874 -37
rect -2790 -71 -2756 -37
rect -2672 -71 -2638 -37
rect -2554 -71 -2520 -37
rect -2436 -71 -2402 -37
rect -2318 -71 -2284 -37
rect -2200 -71 -2166 -37
rect -2082 -71 -2048 -37
rect -1964 -71 -1930 -37
rect -1846 -71 -1812 -37
rect -1728 -71 -1694 -37
rect -1610 -71 -1576 -37
rect -1492 -71 -1458 -37
rect -1374 -71 -1340 -37
rect -1256 -71 -1222 -37
rect -1138 -71 -1104 -37
rect -1020 -71 -986 -37
rect -902 -71 -868 -37
rect -784 -71 -750 -37
rect -666 -71 -632 -37
rect -548 -71 -514 -37
rect -430 -71 -396 -37
rect -312 -71 -278 -37
rect -194 -71 -160 -37
rect -76 -71 -42 -37
rect 42 -71 76 -37
rect 160 -71 194 -37
rect 278 -71 312 -37
rect 396 -71 430 -37
rect 514 -71 548 -37
rect 632 -71 666 -37
rect 750 -71 784 -37
rect 868 -71 902 -37
rect 986 -71 1020 -37
rect 1104 -71 1138 -37
rect 1222 -71 1256 -37
rect 1340 -71 1374 -37
rect 1458 -71 1492 -37
rect 1576 -71 1610 -37
rect 1694 -71 1728 -37
rect 1812 -71 1846 -37
rect 1930 -71 1964 -37
rect 2048 -71 2082 -37
rect 2166 -71 2200 -37
rect 2284 -71 2318 -37
rect 2402 -71 2436 -37
rect 2520 -71 2554 -37
rect 2638 -71 2672 -37
rect 2756 -71 2790 -37
rect 2874 -71 2908 -37
rect 2992 -71 3026 -37
rect 3110 -71 3144 -37
rect 3228 -71 3262 -37
rect 3346 -71 3380 -37
rect 3464 -71 3498 -37
rect -3498 -799 -3464 -765
rect -3380 -799 -3346 -765
rect -3262 -799 -3228 -765
rect -3144 -799 -3110 -765
rect -3026 -799 -2992 -765
rect -2908 -799 -2874 -765
rect -2790 -799 -2756 -765
rect -2672 -799 -2638 -765
rect -2554 -799 -2520 -765
rect -2436 -799 -2402 -765
rect -2318 -799 -2284 -765
rect -2200 -799 -2166 -765
rect -2082 -799 -2048 -765
rect -1964 -799 -1930 -765
rect -1846 -799 -1812 -765
rect -1728 -799 -1694 -765
rect -1610 -799 -1576 -765
rect -1492 -799 -1458 -765
rect -1374 -799 -1340 -765
rect -1256 -799 -1222 -765
rect -1138 -799 -1104 -765
rect -1020 -799 -986 -765
rect -902 -799 -868 -765
rect -784 -799 -750 -765
rect -666 -799 -632 -765
rect -548 -799 -514 -765
rect -430 -799 -396 -765
rect -312 -799 -278 -765
rect -194 -799 -160 -765
rect -76 -799 -42 -765
rect 42 -799 76 -765
rect 160 -799 194 -765
rect 278 -799 312 -765
rect 396 -799 430 -765
rect 514 -799 548 -765
rect 632 -799 666 -765
rect 750 -799 784 -765
rect 868 -799 902 -765
rect 986 -799 1020 -765
rect 1104 -799 1138 -765
rect 1222 -799 1256 -765
rect 1340 -799 1374 -765
rect 1458 -799 1492 -765
rect 1576 -799 1610 -765
rect 1694 -799 1728 -765
rect 1812 -799 1846 -765
rect 1930 -799 1964 -765
rect 2048 -799 2082 -765
rect 2166 -799 2200 -765
rect 2284 -799 2318 -765
rect 2402 -799 2436 -765
rect 2520 -799 2554 -765
rect 2638 -799 2672 -765
rect 2756 -799 2790 -765
rect 2874 -799 2908 -765
rect 2992 -799 3026 -765
rect 3110 -799 3144 -765
rect 3228 -799 3262 -765
rect 3346 -799 3380 -765
rect 3464 -799 3498 -765
<< locali >>
rect -3671 867 -3575 901
rect 3575 867 3671 901
rect -3671 805 -3637 867
rect 3637 805 3671 867
rect -3514 765 -3498 799
rect -3464 765 -3448 799
rect -3396 765 -3380 799
rect -3346 765 -3330 799
rect -3278 765 -3262 799
rect -3228 765 -3212 799
rect -3160 765 -3144 799
rect -3110 765 -3094 799
rect -3042 765 -3026 799
rect -2992 765 -2976 799
rect -2924 765 -2908 799
rect -2874 765 -2858 799
rect -2806 765 -2790 799
rect -2756 765 -2740 799
rect -2688 765 -2672 799
rect -2638 765 -2622 799
rect -2570 765 -2554 799
rect -2520 765 -2504 799
rect -2452 765 -2436 799
rect -2402 765 -2386 799
rect -2334 765 -2318 799
rect -2284 765 -2268 799
rect -2216 765 -2200 799
rect -2166 765 -2150 799
rect -2098 765 -2082 799
rect -2048 765 -2032 799
rect -1980 765 -1964 799
rect -1930 765 -1914 799
rect -1862 765 -1846 799
rect -1812 765 -1796 799
rect -1744 765 -1728 799
rect -1694 765 -1678 799
rect -1626 765 -1610 799
rect -1576 765 -1560 799
rect -1508 765 -1492 799
rect -1458 765 -1442 799
rect -1390 765 -1374 799
rect -1340 765 -1324 799
rect -1272 765 -1256 799
rect -1222 765 -1206 799
rect -1154 765 -1138 799
rect -1104 765 -1088 799
rect -1036 765 -1020 799
rect -986 765 -970 799
rect -918 765 -902 799
rect -868 765 -852 799
rect -800 765 -784 799
rect -750 765 -734 799
rect -682 765 -666 799
rect -632 765 -616 799
rect -564 765 -548 799
rect -514 765 -498 799
rect -446 765 -430 799
rect -396 765 -380 799
rect -328 765 -312 799
rect -278 765 -262 799
rect -210 765 -194 799
rect -160 765 -144 799
rect -92 765 -76 799
rect -42 765 -26 799
rect 26 765 42 799
rect 76 765 92 799
rect 144 765 160 799
rect 194 765 210 799
rect 262 765 278 799
rect 312 765 328 799
rect 380 765 396 799
rect 430 765 446 799
rect 498 765 514 799
rect 548 765 564 799
rect 616 765 632 799
rect 666 765 682 799
rect 734 765 750 799
rect 784 765 800 799
rect 852 765 868 799
rect 902 765 918 799
rect 970 765 986 799
rect 1020 765 1036 799
rect 1088 765 1104 799
rect 1138 765 1154 799
rect 1206 765 1222 799
rect 1256 765 1272 799
rect 1324 765 1340 799
rect 1374 765 1390 799
rect 1442 765 1458 799
rect 1492 765 1508 799
rect 1560 765 1576 799
rect 1610 765 1626 799
rect 1678 765 1694 799
rect 1728 765 1744 799
rect 1796 765 1812 799
rect 1846 765 1862 799
rect 1914 765 1930 799
rect 1964 765 1980 799
rect 2032 765 2048 799
rect 2082 765 2098 799
rect 2150 765 2166 799
rect 2200 765 2216 799
rect 2268 765 2284 799
rect 2318 765 2334 799
rect 2386 765 2402 799
rect 2436 765 2452 799
rect 2504 765 2520 799
rect 2554 765 2570 799
rect 2622 765 2638 799
rect 2672 765 2688 799
rect 2740 765 2756 799
rect 2790 765 2806 799
rect 2858 765 2874 799
rect 2908 765 2924 799
rect 2976 765 2992 799
rect 3026 765 3042 799
rect 3094 765 3110 799
rect 3144 765 3160 799
rect 3212 765 3228 799
rect 3262 765 3278 799
rect 3330 765 3346 799
rect 3380 765 3396 799
rect 3448 765 3464 799
rect 3498 765 3514 799
rect -3557 706 -3523 722
rect -3557 114 -3523 130
rect -3439 706 -3405 722
rect -3439 114 -3405 130
rect -3321 706 -3287 722
rect -3321 114 -3287 130
rect -3203 706 -3169 722
rect -3203 114 -3169 130
rect -3085 706 -3051 722
rect -3085 114 -3051 130
rect -2967 706 -2933 722
rect -2967 114 -2933 130
rect -2849 706 -2815 722
rect -2849 114 -2815 130
rect -2731 706 -2697 722
rect -2731 114 -2697 130
rect -2613 706 -2579 722
rect -2613 114 -2579 130
rect -2495 706 -2461 722
rect -2495 114 -2461 130
rect -2377 706 -2343 722
rect -2377 114 -2343 130
rect -2259 706 -2225 722
rect -2259 114 -2225 130
rect -2141 706 -2107 722
rect -2141 114 -2107 130
rect -2023 706 -1989 722
rect -2023 114 -1989 130
rect -1905 706 -1871 722
rect -1905 114 -1871 130
rect -1787 706 -1753 722
rect -1787 114 -1753 130
rect -1669 706 -1635 722
rect -1669 114 -1635 130
rect -1551 706 -1517 722
rect -1551 114 -1517 130
rect -1433 706 -1399 722
rect -1433 114 -1399 130
rect -1315 706 -1281 722
rect -1315 114 -1281 130
rect -1197 706 -1163 722
rect -1197 114 -1163 130
rect -1079 706 -1045 722
rect -1079 114 -1045 130
rect -961 706 -927 722
rect -961 114 -927 130
rect -843 706 -809 722
rect -843 114 -809 130
rect -725 706 -691 722
rect -725 114 -691 130
rect -607 706 -573 722
rect -607 114 -573 130
rect -489 706 -455 722
rect -489 114 -455 130
rect -371 706 -337 722
rect -371 114 -337 130
rect -253 706 -219 722
rect -253 114 -219 130
rect -135 706 -101 722
rect -135 114 -101 130
rect -17 706 17 722
rect -17 114 17 130
rect 101 706 135 722
rect 101 114 135 130
rect 219 706 253 722
rect 219 114 253 130
rect 337 706 371 722
rect 337 114 371 130
rect 455 706 489 722
rect 455 114 489 130
rect 573 706 607 722
rect 573 114 607 130
rect 691 706 725 722
rect 691 114 725 130
rect 809 706 843 722
rect 809 114 843 130
rect 927 706 961 722
rect 927 114 961 130
rect 1045 706 1079 722
rect 1045 114 1079 130
rect 1163 706 1197 722
rect 1163 114 1197 130
rect 1281 706 1315 722
rect 1281 114 1315 130
rect 1399 706 1433 722
rect 1399 114 1433 130
rect 1517 706 1551 722
rect 1517 114 1551 130
rect 1635 706 1669 722
rect 1635 114 1669 130
rect 1753 706 1787 722
rect 1753 114 1787 130
rect 1871 706 1905 722
rect 1871 114 1905 130
rect 1989 706 2023 722
rect 1989 114 2023 130
rect 2107 706 2141 722
rect 2107 114 2141 130
rect 2225 706 2259 722
rect 2225 114 2259 130
rect 2343 706 2377 722
rect 2343 114 2377 130
rect 2461 706 2495 722
rect 2461 114 2495 130
rect 2579 706 2613 722
rect 2579 114 2613 130
rect 2697 706 2731 722
rect 2697 114 2731 130
rect 2815 706 2849 722
rect 2815 114 2849 130
rect 2933 706 2967 722
rect 2933 114 2967 130
rect 3051 706 3085 722
rect 3051 114 3085 130
rect 3169 706 3203 722
rect 3169 114 3203 130
rect 3287 706 3321 722
rect 3287 114 3321 130
rect 3405 706 3439 722
rect 3405 114 3439 130
rect 3523 706 3557 722
rect 3523 114 3557 130
rect -3514 37 -3498 71
rect -3464 37 -3448 71
rect -3396 37 -3380 71
rect -3346 37 -3330 71
rect -3278 37 -3262 71
rect -3228 37 -3212 71
rect -3160 37 -3144 71
rect -3110 37 -3094 71
rect -3042 37 -3026 71
rect -2992 37 -2976 71
rect -2924 37 -2908 71
rect -2874 37 -2858 71
rect -2806 37 -2790 71
rect -2756 37 -2740 71
rect -2688 37 -2672 71
rect -2638 37 -2622 71
rect -2570 37 -2554 71
rect -2520 37 -2504 71
rect -2452 37 -2436 71
rect -2402 37 -2386 71
rect -2334 37 -2318 71
rect -2284 37 -2268 71
rect -2216 37 -2200 71
rect -2166 37 -2150 71
rect -2098 37 -2082 71
rect -2048 37 -2032 71
rect -1980 37 -1964 71
rect -1930 37 -1914 71
rect -1862 37 -1846 71
rect -1812 37 -1796 71
rect -1744 37 -1728 71
rect -1694 37 -1678 71
rect -1626 37 -1610 71
rect -1576 37 -1560 71
rect -1508 37 -1492 71
rect -1458 37 -1442 71
rect -1390 37 -1374 71
rect -1340 37 -1324 71
rect -1272 37 -1256 71
rect -1222 37 -1206 71
rect -1154 37 -1138 71
rect -1104 37 -1088 71
rect -1036 37 -1020 71
rect -986 37 -970 71
rect -918 37 -902 71
rect -868 37 -852 71
rect -800 37 -784 71
rect -750 37 -734 71
rect -682 37 -666 71
rect -632 37 -616 71
rect -564 37 -548 71
rect -514 37 -498 71
rect -446 37 -430 71
rect -396 37 -380 71
rect -328 37 -312 71
rect -278 37 -262 71
rect -210 37 -194 71
rect -160 37 -144 71
rect -92 37 -76 71
rect -42 37 -26 71
rect 26 37 42 71
rect 76 37 92 71
rect 144 37 160 71
rect 194 37 210 71
rect 262 37 278 71
rect 312 37 328 71
rect 380 37 396 71
rect 430 37 446 71
rect 498 37 514 71
rect 548 37 564 71
rect 616 37 632 71
rect 666 37 682 71
rect 734 37 750 71
rect 784 37 800 71
rect 852 37 868 71
rect 902 37 918 71
rect 970 37 986 71
rect 1020 37 1036 71
rect 1088 37 1104 71
rect 1138 37 1154 71
rect 1206 37 1222 71
rect 1256 37 1272 71
rect 1324 37 1340 71
rect 1374 37 1390 71
rect 1442 37 1458 71
rect 1492 37 1508 71
rect 1560 37 1576 71
rect 1610 37 1626 71
rect 1678 37 1694 71
rect 1728 37 1744 71
rect 1796 37 1812 71
rect 1846 37 1862 71
rect 1914 37 1930 71
rect 1964 37 1980 71
rect 2032 37 2048 71
rect 2082 37 2098 71
rect 2150 37 2166 71
rect 2200 37 2216 71
rect 2268 37 2284 71
rect 2318 37 2334 71
rect 2386 37 2402 71
rect 2436 37 2452 71
rect 2504 37 2520 71
rect 2554 37 2570 71
rect 2622 37 2638 71
rect 2672 37 2688 71
rect 2740 37 2756 71
rect 2790 37 2806 71
rect 2858 37 2874 71
rect 2908 37 2924 71
rect 2976 37 2992 71
rect 3026 37 3042 71
rect 3094 37 3110 71
rect 3144 37 3160 71
rect 3212 37 3228 71
rect 3262 37 3278 71
rect 3330 37 3346 71
rect 3380 37 3396 71
rect 3448 37 3464 71
rect 3498 37 3514 71
rect -3514 -71 -3498 -37
rect -3464 -71 -3448 -37
rect -3396 -71 -3380 -37
rect -3346 -71 -3330 -37
rect -3278 -71 -3262 -37
rect -3228 -71 -3212 -37
rect -3160 -71 -3144 -37
rect -3110 -71 -3094 -37
rect -3042 -71 -3026 -37
rect -2992 -71 -2976 -37
rect -2924 -71 -2908 -37
rect -2874 -71 -2858 -37
rect -2806 -71 -2790 -37
rect -2756 -71 -2740 -37
rect -2688 -71 -2672 -37
rect -2638 -71 -2622 -37
rect -2570 -71 -2554 -37
rect -2520 -71 -2504 -37
rect -2452 -71 -2436 -37
rect -2402 -71 -2386 -37
rect -2334 -71 -2318 -37
rect -2284 -71 -2268 -37
rect -2216 -71 -2200 -37
rect -2166 -71 -2150 -37
rect -2098 -71 -2082 -37
rect -2048 -71 -2032 -37
rect -1980 -71 -1964 -37
rect -1930 -71 -1914 -37
rect -1862 -71 -1846 -37
rect -1812 -71 -1796 -37
rect -1744 -71 -1728 -37
rect -1694 -71 -1678 -37
rect -1626 -71 -1610 -37
rect -1576 -71 -1560 -37
rect -1508 -71 -1492 -37
rect -1458 -71 -1442 -37
rect -1390 -71 -1374 -37
rect -1340 -71 -1324 -37
rect -1272 -71 -1256 -37
rect -1222 -71 -1206 -37
rect -1154 -71 -1138 -37
rect -1104 -71 -1088 -37
rect -1036 -71 -1020 -37
rect -986 -71 -970 -37
rect -918 -71 -902 -37
rect -868 -71 -852 -37
rect -800 -71 -784 -37
rect -750 -71 -734 -37
rect -682 -71 -666 -37
rect -632 -71 -616 -37
rect -564 -71 -548 -37
rect -514 -71 -498 -37
rect -446 -71 -430 -37
rect -396 -71 -380 -37
rect -328 -71 -312 -37
rect -278 -71 -262 -37
rect -210 -71 -194 -37
rect -160 -71 -144 -37
rect -92 -71 -76 -37
rect -42 -71 -26 -37
rect 26 -71 42 -37
rect 76 -71 92 -37
rect 144 -71 160 -37
rect 194 -71 210 -37
rect 262 -71 278 -37
rect 312 -71 328 -37
rect 380 -71 396 -37
rect 430 -71 446 -37
rect 498 -71 514 -37
rect 548 -71 564 -37
rect 616 -71 632 -37
rect 666 -71 682 -37
rect 734 -71 750 -37
rect 784 -71 800 -37
rect 852 -71 868 -37
rect 902 -71 918 -37
rect 970 -71 986 -37
rect 1020 -71 1036 -37
rect 1088 -71 1104 -37
rect 1138 -71 1154 -37
rect 1206 -71 1222 -37
rect 1256 -71 1272 -37
rect 1324 -71 1340 -37
rect 1374 -71 1390 -37
rect 1442 -71 1458 -37
rect 1492 -71 1508 -37
rect 1560 -71 1576 -37
rect 1610 -71 1626 -37
rect 1678 -71 1694 -37
rect 1728 -71 1744 -37
rect 1796 -71 1812 -37
rect 1846 -71 1862 -37
rect 1914 -71 1930 -37
rect 1964 -71 1980 -37
rect 2032 -71 2048 -37
rect 2082 -71 2098 -37
rect 2150 -71 2166 -37
rect 2200 -71 2216 -37
rect 2268 -71 2284 -37
rect 2318 -71 2334 -37
rect 2386 -71 2402 -37
rect 2436 -71 2452 -37
rect 2504 -71 2520 -37
rect 2554 -71 2570 -37
rect 2622 -71 2638 -37
rect 2672 -71 2688 -37
rect 2740 -71 2756 -37
rect 2790 -71 2806 -37
rect 2858 -71 2874 -37
rect 2908 -71 2924 -37
rect 2976 -71 2992 -37
rect 3026 -71 3042 -37
rect 3094 -71 3110 -37
rect 3144 -71 3160 -37
rect 3212 -71 3228 -37
rect 3262 -71 3278 -37
rect 3330 -71 3346 -37
rect 3380 -71 3396 -37
rect 3448 -71 3464 -37
rect 3498 -71 3514 -37
rect -3557 -130 -3523 -114
rect -3557 -722 -3523 -706
rect -3439 -130 -3405 -114
rect -3439 -722 -3405 -706
rect -3321 -130 -3287 -114
rect -3321 -722 -3287 -706
rect -3203 -130 -3169 -114
rect -3203 -722 -3169 -706
rect -3085 -130 -3051 -114
rect -3085 -722 -3051 -706
rect -2967 -130 -2933 -114
rect -2967 -722 -2933 -706
rect -2849 -130 -2815 -114
rect -2849 -722 -2815 -706
rect -2731 -130 -2697 -114
rect -2731 -722 -2697 -706
rect -2613 -130 -2579 -114
rect -2613 -722 -2579 -706
rect -2495 -130 -2461 -114
rect -2495 -722 -2461 -706
rect -2377 -130 -2343 -114
rect -2377 -722 -2343 -706
rect -2259 -130 -2225 -114
rect -2259 -722 -2225 -706
rect -2141 -130 -2107 -114
rect -2141 -722 -2107 -706
rect -2023 -130 -1989 -114
rect -2023 -722 -1989 -706
rect -1905 -130 -1871 -114
rect -1905 -722 -1871 -706
rect -1787 -130 -1753 -114
rect -1787 -722 -1753 -706
rect -1669 -130 -1635 -114
rect -1669 -722 -1635 -706
rect -1551 -130 -1517 -114
rect -1551 -722 -1517 -706
rect -1433 -130 -1399 -114
rect -1433 -722 -1399 -706
rect -1315 -130 -1281 -114
rect -1315 -722 -1281 -706
rect -1197 -130 -1163 -114
rect -1197 -722 -1163 -706
rect -1079 -130 -1045 -114
rect -1079 -722 -1045 -706
rect -961 -130 -927 -114
rect -961 -722 -927 -706
rect -843 -130 -809 -114
rect -843 -722 -809 -706
rect -725 -130 -691 -114
rect -725 -722 -691 -706
rect -607 -130 -573 -114
rect -607 -722 -573 -706
rect -489 -130 -455 -114
rect -489 -722 -455 -706
rect -371 -130 -337 -114
rect -371 -722 -337 -706
rect -253 -130 -219 -114
rect -253 -722 -219 -706
rect -135 -130 -101 -114
rect -135 -722 -101 -706
rect -17 -130 17 -114
rect -17 -722 17 -706
rect 101 -130 135 -114
rect 101 -722 135 -706
rect 219 -130 253 -114
rect 219 -722 253 -706
rect 337 -130 371 -114
rect 337 -722 371 -706
rect 455 -130 489 -114
rect 455 -722 489 -706
rect 573 -130 607 -114
rect 573 -722 607 -706
rect 691 -130 725 -114
rect 691 -722 725 -706
rect 809 -130 843 -114
rect 809 -722 843 -706
rect 927 -130 961 -114
rect 927 -722 961 -706
rect 1045 -130 1079 -114
rect 1045 -722 1079 -706
rect 1163 -130 1197 -114
rect 1163 -722 1197 -706
rect 1281 -130 1315 -114
rect 1281 -722 1315 -706
rect 1399 -130 1433 -114
rect 1399 -722 1433 -706
rect 1517 -130 1551 -114
rect 1517 -722 1551 -706
rect 1635 -130 1669 -114
rect 1635 -722 1669 -706
rect 1753 -130 1787 -114
rect 1753 -722 1787 -706
rect 1871 -130 1905 -114
rect 1871 -722 1905 -706
rect 1989 -130 2023 -114
rect 1989 -722 2023 -706
rect 2107 -130 2141 -114
rect 2107 -722 2141 -706
rect 2225 -130 2259 -114
rect 2225 -722 2259 -706
rect 2343 -130 2377 -114
rect 2343 -722 2377 -706
rect 2461 -130 2495 -114
rect 2461 -722 2495 -706
rect 2579 -130 2613 -114
rect 2579 -722 2613 -706
rect 2697 -130 2731 -114
rect 2697 -722 2731 -706
rect 2815 -130 2849 -114
rect 2815 -722 2849 -706
rect 2933 -130 2967 -114
rect 2933 -722 2967 -706
rect 3051 -130 3085 -114
rect 3051 -722 3085 -706
rect 3169 -130 3203 -114
rect 3169 -722 3203 -706
rect 3287 -130 3321 -114
rect 3287 -722 3321 -706
rect 3405 -130 3439 -114
rect 3405 -722 3439 -706
rect 3523 -130 3557 -114
rect 3523 -722 3557 -706
rect -3514 -799 -3498 -765
rect -3464 -799 -3448 -765
rect -3396 -799 -3380 -765
rect -3346 -799 -3330 -765
rect -3278 -799 -3262 -765
rect -3228 -799 -3212 -765
rect -3160 -799 -3144 -765
rect -3110 -799 -3094 -765
rect -3042 -799 -3026 -765
rect -2992 -799 -2976 -765
rect -2924 -799 -2908 -765
rect -2874 -799 -2858 -765
rect -2806 -799 -2790 -765
rect -2756 -799 -2740 -765
rect -2688 -799 -2672 -765
rect -2638 -799 -2622 -765
rect -2570 -799 -2554 -765
rect -2520 -799 -2504 -765
rect -2452 -799 -2436 -765
rect -2402 -799 -2386 -765
rect -2334 -799 -2318 -765
rect -2284 -799 -2268 -765
rect -2216 -799 -2200 -765
rect -2166 -799 -2150 -765
rect -2098 -799 -2082 -765
rect -2048 -799 -2032 -765
rect -1980 -799 -1964 -765
rect -1930 -799 -1914 -765
rect -1862 -799 -1846 -765
rect -1812 -799 -1796 -765
rect -1744 -799 -1728 -765
rect -1694 -799 -1678 -765
rect -1626 -799 -1610 -765
rect -1576 -799 -1560 -765
rect -1508 -799 -1492 -765
rect -1458 -799 -1442 -765
rect -1390 -799 -1374 -765
rect -1340 -799 -1324 -765
rect -1272 -799 -1256 -765
rect -1222 -799 -1206 -765
rect -1154 -799 -1138 -765
rect -1104 -799 -1088 -765
rect -1036 -799 -1020 -765
rect -986 -799 -970 -765
rect -918 -799 -902 -765
rect -868 -799 -852 -765
rect -800 -799 -784 -765
rect -750 -799 -734 -765
rect -682 -799 -666 -765
rect -632 -799 -616 -765
rect -564 -799 -548 -765
rect -514 -799 -498 -765
rect -446 -799 -430 -765
rect -396 -799 -380 -765
rect -328 -799 -312 -765
rect -278 -799 -262 -765
rect -210 -799 -194 -765
rect -160 -799 -144 -765
rect -92 -799 -76 -765
rect -42 -799 -26 -765
rect 26 -799 42 -765
rect 76 -799 92 -765
rect 144 -799 160 -765
rect 194 -799 210 -765
rect 262 -799 278 -765
rect 312 -799 328 -765
rect 380 -799 396 -765
rect 430 -799 446 -765
rect 498 -799 514 -765
rect 548 -799 564 -765
rect 616 -799 632 -765
rect 666 -799 682 -765
rect 734 -799 750 -765
rect 784 -799 800 -765
rect 852 -799 868 -765
rect 902 -799 918 -765
rect 970 -799 986 -765
rect 1020 -799 1036 -765
rect 1088 -799 1104 -765
rect 1138 -799 1154 -765
rect 1206 -799 1222 -765
rect 1256 -799 1272 -765
rect 1324 -799 1340 -765
rect 1374 -799 1390 -765
rect 1442 -799 1458 -765
rect 1492 -799 1508 -765
rect 1560 -799 1576 -765
rect 1610 -799 1626 -765
rect 1678 -799 1694 -765
rect 1728 -799 1744 -765
rect 1796 -799 1812 -765
rect 1846 -799 1862 -765
rect 1914 -799 1930 -765
rect 1964 -799 1980 -765
rect 2032 -799 2048 -765
rect 2082 -799 2098 -765
rect 2150 -799 2166 -765
rect 2200 -799 2216 -765
rect 2268 -799 2284 -765
rect 2318 -799 2334 -765
rect 2386 -799 2402 -765
rect 2436 -799 2452 -765
rect 2504 -799 2520 -765
rect 2554 -799 2570 -765
rect 2622 -799 2638 -765
rect 2672 -799 2688 -765
rect 2740 -799 2756 -765
rect 2790 -799 2806 -765
rect 2858 -799 2874 -765
rect 2908 -799 2924 -765
rect 2976 -799 2992 -765
rect 3026 -799 3042 -765
rect 3094 -799 3110 -765
rect 3144 -799 3160 -765
rect 3212 -799 3228 -765
rect 3262 -799 3278 -765
rect 3330 -799 3346 -765
rect 3380 -799 3396 -765
rect 3448 -799 3464 -765
rect 3498 -799 3514 -765
rect -3671 -867 -3637 -805
rect 3637 -867 3671 -805
rect -3671 -901 -3575 -867
rect 3575 -901 3671 -867
<< viali >>
rect -3498 765 -3464 799
rect -3380 765 -3346 799
rect -3262 765 -3228 799
rect -3144 765 -3110 799
rect -3026 765 -2992 799
rect -2908 765 -2874 799
rect -2790 765 -2756 799
rect -2672 765 -2638 799
rect -2554 765 -2520 799
rect -2436 765 -2402 799
rect -2318 765 -2284 799
rect -2200 765 -2166 799
rect -2082 765 -2048 799
rect -1964 765 -1930 799
rect -1846 765 -1812 799
rect -1728 765 -1694 799
rect -1610 765 -1576 799
rect -1492 765 -1458 799
rect -1374 765 -1340 799
rect -1256 765 -1222 799
rect -1138 765 -1104 799
rect -1020 765 -986 799
rect -902 765 -868 799
rect -784 765 -750 799
rect -666 765 -632 799
rect -548 765 -514 799
rect -430 765 -396 799
rect -312 765 -278 799
rect -194 765 -160 799
rect -76 765 -42 799
rect 42 765 76 799
rect 160 765 194 799
rect 278 765 312 799
rect 396 765 430 799
rect 514 765 548 799
rect 632 765 666 799
rect 750 765 784 799
rect 868 765 902 799
rect 986 765 1020 799
rect 1104 765 1138 799
rect 1222 765 1256 799
rect 1340 765 1374 799
rect 1458 765 1492 799
rect 1576 765 1610 799
rect 1694 765 1728 799
rect 1812 765 1846 799
rect 1930 765 1964 799
rect 2048 765 2082 799
rect 2166 765 2200 799
rect 2284 765 2318 799
rect 2402 765 2436 799
rect 2520 765 2554 799
rect 2638 765 2672 799
rect 2756 765 2790 799
rect 2874 765 2908 799
rect 2992 765 3026 799
rect 3110 765 3144 799
rect 3228 765 3262 799
rect 3346 765 3380 799
rect 3464 765 3498 799
rect -3557 130 -3523 706
rect -3439 130 -3405 706
rect -3321 130 -3287 706
rect -3203 130 -3169 706
rect -3085 130 -3051 706
rect -2967 130 -2933 706
rect -2849 130 -2815 706
rect -2731 130 -2697 706
rect -2613 130 -2579 706
rect -2495 130 -2461 706
rect -2377 130 -2343 706
rect -2259 130 -2225 706
rect -2141 130 -2107 706
rect -2023 130 -1989 706
rect -1905 130 -1871 706
rect -1787 130 -1753 706
rect -1669 130 -1635 706
rect -1551 130 -1517 706
rect -1433 130 -1399 706
rect -1315 130 -1281 706
rect -1197 130 -1163 706
rect -1079 130 -1045 706
rect -961 130 -927 706
rect -843 130 -809 706
rect -725 130 -691 706
rect -607 130 -573 706
rect -489 130 -455 706
rect -371 130 -337 706
rect -253 130 -219 706
rect -135 130 -101 706
rect -17 130 17 706
rect 101 130 135 706
rect 219 130 253 706
rect 337 130 371 706
rect 455 130 489 706
rect 573 130 607 706
rect 691 130 725 706
rect 809 130 843 706
rect 927 130 961 706
rect 1045 130 1079 706
rect 1163 130 1197 706
rect 1281 130 1315 706
rect 1399 130 1433 706
rect 1517 130 1551 706
rect 1635 130 1669 706
rect 1753 130 1787 706
rect 1871 130 1905 706
rect 1989 130 2023 706
rect 2107 130 2141 706
rect 2225 130 2259 706
rect 2343 130 2377 706
rect 2461 130 2495 706
rect 2579 130 2613 706
rect 2697 130 2731 706
rect 2815 130 2849 706
rect 2933 130 2967 706
rect 3051 130 3085 706
rect 3169 130 3203 706
rect 3287 130 3321 706
rect 3405 130 3439 706
rect 3523 130 3557 706
rect -3498 37 -3464 71
rect -3380 37 -3346 71
rect -3262 37 -3228 71
rect -3144 37 -3110 71
rect -3026 37 -2992 71
rect -2908 37 -2874 71
rect -2790 37 -2756 71
rect -2672 37 -2638 71
rect -2554 37 -2520 71
rect -2436 37 -2402 71
rect -2318 37 -2284 71
rect -2200 37 -2166 71
rect -2082 37 -2048 71
rect -1964 37 -1930 71
rect -1846 37 -1812 71
rect -1728 37 -1694 71
rect -1610 37 -1576 71
rect -1492 37 -1458 71
rect -1374 37 -1340 71
rect -1256 37 -1222 71
rect -1138 37 -1104 71
rect -1020 37 -986 71
rect -902 37 -868 71
rect -784 37 -750 71
rect -666 37 -632 71
rect -548 37 -514 71
rect -430 37 -396 71
rect -312 37 -278 71
rect -194 37 -160 71
rect -76 37 -42 71
rect 42 37 76 71
rect 160 37 194 71
rect 278 37 312 71
rect 396 37 430 71
rect 514 37 548 71
rect 632 37 666 71
rect 750 37 784 71
rect 868 37 902 71
rect 986 37 1020 71
rect 1104 37 1138 71
rect 1222 37 1256 71
rect 1340 37 1374 71
rect 1458 37 1492 71
rect 1576 37 1610 71
rect 1694 37 1728 71
rect 1812 37 1846 71
rect 1930 37 1964 71
rect 2048 37 2082 71
rect 2166 37 2200 71
rect 2284 37 2318 71
rect 2402 37 2436 71
rect 2520 37 2554 71
rect 2638 37 2672 71
rect 2756 37 2790 71
rect 2874 37 2908 71
rect 2992 37 3026 71
rect 3110 37 3144 71
rect 3228 37 3262 71
rect 3346 37 3380 71
rect 3464 37 3498 71
rect -3498 -71 -3464 -37
rect -3380 -71 -3346 -37
rect -3262 -71 -3228 -37
rect -3144 -71 -3110 -37
rect -3026 -71 -2992 -37
rect -2908 -71 -2874 -37
rect -2790 -71 -2756 -37
rect -2672 -71 -2638 -37
rect -2554 -71 -2520 -37
rect -2436 -71 -2402 -37
rect -2318 -71 -2284 -37
rect -2200 -71 -2166 -37
rect -2082 -71 -2048 -37
rect -1964 -71 -1930 -37
rect -1846 -71 -1812 -37
rect -1728 -71 -1694 -37
rect -1610 -71 -1576 -37
rect -1492 -71 -1458 -37
rect -1374 -71 -1340 -37
rect -1256 -71 -1222 -37
rect -1138 -71 -1104 -37
rect -1020 -71 -986 -37
rect -902 -71 -868 -37
rect -784 -71 -750 -37
rect -666 -71 -632 -37
rect -548 -71 -514 -37
rect -430 -71 -396 -37
rect -312 -71 -278 -37
rect -194 -71 -160 -37
rect -76 -71 -42 -37
rect 42 -71 76 -37
rect 160 -71 194 -37
rect 278 -71 312 -37
rect 396 -71 430 -37
rect 514 -71 548 -37
rect 632 -71 666 -37
rect 750 -71 784 -37
rect 868 -71 902 -37
rect 986 -71 1020 -37
rect 1104 -71 1138 -37
rect 1222 -71 1256 -37
rect 1340 -71 1374 -37
rect 1458 -71 1492 -37
rect 1576 -71 1610 -37
rect 1694 -71 1728 -37
rect 1812 -71 1846 -37
rect 1930 -71 1964 -37
rect 2048 -71 2082 -37
rect 2166 -71 2200 -37
rect 2284 -71 2318 -37
rect 2402 -71 2436 -37
rect 2520 -71 2554 -37
rect 2638 -71 2672 -37
rect 2756 -71 2790 -37
rect 2874 -71 2908 -37
rect 2992 -71 3026 -37
rect 3110 -71 3144 -37
rect 3228 -71 3262 -37
rect 3346 -71 3380 -37
rect 3464 -71 3498 -37
rect -3557 -706 -3523 -130
rect -3439 -706 -3405 -130
rect -3321 -706 -3287 -130
rect -3203 -706 -3169 -130
rect -3085 -706 -3051 -130
rect -2967 -706 -2933 -130
rect -2849 -706 -2815 -130
rect -2731 -706 -2697 -130
rect -2613 -706 -2579 -130
rect -2495 -706 -2461 -130
rect -2377 -706 -2343 -130
rect -2259 -706 -2225 -130
rect -2141 -706 -2107 -130
rect -2023 -706 -1989 -130
rect -1905 -706 -1871 -130
rect -1787 -706 -1753 -130
rect -1669 -706 -1635 -130
rect -1551 -706 -1517 -130
rect -1433 -706 -1399 -130
rect -1315 -706 -1281 -130
rect -1197 -706 -1163 -130
rect -1079 -706 -1045 -130
rect -961 -706 -927 -130
rect -843 -706 -809 -130
rect -725 -706 -691 -130
rect -607 -706 -573 -130
rect -489 -706 -455 -130
rect -371 -706 -337 -130
rect -253 -706 -219 -130
rect -135 -706 -101 -130
rect -17 -706 17 -130
rect 101 -706 135 -130
rect 219 -706 253 -130
rect 337 -706 371 -130
rect 455 -706 489 -130
rect 573 -706 607 -130
rect 691 -706 725 -130
rect 809 -706 843 -130
rect 927 -706 961 -130
rect 1045 -706 1079 -130
rect 1163 -706 1197 -130
rect 1281 -706 1315 -130
rect 1399 -706 1433 -130
rect 1517 -706 1551 -130
rect 1635 -706 1669 -130
rect 1753 -706 1787 -130
rect 1871 -706 1905 -130
rect 1989 -706 2023 -130
rect 2107 -706 2141 -130
rect 2225 -706 2259 -130
rect 2343 -706 2377 -130
rect 2461 -706 2495 -130
rect 2579 -706 2613 -130
rect 2697 -706 2731 -130
rect 2815 -706 2849 -130
rect 2933 -706 2967 -130
rect 3051 -706 3085 -130
rect 3169 -706 3203 -130
rect 3287 -706 3321 -130
rect 3405 -706 3439 -130
rect 3523 -706 3557 -130
rect -3498 -799 -3464 -765
rect -3380 -799 -3346 -765
rect -3262 -799 -3228 -765
rect -3144 -799 -3110 -765
rect -3026 -799 -2992 -765
rect -2908 -799 -2874 -765
rect -2790 -799 -2756 -765
rect -2672 -799 -2638 -765
rect -2554 -799 -2520 -765
rect -2436 -799 -2402 -765
rect -2318 -799 -2284 -765
rect -2200 -799 -2166 -765
rect -2082 -799 -2048 -765
rect -1964 -799 -1930 -765
rect -1846 -799 -1812 -765
rect -1728 -799 -1694 -765
rect -1610 -799 -1576 -765
rect -1492 -799 -1458 -765
rect -1374 -799 -1340 -765
rect -1256 -799 -1222 -765
rect -1138 -799 -1104 -765
rect -1020 -799 -986 -765
rect -902 -799 -868 -765
rect -784 -799 -750 -765
rect -666 -799 -632 -765
rect -548 -799 -514 -765
rect -430 -799 -396 -765
rect -312 -799 -278 -765
rect -194 -799 -160 -765
rect -76 -799 -42 -765
rect 42 -799 76 -765
rect 160 -799 194 -765
rect 278 -799 312 -765
rect 396 -799 430 -765
rect 514 -799 548 -765
rect 632 -799 666 -765
rect 750 -799 784 -765
rect 868 -799 902 -765
rect 986 -799 1020 -765
rect 1104 -799 1138 -765
rect 1222 -799 1256 -765
rect 1340 -799 1374 -765
rect 1458 -799 1492 -765
rect 1576 -799 1610 -765
rect 1694 -799 1728 -765
rect 1812 -799 1846 -765
rect 1930 -799 1964 -765
rect 2048 -799 2082 -765
rect 2166 -799 2200 -765
rect 2284 -799 2318 -765
rect 2402 -799 2436 -765
rect 2520 -799 2554 -765
rect 2638 -799 2672 -765
rect 2756 -799 2790 -765
rect 2874 -799 2908 -765
rect 2992 -799 3026 -765
rect 3110 -799 3144 -765
rect 3228 -799 3262 -765
rect 3346 -799 3380 -765
rect 3464 -799 3498 -765
<< metal1 >>
rect -3510 799 -3452 805
rect -3510 765 -3498 799
rect -3464 765 -3452 799
rect -3510 759 -3452 765
rect -3392 799 -3334 805
rect -3392 765 -3380 799
rect -3346 765 -3334 799
rect -3392 759 -3334 765
rect -3274 799 -3216 805
rect -3274 765 -3262 799
rect -3228 765 -3216 799
rect -3274 759 -3216 765
rect -3156 799 -3098 805
rect -3156 765 -3144 799
rect -3110 765 -3098 799
rect -3156 759 -3098 765
rect -3038 799 -2980 805
rect -3038 765 -3026 799
rect -2992 765 -2980 799
rect -3038 759 -2980 765
rect -2920 799 -2862 805
rect -2920 765 -2908 799
rect -2874 765 -2862 799
rect -2920 759 -2862 765
rect -2802 799 -2744 805
rect -2802 765 -2790 799
rect -2756 765 -2744 799
rect -2802 759 -2744 765
rect -2684 799 -2626 805
rect -2684 765 -2672 799
rect -2638 765 -2626 799
rect -2684 759 -2626 765
rect -2566 799 -2508 805
rect -2566 765 -2554 799
rect -2520 765 -2508 799
rect -2566 759 -2508 765
rect -2448 799 -2390 805
rect -2448 765 -2436 799
rect -2402 765 -2390 799
rect -2448 759 -2390 765
rect -2330 799 -2272 805
rect -2330 765 -2318 799
rect -2284 765 -2272 799
rect -2330 759 -2272 765
rect -2212 799 -2154 805
rect -2212 765 -2200 799
rect -2166 765 -2154 799
rect -2212 759 -2154 765
rect -2094 799 -2036 805
rect -2094 765 -2082 799
rect -2048 765 -2036 799
rect -2094 759 -2036 765
rect -1976 799 -1918 805
rect -1976 765 -1964 799
rect -1930 765 -1918 799
rect -1976 759 -1918 765
rect -1858 799 -1800 805
rect -1858 765 -1846 799
rect -1812 765 -1800 799
rect -1858 759 -1800 765
rect -1740 799 -1682 805
rect -1740 765 -1728 799
rect -1694 765 -1682 799
rect -1740 759 -1682 765
rect -1622 799 -1564 805
rect -1622 765 -1610 799
rect -1576 765 -1564 799
rect -1622 759 -1564 765
rect -1504 799 -1446 805
rect -1504 765 -1492 799
rect -1458 765 -1446 799
rect -1504 759 -1446 765
rect -1386 799 -1328 805
rect -1386 765 -1374 799
rect -1340 765 -1328 799
rect -1386 759 -1328 765
rect -1268 799 -1210 805
rect -1268 765 -1256 799
rect -1222 765 -1210 799
rect -1268 759 -1210 765
rect -1150 799 -1092 805
rect -1150 765 -1138 799
rect -1104 765 -1092 799
rect -1150 759 -1092 765
rect -1032 799 -974 805
rect -1032 765 -1020 799
rect -986 765 -974 799
rect -1032 759 -974 765
rect -914 799 -856 805
rect -914 765 -902 799
rect -868 765 -856 799
rect -914 759 -856 765
rect -796 799 -738 805
rect -796 765 -784 799
rect -750 765 -738 799
rect -796 759 -738 765
rect -678 799 -620 805
rect -678 765 -666 799
rect -632 765 -620 799
rect -678 759 -620 765
rect -560 799 -502 805
rect -560 765 -548 799
rect -514 765 -502 799
rect -560 759 -502 765
rect -442 799 -384 805
rect -442 765 -430 799
rect -396 765 -384 799
rect -442 759 -384 765
rect -324 799 -266 805
rect -324 765 -312 799
rect -278 765 -266 799
rect -324 759 -266 765
rect -206 799 -148 805
rect -206 765 -194 799
rect -160 765 -148 799
rect -206 759 -148 765
rect -88 799 -30 805
rect -88 765 -76 799
rect -42 765 -30 799
rect -88 759 -30 765
rect 30 799 88 805
rect 30 765 42 799
rect 76 765 88 799
rect 30 759 88 765
rect 148 799 206 805
rect 148 765 160 799
rect 194 765 206 799
rect 148 759 206 765
rect 266 799 324 805
rect 266 765 278 799
rect 312 765 324 799
rect 266 759 324 765
rect 384 799 442 805
rect 384 765 396 799
rect 430 765 442 799
rect 384 759 442 765
rect 502 799 560 805
rect 502 765 514 799
rect 548 765 560 799
rect 502 759 560 765
rect 620 799 678 805
rect 620 765 632 799
rect 666 765 678 799
rect 620 759 678 765
rect 738 799 796 805
rect 738 765 750 799
rect 784 765 796 799
rect 738 759 796 765
rect 856 799 914 805
rect 856 765 868 799
rect 902 765 914 799
rect 856 759 914 765
rect 974 799 1032 805
rect 974 765 986 799
rect 1020 765 1032 799
rect 974 759 1032 765
rect 1092 799 1150 805
rect 1092 765 1104 799
rect 1138 765 1150 799
rect 1092 759 1150 765
rect 1210 799 1268 805
rect 1210 765 1222 799
rect 1256 765 1268 799
rect 1210 759 1268 765
rect 1328 799 1386 805
rect 1328 765 1340 799
rect 1374 765 1386 799
rect 1328 759 1386 765
rect 1446 799 1504 805
rect 1446 765 1458 799
rect 1492 765 1504 799
rect 1446 759 1504 765
rect 1564 799 1622 805
rect 1564 765 1576 799
rect 1610 765 1622 799
rect 1564 759 1622 765
rect 1682 799 1740 805
rect 1682 765 1694 799
rect 1728 765 1740 799
rect 1682 759 1740 765
rect 1800 799 1858 805
rect 1800 765 1812 799
rect 1846 765 1858 799
rect 1800 759 1858 765
rect 1918 799 1976 805
rect 1918 765 1930 799
rect 1964 765 1976 799
rect 1918 759 1976 765
rect 2036 799 2094 805
rect 2036 765 2048 799
rect 2082 765 2094 799
rect 2036 759 2094 765
rect 2154 799 2212 805
rect 2154 765 2166 799
rect 2200 765 2212 799
rect 2154 759 2212 765
rect 2272 799 2330 805
rect 2272 765 2284 799
rect 2318 765 2330 799
rect 2272 759 2330 765
rect 2390 799 2448 805
rect 2390 765 2402 799
rect 2436 765 2448 799
rect 2390 759 2448 765
rect 2508 799 2566 805
rect 2508 765 2520 799
rect 2554 765 2566 799
rect 2508 759 2566 765
rect 2626 799 2684 805
rect 2626 765 2638 799
rect 2672 765 2684 799
rect 2626 759 2684 765
rect 2744 799 2802 805
rect 2744 765 2756 799
rect 2790 765 2802 799
rect 2744 759 2802 765
rect 2862 799 2920 805
rect 2862 765 2874 799
rect 2908 765 2920 799
rect 2862 759 2920 765
rect 2980 799 3038 805
rect 2980 765 2992 799
rect 3026 765 3038 799
rect 2980 759 3038 765
rect 3098 799 3156 805
rect 3098 765 3110 799
rect 3144 765 3156 799
rect 3098 759 3156 765
rect 3216 799 3274 805
rect 3216 765 3228 799
rect 3262 765 3274 799
rect 3216 759 3274 765
rect 3334 799 3392 805
rect 3334 765 3346 799
rect 3380 765 3392 799
rect 3334 759 3392 765
rect 3452 799 3510 805
rect 3452 765 3464 799
rect 3498 765 3510 799
rect 3452 759 3510 765
rect -3563 706 -3517 718
rect -3563 130 -3557 706
rect -3523 130 -3517 706
rect -3563 118 -3517 130
rect -3445 706 -3399 718
rect -3445 130 -3439 706
rect -3405 130 -3399 706
rect -3445 118 -3399 130
rect -3327 706 -3281 718
rect -3327 130 -3321 706
rect -3287 130 -3281 706
rect -3327 118 -3281 130
rect -3209 706 -3163 718
rect -3209 130 -3203 706
rect -3169 130 -3163 706
rect -3209 118 -3163 130
rect -3091 706 -3045 718
rect -3091 130 -3085 706
rect -3051 130 -3045 706
rect -3091 118 -3045 130
rect -2973 706 -2927 718
rect -2973 130 -2967 706
rect -2933 130 -2927 706
rect -2973 118 -2927 130
rect -2855 706 -2809 718
rect -2855 130 -2849 706
rect -2815 130 -2809 706
rect -2855 118 -2809 130
rect -2737 706 -2691 718
rect -2737 130 -2731 706
rect -2697 130 -2691 706
rect -2737 118 -2691 130
rect -2619 706 -2573 718
rect -2619 130 -2613 706
rect -2579 130 -2573 706
rect -2619 118 -2573 130
rect -2501 706 -2455 718
rect -2501 130 -2495 706
rect -2461 130 -2455 706
rect -2501 118 -2455 130
rect -2383 706 -2337 718
rect -2383 130 -2377 706
rect -2343 130 -2337 706
rect -2383 118 -2337 130
rect -2265 706 -2219 718
rect -2265 130 -2259 706
rect -2225 130 -2219 706
rect -2265 118 -2219 130
rect -2147 706 -2101 718
rect -2147 130 -2141 706
rect -2107 130 -2101 706
rect -2147 118 -2101 130
rect -2029 706 -1983 718
rect -2029 130 -2023 706
rect -1989 130 -1983 706
rect -2029 118 -1983 130
rect -1911 706 -1865 718
rect -1911 130 -1905 706
rect -1871 130 -1865 706
rect -1911 118 -1865 130
rect -1793 706 -1747 718
rect -1793 130 -1787 706
rect -1753 130 -1747 706
rect -1793 118 -1747 130
rect -1675 706 -1629 718
rect -1675 130 -1669 706
rect -1635 130 -1629 706
rect -1675 118 -1629 130
rect -1557 706 -1511 718
rect -1557 130 -1551 706
rect -1517 130 -1511 706
rect -1557 118 -1511 130
rect -1439 706 -1393 718
rect -1439 130 -1433 706
rect -1399 130 -1393 706
rect -1439 118 -1393 130
rect -1321 706 -1275 718
rect -1321 130 -1315 706
rect -1281 130 -1275 706
rect -1321 118 -1275 130
rect -1203 706 -1157 718
rect -1203 130 -1197 706
rect -1163 130 -1157 706
rect -1203 118 -1157 130
rect -1085 706 -1039 718
rect -1085 130 -1079 706
rect -1045 130 -1039 706
rect -1085 118 -1039 130
rect -967 706 -921 718
rect -967 130 -961 706
rect -927 130 -921 706
rect -967 118 -921 130
rect -849 706 -803 718
rect -849 130 -843 706
rect -809 130 -803 706
rect -849 118 -803 130
rect -731 706 -685 718
rect -731 130 -725 706
rect -691 130 -685 706
rect -731 118 -685 130
rect -613 706 -567 718
rect -613 130 -607 706
rect -573 130 -567 706
rect -613 118 -567 130
rect -495 706 -449 718
rect -495 130 -489 706
rect -455 130 -449 706
rect -495 118 -449 130
rect -377 706 -331 718
rect -377 130 -371 706
rect -337 130 -331 706
rect -377 118 -331 130
rect -259 706 -213 718
rect -259 130 -253 706
rect -219 130 -213 706
rect -259 118 -213 130
rect -141 706 -95 718
rect -141 130 -135 706
rect -101 130 -95 706
rect -141 118 -95 130
rect -23 706 23 718
rect -23 130 -17 706
rect 17 130 23 706
rect -23 118 23 130
rect 95 706 141 718
rect 95 130 101 706
rect 135 130 141 706
rect 95 118 141 130
rect 213 706 259 718
rect 213 130 219 706
rect 253 130 259 706
rect 213 118 259 130
rect 331 706 377 718
rect 331 130 337 706
rect 371 130 377 706
rect 331 118 377 130
rect 449 706 495 718
rect 449 130 455 706
rect 489 130 495 706
rect 449 118 495 130
rect 567 706 613 718
rect 567 130 573 706
rect 607 130 613 706
rect 567 118 613 130
rect 685 706 731 718
rect 685 130 691 706
rect 725 130 731 706
rect 685 118 731 130
rect 803 706 849 718
rect 803 130 809 706
rect 843 130 849 706
rect 803 118 849 130
rect 921 706 967 718
rect 921 130 927 706
rect 961 130 967 706
rect 921 118 967 130
rect 1039 706 1085 718
rect 1039 130 1045 706
rect 1079 130 1085 706
rect 1039 118 1085 130
rect 1157 706 1203 718
rect 1157 130 1163 706
rect 1197 130 1203 706
rect 1157 118 1203 130
rect 1275 706 1321 718
rect 1275 130 1281 706
rect 1315 130 1321 706
rect 1275 118 1321 130
rect 1393 706 1439 718
rect 1393 130 1399 706
rect 1433 130 1439 706
rect 1393 118 1439 130
rect 1511 706 1557 718
rect 1511 130 1517 706
rect 1551 130 1557 706
rect 1511 118 1557 130
rect 1629 706 1675 718
rect 1629 130 1635 706
rect 1669 130 1675 706
rect 1629 118 1675 130
rect 1747 706 1793 718
rect 1747 130 1753 706
rect 1787 130 1793 706
rect 1747 118 1793 130
rect 1865 706 1911 718
rect 1865 130 1871 706
rect 1905 130 1911 706
rect 1865 118 1911 130
rect 1983 706 2029 718
rect 1983 130 1989 706
rect 2023 130 2029 706
rect 1983 118 2029 130
rect 2101 706 2147 718
rect 2101 130 2107 706
rect 2141 130 2147 706
rect 2101 118 2147 130
rect 2219 706 2265 718
rect 2219 130 2225 706
rect 2259 130 2265 706
rect 2219 118 2265 130
rect 2337 706 2383 718
rect 2337 130 2343 706
rect 2377 130 2383 706
rect 2337 118 2383 130
rect 2455 706 2501 718
rect 2455 130 2461 706
rect 2495 130 2501 706
rect 2455 118 2501 130
rect 2573 706 2619 718
rect 2573 130 2579 706
rect 2613 130 2619 706
rect 2573 118 2619 130
rect 2691 706 2737 718
rect 2691 130 2697 706
rect 2731 130 2737 706
rect 2691 118 2737 130
rect 2809 706 2855 718
rect 2809 130 2815 706
rect 2849 130 2855 706
rect 2809 118 2855 130
rect 2927 706 2973 718
rect 2927 130 2933 706
rect 2967 130 2973 706
rect 2927 118 2973 130
rect 3045 706 3091 718
rect 3045 130 3051 706
rect 3085 130 3091 706
rect 3045 118 3091 130
rect 3163 706 3209 718
rect 3163 130 3169 706
rect 3203 130 3209 706
rect 3163 118 3209 130
rect 3281 706 3327 718
rect 3281 130 3287 706
rect 3321 130 3327 706
rect 3281 118 3327 130
rect 3399 706 3445 718
rect 3399 130 3405 706
rect 3439 130 3445 706
rect 3399 118 3445 130
rect 3517 706 3563 718
rect 3517 130 3523 706
rect 3557 130 3563 706
rect 3517 118 3563 130
rect -3510 71 -3452 77
rect -3510 37 -3498 71
rect -3464 37 -3452 71
rect -3510 31 -3452 37
rect -3392 71 -3334 77
rect -3392 37 -3380 71
rect -3346 37 -3334 71
rect -3392 31 -3334 37
rect -3274 71 -3216 77
rect -3274 37 -3262 71
rect -3228 37 -3216 71
rect -3274 31 -3216 37
rect -3156 71 -3098 77
rect -3156 37 -3144 71
rect -3110 37 -3098 71
rect -3156 31 -3098 37
rect -3038 71 -2980 77
rect -3038 37 -3026 71
rect -2992 37 -2980 71
rect -3038 31 -2980 37
rect -2920 71 -2862 77
rect -2920 37 -2908 71
rect -2874 37 -2862 71
rect -2920 31 -2862 37
rect -2802 71 -2744 77
rect -2802 37 -2790 71
rect -2756 37 -2744 71
rect -2802 31 -2744 37
rect -2684 71 -2626 77
rect -2684 37 -2672 71
rect -2638 37 -2626 71
rect -2684 31 -2626 37
rect -2566 71 -2508 77
rect -2566 37 -2554 71
rect -2520 37 -2508 71
rect -2566 31 -2508 37
rect -2448 71 -2390 77
rect -2448 37 -2436 71
rect -2402 37 -2390 71
rect -2448 31 -2390 37
rect -2330 71 -2272 77
rect -2330 37 -2318 71
rect -2284 37 -2272 71
rect -2330 31 -2272 37
rect -2212 71 -2154 77
rect -2212 37 -2200 71
rect -2166 37 -2154 71
rect -2212 31 -2154 37
rect -2094 71 -2036 77
rect -2094 37 -2082 71
rect -2048 37 -2036 71
rect -2094 31 -2036 37
rect -1976 71 -1918 77
rect -1976 37 -1964 71
rect -1930 37 -1918 71
rect -1976 31 -1918 37
rect -1858 71 -1800 77
rect -1858 37 -1846 71
rect -1812 37 -1800 71
rect -1858 31 -1800 37
rect -1740 71 -1682 77
rect -1740 37 -1728 71
rect -1694 37 -1682 71
rect -1740 31 -1682 37
rect -1622 71 -1564 77
rect -1622 37 -1610 71
rect -1576 37 -1564 71
rect -1622 31 -1564 37
rect -1504 71 -1446 77
rect -1504 37 -1492 71
rect -1458 37 -1446 71
rect -1504 31 -1446 37
rect -1386 71 -1328 77
rect -1386 37 -1374 71
rect -1340 37 -1328 71
rect -1386 31 -1328 37
rect -1268 71 -1210 77
rect -1268 37 -1256 71
rect -1222 37 -1210 71
rect -1268 31 -1210 37
rect -1150 71 -1092 77
rect -1150 37 -1138 71
rect -1104 37 -1092 71
rect -1150 31 -1092 37
rect -1032 71 -974 77
rect -1032 37 -1020 71
rect -986 37 -974 71
rect -1032 31 -974 37
rect -914 71 -856 77
rect -914 37 -902 71
rect -868 37 -856 71
rect -914 31 -856 37
rect -796 71 -738 77
rect -796 37 -784 71
rect -750 37 -738 71
rect -796 31 -738 37
rect -678 71 -620 77
rect -678 37 -666 71
rect -632 37 -620 71
rect -678 31 -620 37
rect -560 71 -502 77
rect -560 37 -548 71
rect -514 37 -502 71
rect -560 31 -502 37
rect -442 71 -384 77
rect -442 37 -430 71
rect -396 37 -384 71
rect -442 31 -384 37
rect -324 71 -266 77
rect -324 37 -312 71
rect -278 37 -266 71
rect -324 31 -266 37
rect -206 71 -148 77
rect -206 37 -194 71
rect -160 37 -148 71
rect -206 31 -148 37
rect -88 71 -30 77
rect -88 37 -76 71
rect -42 37 -30 71
rect -88 31 -30 37
rect 30 71 88 77
rect 30 37 42 71
rect 76 37 88 71
rect 30 31 88 37
rect 148 71 206 77
rect 148 37 160 71
rect 194 37 206 71
rect 148 31 206 37
rect 266 71 324 77
rect 266 37 278 71
rect 312 37 324 71
rect 266 31 324 37
rect 384 71 442 77
rect 384 37 396 71
rect 430 37 442 71
rect 384 31 442 37
rect 502 71 560 77
rect 502 37 514 71
rect 548 37 560 71
rect 502 31 560 37
rect 620 71 678 77
rect 620 37 632 71
rect 666 37 678 71
rect 620 31 678 37
rect 738 71 796 77
rect 738 37 750 71
rect 784 37 796 71
rect 738 31 796 37
rect 856 71 914 77
rect 856 37 868 71
rect 902 37 914 71
rect 856 31 914 37
rect 974 71 1032 77
rect 974 37 986 71
rect 1020 37 1032 71
rect 974 31 1032 37
rect 1092 71 1150 77
rect 1092 37 1104 71
rect 1138 37 1150 71
rect 1092 31 1150 37
rect 1210 71 1268 77
rect 1210 37 1222 71
rect 1256 37 1268 71
rect 1210 31 1268 37
rect 1328 71 1386 77
rect 1328 37 1340 71
rect 1374 37 1386 71
rect 1328 31 1386 37
rect 1446 71 1504 77
rect 1446 37 1458 71
rect 1492 37 1504 71
rect 1446 31 1504 37
rect 1564 71 1622 77
rect 1564 37 1576 71
rect 1610 37 1622 71
rect 1564 31 1622 37
rect 1682 71 1740 77
rect 1682 37 1694 71
rect 1728 37 1740 71
rect 1682 31 1740 37
rect 1800 71 1858 77
rect 1800 37 1812 71
rect 1846 37 1858 71
rect 1800 31 1858 37
rect 1918 71 1976 77
rect 1918 37 1930 71
rect 1964 37 1976 71
rect 1918 31 1976 37
rect 2036 71 2094 77
rect 2036 37 2048 71
rect 2082 37 2094 71
rect 2036 31 2094 37
rect 2154 71 2212 77
rect 2154 37 2166 71
rect 2200 37 2212 71
rect 2154 31 2212 37
rect 2272 71 2330 77
rect 2272 37 2284 71
rect 2318 37 2330 71
rect 2272 31 2330 37
rect 2390 71 2448 77
rect 2390 37 2402 71
rect 2436 37 2448 71
rect 2390 31 2448 37
rect 2508 71 2566 77
rect 2508 37 2520 71
rect 2554 37 2566 71
rect 2508 31 2566 37
rect 2626 71 2684 77
rect 2626 37 2638 71
rect 2672 37 2684 71
rect 2626 31 2684 37
rect 2744 71 2802 77
rect 2744 37 2756 71
rect 2790 37 2802 71
rect 2744 31 2802 37
rect 2862 71 2920 77
rect 2862 37 2874 71
rect 2908 37 2920 71
rect 2862 31 2920 37
rect 2980 71 3038 77
rect 2980 37 2992 71
rect 3026 37 3038 71
rect 2980 31 3038 37
rect 3098 71 3156 77
rect 3098 37 3110 71
rect 3144 37 3156 71
rect 3098 31 3156 37
rect 3216 71 3274 77
rect 3216 37 3228 71
rect 3262 37 3274 71
rect 3216 31 3274 37
rect 3334 71 3392 77
rect 3334 37 3346 71
rect 3380 37 3392 71
rect 3334 31 3392 37
rect 3452 71 3510 77
rect 3452 37 3464 71
rect 3498 37 3510 71
rect 3452 31 3510 37
rect -3510 -37 -3452 -31
rect -3510 -71 -3498 -37
rect -3464 -71 -3452 -37
rect -3510 -77 -3452 -71
rect -3392 -37 -3334 -31
rect -3392 -71 -3380 -37
rect -3346 -71 -3334 -37
rect -3392 -77 -3334 -71
rect -3274 -37 -3216 -31
rect -3274 -71 -3262 -37
rect -3228 -71 -3216 -37
rect -3274 -77 -3216 -71
rect -3156 -37 -3098 -31
rect -3156 -71 -3144 -37
rect -3110 -71 -3098 -37
rect -3156 -77 -3098 -71
rect -3038 -37 -2980 -31
rect -3038 -71 -3026 -37
rect -2992 -71 -2980 -37
rect -3038 -77 -2980 -71
rect -2920 -37 -2862 -31
rect -2920 -71 -2908 -37
rect -2874 -71 -2862 -37
rect -2920 -77 -2862 -71
rect -2802 -37 -2744 -31
rect -2802 -71 -2790 -37
rect -2756 -71 -2744 -37
rect -2802 -77 -2744 -71
rect -2684 -37 -2626 -31
rect -2684 -71 -2672 -37
rect -2638 -71 -2626 -37
rect -2684 -77 -2626 -71
rect -2566 -37 -2508 -31
rect -2566 -71 -2554 -37
rect -2520 -71 -2508 -37
rect -2566 -77 -2508 -71
rect -2448 -37 -2390 -31
rect -2448 -71 -2436 -37
rect -2402 -71 -2390 -37
rect -2448 -77 -2390 -71
rect -2330 -37 -2272 -31
rect -2330 -71 -2318 -37
rect -2284 -71 -2272 -37
rect -2330 -77 -2272 -71
rect -2212 -37 -2154 -31
rect -2212 -71 -2200 -37
rect -2166 -71 -2154 -37
rect -2212 -77 -2154 -71
rect -2094 -37 -2036 -31
rect -2094 -71 -2082 -37
rect -2048 -71 -2036 -37
rect -2094 -77 -2036 -71
rect -1976 -37 -1918 -31
rect -1976 -71 -1964 -37
rect -1930 -71 -1918 -37
rect -1976 -77 -1918 -71
rect -1858 -37 -1800 -31
rect -1858 -71 -1846 -37
rect -1812 -71 -1800 -37
rect -1858 -77 -1800 -71
rect -1740 -37 -1682 -31
rect -1740 -71 -1728 -37
rect -1694 -71 -1682 -37
rect -1740 -77 -1682 -71
rect -1622 -37 -1564 -31
rect -1622 -71 -1610 -37
rect -1576 -71 -1564 -37
rect -1622 -77 -1564 -71
rect -1504 -37 -1446 -31
rect -1504 -71 -1492 -37
rect -1458 -71 -1446 -37
rect -1504 -77 -1446 -71
rect -1386 -37 -1328 -31
rect -1386 -71 -1374 -37
rect -1340 -71 -1328 -37
rect -1386 -77 -1328 -71
rect -1268 -37 -1210 -31
rect -1268 -71 -1256 -37
rect -1222 -71 -1210 -37
rect -1268 -77 -1210 -71
rect -1150 -37 -1092 -31
rect -1150 -71 -1138 -37
rect -1104 -71 -1092 -37
rect -1150 -77 -1092 -71
rect -1032 -37 -974 -31
rect -1032 -71 -1020 -37
rect -986 -71 -974 -37
rect -1032 -77 -974 -71
rect -914 -37 -856 -31
rect -914 -71 -902 -37
rect -868 -71 -856 -37
rect -914 -77 -856 -71
rect -796 -37 -738 -31
rect -796 -71 -784 -37
rect -750 -71 -738 -37
rect -796 -77 -738 -71
rect -678 -37 -620 -31
rect -678 -71 -666 -37
rect -632 -71 -620 -37
rect -678 -77 -620 -71
rect -560 -37 -502 -31
rect -560 -71 -548 -37
rect -514 -71 -502 -37
rect -560 -77 -502 -71
rect -442 -37 -384 -31
rect -442 -71 -430 -37
rect -396 -71 -384 -37
rect -442 -77 -384 -71
rect -324 -37 -266 -31
rect -324 -71 -312 -37
rect -278 -71 -266 -37
rect -324 -77 -266 -71
rect -206 -37 -148 -31
rect -206 -71 -194 -37
rect -160 -71 -148 -37
rect -206 -77 -148 -71
rect -88 -37 -30 -31
rect -88 -71 -76 -37
rect -42 -71 -30 -37
rect -88 -77 -30 -71
rect 30 -37 88 -31
rect 30 -71 42 -37
rect 76 -71 88 -37
rect 30 -77 88 -71
rect 148 -37 206 -31
rect 148 -71 160 -37
rect 194 -71 206 -37
rect 148 -77 206 -71
rect 266 -37 324 -31
rect 266 -71 278 -37
rect 312 -71 324 -37
rect 266 -77 324 -71
rect 384 -37 442 -31
rect 384 -71 396 -37
rect 430 -71 442 -37
rect 384 -77 442 -71
rect 502 -37 560 -31
rect 502 -71 514 -37
rect 548 -71 560 -37
rect 502 -77 560 -71
rect 620 -37 678 -31
rect 620 -71 632 -37
rect 666 -71 678 -37
rect 620 -77 678 -71
rect 738 -37 796 -31
rect 738 -71 750 -37
rect 784 -71 796 -37
rect 738 -77 796 -71
rect 856 -37 914 -31
rect 856 -71 868 -37
rect 902 -71 914 -37
rect 856 -77 914 -71
rect 974 -37 1032 -31
rect 974 -71 986 -37
rect 1020 -71 1032 -37
rect 974 -77 1032 -71
rect 1092 -37 1150 -31
rect 1092 -71 1104 -37
rect 1138 -71 1150 -37
rect 1092 -77 1150 -71
rect 1210 -37 1268 -31
rect 1210 -71 1222 -37
rect 1256 -71 1268 -37
rect 1210 -77 1268 -71
rect 1328 -37 1386 -31
rect 1328 -71 1340 -37
rect 1374 -71 1386 -37
rect 1328 -77 1386 -71
rect 1446 -37 1504 -31
rect 1446 -71 1458 -37
rect 1492 -71 1504 -37
rect 1446 -77 1504 -71
rect 1564 -37 1622 -31
rect 1564 -71 1576 -37
rect 1610 -71 1622 -37
rect 1564 -77 1622 -71
rect 1682 -37 1740 -31
rect 1682 -71 1694 -37
rect 1728 -71 1740 -37
rect 1682 -77 1740 -71
rect 1800 -37 1858 -31
rect 1800 -71 1812 -37
rect 1846 -71 1858 -37
rect 1800 -77 1858 -71
rect 1918 -37 1976 -31
rect 1918 -71 1930 -37
rect 1964 -71 1976 -37
rect 1918 -77 1976 -71
rect 2036 -37 2094 -31
rect 2036 -71 2048 -37
rect 2082 -71 2094 -37
rect 2036 -77 2094 -71
rect 2154 -37 2212 -31
rect 2154 -71 2166 -37
rect 2200 -71 2212 -37
rect 2154 -77 2212 -71
rect 2272 -37 2330 -31
rect 2272 -71 2284 -37
rect 2318 -71 2330 -37
rect 2272 -77 2330 -71
rect 2390 -37 2448 -31
rect 2390 -71 2402 -37
rect 2436 -71 2448 -37
rect 2390 -77 2448 -71
rect 2508 -37 2566 -31
rect 2508 -71 2520 -37
rect 2554 -71 2566 -37
rect 2508 -77 2566 -71
rect 2626 -37 2684 -31
rect 2626 -71 2638 -37
rect 2672 -71 2684 -37
rect 2626 -77 2684 -71
rect 2744 -37 2802 -31
rect 2744 -71 2756 -37
rect 2790 -71 2802 -37
rect 2744 -77 2802 -71
rect 2862 -37 2920 -31
rect 2862 -71 2874 -37
rect 2908 -71 2920 -37
rect 2862 -77 2920 -71
rect 2980 -37 3038 -31
rect 2980 -71 2992 -37
rect 3026 -71 3038 -37
rect 2980 -77 3038 -71
rect 3098 -37 3156 -31
rect 3098 -71 3110 -37
rect 3144 -71 3156 -37
rect 3098 -77 3156 -71
rect 3216 -37 3274 -31
rect 3216 -71 3228 -37
rect 3262 -71 3274 -37
rect 3216 -77 3274 -71
rect 3334 -37 3392 -31
rect 3334 -71 3346 -37
rect 3380 -71 3392 -37
rect 3334 -77 3392 -71
rect 3452 -37 3510 -31
rect 3452 -71 3464 -37
rect 3498 -71 3510 -37
rect 3452 -77 3510 -71
rect -3563 -130 -3517 -118
rect -3563 -706 -3557 -130
rect -3523 -706 -3517 -130
rect -3563 -718 -3517 -706
rect -3445 -130 -3399 -118
rect -3445 -706 -3439 -130
rect -3405 -706 -3399 -130
rect -3445 -718 -3399 -706
rect -3327 -130 -3281 -118
rect -3327 -706 -3321 -130
rect -3287 -706 -3281 -130
rect -3327 -718 -3281 -706
rect -3209 -130 -3163 -118
rect -3209 -706 -3203 -130
rect -3169 -706 -3163 -130
rect -3209 -718 -3163 -706
rect -3091 -130 -3045 -118
rect -3091 -706 -3085 -130
rect -3051 -706 -3045 -130
rect -3091 -718 -3045 -706
rect -2973 -130 -2927 -118
rect -2973 -706 -2967 -130
rect -2933 -706 -2927 -130
rect -2973 -718 -2927 -706
rect -2855 -130 -2809 -118
rect -2855 -706 -2849 -130
rect -2815 -706 -2809 -130
rect -2855 -718 -2809 -706
rect -2737 -130 -2691 -118
rect -2737 -706 -2731 -130
rect -2697 -706 -2691 -130
rect -2737 -718 -2691 -706
rect -2619 -130 -2573 -118
rect -2619 -706 -2613 -130
rect -2579 -706 -2573 -130
rect -2619 -718 -2573 -706
rect -2501 -130 -2455 -118
rect -2501 -706 -2495 -130
rect -2461 -706 -2455 -130
rect -2501 -718 -2455 -706
rect -2383 -130 -2337 -118
rect -2383 -706 -2377 -130
rect -2343 -706 -2337 -130
rect -2383 -718 -2337 -706
rect -2265 -130 -2219 -118
rect -2265 -706 -2259 -130
rect -2225 -706 -2219 -130
rect -2265 -718 -2219 -706
rect -2147 -130 -2101 -118
rect -2147 -706 -2141 -130
rect -2107 -706 -2101 -130
rect -2147 -718 -2101 -706
rect -2029 -130 -1983 -118
rect -2029 -706 -2023 -130
rect -1989 -706 -1983 -130
rect -2029 -718 -1983 -706
rect -1911 -130 -1865 -118
rect -1911 -706 -1905 -130
rect -1871 -706 -1865 -130
rect -1911 -718 -1865 -706
rect -1793 -130 -1747 -118
rect -1793 -706 -1787 -130
rect -1753 -706 -1747 -130
rect -1793 -718 -1747 -706
rect -1675 -130 -1629 -118
rect -1675 -706 -1669 -130
rect -1635 -706 -1629 -130
rect -1675 -718 -1629 -706
rect -1557 -130 -1511 -118
rect -1557 -706 -1551 -130
rect -1517 -706 -1511 -130
rect -1557 -718 -1511 -706
rect -1439 -130 -1393 -118
rect -1439 -706 -1433 -130
rect -1399 -706 -1393 -130
rect -1439 -718 -1393 -706
rect -1321 -130 -1275 -118
rect -1321 -706 -1315 -130
rect -1281 -706 -1275 -130
rect -1321 -718 -1275 -706
rect -1203 -130 -1157 -118
rect -1203 -706 -1197 -130
rect -1163 -706 -1157 -130
rect -1203 -718 -1157 -706
rect -1085 -130 -1039 -118
rect -1085 -706 -1079 -130
rect -1045 -706 -1039 -130
rect -1085 -718 -1039 -706
rect -967 -130 -921 -118
rect -967 -706 -961 -130
rect -927 -706 -921 -130
rect -967 -718 -921 -706
rect -849 -130 -803 -118
rect -849 -706 -843 -130
rect -809 -706 -803 -130
rect -849 -718 -803 -706
rect -731 -130 -685 -118
rect -731 -706 -725 -130
rect -691 -706 -685 -130
rect -731 -718 -685 -706
rect -613 -130 -567 -118
rect -613 -706 -607 -130
rect -573 -706 -567 -130
rect -613 -718 -567 -706
rect -495 -130 -449 -118
rect -495 -706 -489 -130
rect -455 -706 -449 -130
rect -495 -718 -449 -706
rect -377 -130 -331 -118
rect -377 -706 -371 -130
rect -337 -706 -331 -130
rect -377 -718 -331 -706
rect -259 -130 -213 -118
rect -259 -706 -253 -130
rect -219 -706 -213 -130
rect -259 -718 -213 -706
rect -141 -130 -95 -118
rect -141 -706 -135 -130
rect -101 -706 -95 -130
rect -141 -718 -95 -706
rect -23 -130 23 -118
rect -23 -706 -17 -130
rect 17 -706 23 -130
rect -23 -718 23 -706
rect 95 -130 141 -118
rect 95 -706 101 -130
rect 135 -706 141 -130
rect 95 -718 141 -706
rect 213 -130 259 -118
rect 213 -706 219 -130
rect 253 -706 259 -130
rect 213 -718 259 -706
rect 331 -130 377 -118
rect 331 -706 337 -130
rect 371 -706 377 -130
rect 331 -718 377 -706
rect 449 -130 495 -118
rect 449 -706 455 -130
rect 489 -706 495 -130
rect 449 -718 495 -706
rect 567 -130 613 -118
rect 567 -706 573 -130
rect 607 -706 613 -130
rect 567 -718 613 -706
rect 685 -130 731 -118
rect 685 -706 691 -130
rect 725 -706 731 -130
rect 685 -718 731 -706
rect 803 -130 849 -118
rect 803 -706 809 -130
rect 843 -706 849 -130
rect 803 -718 849 -706
rect 921 -130 967 -118
rect 921 -706 927 -130
rect 961 -706 967 -130
rect 921 -718 967 -706
rect 1039 -130 1085 -118
rect 1039 -706 1045 -130
rect 1079 -706 1085 -130
rect 1039 -718 1085 -706
rect 1157 -130 1203 -118
rect 1157 -706 1163 -130
rect 1197 -706 1203 -130
rect 1157 -718 1203 -706
rect 1275 -130 1321 -118
rect 1275 -706 1281 -130
rect 1315 -706 1321 -130
rect 1275 -718 1321 -706
rect 1393 -130 1439 -118
rect 1393 -706 1399 -130
rect 1433 -706 1439 -130
rect 1393 -718 1439 -706
rect 1511 -130 1557 -118
rect 1511 -706 1517 -130
rect 1551 -706 1557 -130
rect 1511 -718 1557 -706
rect 1629 -130 1675 -118
rect 1629 -706 1635 -130
rect 1669 -706 1675 -130
rect 1629 -718 1675 -706
rect 1747 -130 1793 -118
rect 1747 -706 1753 -130
rect 1787 -706 1793 -130
rect 1747 -718 1793 -706
rect 1865 -130 1911 -118
rect 1865 -706 1871 -130
rect 1905 -706 1911 -130
rect 1865 -718 1911 -706
rect 1983 -130 2029 -118
rect 1983 -706 1989 -130
rect 2023 -706 2029 -130
rect 1983 -718 2029 -706
rect 2101 -130 2147 -118
rect 2101 -706 2107 -130
rect 2141 -706 2147 -130
rect 2101 -718 2147 -706
rect 2219 -130 2265 -118
rect 2219 -706 2225 -130
rect 2259 -706 2265 -130
rect 2219 -718 2265 -706
rect 2337 -130 2383 -118
rect 2337 -706 2343 -130
rect 2377 -706 2383 -130
rect 2337 -718 2383 -706
rect 2455 -130 2501 -118
rect 2455 -706 2461 -130
rect 2495 -706 2501 -130
rect 2455 -718 2501 -706
rect 2573 -130 2619 -118
rect 2573 -706 2579 -130
rect 2613 -706 2619 -130
rect 2573 -718 2619 -706
rect 2691 -130 2737 -118
rect 2691 -706 2697 -130
rect 2731 -706 2737 -130
rect 2691 -718 2737 -706
rect 2809 -130 2855 -118
rect 2809 -706 2815 -130
rect 2849 -706 2855 -130
rect 2809 -718 2855 -706
rect 2927 -130 2973 -118
rect 2927 -706 2933 -130
rect 2967 -706 2973 -130
rect 2927 -718 2973 -706
rect 3045 -130 3091 -118
rect 3045 -706 3051 -130
rect 3085 -706 3091 -130
rect 3045 -718 3091 -706
rect 3163 -130 3209 -118
rect 3163 -706 3169 -130
rect 3203 -706 3209 -130
rect 3163 -718 3209 -706
rect 3281 -130 3327 -118
rect 3281 -706 3287 -130
rect 3321 -706 3327 -130
rect 3281 -718 3327 -706
rect 3399 -130 3445 -118
rect 3399 -706 3405 -130
rect 3439 -706 3445 -130
rect 3399 -718 3445 -706
rect 3517 -130 3563 -118
rect 3517 -706 3523 -130
rect 3557 -706 3563 -130
rect 3517 -718 3563 -706
rect -3510 -765 -3452 -759
rect -3510 -799 -3498 -765
rect -3464 -799 -3452 -765
rect -3510 -805 -3452 -799
rect -3392 -765 -3334 -759
rect -3392 -799 -3380 -765
rect -3346 -799 -3334 -765
rect -3392 -805 -3334 -799
rect -3274 -765 -3216 -759
rect -3274 -799 -3262 -765
rect -3228 -799 -3216 -765
rect -3274 -805 -3216 -799
rect -3156 -765 -3098 -759
rect -3156 -799 -3144 -765
rect -3110 -799 -3098 -765
rect -3156 -805 -3098 -799
rect -3038 -765 -2980 -759
rect -3038 -799 -3026 -765
rect -2992 -799 -2980 -765
rect -3038 -805 -2980 -799
rect -2920 -765 -2862 -759
rect -2920 -799 -2908 -765
rect -2874 -799 -2862 -765
rect -2920 -805 -2862 -799
rect -2802 -765 -2744 -759
rect -2802 -799 -2790 -765
rect -2756 -799 -2744 -765
rect -2802 -805 -2744 -799
rect -2684 -765 -2626 -759
rect -2684 -799 -2672 -765
rect -2638 -799 -2626 -765
rect -2684 -805 -2626 -799
rect -2566 -765 -2508 -759
rect -2566 -799 -2554 -765
rect -2520 -799 -2508 -765
rect -2566 -805 -2508 -799
rect -2448 -765 -2390 -759
rect -2448 -799 -2436 -765
rect -2402 -799 -2390 -765
rect -2448 -805 -2390 -799
rect -2330 -765 -2272 -759
rect -2330 -799 -2318 -765
rect -2284 -799 -2272 -765
rect -2330 -805 -2272 -799
rect -2212 -765 -2154 -759
rect -2212 -799 -2200 -765
rect -2166 -799 -2154 -765
rect -2212 -805 -2154 -799
rect -2094 -765 -2036 -759
rect -2094 -799 -2082 -765
rect -2048 -799 -2036 -765
rect -2094 -805 -2036 -799
rect -1976 -765 -1918 -759
rect -1976 -799 -1964 -765
rect -1930 -799 -1918 -765
rect -1976 -805 -1918 -799
rect -1858 -765 -1800 -759
rect -1858 -799 -1846 -765
rect -1812 -799 -1800 -765
rect -1858 -805 -1800 -799
rect -1740 -765 -1682 -759
rect -1740 -799 -1728 -765
rect -1694 -799 -1682 -765
rect -1740 -805 -1682 -799
rect -1622 -765 -1564 -759
rect -1622 -799 -1610 -765
rect -1576 -799 -1564 -765
rect -1622 -805 -1564 -799
rect -1504 -765 -1446 -759
rect -1504 -799 -1492 -765
rect -1458 -799 -1446 -765
rect -1504 -805 -1446 -799
rect -1386 -765 -1328 -759
rect -1386 -799 -1374 -765
rect -1340 -799 -1328 -765
rect -1386 -805 -1328 -799
rect -1268 -765 -1210 -759
rect -1268 -799 -1256 -765
rect -1222 -799 -1210 -765
rect -1268 -805 -1210 -799
rect -1150 -765 -1092 -759
rect -1150 -799 -1138 -765
rect -1104 -799 -1092 -765
rect -1150 -805 -1092 -799
rect -1032 -765 -974 -759
rect -1032 -799 -1020 -765
rect -986 -799 -974 -765
rect -1032 -805 -974 -799
rect -914 -765 -856 -759
rect -914 -799 -902 -765
rect -868 -799 -856 -765
rect -914 -805 -856 -799
rect -796 -765 -738 -759
rect -796 -799 -784 -765
rect -750 -799 -738 -765
rect -796 -805 -738 -799
rect -678 -765 -620 -759
rect -678 -799 -666 -765
rect -632 -799 -620 -765
rect -678 -805 -620 -799
rect -560 -765 -502 -759
rect -560 -799 -548 -765
rect -514 -799 -502 -765
rect -560 -805 -502 -799
rect -442 -765 -384 -759
rect -442 -799 -430 -765
rect -396 -799 -384 -765
rect -442 -805 -384 -799
rect -324 -765 -266 -759
rect -324 -799 -312 -765
rect -278 -799 -266 -765
rect -324 -805 -266 -799
rect -206 -765 -148 -759
rect -206 -799 -194 -765
rect -160 -799 -148 -765
rect -206 -805 -148 -799
rect -88 -765 -30 -759
rect -88 -799 -76 -765
rect -42 -799 -30 -765
rect -88 -805 -30 -799
rect 30 -765 88 -759
rect 30 -799 42 -765
rect 76 -799 88 -765
rect 30 -805 88 -799
rect 148 -765 206 -759
rect 148 -799 160 -765
rect 194 -799 206 -765
rect 148 -805 206 -799
rect 266 -765 324 -759
rect 266 -799 278 -765
rect 312 -799 324 -765
rect 266 -805 324 -799
rect 384 -765 442 -759
rect 384 -799 396 -765
rect 430 -799 442 -765
rect 384 -805 442 -799
rect 502 -765 560 -759
rect 502 -799 514 -765
rect 548 -799 560 -765
rect 502 -805 560 -799
rect 620 -765 678 -759
rect 620 -799 632 -765
rect 666 -799 678 -765
rect 620 -805 678 -799
rect 738 -765 796 -759
rect 738 -799 750 -765
rect 784 -799 796 -765
rect 738 -805 796 -799
rect 856 -765 914 -759
rect 856 -799 868 -765
rect 902 -799 914 -765
rect 856 -805 914 -799
rect 974 -765 1032 -759
rect 974 -799 986 -765
rect 1020 -799 1032 -765
rect 974 -805 1032 -799
rect 1092 -765 1150 -759
rect 1092 -799 1104 -765
rect 1138 -799 1150 -765
rect 1092 -805 1150 -799
rect 1210 -765 1268 -759
rect 1210 -799 1222 -765
rect 1256 -799 1268 -765
rect 1210 -805 1268 -799
rect 1328 -765 1386 -759
rect 1328 -799 1340 -765
rect 1374 -799 1386 -765
rect 1328 -805 1386 -799
rect 1446 -765 1504 -759
rect 1446 -799 1458 -765
rect 1492 -799 1504 -765
rect 1446 -805 1504 -799
rect 1564 -765 1622 -759
rect 1564 -799 1576 -765
rect 1610 -799 1622 -765
rect 1564 -805 1622 -799
rect 1682 -765 1740 -759
rect 1682 -799 1694 -765
rect 1728 -799 1740 -765
rect 1682 -805 1740 -799
rect 1800 -765 1858 -759
rect 1800 -799 1812 -765
rect 1846 -799 1858 -765
rect 1800 -805 1858 -799
rect 1918 -765 1976 -759
rect 1918 -799 1930 -765
rect 1964 -799 1976 -765
rect 1918 -805 1976 -799
rect 2036 -765 2094 -759
rect 2036 -799 2048 -765
rect 2082 -799 2094 -765
rect 2036 -805 2094 -799
rect 2154 -765 2212 -759
rect 2154 -799 2166 -765
rect 2200 -799 2212 -765
rect 2154 -805 2212 -799
rect 2272 -765 2330 -759
rect 2272 -799 2284 -765
rect 2318 -799 2330 -765
rect 2272 -805 2330 -799
rect 2390 -765 2448 -759
rect 2390 -799 2402 -765
rect 2436 -799 2448 -765
rect 2390 -805 2448 -799
rect 2508 -765 2566 -759
rect 2508 -799 2520 -765
rect 2554 -799 2566 -765
rect 2508 -805 2566 -799
rect 2626 -765 2684 -759
rect 2626 -799 2638 -765
rect 2672 -799 2684 -765
rect 2626 -805 2684 -799
rect 2744 -765 2802 -759
rect 2744 -799 2756 -765
rect 2790 -799 2802 -765
rect 2744 -805 2802 -799
rect 2862 -765 2920 -759
rect 2862 -799 2874 -765
rect 2908 -799 2920 -765
rect 2862 -805 2920 -799
rect 2980 -765 3038 -759
rect 2980 -799 2992 -765
rect 3026 -799 3038 -765
rect 2980 -805 3038 -799
rect 3098 -765 3156 -759
rect 3098 -799 3110 -765
rect 3144 -799 3156 -765
rect 3098 -805 3156 -799
rect 3216 -765 3274 -759
rect 3216 -799 3228 -765
rect 3262 -799 3274 -765
rect 3216 -805 3274 -799
rect 3334 -765 3392 -759
rect 3334 -799 3346 -765
rect 3380 -799 3392 -765
rect 3334 -805 3392 -799
rect 3452 -765 3510 -759
rect 3452 -799 3464 -765
rect 3498 -799 3510 -765
rect 3452 -805 3510 -799
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -3654 -884 3654 884
string parameters w 3 l 0.3 m 2 nf 60 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
