magic
tech sky130A
magscale 1 2
timestamp 1605995445
<< error_s >>
rect -4389 9085 -4379 9131
rect -4361 9057 -4351 9159
rect -4073 9057 -4066 9159
rect -4045 9085 -4038 9131
rect -1626 9085 -1613 9131
rect -1598 9057 -1585 9159
rect -592 8620 -576 8678
rect 26 8666 30 8678
rect 38 8632 42 8666
rect -5119 8532 -5112 8578
rect -5091 8504 -5084 8605
rect -404 8054 -392 8100
rect -125 8074 -121 8108
<< pwell >>
rect -7384 8100 -7328 8110
rect -5312 7347 -5094 7557
<< locali >>
rect -7906 8982 -7699 9791
rect -1438 8986 -1313 9791
rect -4804 8982 -1313 8986
rect -7906 8906 -1313 8982
rect -7906 8836 -787 8906
rect -4804 8732 -787 8836
rect -7912 7919 -7726 8710
rect -4804 8536 -1313 8732
rect -4940 7919 -1313 8369
rect -7912 7674 2913 7919
rect -7912 7344 -7258 7674
rect -6941 7344 -6554 7560
rect -6169 7344 -5782 7560
rect -5397 7546 -5010 7560
rect -5397 7360 -5299 7546
rect -5107 7360 -5010 7546
rect -5397 7344 -5010 7360
rect -4625 7344 -4238 7560
rect -3853 7344 -3466 7560
rect -3081 7344 -2694 7560
rect -2309 7344 -1922 7560
rect -1537 7344 -1150 7560
rect -765 7344 -378 7560
rect 7 7344 394 7560
rect 779 7344 1166 7560
rect 1551 7344 1938 7560
rect 2709 7344 2890 7560
rect -7896 1696 -7713 1912
rect -7328 1696 -6941 1912
rect -6556 1696 -6169 1912
rect -5784 1696 -5397 1912
rect -5012 1696 -4625 1912
rect -4240 1696 -3853 1912
rect -3468 1696 -3081 1912
rect -2696 1696 -2309 1912
rect -1924 1696 -1537 1912
rect -1152 1696 -765 1912
rect -380 1696 7 1912
rect 392 1696 779 1912
rect 1164 1696 1551 1912
rect 1936 1696 2323 1912
rect 2708 1696 2888 1912
<< viali >>
rect -5299 7360 -5107 7546
rect 2254 7128 2392 7560
<< metal1 >>
rect -7034 9616 -5348 9660
rect -3564 9612 -2090 9656
rect -1167 9603 2564 9740
rect -1167 9579 -783 9603
rect -7662 9555 -7565 9557
rect -7662 9170 -7534 9555
rect -7220 9423 -5026 9559
rect -7345 9184 -5310 9319
rect -4854 9189 -4547 9335
rect -7662 8652 -7565 9170
rect -7034 9084 -5348 9128
rect -4361 8875 -4291 9566
rect -5465 8805 -4291 8875
rect -7662 8500 -7584 8652
rect -7662 8104 -7565 8500
rect -7502 7475 -7448 8564
rect -7066 8534 -5592 8578
rect -7384 8276 -7213 8503
rect -5465 8483 -5395 8805
rect -4361 8804 -4291 8805
rect -7126 8346 -5395 8483
rect -5091 8696 -5021 8704
rect -4148 8696 -4066 9575
rect -3738 9403 -1776 9564
rect -3881 9176 -2045 9336
rect -3568 9084 -2094 9128
rect -5091 8605 -4066 8696
rect -7384 8110 -5287 8276
rect -7384 8100 -7213 8110
rect -5091 8104 -5005 8605
rect -1598 8249 -1516 9575
rect -7342 7864 -7213 8100
rect -7066 8020 -5592 8064
rect -1167 7664 -943 9579
rect -789 8765 2570 9020
rect -789 8632 2734 8765
rect 2569 8624 2734 8632
rect -794 7916 2562 8053
rect 2274 7801 2368 7805
rect 2640 7801 2734 8624
rect 2274 7707 2734 7801
rect 2274 7576 2368 7707
rect 2240 7560 2406 7576
rect -5312 7546 -5094 7557
rect -5312 7475 -5299 7546
rect -7502 7421 -5299 7475
rect -5312 7360 -5299 7421
rect -5107 7360 -5094 7546
rect -5312 7347 -5094 7360
rect 2240 7128 2254 7560
rect 2392 7128 2406 7560
rect 2240 7113 2406 7128
<< metal2 >>
rect 2824 8538 2880 9338
rect 3028 8538 3084 9338
rect 3232 8538 3288 9338
rect 2838 8440 2866 8538
rect 3042 8440 3070 8538
rect 3246 8440 3274 8538
rect 15 581 71 1381
rect 219 581 275 1381
<< metal3 >>
rect 3560 3862 4360 3982
use sky130_fd_pr__pfet_g5v0d10v5_6UDFJU  sky130_fd_pr__pfet_g5v0d10v5_6UDFJU_0
timestamp 1605994897
transform 1 0 -6190 0 1 9372
box -1101 -497 1101 497
use sky130_fd_pr__pfet_g5v0d10v5_6E4TNU  sky130_fd_pr__pfet_g5v0d10v5_6E4TNU_0
timestamp 1605994897
transform 1 0 -7439 0 1 9372
box -338 -497 338 497
use sky130_fd_pr__nfet_g5v0d10v5_CWNXJM  sky130_fd_pr__nfet_g5v0d10v5_CWNXJM_0
timestamp 1605994897
transform 1 0 -6332 0 1 8300
box -962 -458 962 458
use sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC  sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC_1
timestamp 1605994897
transform -1 0 -7476 0 1 8300
box -308 -458 308 458
use sky130_fd_pr__pfet_g5v0d10v5_ZPXEXA  sky130_fd_pr__pfet_g5v0d10v5_ZPXEXA_0
timestamp 1605995445
transform 1 0 -2829 0 1 9372
box -992 -497 992 497
use sky130_fd_pr__pfet_g5v0d10v5_Z95PRA  sky130_fd_pr__pfet_g5v0d10v5_Z95PRA_0
timestamp 1605995445
transform 1 0 -4941 0 1 9372
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_6E4TNU  sky130_fd_pr__pfet_g5v0d10v5_6E4TNU_2
timestamp 1605994897
transform 1 0 -4455 0 1 9372
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_6E4TNU  sky130_fd_pr__pfet_g5v0d10v5_6E4TNU_3
timestamp 1605994897
transform 1 0 -3969 0 1 9372
box -338 -497 338 497
use sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC  sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC_0
timestamp 1605994897
transform 1 0 -5188 0 1 8300
box -308 -458 308 458
use sky130_fd_pr__pfet_g5v0d10v5_6E4TNU  sky130_fd_pr__pfet_g5v0d10v5_6E4TNU_4
timestamp 1605994897
transform 1 0 -1689 0 1 9372
box -338 -497 338 497
use sky130_fd_sc_hvl__schmittbuf_1  sky130_fd_sc_hvl__schmittbuf_1_0 ~/projects/efabless/tech/SW/sky130A/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1605995445
transform 1 0 -790 0 1 7935
box -66 -23 1122 897
use sky130_fd_sc_hvl__buf_8  sky130_fd_sc_hvl__buf_8_0 ~/projects/efabless/tech/SW/sky130A/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1605995445
transform 1 0 266 0 1 7935
box -66 -23 1986 897
use sky130_fd_sc_hvl__buf_8  sky130_fd_sc_hvl__buf_8_1
timestamp 1605995445
transform 1 0 -790 0 -1 9703
box -66 -23 1986 897
use sky130_fd_sc_hvl__fill_4  sky130_fd_sc_hvl__fill_4_0 ~/projects/efabless/tech/SW/sky130A/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1605995445
transform 1 0 2186 0 1 7935
box -66 -23 450 897
use sky130_fd_sc_hvl__inv_8  sky130_fd_sc_hvl__inv_8_0 ~/projects/efabless/tech/SW/sky130A/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1605995445
transform 1 0 1130 0 -1 9703
box -66 -23 1506 897
use sky130_fd_pr__res_xhigh_po_0p69_LV2JUS  sky130_fd_pr__res_xhigh_po_0p69_LV2JUS_0
timestamp 1605923309
transform 1 0 -2502 0 1 4628
box -5446 -3098 5446 3098
use sky130_fd_pr__cap_mim_m3_2_N249RX  sky130_fd_pr__cap_mim_m3_2_N249RX_0
timestamp 1605923309
transform 1 0 -77 0 1 4682
box -3379 -3101 3401 3101
use sky130_fd_pr__cap_mim_m3_1_N249RX  sky130_fd_pr__cap_mim_m3_1_N249RX_0
timestamp 1605923309
transform -1 0 -450 0 1 4682
box -3186 -3100 3186 3100
<< labels >>
rlabel metal3 s 3560 3862 4360 3982 6 vss
port 2 nsew default input
rlabel metal2 s 2824 8538 2880 9338 6 porb_h
port 0 nsew default tristate
rlabel metal2 s 3028 8538 3084 9338 6 porb_l
port 0 nsew default tristate
rlabel metal2 s 3232 8538 3288 9338 6 por_l
port 0 nsew default tristate
rlabel metal2 s 15 581 71 1381 6 vdd3v3
port 1 nsew default input
rlabel metal2 s 219 581 275 1381 6 vdd1v8
port 1 nsew default input
<< properties >>
string FIXED_BBOX 0 0 4360 9164
<< end >>
