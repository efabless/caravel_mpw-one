magic
tech sky130A
timestamp 1606369131
<< checkpaint >>
rect -630 -630 300088 359022
<< metal2 >>
rect 7805 354972 7833 355212
rect 15901 354972 15929 355212
rect 23997 354972 24025 355212
rect 32139 354972 32167 355212
rect 40235 354972 40263 355212
rect 48331 354972 48359 355212
rect 56473 354972 56501 355212
rect 64569 354972 64597 355212
rect 72665 354972 72693 355212
rect 80807 354972 80835 355212
rect 88903 354972 88931 355212
rect 96999 354972 97027 355212
rect 105141 354972 105169 355212
rect 113237 354972 113265 355212
rect 121333 354972 121361 355212
rect 129475 354972 129503 355212
rect 137571 354972 137599 355212
rect 145667 354972 145695 355212
rect 153809 354972 153837 355212
rect 161905 354972 161933 355212
rect 170001 354972 170029 355212
rect 178143 354972 178171 355212
rect 186239 354972 186267 355212
rect 194335 354972 194363 355212
rect 202477 354972 202505 355212
rect 210573 354972 210601 355212
rect 218669 354972 218697 355212
rect 226811 354972 226839 355212
rect 234907 354972 234935 355212
rect 243003 354972 243031 355212
rect 251145 354972 251173 355212
rect 259241 354972 259269 355212
rect 267337 354972 267365 355212
rect 275479 354972 275507 355212
rect 283575 354972 283603 355212
rect 291671 354972 291699 355212
rect 4033 3212 4061 3452
rect 4585 3212 4613 3452
rect 5183 3212 5211 3452
rect 5781 3212 5809 3452
rect 6379 3212 6407 3452
rect 6977 3212 7005 3452
rect 7575 3212 7603 3452
rect 8173 3212 8201 3452
rect 8771 3212 8799 3452
rect 9369 3212 9397 3452
rect 9967 3212 9995 3452
rect 10565 3212 10593 3452
rect 11163 3212 11191 3452
rect 11761 3212 11789 3452
rect 12359 3212 12387 3452
rect 12911 3212 12939 3452
rect 13509 3212 13537 3452
rect 14107 3212 14135 3452
rect 14705 3212 14733 3452
rect 15303 3212 15331 3452
rect 15901 3212 15929 3452
rect 16499 3212 16527 3452
rect 17097 3212 17125 3452
rect 17695 3212 17723 3452
rect 18293 3212 18321 3452
rect 18891 3212 18919 3452
rect 19489 3212 19517 3452
rect 20087 3212 20115 3452
rect 20685 3212 20713 3452
rect 21237 3212 21265 3452
rect 21835 3212 21863 3452
rect 22433 3212 22461 3452
rect 23031 3212 23059 3452
rect 23629 3212 23657 3452
rect 24227 3212 24255 3452
rect 24825 3212 24853 3452
rect 25423 3212 25451 3452
rect 26021 3212 26049 3452
rect 26619 3212 26647 3452
rect 27217 3212 27245 3452
rect 27815 3212 27843 3452
rect 28413 3212 28441 3452
rect 29011 3212 29039 3452
rect 29563 3212 29591 3452
rect 30161 3212 30189 3452
rect 30759 3212 30787 3452
rect 31357 3212 31385 3452
rect 31955 3212 31983 3452
rect 32553 3212 32581 3452
rect 33151 3212 33179 3452
rect 33749 3212 33777 3452
rect 34347 3212 34375 3452
rect 34945 3212 34973 3452
rect 35543 3212 35571 3452
rect 36141 3212 36169 3452
rect 36739 3212 36767 3452
rect 37337 3212 37365 3452
rect 37889 3212 37917 3452
rect 38487 3212 38515 3452
rect 39085 3212 39113 3452
rect 39683 3212 39711 3452
rect 40281 3212 40309 3452
rect 40879 3212 40907 3452
rect 41477 3212 41505 3452
rect 42075 3212 42103 3452
rect 42673 3212 42701 3452
rect 43271 3212 43299 3452
rect 43869 3212 43897 3452
rect 44467 3212 44495 3452
rect 45065 3212 45093 3452
rect 45663 3212 45691 3452
rect 46215 3212 46243 3452
rect 46813 3212 46841 3452
rect 47411 3212 47439 3452
rect 48009 3212 48037 3452
rect 48607 3212 48635 3452
rect 49205 3212 49233 3452
rect 49803 3212 49831 3452
rect 50401 3212 50429 3452
rect 50999 3212 51027 3452
rect 51597 3212 51625 3452
rect 52195 3212 52223 3452
rect 52793 3212 52821 3452
rect 53391 3212 53419 3452
rect 53989 3212 54017 3452
rect 54541 3212 54569 3452
rect 55139 3212 55167 3452
rect 55737 3212 55765 3452
rect 56335 3212 56363 3452
rect 56933 3212 56961 3452
rect 57531 3212 57559 3452
rect 58129 3212 58157 3452
rect 58727 3212 58755 3452
rect 59325 3212 59353 3452
rect 59923 3212 59951 3452
rect 60521 3212 60549 3452
rect 61119 3212 61147 3452
rect 61717 3212 61745 3452
rect 62315 3212 62343 3452
rect 62867 3212 62895 3452
rect 63465 3212 63493 3452
rect 64063 3212 64091 3452
rect 64661 3212 64689 3452
rect 65259 3212 65287 3452
rect 65857 3212 65885 3452
rect 66455 3212 66483 3452
rect 67053 3212 67081 3452
rect 67651 3212 67679 3452
rect 68249 3212 68277 3452
rect 68847 3212 68875 3452
rect 69445 3212 69473 3452
rect 70043 3212 70071 3452
rect 70641 3212 70669 3452
rect 71193 3212 71221 3452
rect 71791 3212 71819 3452
rect 72389 3212 72417 3452
rect 72987 3212 73015 3452
rect 73585 3212 73613 3452
rect 74183 3212 74211 3452
rect 74781 3212 74809 3452
rect 75379 3212 75407 3452
rect 75977 3212 76005 3452
rect 76575 3212 76603 3452
rect 77173 3212 77201 3452
rect 77771 3212 77799 3452
rect 78369 3212 78397 3452
rect 78967 3212 78995 3452
rect 79519 3212 79547 3452
rect 80117 3212 80145 3452
rect 80715 3212 80743 3452
rect 81313 3212 81341 3452
rect 81911 3212 81939 3452
rect 82509 3212 82537 3452
rect 83107 3212 83135 3452
rect 83705 3212 83733 3452
rect 84303 3212 84331 3452
rect 84901 3212 84929 3452
rect 85499 3212 85527 3452
rect 86097 3212 86125 3452
rect 86695 3212 86723 3452
rect 87293 3212 87321 3452
rect 87845 3212 87873 3452
rect 88443 3212 88471 3452
rect 89041 3212 89069 3452
rect 89639 3212 89667 3452
rect 90237 3212 90265 3452
rect 90835 3212 90863 3452
rect 91433 3212 91461 3452
rect 92031 3212 92059 3452
rect 92629 3212 92657 3452
rect 93227 3212 93255 3452
rect 93825 3212 93853 3452
rect 94423 3212 94451 3452
rect 95021 3212 95049 3452
rect 95619 3212 95647 3452
rect 96171 3212 96199 3452
rect 96769 3212 96797 3452
rect 97367 3212 97395 3452
rect 97965 3212 97993 3452
rect 98563 3212 98591 3452
rect 99161 3212 99189 3452
rect 99759 3212 99787 3452
rect 100357 3212 100385 3452
rect 100955 3212 100983 3452
rect 101553 3212 101581 3452
rect 102151 3212 102179 3452
rect 102749 3212 102777 3452
rect 103347 3212 103375 3452
rect 103945 3212 103973 3452
rect 104497 3212 104525 3452
rect 105095 3212 105123 3452
rect 105693 3212 105721 3452
rect 106291 3212 106319 3452
rect 106889 3212 106917 3452
rect 107487 3212 107515 3452
rect 108085 3212 108113 3452
rect 108683 3212 108711 3452
rect 109281 3212 109309 3452
rect 109879 3212 109907 3452
rect 110477 3212 110505 3452
rect 111075 3212 111103 3452
rect 111673 3212 111701 3452
rect 112271 3212 112299 3452
rect 112823 3212 112851 3452
rect 113421 3212 113449 3452
rect 114019 3212 114047 3452
rect 114617 3212 114645 3452
rect 115215 3212 115243 3452
rect 115813 3212 115841 3452
rect 116411 3212 116439 3452
rect 117009 3212 117037 3452
rect 117607 3212 117635 3452
rect 118205 3212 118233 3452
rect 118803 3212 118831 3452
rect 119401 3212 119429 3452
rect 119999 3212 120027 3452
rect 120597 3212 120625 3452
rect 121149 3212 121177 3452
rect 121747 3212 121775 3452
rect 122345 3212 122373 3452
rect 122943 3212 122971 3452
rect 123541 3212 123569 3452
rect 124139 3212 124167 3452
rect 124737 3212 124765 3452
rect 125335 3212 125363 3452
rect 125933 3212 125961 3452
rect 126531 3212 126559 3452
rect 127129 3212 127157 3452
rect 127727 3212 127755 3452
rect 128325 3212 128353 3452
rect 128923 3212 128951 3452
rect 129475 3212 129503 3452
rect 130073 3212 130101 3452
rect 130671 3212 130699 3452
rect 131269 3212 131297 3452
rect 131867 3212 131895 3452
rect 132465 3212 132493 3452
rect 133063 3212 133091 3452
rect 133661 3212 133689 3452
rect 134259 3212 134287 3452
rect 134857 3212 134885 3452
rect 135455 3212 135483 3452
rect 136053 3212 136081 3452
rect 136651 3212 136679 3452
rect 137249 3212 137277 3452
rect 137801 3212 137829 3452
rect 138399 3212 138427 3452
rect 138997 3212 139025 3452
rect 139595 3212 139623 3452
rect 140193 3212 140221 3452
rect 140791 3212 140819 3452
rect 141389 3212 141417 3452
rect 141987 3212 142015 3452
rect 142585 3212 142613 3452
rect 143183 3212 143211 3452
rect 143781 3212 143809 3452
rect 144379 3212 144407 3452
rect 144977 3212 145005 3452
rect 145575 3212 145603 3452
rect 146127 3212 146155 3452
rect 146725 3212 146753 3452
rect 147323 3212 147351 3452
rect 147921 3212 147949 3452
rect 148519 3212 148547 3452
rect 149117 3212 149145 3452
rect 149715 3212 149743 3452
rect 150313 3212 150341 3452
rect 150911 3212 150939 3452
rect 151509 3212 151537 3452
rect 152107 3212 152135 3452
rect 152705 3212 152733 3452
rect 153303 3212 153331 3452
rect 153901 3212 153929 3452
rect 154453 3212 154481 3452
rect 155051 3212 155079 3452
rect 155649 3212 155677 3452
rect 156247 3212 156275 3452
rect 156845 3212 156873 3452
rect 157443 3212 157471 3452
rect 158041 3212 158069 3452
rect 158639 3212 158667 3452
rect 159237 3212 159265 3452
rect 159835 3212 159863 3452
rect 160433 3212 160461 3452
rect 161031 3212 161059 3452
rect 161629 3212 161657 3452
rect 162227 3212 162255 3452
rect 162779 3212 162807 3452
rect 163377 3212 163405 3452
rect 163975 3212 164003 3452
rect 164573 3212 164601 3452
rect 165171 3212 165199 3452
rect 165769 3212 165797 3452
rect 166367 3212 166395 3452
rect 166965 3212 166993 3452
rect 167563 3212 167591 3452
rect 168161 3212 168189 3452
rect 168759 3212 168787 3452
rect 169357 3212 169385 3452
rect 169955 3212 169983 3452
rect 170553 3212 170581 3452
rect 171105 3212 171133 3452
rect 171703 3212 171731 3452
rect 172301 3212 172329 3452
rect 172899 3212 172927 3452
rect 173497 3212 173525 3452
rect 174095 3212 174123 3452
rect 174693 3212 174721 3452
rect 175291 3212 175319 3452
rect 175889 3212 175917 3452
rect 176487 3212 176515 3452
rect 177085 3212 177113 3452
rect 177683 3212 177711 3452
rect 178281 3212 178309 3452
rect 178879 3212 178907 3452
rect 179431 3212 179459 3452
rect 180029 3212 180057 3452
rect 180627 3212 180655 3452
rect 181225 3212 181253 3452
rect 181823 3212 181851 3452
rect 182421 3212 182449 3452
rect 183019 3212 183047 3452
rect 183617 3212 183645 3452
rect 184215 3212 184243 3452
rect 184813 3212 184841 3452
rect 185411 3212 185439 3452
rect 186009 3212 186037 3452
rect 186607 3212 186635 3452
rect 187205 3212 187233 3452
rect 187757 3212 187785 3452
rect 188355 3212 188383 3452
rect 188953 3212 188981 3452
rect 189551 3212 189579 3452
rect 190149 3212 190177 3452
rect 190747 3212 190775 3452
rect 191345 3212 191373 3452
rect 191943 3212 191971 3452
rect 192541 3212 192569 3452
rect 193139 3212 193167 3452
rect 193737 3212 193765 3452
rect 194335 3212 194363 3452
rect 194933 3212 194961 3452
rect 195531 3212 195559 3452
rect 196083 3212 196111 3452
rect 196681 3212 196709 3452
rect 197279 3212 197307 3452
rect 197877 3212 197905 3452
rect 198475 3212 198503 3452
rect 199073 3212 199101 3452
rect 199671 3212 199699 3452
rect 200269 3212 200297 3452
rect 200867 3212 200895 3452
rect 201465 3212 201493 3452
rect 202063 3212 202091 3452
rect 202661 3212 202689 3452
rect 203259 3212 203287 3452
rect 203857 3212 203885 3452
rect 204409 3212 204437 3452
rect 205007 3212 205035 3452
rect 205605 3212 205633 3452
rect 206203 3212 206231 3452
rect 206801 3212 206829 3452
rect 207399 3212 207427 3452
rect 207997 3212 208025 3452
rect 208595 3212 208623 3452
rect 209193 3212 209221 3452
rect 209791 3212 209819 3452
rect 210389 3212 210417 3452
rect 210987 3212 211015 3452
rect 211585 3212 211613 3452
rect 212183 3212 212211 3452
rect 212735 3212 212763 3452
rect 213333 3212 213361 3452
rect 213931 3212 213959 3452
rect 214529 3212 214557 3452
rect 215127 3212 215155 3452
rect 215725 3212 215753 3452
rect 216323 3212 216351 3452
rect 216921 3212 216949 3452
rect 217519 3212 217547 3452
rect 218117 3212 218145 3452
rect 218715 3212 218743 3452
rect 219313 3212 219341 3452
rect 219911 3212 219939 3452
rect 220509 3212 220537 3452
rect 221061 3212 221089 3452
rect 221659 3212 221687 3452
rect 222257 3212 222285 3452
rect 222855 3212 222883 3452
rect 223453 3212 223481 3452
rect 224051 3212 224079 3452
rect 224649 3212 224677 3452
rect 225247 3212 225275 3452
rect 225845 3212 225873 3452
rect 226443 3212 226471 3452
rect 227041 3212 227069 3452
rect 227639 3212 227667 3452
rect 228237 3212 228265 3452
rect 228835 3212 228863 3452
rect 229387 3212 229415 3452
rect 229985 3212 230013 3452
rect 230583 3212 230611 3452
rect 231181 3212 231209 3452
rect 231779 3212 231807 3452
rect 232377 3212 232405 3452
rect 232975 3212 233003 3452
rect 233573 3212 233601 3452
rect 234171 3212 234199 3452
rect 234769 3212 234797 3452
rect 235367 3212 235395 3452
rect 235965 3212 235993 3452
rect 236563 3212 236591 3452
rect 237161 3212 237189 3452
rect 237713 3212 237741 3452
rect 238311 3212 238339 3452
rect 238909 3212 238937 3452
rect 239507 3212 239535 3452
rect 240105 3212 240133 3452
rect 240703 3212 240731 3452
rect 241301 3212 241329 3452
rect 241899 3212 241927 3452
rect 242497 3212 242525 3452
rect 243095 3212 243123 3452
rect 243693 3212 243721 3452
rect 244291 3212 244319 3452
rect 244889 3212 244917 3452
rect 245487 3212 245515 3452
rect 246039 3212 246067 3452
rect 246637 3212 246665 3452
rect 247235 3212 247263 3452
rect 247833 3212 247861 3452
rect 248431 3212 248459 3452
rect 249029 3212 249057 3452
rect 249627 3212 249655 3452
rect 250225 3212 250253 3452
rect 250823 3212 250851 3452
rect 251421 3212 251449 3452
rect 252019 3212 252047 3452
rect 252617 3212 252645 3452
rect 253215 3212 253243 3452
rect 253813 3212 253841 3452
rect 254365 3212 254393 3452
rect 254963 3212 254991 3452
rect 255561 3212 255589 3452
rect 256159 3212 256187 3452
rect 256757 3212 256785 3452
rect 257355 3212 257383 3452
rect 257953 3212 257981 3452
rect 258551 3212 258579 3452
rect 259149 3212 259177 3452
rect 259747 3212 259775 3452
rect 260345 3212 260373 3452
rect 260943 3212 260971 3452
rect 261541 3212 261569 3452
rect 262139 3212 262167 3452
rect 262691 3212 262719 3452
rect 263289 3212 263317 3452
rect 263887 3212 263915 3452
rect 264485 3212 264513 3452
rect 265083 3212 265111 3452
rect 265681 3212 265709 3452
rect 266279 3212 266307 3452
rect 266877 3212 266905 3452
rect 267475 3212 267503 3452
rect 268073 3212 268101 3452
rect 268671 3212 268699 3452
rect 269269 3212 269297 3452
rect 269867 3212 269895 3452
rect 270465 3212 270493 3452
rect 271017 3212 271045 3452
rect 271615 3212 271643 3452
rect 272213 3212 272241 3452
rect 272811 3212 272839 3452
rect 273409 3212 273437 3452
rect 274007 3212 274035 3452
rect 274605 3212 274633 3452
rect 275203 3212 275231 3452
rect 275801 3212 275829 3452
rect 276399 3212 276427 3452
rect 276997 3212 277025 3452
rect 277595 3212 277623 3452
rect 278193 3212 278221 3452
rect 278791 3212 278819 3452
rect 279343 3212 279371 3452
rect 279941 3212 279969 3452
rect 280539 3212 280567 3452
rect 281137 3212 281165 3452
rect 281735 3212 281763 3452
rect 282333 3212 282361 3452
rect 282931 3212 282959 3452
rect 283529 3212 283557 3452
rect 284127 3212 284155 3452
rect 284725 3212 284753 3452
rect 285323 3212 285351 3452
rect 285921 3212 285949 3452
rect 286519 3212 286547 3452
rect 287117 3212 287145 3452
rect 287669 3212 287697 3452
rect 288267 3212 288295 3452
rect 288865 3212 288893 3452
rect 289463 3212 289491 3452
rect 290061 3212 290089 3452
rect 290659 3212 290687 3452
rect 291257 3212 291285 3452
rect 291855 3212 291883 3452
rect 292453 3212 292481 3452
rect 293051 3212 293079 3452
rect 293649 3212 293677 3452
rect 294247 3212 294275 3452
rect 294845 3212 294873 3452
rect 295443 3212 295471 3452
<< metal3 >>
rect 295508 352192 295748 352252
rect 3748 351512 3988 351572
rect 295508 346344 295748 346404
rect 3748 344304 3988 344364
rect 295508 340496 295748 340556
rect 3748 337164 3988 337224
rect 295508 334580 295748 334640
rect 3748 329956 3988 330016
rect 295508 328732 295748 328792
rect 295508 322884 295748 322944
rect 3748 322748 3988 322808
rect 295508 317036 295748 317096
rect 3748 315608 3988 315668
rect 295508 311120 295748 311180
rect 3748 308400 3988 308460
rect 295508 305272 295748 305332
rect 3748 301192 3988 301252
rect 295508 299424 295748 299484
rect 3748 294052 3988 294112
rect 295508 293576 295748 293636
rect 295508 287660 295748 287720
rect 3748 286844 3988 286904
rect 295508 281812 295748 281872
rect 3748 279704 3988 279764
rect 295508 275964 295748 276024
rect 3748 272496 3988 272556
rect 295508 270116 295748 270176
rect 3748 265288 3988 265348
rect 295508 264200 295748 264260
rect 295508 258352 295748 258412
rect 3748 258148 3988 258208
rect 295508 252504 295748 252564
rect 3748 250940 3988 251000
rect 295508 246588 295748 246648
rect 3748 243732 3988 243792
rect 295508 240740 295748 240800
rect 3748 236592 3988 236652
rect 295508 234892 295748 234952
rect 3748 229384 3988 229444
rect 295508 229044 295748 229104
rect 295508 223128 295748 223188
rect 3748 222176 3988 222236
rect 295508 217280 295748 217340
rect 3748 215036 3988 215096
rect 295508 211432 295748 211492
rect 3748 207828 3988 207888
rect 295508 205584 295748 205644
rect 3748 200688 3988 200748
rect 295508 199668 295748 199728
rect 295508 193820 295748 193880
rect 3748 193480 3988 193540
rect 295508 187972 295748 188032
rect 3748 186272 3988 186332
rect 295508 182124 295748 182184
rect 3748 179132 3988 179192
rect 295508 176208 295748 176268
rect 3748 171924 3988 171984
rect 295508 170360 295748 170420
rect 3748 164716 3988 164776
rect 295508 164512 295748 164572
rect 295508 158596 295748 158656
rect 3748 157576 3988 157636
rect 295508 152748 295748 152808
rect 3748 150368 3988 150428
rect 295508 146900 295748 146960
rect 3748 143228 3988 143288
rect 295508 141052 295748 141112
rect 3748 136020 3988 136080
rect 295508 135136 295748 135196
rect 295508 129288 295748 129348
rect 3748 128812 3988 128872
rect 295508 123440 295748 123500
rect 3748 121672 3988 121732
rect 295508 117592 295748 117652
rect 3748 114464 3988 114524
rect 295508 111676 295748 111736
rect 3748 107256 3988 107316
rect 295508 105828 295748 105888
rect 3748 100116 3988 100176
rect 295508 99980 295748 100040
rect 295508 94132 295748 94192
rect 3748 92908 3988 92968
rect 295508 88216 295748 88276
rect 3748 85700 3988 85760
rect 295508 82368 295748 82428
rect 3748 78560 3988 78620
rect 295508 76520 295748 76580
rect 3748 71352 3988 71412
rect 295508 70604 295748 70664
rect 295508 64756 295748 64816
rect 3748 64212 3988 64272
rect 295508 58908 295748 58968
rect 3748 57004 3988 57064
rect 295508 53060 295748 53120
rect 3748 49796 3988 49856
rect 295508 47144 295748 47204
rect 3748 42656 3988 42716
rect 295508 41296 295748 41356
rect 3748 35448 3988 35508
rect 295508 35448 295748 35508
rect 295508 29600 295748 29660
rect 3748 28240 3988 28300
rect 295508 23684 295748 23744
rect 3748 21100 3988 21160
rect 295508 17836 295748 17896
rect 3748 13892 3988 13952
rect 295508 11988 295748 12048
rect 3748 6752 3988 6812
rect 295508 6140 295748 6200
<< metal4 >>
rect 0 358351 200 358392
rect 0 358233 41 358351
rect 159 358233 200 358351
rect 0 352239 200 358233
rect 0 352121 41 352239
rect 159 352121 200 352239
rect 0 342239 200 352121
rect 0 342121 41 342239
rect 159 342121 200 342239
rect 0 332239 200 342121
rect 0 332121 41 332239
rect 159 332121 200 332239
rect 0 322239 200 332121
rect 0 322121 41 322239
rect 159 322121 200 322239
rect 0 312239 200 322121
rect 0 312121 41 312239
rect 159 312121 200 312239
rect 0 302239 200 312121
rect 0 302121 41 302239
rect 159 302121 200 302239
rect 0 292239 200 302121
rect 0 292121 41 292239
rect 159 292121 200 292239
rect 0 282239 200 292121
rect 0 282121 41 282239
rect 159 282121 200 282239
rect 0 272239 200 282121
rect 0 272121 41 272239
rect 159 272121 200 272239
rect 0 262239 200 272121
rect 0 262121 41 262239
rect 159 262121 200 262239
rect 0 252239 200 262121
rect 0 252121 41 252239
rect 159 252121 200 252239
rect 0 242239 200 252121
rect 0 242121 41 242239
rect 159 242121 200 242239
rect 0 232239 200 242121
rect 0 232121 41 232239
rect 159 232121 200 232239
rect 0 222239 200 232121
rect 0 222121 41 222239
rect 159 222121 200 222239
rect 0 212239 200 222121
rect 0 212121 41 212239
rect 159 212121 200 212239
rect 0 202239 200 212121
rect 0 202121 41 202239
rect 159 202121 200 202239
rect 0 192239 200 202121
rect 0 192121 41 192239
rect 159 192121 200 192239
rect 0 182239 200 192121
rect 0 182121 41 182239
rect 159 182121 200 182239
rect 0 172239 200 182121
rect 0 172121 41 172239
rect 159 172121 200 172239
rect 0 162239 200 172121
rect 0 162121 41 162239
rect 159 162121 200 162239
rect 0 152239 200 162121
rect 0 152121 41 152239
rect 159 152121 200 152239
rect 0 142239 200 152121
rect 0 142121 41 142239
rect 159 142121 200 142239
rect 0 132239 200 142121
rect 0 132121 41 132239
rect 159 132121 200 132239
rect 0 122239 200 132121
rect 0 122121 41 122239
rect 159 122121 200 122239
rect 0 112239 200 122121
rect 0 112121 41 112239
rect 159 112121 200 112239
rect 0 102239 200 112121
rect 0 102121 41 102239
rect 159 102121 200 102239
rect 0 92239 200 102121
rect 0 92121 41 92239
rect 159 92121 200 92239
rect 0 82239 200 92121
rect 0 82121 41 82239
rect 159 82121 200 82239
rect 0 72239 200 82121
rect 0 72121 41 72239
rect 159 72121 200 72239
rect 0 62239 200 72121
rect 0 62121 41 62239
rect 159 62121 200 62239
rect 0 52239 200 62121
rect 0 52121 41 52239
rect 159 52121 200 52239
rect 0 42239 200 52121
rect 0 42121 41 42239
rect 159 42121 200 42239
rect 0 32239 200 42121
rect 0 32121 41 32239
rect 159 32121 200 32239
rect 0 22239 200 32121
rect 0 22121 41 22239
rect 159 22121 200 22239
rect 0 12239 200 22121
rect 0 12121 41 12239
rect 159 12121 200 12239
rect 0 159 200 12121
rect 400 357951 600 357992
rect 400 357833 441 357951
rect 559 357833 600 357951
rect 400 347239 600 357833
rect 7080 357951 7280 358392
rect 7080 357833 7121 357951
rect 7239 357833 7280 357951
rect 400 347121 441 347239
rect 559 347121 600 347239
rect 400 337239 600 347121
rect 400 337121 441 337239
rect 559 337121 600 337239
rect 400 327239 600 337121
rect 400 327121 441 327239
rect 559 327121 600 327239
rect 400 317239 600 327121
rect 400 317121 441 317239
rect 559 317121 600 317239
rect 400 307239 600 317121
rect 400 307121 441 307239
rect 559 307121 600 307239
rect 400 297239 600 307121
rect 400 297121 441 297239
rect 559 297121 600 297239
rect 400 287239 600 297121
rect 400 287121 441 287239
rect 559 287121 600 287239
rect 400 277239 600 287121
rect 400 277121 441 277239
rect 559 277121 600 277239
rect 400 267239 600 277121
rect 400 267121 441 267239
rect 559 267121 600 267239
rect 400 257239 600 267121
rect 400 257121 441 257239
rect 559 257121 600 257239
rect 400 247239 600 257121
rect 400 247121 441 247239
rect 559 247121 600 247239
rect 400 237239 600 247121
rect 400 237121 441 237239
rect 559 237121 600 237239
rect 400 227239 600 237121
rect 400 227121 441 227239
rect 559 227121 600 227239
rect 400 217239 600 227121
rect 400 217121 441 217239
rect 559 217121 600 217239
rect 400 207239 600 217121
rect 400 207121 441 207239
rect 559 207121 600 207239
rect 400 197239 600 207121
rect 400 197121 441 197239
rect 559 197121 600 197239
rect 400 187239 600 197121
rect 400 187121 441 187239
rect 559 187121 600 187239
rect 400 177239 600 187121
rect 400 177121 441 177239
rect 559 177121 600 177239
rect 400 167239 600 177121
rect 400 167121 441 167239
rect 559 167121 600 167239
rect 400 157239 600 167121
rect 400 157121 441 157239
rect 559 157121 600 157239
rect 400 147239 600 157121
rect 400 147121 441 147239
rect 559 147121 600 147239
rect 400 137239 600 147121
rect 400 137121 441 137239
rect 559 137121 600 137239
rect 400 127239 600 137121
rect 400 127121 441 127239
rect 559 127121 600 127239
rect 400 117239 600 127121
rect 400 117121 441 117239
rect 559 117121 600 117239
rect 400 107239 600 117121
rect 400 107121 441 107239
rect 559 107121 600 107239
rect 400 97239 600 107121
rect 400 97121 441 97239
rect 559 97121 600 97239
rect 400 87239 600 97121
rect 400 87121 441 87239
rect 559 87121 600 87239
rect 400 77239 600 87121
rect 400 77121 441 77239
rect 559 77121 600 77239
rect 400 67239 600 77121
rect 400 67121 441 67239
rect 559 67121 600 67239
rect 400 57239 600 67121
rect 400 57121 441 57239
rect 559 57121 600 57239
rect 400 47239 600 57121
rect 400 47121 441 47239
rect 559 47121 600 47239
rect 400 37239 600 47121
rect 400 37121 441 37239
rect 559 37121 600 37239
rect 400 27239 600 37121
rect 400 27121 441 27239
rect 559 27121 600 27239
rect 400 17239 600 27121
rect 400 17121 441 17239
rect 559 17121 600 17239
rect 400 7239 600 17121
rect 400 7121 441 7239
rect 559 7121 600 7239
rect 400 559 600 7121
rect 800 357551 1000 357592
rect 800 357433 841 357551
rect 959 357433 1000 357551
rect 800 351279 1000 357433
rect 800 351161 841 351279
rect 959 351161 1000 351279
rect 800 341279 1000 351161
rect 800 341161 841 341279
rect 959 341161 1000 341279
rect 800 331279 1000 341161
rect 800 331161 841 331279
rect 959 331161 1000 331279
rect 800 321279 1000 331161
rect 800 321161 841 321279
rect 959 321161 1000 321279
rect 800 311279 1000 321161
rect 800 311161 841 311279
rect 959 311161 1000 311279
rect 800 301279 1000 311161
rect 800 301161 841 301279
rect 959 301161 1000 301279
rect 800 291279 1000 301161
rect 800 291161 841 291279
rect 959 291161 1000 291279
rect 800 281279 1000 291161
rect 800 281161 841 281279
rect 959 281161 1000 281279
rect 800 271279 1000 281161
rect 800 271161 841 271279
rect 959 271161 1000 271279
rect 800 261279 1000 271161
rect 800 261161 841 261279
rect 959 261161 1000 261279
rect 800 251279 1000 261161
rect 800 251161 841 251279
rect 959 251161 1000 251279
rect 800 241279 1000 251161
rect 800 241161 841 241279
rect 959 241161 1000 241279
rect 800 231279 1000 241161
rect 800 231161 841 231279
rect 959 231161 1000 231279
rect 800 221279 1000 231161
rect 800 221161 841 221279
rect 959 221161 1000 221279
rect 800 211279 1000 221161
rect 800 211161 841 211279
rect 959 211161 1000 211279
rect 800 201279 1000 211161
rect 800 201161 841 201279
rect 959 201161 1000 201279
rect 800 191279 1000 201161
rect 800 191161 841 191279
rect 959 191161 1000 191279
rect 800 181279 1000 191161
rect 800 181161 841 181279
rect 959 181161 1000 181279
rect 800 171279 1000 181161
rect 800 171161 841 171279
rect 959 171161 1000 171279
rect 800 161279 1000 171161
rect 800 161161 841 161279
rect 959 161161 1000 161279
rect 800 151279 1000 161161
rect 800 151161 841 151279
rect 959 151161 1000 151279
rect 800 141279 1000 151161
rect 800 141161 841 141279
rect 959 141161 1000 141279
rect 800 131279 1000 141161
rect 800 131161 841 131279
rect 959 131161 1000 131279
rect 800 121279 1000 131161
rect 800 121161 841 121279
rect 959 121161 1000 121279
rect 800 111279 1000 121161
rect 800 111161 841 111279
rect 959 111161 1000 111279
rect 800 101279 1000 111161
rect 800 101161 841 101279
rect 959 101161 1000 101279
rect 800 91279 1000 101161
rect 800 91161 841 91279
rect 959 91161 1000 91279
rect 800 81279 1000 91161
rect 800 81161 841 81279
rect 959 81161 1000 81279
rect 800 71279 1000 81161
rect 800 71161 841 71279
rect 959 71161 1000 71279
rect 800 61279 1000 71161
rect 800 61161 841 61279
rect 959 61161 1000 61279
rect 800 51279 1000 61161
rect 800 51161 841 51279
rect 959 51161 1000 51279
rect 800 41279 1000 51161
rect 800 41161 841 41279
rect 959 41161 1000 41279
rect 800 31279 1000 41161
rect 800 31161 841 31279
rect 959 31161 1000 31279
rect 800 21279 1000 31161
rect 800 21161 841 21279
rect 959 21161 1000 21279
rect 800 11279 1000 21161
rect 800 11161 841 11279
rect 959 11161 1000 11279
rect 800 959 1000 11161
rect 1200 357151 1400 357192
rect 1200 357033 1241 357151
rect 1359 357033 1400 357151
rect 1200 346279 1400 357033
rect 6120 357151 6320 357592
rect 6120 357033 6161 357151
rect 6279 357033 6320 357151
rect 1200 346161 1241 346279
rect 1359 346161 1400 346279
rect 1200 336279 1400 346161
rect 1200 336161 1241 336279
rect 1359 336161 1400 336279
rect 1200 326279 1400 336161
rect 1200 326161 1241 326279
rect 1359 326161 1400 326279
rect 1200 316279 1400 326161
rect 1200 316161 1241 316279
rect 1359 316161 1400 316279
rect 1200 306279 1400 316161
rect 1200 306161 1241 306279
rect 1359 306161 1400 306279
rect 1200 296279 1400 306161
rect 1200 296161 1241 296279
rect 1359 296161 1400 296279
rect 1200 286279 1400 296161
rect 1200 286161 1241 286279
rect 1359 286161 1400 286279
rect 1200 276279 1400 286161
rect 1200 276161 1241 276279
rect 1359 276161 1400 276279
rect 1200 266279 1400 276161
rect 1200 266161 1241 266279
rect 1359 266161 1400 266279
rect 1200 256279 1400 266161
rect 1200 256161 1241 256279
rect 1359 256161 1400 256279
rect 1200 246279 1400 256161
rect 1200 246161 1241 246279
rect 1359 246161 1400 246279
rect 1200 236279 1400 246161
rect 1200 236161 1241 236279
rect 1359 236161 1400 236279
rect 1200 226279 1400 236161
rect 1200 226161 1241 226279
rect 1359 226161 1400 226279
rect 1200 216279 1400 226161
rect 1200 216161 1241 216279
rect 1359 216161 1400 216279
rect 1200 206279 1400 216161
rect 1200 206161 1241 206279
rect 1359 206161 1400 206279
rect 1200 196279 1400 206161
rect 1200 196161 1241 196279
rect 1359 196161 1400 196279
rect 1200 186279 1400 196161
rect 1200 186161 1241 186279
rect 1359 186161 1400 186279
rect 1200 176279 1400 186161
rect 1200 176161 1241 176279
rect 1359 176161 1400 176279
rect 1200 166279 1400 176161
rect 1200 166161 1241 166279
rect 1359 166161 1400 166279
rect 1200 156279 1400 166161
rect 1200 156161 1241 156279
rect 1359 156161 1400 156279
rect 1200 146279 1400 156161
rect 1200 146161 1241 146279
rect 1359 146161 1400 146279
rect 1200 136279 1400 146161
rect 1200 136161 1241 136279
rect 1359 136161 1400 136279
rect 1200 126279 1400 136161
rect 1200 126161 1241 126279
rect 1359 126161 1400 126279
rect 1200 116279 1400 126161
rect 1200 116161 1241 116279
rect 1359 116161 1400 116279
rect 1200 106279 1400 116161
rect 1200 106161 1241 106279
rect 1359 106161 1400 106279
rect 1200 96279 1400 106161
rect 1200 96161 1241 96279
rect 1359 96161 1400 96279
rect 1200 86279 1400 96161
rect 1200 86161 1241 86279
rect 1359 86161 1400 86279
rect 1200 76279 1400 86161
rect 1200 76161 1241 76279
rect 1359 76161 1400 76279
rect 1200 66279 1400 76161
rect 1200 66161 1241 66279
rect 1359 66161 1400 66279
rect 1200 56279 1400 66161
rect 1200 56161 1241 56279
rect 1359 56161 1400 56279
rect 1200 46279 1400 56161
rect 1200 46161 1241 46279
rect 1359 46161 1400 46279
rect 1200 36279 1400 46161
rect 1200 36161 1241 36279
rect 1359 36161 1400 36279
rect 1200 26279 1400 36161
rect 1200 26161 1241 26279
rect 1359 26161 1400 26279
rect 1200 16279 1400 26161
rect 1200 16161 1241 16279
rect 1359 16161 1400 16279
rect 1200 6279 1400 16161
rect 1200 6161 1241 6279
rect 1359 6161 1400 6279
rect 1200 1359 1400 6161
rect 1600 356751 1800 356792
rect 1600 356633 1641 356751
rect 1759 356633 1800 356751
rect 1600 350319 1800 356633
rect 1600 350201 1641 350319
rect 1759 350201 1800 350319
rect 1600 340319 1800 350201
rect 1600 340201 1641 340319
rect 1759 340201 1800 340319
rect 1600 330319 1800 340201
rect 1600 330201 1641 330319
rect 1759 330201 1800 330319
rect 1600 320319 1800 330201
rect 1600 320201 1641 320319
rect 1759 320201 1800 320319
rect 1600 310319 1800 320201
rect 1600 310201 1641 310319
rect 1759 310201 1800 310319
rect 1600 300319 1800 310201
rect 1600 300201 1641 300319
rect 1759 300201 1800 300319
rect 1600 290319 1800 300201
rect 1600 290201 1641 290319
rect 1759 290201 1800 290319
rect 1600 280319 1800 290201
rect 1600 280201 1641 280319
rect 1759 280201 1800 280319
rect 1600 270319 1800 280201
rect 1600 270201 1641 270319
rect 1759 270201 1800 270319
rect 1600 260319 1800 270201
rect 1600 260201 1641 260319
rect 1759 260201 1800 260319
rect 1600 250319 1800 260201
rect 1600 250201 1641 250319
rect 1759 250201 1800 250319
rect 1600 240319 1800 250201
rect 1600 240201 1641 240319
rect 1759 240201 1800 240319
rect 1600 230319 1800 240201
rect 1600 230201 1641 230319
rect 1759 230201 1800 230319
rect 1600 220319 1800 230201
rect 1600 220201 1641 220319
rect 1759 220201 1800 220319
rect 1600 210319 1800 220201
rect 1600 210201 1641 210319
rect 1759 210201 1800 210319
rect 1600 200319 1800 210201
rect 1600 200201 1641 200319
rect 1759 200201 1800 200319
rect 1600 190319 1800 200201
rect 1600 190201 1641 190319
rect 1759 190201 1800 190319
rect 1600 180319 1800 190201
rect 1600 180201 1641 180319
rect 1759 180201 1800 180319
rect 1600 170319 1800 180201
rect 1600 170201 1641 170319
rect 1759 170201 1800 170319
rect 1600 160319 1800 170201
rect 1600 160201 1641 160319
rect 1759 160201 1800 160319
rect 1600 150319 1800 160201
rect 1600 150201 1641 150319
rect 1759 150201 1800 150319
rect 1600 140319 1800 150201
rect 1600 140201 1641 140319
rect 1759 140201 1800 140319
rect 1600 130319 1800 140201
rect 1600 130201 1641 130319
rect 1759 130201 1800 130319
rect 1600 120319 1800 130201
rect 1600 120201 1641 120319
rect 1759 120201 1800 120319
rect 1600 110319 1800 120201
rect 1600 110201 1641 110319
rect 1759 110201 1800 110319
rect 1600 100319 1800 110201
rect 1600 100201 1641 100319
rect 1759 100201 1800 100319
rect 1600 90319 1800 100201
rect 1600 90201 1641 90319
rect 1759 90201 1800 90319
rect 1600 80319 1800 90201
rect 1600 80201 1641 80319
rect 1759 80201 1800 80319
rect 1600 70319 1800 80201
rect 1600 70201 1641 70319
rect 1759 70201 1800 70319
rect 1600 60319 1800 70201
rect 1600 60201 1641 60319
rect 1759 60201 1800 60319
rect 1600 50319 1800 60201
rect 1600 50201 1641 50319
rect 1759 50201 1800 50319
rect 1600 40319 1800 50201
rect 1600 40201 1641 40319
rect 1759 40201 1800 40319
rect 1600 30319 1800 40201
rect 1600 30201 1641 30319
rect 1759 30201 1800 30319
rect 1600 20319 1800 30201
rect 1600 20201 1641 20319
rect 1759 20201 1800 20319
rect 1600 10319 1800 20201
rect 1600 10201 1641 10319
rect 1759 10201 1800 10319
rect 1600 1759 1800 10201
rect 2000 356351 2200 356392
rect 2000 356233 2041 356351
rect 2159 356233 2200 356351
rect 2000 345319 2200 356233
rect 5160 356351 5360 356792
rect 5160 356233 5201 356351
rect 5319 356233 5360 356351
rect 2000 345201 2041 345319
rect 2159 345201 2200 345319
rect 2000 335319 2200 345201
rect 2000 335201 2041 335319
rect 2159 335201 2200 335319
rect 2000 325319 2200 335201
rect 2000 325201 2041 325319
rect 2159 325201 2200 325319
rect 2000 315319 2200 325201
rect 2000 315201 2041 315319
rect 2159 315201 2200 315319
rect 2000 305319 2200 315201
rect 2000 305201 2041 305319
rect 2159 305201 2200 305319
rect 2000 295319 2200 305201
rect 2000 295201 2041 295319
rect 2159 295201 2200 295319
rect 2000 285319 2200 295201
rect 2000 285201 2041 285319
rect 2159 285201 2200 285319
rect 2000 275319 2200 285201
rect 2000 275201 2041 275319
rect 2159 275201 2200 275319
rect 2000 265319 2200 275201
rect 2000 265201 2041 265319
rect 2159 265201 2200 265319
rect 2000 255319 2200 265201
rect 2000 255201 2041 255319
rect 2159 255201 2200 255319
rect 2000 245319 2200 255201
rect 2000 245201 2041 245319
rect 2159 245201 2200 245319
rect 2000 235319 2200 245201
rect 2000 235201 2041 235319
rect 2159 235201 2200 235319
rect 2000 225319 2200 235201
rect 2000 225201 2041 225319
rect 2159 225201 2200 225319
rect 2000 215319 2200 225201
rect 2000 215201 2041 215319
rect 2159 215201 2200 215319
rect 2000 205319 2200 215201
rect 2000 205201 2041 205319
rect 2159 205201 2200 205319
rect 2000 195319 2200 205201
rect 2000 195201 2041 195319
rect 2159 195201 2200 195319
rect 2000 185319 2200 195201
rect 2000 185201 2041 185319
rect 2159 185201 2200 185319
rect 2000 175319 2200 185201
rect 2000 175201 2041 175319
rect 2159 175201 2200 175319
rect 2000 165319 2200 175201
rect 2000 165201 2041 165319
rect 2159 165201 2200 165319
rect 2000 155319 2200 165201
rect 2000 155201 2041 155319
rect 2159 155201 2200 155319
rect 2000 145319 2200 155201
rect 2000 145201 2041 145319
rect 2159 145201 2200 145319
rect 2000 135319 2200 145201
rect 2000 135201 2041 135319
rect 2159 135201 2200 135319
rect 2000 125319 2200 135201
rect 2000 125201 2041 125319
rect 2159 125201 2200 125319
rect 2000 115319 2200 125201
rect 2000 115201 2041 115319
rect 2159 115201 2200 115319
rect 2000 105319 2200 115201
rect 2000 105201 2041 105319
rect 2159 105201 2200 105319
rect 2000 95319 2200 105201
rect 2000 95201 2041 95319
rect 2159 95201 2200 95319
rect 2000 85319 2200 95201
rect 2000 85201 2041 85319
rect 2159 85201 2200 85319
rect 2000 75319 2200 85201
rect 2000 75201 2041 75319
rect 2159 75201 2200 75319
rect 2000 65319 2200 75201
rect 2000 65201 2041 65319
rect 2159 65201 2200 65319
rect 2000 55319 2200 65201
rect 2000 55201 2041 55319
rect 2159 55201 2200 55319
rect 2000 45319 2200 55201
rect 2000 45201 2041 45319
rect 2159 45201 2200 45319
rect 2000 35319 2200 45201
rect 2000 35201 2041 35319
rect 2159 35201 2200 35319
rect 2000 25319 2200 35201
rect 2000 25201 2041 25319
rect 2159 25201 2200 25319
rect 2000 15319 2200 25201
rect 2000 15201 2041 15319
rect 2159 15201 2200 15319
rect 2000 5319 2200 15201
rect 2000 5201 2041 5319
rect 2159 5201 2200 5319
rect 2000 2159 2200 5201
rect 2400 355951 2600 355992
rect 2400 355833 2441 355951
rect 2559 355833 2600 355951
rect 2400 349359 2600 355833
rect 2400 349241 2441 349359
rect 2559 349241 2600 349359
rect 2400 339359 2600 349241
rect 2400 339241 2441 339359
rect 2559 339241 2600 339359
rect 2400 329359 2600 339241
rect 2400 329241 2441 329359
rect 2559 329241 2600 329359
rect 2400 319359 2600 329241
rect 2400 319241 2441 319359
rect 2559 319241 2600 319359
rect 2400 309359 2600 319241
rect 2400 309241 2441 309359
rect 2559 309241 2600 309359
rect 2400 299359 2600 309241
rect 2400 299241 2441 299359
rect 2559 299241 2600 299359
rect 2400 289359 2600 299241
rect 2400 289241 2441 289359
rect 2559 289241 2600 289359
rect 2400 279359 2600 289241
rect 2400 279241 2441 279359
rect 2559 279241 2600 279359
rect 2400 269359 2600 279241
rect 2400 269241 2441 269359
rect 2559 269241 2600 269359
rect 2400 259359 2600 269241
rect 2400 259241 2441 259359
rect 2559 259241 2600 259359
rect 2400 249359 2600 259241
rect 2400 249241 2441 249359
rect 2559 249241 2600 249359
rect 2400 239359 2600 249241
rect 2400 239241 2441 239359
rect 2559 239241 2600 239359
rect 2400 229359 2600 239241
rect 2400 229241 2441 229359
rect 2559 229241 2600 229359
rect 2400 219359 2600 229241
rect 2400 219241 2441 219359
rect 2559 219241 2600 219359
rect 2400 209359 2600 219241
rect 2400 209241 2441 209359
rect 2559 209241 2600 209359
rect 2400 199359 2600 209241
rect 2400 199241 2441 199359
rect 2559 199241 2600 199359
rect 2400 189359 2600 199241
rect 2400 189241 2441 189359
rect 2559 189241 2600 189359
rect 2400 179359 2600 189241
rect 2400 179241 2441 179359
rect 2559 179241 2600 179359
rect 2400 169359 2600 179241
rect 2400 169241 2441 169359
rect 2559 169241 2600 169359
rect 2400 159359 2600 169241
rect 2400 159241 2441 159359
rect 2559 159241 2600 159359
rect 2400 149359 2600 159241
rect 2400 149241 2441 149359
rect 2559 149241 2600 149359
rect 2400 139359 2600 149241
rect 2400 139241 2441 139359
rect 2559 139241 2600 139359
rect 2400 129359 2600 139241
rect 2400 129241 2441 129359
rect 2559 129241 2600 129359
rect 2400 119359 2600 129241
rect 2400 119241 2441 119359
rect 2559 119241 2600 119359
rect 2400 109359 2600 119241
rect 2400 109241 2441 109359
rect 2559 109241 2600 109359
rect 2400 99359 2600 109241
rect 2400 99241 2441 99359
rect 2559 99241 2600 99359
rect 2400 89359 2600 99241
rect 2400 89241 2441 89359
rect 2559 89241 2600 89359
rect 2400 79359 2600 89241
rect 2400 79241 2441 79359
rect 2559 79241 2600 79359
rect 2400 69359 2600 79241
rect 2400 69241 2441 69359
rect 2559 69241 2600 69359
rect 2400 59359 2600 69241
rect 2400 59241 2441 59359
rect 2559 59241 2600 59359
rect 2400 49359 2600 59241
rect 2400 49241 2441 49359
rect 2559 49241 2600 49359
rect 2400 39359 2600 49241
rect 2400 39241 2441 39359
rect 2559 39241 2600 39359
rect 2400 29359 2600 39241
rect 2400 29241 2441 29359
rect 2559 29241 2600 29359
rect 2400 19359 2600 29241
rect 2400 19241 2441 19359
rect 2559 19241 2600 19359
rect 2400 9359 2600 19241
rect 2400 9241 2441 9359
rect 2559 9241 2600 9359
rect 2400 2559 2600 9241
rect 2800 355551 3000 355592
rect 2800 355433 2841 355551
rect 2959 355433 3000 355551
rect 2800 344359 3000 355433
rect 4200 355551 4400 355992
rect 4200 355433 4241 355551
rect 4359 355433 4400 355551
rect 4200 354972 4400 355433
rect 5160 354972 5360 356233
rect 6120 354972 6320 357033
rect 7080 354972 7280 357833
rect 12080 358351 12280 358392
rect 12080 358233 12121 358351
rect 12239 358233 12280 358351
rect 11120 357551 11320 357592
rect 11120 357433 11161 357551
rect 11279 357433 11320 357551
rect 10160 356751 10360 356792
rect 10160 356633 10201 356751
rect 10319 356633 10360 356751
rect 9200 355951 9400 355992
rect 9200 355833 9241 355951
rect 9359 355833 9400 355951
rect 9200 354972 9400 355833
rect 10160 354972 10360 356633
rect 11120 354972 11320 357433
rect 12080 354972 12280 358233
rect 17080 357951 17280 358392
rect 17080 357833 17121 357951
rect 17239 357833 17280 357951
rect 16120 357151 16320 357592
rect 16120 357033 16161 357151
rect 16279 357033 16320 357151
rect 15160 356351 15360 356792
rect 15160 356233 15201 356351
rect 15319 356233 15360 356351
rect 14200 355551 14400 355992
rect 14200 355433 14241 355551
rect 14359 355433 14400 355551
rect 14200 354972 14400 355433
rect 15160 354972 15360 356233
rect 16120 354972 16320 357033
rect 17080 354972 17280 357833
rect 22080 358351 22280 358392
rect 22080 358233 22121 358351
rect 22239 358233 22280 358351
rect 21120 357551 21320 357592
rect 21120 357433 21161 357551
rect 21279 357433 21320 357551
rect 20160 356751 20360 356792
rect 20160 356633 20201 356751
rect 20319 356633 20360 356751
rect 19200 355951 19400 355992
rect 19200 355833 19241 355951
rect 19359 355833 19400 355951
rect 19200 354972 19400 355833
rect 20160 354972 20360 356633
rect 21120 354972 21320 357433
rect 22080 354972 22280 358233
rect 27080 357951 27280 358392
rect 27080 357833 27121 357951
rect 27239 357833 27280 357951
rect 26120 357151 26320 357592
rect 26120 357033 26161 357151
rect 26279 357033 26320 357151
rect 25160 356351 25360 356792
rect 25160 356233 25201 356351
rect 25319 356233 25360 356351
rect 24200 355551 24400 355992
rect 24200 355433 24241 355551
rect 24359 355433 24400 355551
rect 24200 354972 24400 355433
rect 25160 354972 25360 356233
rect 26120 354972 26320 357033
rect 27080 354972 27280 357833
rect 32080 358351 32280 358392
rect 32080 358233 32121 358351
rect 32239 358233 32280 358351
rect 31120 357551 31320 357592
rect 31120 357433 31161 357551
rect 31279 357433 31320 357551
rect 30160 356751 30360 356792
rect 30160 356633 30201 356751
rect 30319 356633 30360 356751
rect 29200 355951 29400 355992
rect 29200 355833 29241 355951
rect 29359 355833 29400 355951
rect 29200 354972 29400 355833
rect 30160 354972 30360 356633
rect 31120 354972 31320 357433
rect 32080 354972 32280 358233
rect 37080 357951 37280 358392
rect 37080 357833 37121 357951
rect 37239 357833 37280 357951
rect 36120 357151 36320 357592
rect 36120 357033 36161 357151
rect 36279 357033 36320 357151
rect 35160 356351 35360 356792
rect 35160 356233 35201 356351
rect 35319 356233 35360 356351
rect 34200 355551 34400 355992
rect 34200 355433 34241 355551
rect 34359 355433 34400 355551
rect 34200 354972 34400 355433
rect 35160 354972 35360 356233
rect 36120 354972 36320 357033
rect 37080 354972 37280 357833
rect 42080 358351 42280 358392
rect 42080 358233 42121 358351
rect 42239 358233 42280 358351
rect 41120 357551 41320 357592
rect 41120 357433 41161 357551
rect 41279 357433 41320 357551
rect 40160 356751 40360 356792
rect 40160 356633 40201 356751
rect 40319 356633 40360 356751
rect 39200 355951 39400 355992
rect 39200 355833 39241 355951
rect 39359 355833 39400 355951
rect 39200 354972 39400 355833
rect 40160 354972 40360 356633
rect 41120 354972 41320 357433
rect 42080 354972 42280 358233
rect 47080 357951 47280 358392
rect 47080 357833 47121 357951
rect 47239 357833 47280 357951
rect 46120 357151 46320 357592
rect 46120 357033 46161 357151
rect 46279 357033 46320 357151
rect 45160 356351 45360 356792
rect 45160 356233 45201 356351
rect 45319 356233 45360 356351
rect 44200 355551 44400 355992
rect 44200 355433 44241 355551
rect 44359 355433 44400 355551
rect 44200 354972 44400 355433
rect 45160 354972 45360 356233
rect 46120 354972 46320 357033
rect 47080 354972 47280 357833
rect 52080 358351 52280 358392
rect 52080 358233 52121 358351
rect 52239 358233 52280 358351
rect 51120 357551 51320 357592
rect 51120 357433 51161 357551
rect 51279 357433 51320 357551
rect 50160 356751 50360 356792
rect 50160 356633 50201 356751
rect 50319 356633 50360 356751
rect 49200 355951 49400 355992
rect 49200 355833 49241 355951
rect 49359 355833 49400 355951
rect 49200 354972 49400 355833
rect 50160 354972 50360 356633
rect 51120 354972 51320 357433
rect 52080 354972 52280 358233
rect 57080 357951 57280 358392
rect 57080 357833 57121 357951
rect 57239 357833 57280 357951
rect 56120 357151 56320 357592
rect 56120 357033 56161 357151
rect 56279 357033 56320 357151
rect 55160 356351 55360 356792
rect 55160 356233 55201 356351
rect 55319 356233 55360 356351
rect 54200 355551 54400 355992
rect 54200 355433 54241 355551
rect 54359 355433 54400 355551
rect 54200 354972 54400 355433
rect 55160 354972 55360 356233
rect 56120 354972 56320 357033
rect 57080 354972 57280 357833
rect 62080 358351 62280 358392
rect 62080 358233 62121 358351
rect 62239 358233 62280 358351
rect 61120 357551 61320 357592
rect 61120 357433 61161 357551
rect 61279 357433 61320 357551
rect 60160 356751 60360 356792
rect 60160 356633 60201 356751
rect 60319 356633 60360 356751
rect 59200 355951 59400 355992
rect 59200 355833 59241 355951
rect 59359 355833 59400 355951
rect 59200 354972 59400 355833
rect 60160 354972 60360 356633
rect 61120 354972 61320 357433
rect 62080 354972 62280 358233
rect 67080 357951 67280 358392
rect 67080 357833 67121 357951
rect 67239 357833 67280 357951
rect 66120 357151 66320 357592
rect 66120 357033 66161 357151
rect 66279 357033 66320 357151
rect 65160 356351 65360 356792
rect 65160 356233 65201 356351
rect 65319 356233 65360 356351
rect 64200 355551 64400 355992
rect 64200 355433 64241 355551
rect 64359 355433 64400 355551
rect 64200 354972 64400 355433
rect 65160 354972 65360 356233
rect 66120 354972 66320 357033
rect 67080 354972 67280 357833
rect 72080 358351 72280 358392
rect 72080 358233 72121 358351
rect 72239 358233 72280 358351
rect 71120 357551 71320 357592
rect 71120 357433 71161 357551
rect 71279 357433 71320 357551
rect 70160 356751 70360 356792
rect 70160 356633 70201 356751
rect 70319 356633 70360 356751
rect 69200 355951 69400 355992
rect 69200 355833 69241 355951
rect 69359 355833 69400 355951
rect 69200 354972 69400 355833
rect 70160 354972 70360 356633
rect 71120 354972 71320 357433
rect 72080 354972 72280 358233
rect 77080 357951 77280 358392
rect 77080 357833 77121 357951
rect 77239 357833 77280 357951
rect 76120 357151 76320 357592
rect 76120 357033 76161 357151
rect 76279 357033 76320 357151
rect 75160 356351 75360 356792
rect 75160 356233 75201 356351
rect 75319 356233 75360 356351
rect 74200 355551 74400 355992
rect 74200 355433 74241 355551
rect 74359 355433 74400 355551
rect 74200 354972 74400 355433
rect 75160 354972 75360 356233
rect 76120 354972 76320 357033
rect 77080 354972 77280 357833
rect 82080 358351 82280 358392
rect 82080 358233 82121 358351
rect 82239 358233 82280 358351
rect 81120 357551 81320 357592
rect 81120 357433 81161 357551
rect 81279 357433 81320 357551
rect 80160 356751 80360 356792
rect 80160 356633 80201 356751
rect 80319 356633 80360 356751
rect 79200 355951 79400 355992
rect 79200 355833 79241 355951
rect 79359 355833 79400 355951
rect 79200 354972 79400 355833
rect 80160 354972 80360 356633
rect 81120 354972 81320 357433
rect 82080 354972 82280 358233
rect 87080 357951 87280 358392
rect 87080 357833 87121 357951
rect 87239 357833 87280 357951
rect 86120 357151 86320 357592
rect 86120 357033 86161 357151
rect 86279 357033 86320 357151
rect 85160 356351 85360 356792
rect 85160 356233 85201 356351
rect 85319 356233 85360 356351
rect 84200 355551 84400 355992
rect 84200 355433 84241 355551
rect 84359 355433 84400 355551
rect 84200 354972 84400 355433
rect 85160 354972 85360 356233
rect 86120 354972 86320 357033
rect 87080 354972 87280 357833
rect 92080 358351 92280 358392
rect 92080 358233 92121 358351
rect 92239 358233 92280 358351
rect 91120 357551 91320 357592
rect 91120 357433 91161 357551
rect 91279 357433 91320 357551
rect 90160 356751 90360 356792
rect 90160 356633 90201 356751
rect 90319 356633 90360 356751
rect 89200 355951 89400 355992
rect 89200 355833 89241 355951
rect 89359 355833 89400 355951
rect 89200 354972 89400 355833
rect 90160 354972 90360 356633
rect 91120 354972 91320 357433
rect 92080 354972 92280 358233
rect 97080 357951 97280 358392
rect 97080 357833 97121 357951
rect 97239 357833 97280 357951
rect 96120 357151 96320 357592
rect 96120 357033 96161 357151
rect 96279 357033 96320 357151
rect 95160 356351 95360 356792
rect 95160 356233 95201 356351
rect 95319 356233 95360 356351
rect 94200 355551 94400 355992
rect 94200 355433 94241 355551
rect 94359 355433 94400 355551
rect 94200 354972 94400 355433
rect 95160 354972 95360 356233
rect 96120 354972 96320 357033
rect 97080 354972 97280 357833
rect 102080 358351 102280 358392
rect 102080 358233 102121 358351
rect 102239 358233 102280 358351
rect 101120 357551 101320 357592
rect 101120 357433 101161 357551
rect 101279 357433 101320 357551
rect 100160 356751 100360 356792
rect 100160 356633 100201 356751
rect 100319 356633 100360 356751
rect 99200 355951 99400 355992
rect 99200 355833 99241 355951
rect 99359 355833 99400 355951
rect 99200 354972 99400 355833
rect 100160 354972 100360 356633
rect 101120 354972 101320 357433
rect 102080 354972 102280 358233
rect 107080 357951 107280 358392
rect 107080 357833 107121 357951
rect 107239 357833 107280 357951
rect 106120 357151 106320 357592
rect 106120 357033 106161 357151
rect 106279 357033 106320 357151
rect 105160 356351 105360 356792
rect 105160 356233 105201 356351
rect 105319 356233 105360 356351
rect 104200 355551 104400 355992
rect 104200 355433 104241 355551
rect 104359 355433 104400 355551
rect 104200 354972 104400 355433
rect 105160 354972 105360 356233
rect 106120 354972 106320 357033
rect 107080 354972 107280 357833
rect 112080 358351 112280 358392
rect 112080 358233 112121 358351
rect 112239 358233 112280 358351
rect 111120 357551 111320 357592
rect 111120 357433 111161 357551
rect 111279 357433 111320 357551
rect 110160 356751 110360 356792
rect 110160 356633 110201 356751
rect 110319 356633 110360 356751
rect 109200 355951 109400 355992
rect 109200 355833 109241 355951
rect 109359 355833 109400 355951
rect 109200 354972 109400 355833
rect 110160 354972 110360 356633
rect 111120 354972 111320 357433
rect 112080 354972 112280 358233
rect 117080 357951 117280 358392
rect 117080 357833 117121 357951
rect 117239 357833 117280 357951
rect 116120 357151 116320 357592
rect 116120 357033 116161 357151
rect 116279 357033 116320 357151
rect 115160 356351 115360 356792
rect 115160 356233 115201 356351
rect 115319 356233 115360 356351
rect 114200 355551 114400 355992
rect 114200 355433 114241 355551
rect 114359 355433 114400 355551
rect 114200 354972 114400 355433
rect 115160 354972 115360 356233
rect 116120 354972 116320 357033
rect 117080 354972 117280 357833
rect 122080 358351 122280 358392
rect 122080 358233 122121 358351
rect 122239 358233 122280 358351
rect 121120 357551 121320 357592
rect 121120 357433 121161 357551
rect 121279 357433 121320 357551
rect 120160 356751 120360 356792
rect 120160 356633 120201 356751
rect 120319 356633 120360 356751
rect 119200 355951 119400 355992
rect 119200 355833 119241 355951
rect 119359 355833 119400 355951
rect 119200 354972 119400 355833
rect 120160 354972 120360 356633
rect 121120 354972 121320 357433
rect 122080 354972 122280 358233
rect 127080 357951 127280 358392
rect 127080 357833 127121 357951
rect 127239 357833 127280 357951
rect 126120 357151 126320 357592
rect 126120 357033 126161 357151
rect 126279 357033 126320 357151
rect 125160 356351 125360 356792
rect 125160 356233 125201 356351
rect 125319 356233 125360 356351
rect 124200 355551 124400 355992
rect 124200 355433 124241 355551
rect 124359 355433 124400 355551
rect 124200 354972 124400 355433
rect 125160 354972 125360 356233
rect 126120 354972 126320 357033
rect 127080 354972 127280 357833
rect 132080 358351 132280 358392
rect 132080 358233 132121 358351
rect 132239 358233 132280 358351
rect 131120 357551 131320 357592
rect 131120 357433 131161 357551
rect 131279 357433 131320 357551
rect 130160 356751 130360 356792
rect 130160 356633 130201 356751
rect 130319 356633 130360 356751
rect 129200 355951 129400 355992
rect 129200 355833 129241 355951
rect 129359 355833 129400 355951
rect 129200 354972 129400 355833
rect 130160 354972 130360 356633
rect 131120 354972 131320 357433
rect 132080 354972 132280 358233
rect 137080 357951 137280 358392
rect 137080 357833 137121 357951
rect 137239 357833 137280 357951
rect 136120 357151 136320 357592
rect 136120 357033 136161 357151
rect 136279 357033 136320 357151
rect 135160 356351 135360 356792
rect 135160 356233 135201 356351
rect 135319 356233 135360 356351
rect 134200 355551 134400 355992
rect 134200 355433 134241 355551
rect 134359 355433 134400 355551
rect 134200 354972 134400 355433
rect 135160 354972 135360 356233
rect 136120 354972 136320 357033
rect 137080 354972 137280 357833
rect 142080 358351 142280 358392
rect 142080 358233 142121 358351
rect 142239 358233 142280 358351
rect 141120 357551 141320 357592
rect 141120 357433 141161 357551
rect 141279 357433 141320 357551
rect 140160 356751 140360 356792
rect 140160 356633 140201 356751
rect 140319 356633 140360 356751
rect 139200 355951 139400 355992
rect 139200 355833 139241 355951
rect 139359 355833 139400 355951
rect 139200 354972 139400 355833
rect 140160 354972 140360 356633
rect 141120 354972 141320 357433
rect 142080 354972 142280 358233
rect 147080 357951 147280 358392
rect 147080 357833 147121 357951
rect 147239 357833 147280 357951
rect 146120 357151 146320 357592
rect 146120 357033 146161 357151
rect 146279 357033 146320 357151
rect 145160 356351 145360 356792
rect 145160 356233 145201 356351
rect 145319 356233 145360 356351
rect 144200 355551 144400 355992
rect 144200 355433 144241 355551
rect 144359 355433 144400 355551
rect 144200 354972 144400 355433
rect 145160 354972 145360 356233
rect 146120 354972 146320 357033
rect 147080 354972 147280 357833
rect 152080 358351 152280 358392
rect 152080 358233 152121 358351
rect 152239 358233 152280 358351
rect 151120 357551 151320 357592
rect 151120 357433 151161 357551
rect 151279 357433 151320 357551
rect 150160 356751 150360 356792
rect 150160 356633 150201 356751
rect 150319 356633 150360 356751
rect 149200 355951 149400 355992
rect 149200 355833 149241 355951
rect 149359 355833 149400 355951
rect 149200 354972 149400 355833
rect 150160 354972 150360 356633
rect 151120 354972 151320 357433
rect 152080 354972 152280 358233
rect 157080 357951 157280 358392
rect 157080 357833 157121 357951
rect 157239 357833 157280 357951
rect 156120 357151 156320 357592
rect 156120 357033 156161 357151
rect 156279 357033 156320 357151
rect 155160 356351 155360 356792
rect 155160 356233 155201 356351
rect 155319 356233 155360 356351
rect 154200 355551 154400 355992
rect 154200 355433 154241 355551
rect 154359 355433 154400 355551
rect 154200 354972 154400 355433
rect 155160 354972 155360 356233
rect 156120 354972 156320 357033
rect 157080 354972 157280 357833
rect 162080 358351 162280 358392
rect 162080 358233 162121 358351
rect 162239 358233 162280 358351
rect 161120 357551 161320 357592
rect 161120 357433 161161 357551
rect 161279 357433 161320 357551
rect 160160 356751 160360 356792
rect 160160 356633 160201 356751
rect 160319 356633 160360 356751
rect 159200 355951 159400 355992
rect 159200 355833 159241 355951
rect 159359 355833 159400 355951
rect 159200 354972 159400 355833
rect 160160 354972 160360 356633
rect 161120 354972 161320 357433
rect 162080 354972 162280 358233
rect 167080 357951 167280 358392
rect 167080 357833 167121 357951
rect 167239 357833 167280 357951
rect 166120 357151 166320 357592
rect 166120 357033 166161 357151
rect 166279 357033 166320 357151
rect 165160 356351 165360 356792
rect 165160 356233 165201 356351
rect 165319 356233 165360 356351
rect 164200 355551 164400 355992
rect 164200 355433 164241 355551
rect 164359 355433 164400 355551
rect 164200 354972 164400 355433
rect 165160 354972 165360 356233
rect 166120 354972 166320 357033
rect 167080 354972 167280 357833
rect 172080 358351 172280 358392
rect 172080 358233 172121 358351
rect 172239 358233 172280 358351
rect 171120 357551 171320 357592
rect 171120 357433 171161 357551
rect 171279 357433 171320 357551
rect 170160 356751 170360 356792
rect 170160 356633 170201 356751
rect 170319 356633 170360 356751
rect 169200 355951 169400 355992
rect 169200 355833 169241 355951
rect 169359 355833 169400 355951
rect 169200 354972 169400 355833
rect 170160 354972 170360 356633
rect 171120 354972 171320 357433
rect 172080 354972 172280 358233
rect 177080 357951 177280 358392
rect 177080 357833 177121 357951
rect 177239 357833 177280 357951
rect 176120 357151 176320 357592
rect 176120 357033 176161 357151
rect 176279 357033 176320 357151
rect 175160 356351 175360 356792
rect 175160 356233 175201 356351
rect 175319 356233 175360 356351
rect 174200 355551 174400 355992
rect 174200 355433 174241 355551
rect 174359 355433 174400 355551
rect 174200 354972 174400 355433
rect 175160 354972 175360 356233
rect 176120 354972 176320 357033
rect 177080 354972 177280 357833
rect 182080 358351 182280 358392
rect 182080 358233 182121 358351
rect 182239 358233 182280 358351
rect 181120 357551 181320 357592
rect 181120 357433 181161 357551
rect 181279 357433 181320 357551
rect 180160 356751 180360 356792
rect 180160 356633 180201 356751
rect 180319 356633 180360 356751
rect 179200 355951 179400 355992
rect 179200 355833 179241 355951
rect 179359 355833 179400 355951
rect 179200 354972 179400 355833
rect 180160 354972 180360 356633
rect 181120 354972 181320 357433
rect 182080 354972 182280 358233
rect 187080 357951 187280 358392
rect 187080 357833 187121 357951
rect 187239 357833 187280 357951
rect 186120 357151 186320 357592
rect 186120 357033 186161 357151
rect 186279 357033 186320 357151
rect 185160 356351 185360 356792
rect 185160 356233 185201 356351
rect 185319 356233 185360 356351
rect 184200 355551 184400 355992
rect 184200 355433 184241 355551
rect 184359 355433 184400 355551
rect 184200 354972 184400 355433
rect 185160 354972 185360 356233
rect 186120 354972 186320 357033
rect 187080 354972 187280 357833
rect 192080 358351 192280 358392
rect 192080 358233 192121 358351
rect 192239 358233 192280 358351
rect 191120 357551 191320 357592
rect 191120 357433 191161 357551
rect 191279 357433 191320 357551
rect 190160 356751 190360 356792
rect 190160 356633 190201 356751
rect 190319 356633 190360 356751
rect 189200 355951 189400 355992
rect 189200 355833 189241 355951
rect 189359 355833 189400 355951
rect 189200 354972 189400 355833
rect 190160 354972 190360 356633
rect 191120 354972 191320 357433
rect 192080 354972 192280 358233
rect 197080 357951 197280 358392
rect 197080 357833 197121 357951
rect 197239 357833 197280 357951
rect 196120 357151 196320 357592
rect 196120 357033 196161 357151
rect 196279 357033 196320 357151
rect 195160 356351 195360 356792
rect 195160 356233 195201 356351
rect 195319 356233 195360 356351
rect 194200 355551 194400 355992
rect 194200 355433 194241 355551
rect 194359 355433 194400 355551
rect 194200 354972 194400 355433
rect 195160 354972 195360 356233
rect 196120 354972 196320 357033
rect 197080 354972 197280 357833
rect 202080 358351 202280 358392
rect 202080 358233 202121 358351
rect 202239 358233 202280 358351
rect 201120 357551 201320 357592
rect 201120 357433 201161 357551
rect 201279 357433 201320 357551
rect 200160 356751 200360 356792
rect 200160 356633 200201 356751
rect 200319 356633 200360 356751
rect 199200 355951 199400 355992
rect 199200 355833 199241 355951
rect 199359 355833 199400 355951
rect 199200 354972 199400 355833
rect 200160 354972 200360 356633
rect 201120 354972 201320 357433
rect 202080 354972 202280 358233
rect 207080 357951 207280 358392
rect 207080 357833 207121 357951
rect 207239 357833 207280 357951
rect 206120 357151 206320 357592
rect 206120 357033 206161 357151
rect 206279 357033 206320 357151
rect 205160 356351 205360 356792
rect 205160 356233 205201 356351
rect 205319 356233 205360 356351
rect 204200 355551 204400 355992
rect 204200 355433 204241 355551
rect 204359 355433 204400 355551
rect 204200 354972 204400 355433
rect 205160 354972 205360 356233
rect 206120 354972 206320 357033
rect 207080 354972 207280 357833
rect 212080 358351 212280 358392
rect 212080 358233 212121 358351
rect 212239 358233 212280 358351
rect 211120 357551 211320 357592
rect 211120 357433 211161 357551
rect 211279 357433 211320 357551
rect 210160 356751 210360 356792
rect 210160 356633 210201 356751
rect 210319 356633 210360 356751
rect 209200 355951 209400 355992
rect 209200 355833 209241 355951
rect 209359 355833 209400 355951
rect 209200 354972 209400 355833
rect 210160 354972 210360 356633
rect 211120 354972 211320 357433
rect 212080 354972 212280 358233
rect 217080 357951 217280 358392
rect 217080 357833 217121 357951
rect 217239 357833 217280 357951
rect 216120 357151 216320 357592
rect 216120 357033 216161 357151
rect 216279 357033 216320 357151
rect 215160 356351 215360 356792
rect 215160 356233 215201 356351
rect 215319 356233 215360 356351
rect 214200 355551 214400 355992
rect 214200 355433 214241 355551
rect 214359 355433 214400 355551
rect 214200 354972 214400 355433
rect 215160 354972 215360 356233
rect 216120 354972 216320 357033
rect 217080 354972 217280 357833
rect 222080 358351 222280 358392
rect 222080 358233 222121 358351
rect 222239 358233 222280 358351
rect 221120 357551 221320 357592
rect 221120 357433 221161 357551
rect 221279 357433 221320 357551
rect 220160 356751 220360 356792
rect 220160 356633 220201 356751
rect 220319 356633 220360 356751
rect 219200 355951 219400 355992
rect 219200 355833 219241 355951
rect 219359 355833 219400 355951
rect 219200 354972 219400 355833
rect 220160 354972 220360 356633
rect 221120 354972 221320 357433
rect 222080 354972 222280 358233
rect 227080 357951 227280 358392
rect 227080 357833 227121 357951
rect 227239 357833 227280 357951
rect 226120 357151 226320 357592
rect 226120 357033 226161 357151
rect 226279 357033 226320 357151
rect 225160 356351 225360 356792
rect 225160 356233 225201 356351
rect 225319 356233 225360 356351
rect 224200 355551 224400 355992
rect 224200 355433 224241 355551
rect 224359 355433 224400 355551
rect 224200 354972 224400 355433
rect 225160 354972 225360 356233
rect 226120 354972 226320 357033
rect 227080 354972 227280 357833
rect 232080 358351 232280 358392
rect 232080 358233 232121 358351
rect 232239 358233 232280 358351
rect 231120 357551 231320 357592
rect 231120 357433 231161 357551
rect 231279 357433 231320 357551
rect 230160 356751 230360 356792
rect 230160 356633 230201 356751
rect 230319 356633 230360 356751
rect 229200 355951 229400 355992
rect 229200 355833 229241 355951
rect 229359 355833 229400 355951
rect 229200 354972 229400 355833
rect 230160 354972 230360 356633
rect 231120 354972 231320 357433
rect 232080 354972 232280 358233
rect 237080 357951 237280 358392
rect 237080 357833 237121 357951
rect 237239 357833 237280 357951
rect 236120 357151 236320 357592
rect 236120 357033 236161 357151
rect 236279 357033 236320 357151
rect 235160 356351 235360 356792
rect 235160 356233 235201 356351
rect 235319 356233 235360 356351
rect 234200 355551 234400 355992
rect 234200 355433 234241 355551
rect 234359 355433 234400 355551
rect 234200 354972 234400 355433
rect 235160 354972 235360 356233
rect 236120 354972 236320 357033
rect 237080 354972 237280 357833
rect 242080 358351 242280 358392
rect 242080 358233 242121 358351
rect 242239 358233 242280 358351
rect 241120 357551 241320 357592
rect 241120 357433 241161 357551
rect 241279 357433 241320 357551
rect 240160 356751 240360 356792
rect 240160 356633 240201 356751
rect 240319 356633 240360 356751
rect 239200 355951 239400 355992
rect 239200 355833 239241 355951
rect 239359 355833 239400 355951
rect 239200 354972 239400 355833
rect 240160 354972 240360 356633
rect 241120 354972 241320 357433
rect 242080 354972 242280 358233
rect 247080 357951 247280 358392
rect 247080 357833 247121 357951
rect 247239 357833 247280 357951
rect 246120 357151 246320 357592
rect 246120 357033 246161 357151
rect 246279 357033 246320 357151
rect 245160 356351 245360 356792
rect 245160 356233 245201 356351
rect 245319 356233 245360 356351
rect 244200 355551 244400 355992
rect 244200 355433 244241 355551
rect 244359 355433 244400 355551
rect 244200 354972 244400 355433
rect 245160 354972 245360 356233
rect 246120 354972 246320 357033
rect 247080 354972 247280 357833
rect 252080 358351 252280 358392
rect 252080 358233 252121 358351
rect 252239 358233 252280 358351
rect 251120 357551 251320 357592
rect 251120 357433 251161 357551
rect 251279 357433 251320 357551
rect 250160 356751 250360 356792
rect 250160 356633 250201 356751
rect 250319 356633 250360 356751
rect 249200 355951 249400 355992
rect 249200 355833 249241 355951
rect 249359 355833 249400 355951
rect 249200 354972 249400 355833
rect 250160 354972 250360 356633
rect 251120 354972 251320 357433
rect 252080 354972 252280 358233
rect 257080 357951 257280 358392
rect 257080 357833 257121 357951
rect 257239 357833 257280 357951
rect 256120 357151 256320 357592
rect 256120 357033 256161 357151
rect 256279 357033 256320 357151
rect 255160 356351 255360 356792
rect 255160 356233 255201 356351
rect 255319 356233 255360 356351
rect 254200 355551 254400 355992
rect 254200 355433 254241 355551
rect 254359 355433 254400 355551
rect 254200 354972 254400 355433
rect 255160 354972 255360 356233
rect 256120 354972 256320 357033
rect 257080 354972 257280 357833
rect 262080 358351 262280 358392
rect 262080 358233 262121 358351
rect 262239 358233 262280 358351
rect 261120 357551 261320 357592
rect 261120 357433 261161 357551
rect 261279 357433 261320 357551
rect 260160 356751 260360 356792
rect 260160 356633 260201 356751
rect 260319 356633 260360 356751
rect 259200 355951 259400 355992
rect 259200 355833 259241 355951
rect 259359 355833 259400 355951
rect 259200 354972 259400 355833
rect 260160 354972 260360 356633
rect 261120 354972 261320 357433
rect 262080 354972 262280 358233
rect 267080 357951 267280 358392
rect 267080 357833 267121 357951
rect 267239 357833 267280 357951
rect 266120 357151 266320 357592
rect 266120 357033 266161 357151
rect 266279 357033 266320 357151
rect 265160 356351 265360 356792
rect 265160 356233 265201 356351
rect 265319 356233 265360 356351
rect 264200 355551 264400 355992
rect 264200 355433 264241 355551
rect 264359 355433 264400 355551
rect 264200 354972 264400 355433
rect 265160 354972 265360 356233
rect 266120 354972 266320 357033
rect 267080 354972 267280 357833
rect 272080 358351 272280 358392
rect 272080 358233 272121 358351
rect 272239 358233 272280 358351
rect 271120 357551 271320 357592
rect 271120 357433 271161 357551
rect 271279 357433 271320 357551
rect 270160 356751 270360 356792
rect 270160 356633 270201 356751
rect 270319 356633 270360 356751
rect 269200 355951 269400 355992
rect 269200 355833 269241 355951
rect 269359 355833 269400 355951
rect 269200 354972 269400 355833
rect 270160 354972 270360 356633
rect 271120 354972 271320 357433
rect 272080 354972 272280 358233
rect 277080 357951 277280 358392
rect 277080 357833 277121 357951
rect 277239 357833 277280 357951
rect 276120 357151 276320 357592
rect 276120 357033 276161 357151
rect 276279 357033 276320 357151
rect 275160 356351 275360 356792
rect 275160 356233 275201 356351
rect 275319 356233 275360 356351
rect 274200 355551 274400 355992
rect 274200 355433 274241 355551
rect 274359 355433 274400 355551
rect 274200 354972 274400 355433
rect 275160 354972 275360 356233
rect 276120 354972 276320 357033
rect 277080 354972 277280 357833
rect 282080 358351 282280 358392
rect 282080 358233 282121 358351
rect 282239 358233 282280 358351
rect 281120 357551 281320 357592
rect 281120 357433 281161 357551
rect 281279 357433 281320 357551
rect 280160 356751 280360 356792
rect 280160 356633 280201 356751
rect 280319 356633 280360 356751
rect 279200 355951 279400 355992
rect 279200 355833 279241 355951
rect 279359 355833 279400 355951
rect 279200 354972 279400 355833
rect 280160 354972 280360 356633
rect 281120 354972 281320 357433
rect 282080 354972 282280 358233
rect 287080 357951 287280 358392
rect 287080 357833 287121 357951
rect 287239 357833 287280 357951
rect 286120 357151 286320 357592
rect 286120 357033 286161 357151
rect 286279 357033 286320 357151
rect 285160 356351 285360 356792
rect 285160 356233 285201 356351
rect 285319 356233 285360 356351
rect 284200 355551 284400 355992
rect 284200 355433 284241 355551
rect 284359 355433 284400 355551
rect 284200 354972 284400 355433
rect 285160 354972 285360 356233
rect 286120 354972 286320 357033
rect 287080 354972 287280 357833
rect 292080 358351 292280 358392
rect 292080 358233 292121 358351
rect 292239 358233 292280 358351
rect 291120 357551 291320 357592
rect 291120 357433 291161 357551
rect 291279 357433 291320 357551
rect 290160 356751 290360 356792
rect 290160 356633 290201 356751
rect 290319 356633 290360 356751
rect 289200 355951 289400 355992
rect 289200 355833 289241 355951
rect 289359 355833 289400 355951
rect 289200 354972 289400 355833
rect 290160 354972 290360 356633
rect 291120 354972 291320 357433
rect 292080 354972 292280 358233
rect 299258 358351 299458 358392
rect 299258 358233 299299 358351
rect 299417 358233 299458 358351
rect 298858 357951 299058 357992
rect 298858 357833 298899 357951
rect 299017 357833 299058 357951
rect 298458 357551 298658 357592
rect 298458 357433 298499 357551
rect 298617 357433 298658 357551
rect 298058 357151 298258 357192
rect 298058 357033 298099 357151
rect 298217 357033 298258 357151
rect 297658 356751 297858 356792
rect 297658 356633 297699 356751
rect 297817 356633 297858 356751
rect 297258 356351 297458 356392
rect 297258 356233 297299 356351
rect 297417 356233 297458 356351
rect 294200 355551 294400 355992
rect 296858 355951 297058 355992
rect 296858 355833 296899 355951
rect 297017 355833 297058 355951
rect 294200 355433 294241 355551
rect 294359 355433 294400 355551
rect 294200 354972 294400 355433
rect 296458 355551 296658 355592
rect 296458 355433 296499 355551
rect 296617 355433 296658 355551
rect 2800 344241 2841 344359
rect 2959 344241 3000 344359
rect 2800 334359 3000 344241
rect 2800 334241 2841 334359
rect 2959 334241 3000 334359
rect 2800 324359 3000 334241
rect 2800 324241 2841 324359
rect 2959 324241 3000 324359
rect 2800 314359 3000 324241
rect 2800 314241 2841 314359
rect 2959 314241 3000 314359
rect 2800 304359 3000 314241
rect 2800 304241 2841 304359
rect 2959 304241 3000 304359
rect 2800 294359 3000 304241
rect 2800 294241 2841 294359
rect 2959 294241 3000 294359
rect 2800 284359 3000 294241
rect 2800 284241 2841 284359
rect 2959 284241 3000 284359
rect 2800 274359 3000 284241
rect 2800 274241 2841 274359
rect 2959 274241 3000 274359
rect 2800 264359 3000 274241
rect 2800 264241 2841 264359
rect 2959 264241 3000 264359
rect 2800 254359 3000 264241
rect 2800 254241 2841 254359
rect 2959 254241 3000 254359
rect 2800 244359 3000 254241
rect 2800 244241 2841 244359
rect 2959 244241 3000 244359
rect 2800 234359 3000 244241
rect 2800 234241 2841 234359
rect 2959 234241 3000 234359
rect 2800 224359 3000 234241
rect 2800 224241 2841 224359
rect 2959 224241 3000 224359
rect 2800 214359 3000 224241
rect 2800 214241 2841 214359
rect 2959 214241 3000 214359
rect 2800 204359 3000 214241
rect 2800 204241 2841 204359
rect 2959 204241 3000 204359
rect 2800 194359 3000 204241
rect 2800 194241 2841 194359
rect 2959 194241 3000 194359
rect 2800 184359 3000 194241
rect 2800 184241 2841 184359
rect 2959 184241 3000 184359
rect 2800 174359 3000 184241
rect 2800 174241 2841 174359
rect 2959 174241 3000 174359
rect 2800 164359 3000 174241
rect 2800 164241 2841 164359
rect 2959 164241 3000 164359
rect 2800 154359 3000 164241
rect 2800 154241 2841 154359
rect 2959 154241 3000 154359
rect 2800 144359 3000 154241
rect 2800 144241 2841 144359
rect 2959 144241 3000 144359
rect 2800 134359 3000 144241
rect 2800 134241 2841 134359
rect 2959 134241 3000 134359
rect 2800 124359 3000 134241
rect 2800 124241 2841 124359
rect 2959 124241 3000 124359
rect 2800 114359 3000 124241
rect 2800 114241 2841 114359
rect 2959 114241 3000 114359
rect 2800 104359 3000 114241
rect 2800 104241 2841 104359
rect 2959 104241 3000 104359
rect 2800 94359 3000 104241
rect 2800 94241 2841 94359
rect 2959 94241 3000 94359
rect 2800 84359 3000 94241
rect 2800 84241 2841 84359
rect 2959 84241 3000 84359
rect 2800 74359 3000 84241
rect 2800 74241 2841 74359
rect 2959 74241 3000 74359
rect 2800 64359 3000 74241
rect 2800 64241 2841 64359
rect 2959 64241 3000 64359
rect 2800 54359 3000 64241
rect 2800 54241 2841 54359
rect 2959 54241 3000 54359
rect 2800 44359 3000 54241
rect 2800 44241 2841 44359
rect 2959 44241 3000 44359
rect 2800 34359 3000 44241
rect 2800 34241 2841 34359
rect 2959 34241 3000 34359
rect 2800 24359 3000 34241
rect 2800 24241 2841 24359
rect 2959 24241 3000 24359
rect 2800 14359 3000 24241
rect 2800 14241 2841 14359
rect 2959 14241 3000 14359
rect 2800 4359 3000 14241
rect 2800 4241 2841 4359
rect 2959 4241 3000 4359
rect 2800 2959 3000 4241
rect 296458 344359 296658 355433
rect 296458 344241 296499 344359
rect 296617 344241 296658 344359
rect 296458 334359 296658 344241
rect 296458 334241 296499 334359
rect 296617 334241 296658 334359
rect 296458 324359 296658 334241
rect 296458 324241 296499 324359
rect 296617 324241 296658 324359
rect 296458 314359 296658 324241
rect 296458 314241 296499 314359
rect 296617 314241 296658 314359
rect 296458 304359 296658 314241
rect 296458 304241 296499 304359
rect 296617 304241 296658 304359
rect 296458 294359 296658 304241
rect 296458 294241 296499 294359
rect 296617 294241 296658 294359
rect 296458 284359 296658 294241
rect 296458 284241 296499 284359
rect 296617 284241 296658 284359
rect 296458 274359 296658 284241
rect 296458 274241 296499 274359
rect 296617 274241 296658 274359
rect 296458 264359 296658 274241
rect 296458 264241 296499 264359
rect 296617 264241 296658 264359
rect 296458 254359 296658 264241
rect 296458 254241 296499 254359
rect 296617 254241 296658 254359
rect 296458 244359 296658 254241
rect 296458 244241 296499 244359
rect 296617 244241 296658 244359
rect 296458 234359 296658 244241
rect 296458 234241 296499 234359
rect 296617 234241 296658 234359
rect 296458 224359 296658 234241
rect 296458 224241 296499 224359
rect 296617 224241 296658 224359
rect 296458 214359 296658 224241
rect 296458 214241 296499 214359
rect 296617 214241 296658 214359
rect 296458 204359 296658 214241
rect 296458 204241 296499 204359
rect 296617 204241 296658 204359
rect 296458 194359 296658 204241
rect 296458 194241 296499 194359
rect 296617 194241 296658 194359
rect 296458 184359 296658 194241
rect 296458 184241 296499 184359
rect 296617 184241 296658 184359
rect 296458 174359 296658 184241
rect 296458 174241 296499 174359
rect 296617 174241 296658 174359
rect 296458 164359 296658 174241
rect 296458 164241 296499 164359
rect 296617 164241 296658 164359
rect 296458 154359 296658 164241
rect 296458 154241 296499 154359
rect 296617 154241 296658 154359
rect 296458 144359 296658 154241
rect 296458 144241 296499 144359
rect 296617 144241 296658 144359
rect 296458 134359 296658 144241
rect 296458 134241 296499 134359
rect 296617 134241 296658 134359
rect 296458 124359 296658 134241
rect 296458 124241 296499 124359
rect 296617 124241 296658 124359
rect 296458 114359 296658 124241
rect 296458 114241 296499 114359
rect 296617 114241 296658 114359
rect 296458 104359 296658 114241
rect 296458 104241 296499 104359
rect 296617 104241 296658 104359
rect 296458 94359 296658 104241
rect 296458 94241 296499 94359
rect 296617 94241 296658 94359
rect 296458 84359 296658 94241
rect 296458 84241 296499 84359
rect 296617 84241 296658 84359
rect 296458 74359 296658 84241
rect 296458 74241 296499 74359
rect 296617 74241 296658 74359
rect 296458 64359 296658 74241
rect 296458 64241 296499 64359
rect 296617 64241 296658 64359
rect 296458 54359 296658 64241
rect 296458 54241 296499 54359
rect 296617 54241 296658 54359
rect 296458 44359 296658 54241
rect 296458 44241 296499 44359
rect 296617 44241 296658 44359
rect 296458 34359 296658 44241
rect 296458 34241 296499 34359
rect 296617 34241 296658 34359
rect 296458 24359 296658 34241
rect 296458 24241 296499 24359
rect 296617 24241 296658 24359
rect 296458 14359 296658 24241
rect 296458 14241 296499 14359
rect 296617 14241 296658 14359
rect 296458 4359 296658 14241
rect 296458 4241 296499 4359
rect 296617 4241 296658 4359
rect 2800 2841 2841 2959
rect 2959 2841 3000 2959
rect 2800 2800 3000 2841
rect 4200 2959 4400 3452
rect 4200 2841 4241 2959
rect 4359 2841 4400 2959
rect 2400 2441 2441 2559
rect 2559 2441 2600 2559
rect 2400 2400 2600 2441
rect 4200 2400 4400 2841
rect 2000 2041 2041 2159
rect 2159 2041 2200 2159
rect 2000 2000 2200 2041
rect 5160 2159 5360 3452
rect 5160 2041 5201 2159
rect 5319 2041 5360 2159
rect 1600 1641 1641 1759
rect 1759 1641 1800 1759
rect 1600 1600 1800 1641
rect 5160 1600 5360 2041
rect 1200 1241 1241 1359
rect 1359 1241 1400 1359
rect 1200 1200 1400 1241
rect 6120 1359 6320 3452
rect 6120 1241 6161 1359
rect 6279 1241 6320 1359
rect 800 841 841 959
rect 959 841 1000 959
rect 800 800 1000 841
rect 6120 800 6320 1241
rect 400 441 441 559
rect 559 441 600 559
rect 400 400 600 441
rect 7080 559 7280 3452
rect 9200 2559 9400 3452
rect 9200 2441 9241 2559
rect 9359 2441 9400 2559
rect 9200 2400 9400 2441
rect 10160 1759 10360 3452
rect 10160 1641 10201 1759
rect 10319 1641 10360 1759
rect 10160 1600 10360 1641
rect 11120 959 11320 3452
rect 11120 841 11161 959
rect 11279 841 11320 959
rect 11120 800 11320 841
rect 7080 441 7121 559
rect 7239 441 7280 559
rect 0 41 41 159
rect 159 41 200 159
rect 0 0 200 41
rect 7080 0 7280 441
rect 12080 159 12280 3452
rect 14200 2959 14400 3452
rect 14200 2841 14241 2959
rect 14359 2841 14400 2959
rect 14200 2400 14400 2841
rect 15160 2159 15360 3452
rect 15160 2041 15201 2159
rect 15319 2041 15360 2159
rect 15160 1600 15360 2041
rect 16120 1359 16320 3452
rect 16120 1241 16161 1359
rect 16279 1241 16320 1359
rect 16120 800 16320 1241
rect 12080 41 12121 159
rect 12239 41 12280 159
rect 12080 0 12280 41
rect 17080 559 17280 3452
rect 19200 2559 19400 3452
rect 19200 2441 19241 2559
rect 19359 2441 19400 2559
rect 19200 2400 19400 2441
rect 20160 1759 20360 3452
rect 20160 1641 20201 1759
rect 20319 1641 20360 1759
rect 20160 1600 20360 1641
rect 21120 959 21320 3452
rect 21120 841 21161 959
rect 21279 841 21320 959
rect 21120 800 21320 841
rect 17080 441 17121 559
rect 17239 441 17280 559
rect 17080 0 17280 441
rect 22080 159 22280 3452
rect 24200 2959 24400 3452
rect 24200 2841 24241 2959
rect 24359 2841 24400 2959
rect 24200 2400 24400 2841
rect 25160 2159 25360 3452
rect 25160 2041 25201 2159
rect 25319 2041 25360 2159
rect 25160 1600 25360 2041
rect 26120 1359 26320 3452
rect 26120 1241 26161 1359
rect 26279 1241 26320 1359
rect 26120 800 26320 1241
rect 22080 41 22121 159
rect 22239 41 22280 159
rect 22080 0 22280 41
rect 27080 559 27280 3452
rect 29200 2559 29400 3452
rect 29200 2441 29241 2559
rect 29359 2441 29400 2559
rect 29200 2400 29400 2441
rect 30160 1759 30360 3452
rect 30160 1641 30201 1759
rect 30319 1641 30360 1759
rect 30160 1600 30360 1641
rect 31120 959 31320 3452
rect 31120 841 31161 959
rect 31279 841 31320 959
rect 31120 800 31320 841
rect 27080 441 27121 559
rect 27239 441 27280 559
rect 27080 0 27280 441
rect 32080 159 32280 3452
rect 34200 2959 34400 3452
rect 34200 2841 34241 2959
rect 34359 2841 34400 2959
rect 34200 2400 34400 2841
rect 35160 2159 35360 3452
rect 35160 2041 35201 2159
rect 35319 2041 35360 2159
rect 35160 1600 35360 2041
rect 36120 1359 36320 3452
rect 36120 1241 36161 1359
rect 36279 1241 36320 1359
rect 36120 800 36320 1241
rect 32080 41 32121 159
rect 32239 41 32280 159
rect 32080 0 32280 41
rect 37080 559 37280 3452
rect 39200 2559 39400 3452
rect 39200 2441 39241 2559
rect 39359 2441 39400 2559
rect 39200 2400 39400 2441
rect 40160 1759 40360 3452
rect 40160 1641 40201 1759
rect 40319 1641 40360 1759
rect 40160 1600 40360 1641
rect 41120 959 41320 3452
rect 41120 841 41161 959
rect 41279 841 41320 959
rect 41120 800 41320 841
rect 37080 441 37121 559
rect 37239 441 37280 559
rect 37080 0 37280 441
rect 42080 159 42280 3452
rect 44200 2959 44400 3452
rect 44200 2841 44241 2959
rect 44359 2841 44400 2959
rect 44200 2400 44400 2841
rect 45160 2159 45360 3452
rect 45160 2041 45201 2159
rect 45319 2041 45360 2159
rect 45160 1600 45360 2041
rect 46120 1359 46320 3452
rect 46120 1241 46161 1359
rect 46279 1241 46320 1359
rect 46120 800 46320 1241
rect 42080 41 42121 159
rect 42239 41 42280 159
rect 42080 0 42280 41
rect 47080 559 47280 3452
rect 49200 2559 49400 3452
rect 49200 2441 49241 2559
rect 49359 2441 49400 2559
rect 49200 2400 49400 2441
rect 50160 1759 50360 3452
rect 50160 1641 50201 1759
rect 50319 1641 50360 1759
rect 50160 1600 50360 1641
rect 51120 959 51320 3452
rect 51120 841 51161 959
rect 51279 841 51320 959
rect 51120 800 51320 841
rect 47080 441 47121 559
rect 47239 441 47280 559
rect 47080 0 47280 441
rect 52080 159 52280 3452
rect 54200 2959 54400 3452
rect 54200 2841 54241 2959
rect 54359 2841 54400 2959
rect 54200 2400 54400 2841
rect 55160 2159 55360 3452
rect 55160 2041 55201 2159
rect 55319 2041 55360 2159
rect 55160 1600 55360 2041
rect 56120 1359 56320 3452
rect 56120 1241 56161 1359
rect 56279 1241 56320 1359
rect 56120 800 56320 1241
rect 52080 41 52121 159
rect 52239 41 52280 159
rect 52080 0 52280 41
rect 57080 559 57280 3452
rect 59200 2559 59400 3452
rect 59200 2441 59241 2559
rect 59359 2441 59400 2559
rect 59200 2400 59400 2441
rect 60160 1759 60360 3452
rect 60160 1641 60201 1759
rect 60319 1641 60360 1759
rect 60160 1600 60360 1641
rect 61120 959 61320 3452
rect 61120 841 61161 959
rect 61279 841 61320 959
rect 61120 800 61320 841
rect 57080 441 57121 559
rect 57239 441 57280 559
rect 57080 0 57280 441
rect 62080 159 62280 3452
rect 64200 2959 64400 3452
rect 64200 2841 64241 2959
rect 64359 2841 64400 2959
rect 64200 2400 64400 2841
rect 65160 2159 65360 3452
rect 65160 2041 65201 2159
rect 65319 2041 65360 2159
rect 65160 1600 65360 2041
rect 66120 1359 66320 3452
rect 66120 1241 66161 1359
rect 66279 1241 66320 1359
rect 66120 800 66320 1241
rect 62080 41 62121 159
rect 62239 41 62280 159
rect 62080 0 62280 41
rect 67080 559 67280 3452
rect 69200 2559 69400 3452
rect 69200 2441 69241 2559
rect 69359 2441 69400 2559
rect 69200 2400 69400 2441
rect 70160 1759 70360 3452
rect 70160 1641 70201 1759
rect 70319 1641 70360 1759
rect 70160 1600 70360 1641
rect 71120 959 71320 3452
rect 71120 841 71161 959
rect 71279 841 71320 959
rect 71120 800 71320 841
rect 67080 441 67121 559
rect 67239 441 67280 559
rect 67080 0 67280 441
rect 72080 159 72280 3452
rect 74200 2959 74400 3452
rect 74200 2841 74241 2959
rect 74359 2841 74400 2959
rect 74200 2400 74400 2841
rect 75160 2159 75360 3452
rect 75160 2041 75201 2159
rect 75319 2041 75360 2159
rect 75160 1600 75360 2041
rect 76120 1359 76320 3452
rect 76120 1241 76161 1359
rect 76279 1241 76320 1359
rect 76120 800 76320 1241
rect 72080 41 72121 159
rect 72239 41 72280 159
rect 72080 0 72280 41
rect 77080 559 77280 3452
rect 79200 2559 79400 3452
rect 79200 2441 79241 2559
rect 79359 2441 79400 2559
rect 79200 2400 79400 2441
rect 80160 1759 80360 3452
rect 80160 1641 80201 1759
rect 80319 1641 80360 1759
rect 80160 1600 80360 1641
rect 81120 959 81320 3452
rect 81120 841 81161 959
rect 81279 841 81320 959
rect 81120 800 81320 841
rect 77080 441 77121 559
rect 77239 441 77280 559
rect 77080 0 77280 441
rect 82080 159 82280 3452
rect 84200 2959 84400 3452
rect 84200 2841 84241 2959
rect 84359 2841 84400 2959
rect 84200 2400 84400 2841
rect 85160 2159 85360 3452
rect 85160 2041 85201 2159
rect 85319 2041 85360 2159
rect 85160 1600 85360 2041
rect 86120 1359 86320 3452
rect 86120 1241 86161 1359
rect 86279 1241 86320 1359
rect 86120 800 86320 1241
rect 82080 41 82121 159
rect 82239 41 82280 159
rect 82080 0 82280 41
rect 87080 559 87280 3452
rect 89200 2559 89400 3452
rect 89200 2441 89241 2559
rect 89359 2441 89400 2559
rect 89200 2400 89400 2441
rect 90160 1759 90360 3452
rect 90160 1641 90201 1759
rect 90319 1641 90360 1759
rect 90160 1600 90360 1641
rect 91120 959 91320 3452
rect 91120 841 91161 959
rect 91279 841 91320 959
rect 91120 800 91320 841
rect 87080 441 87121 559
rect 87239 441 87280 559
rect 87080 0 87280 441
rect 92080 159 92280 3452
rect 94200 2959 94400 3452
rect 94200 2841 94241 2959
rect 94359 2841 94400 2959
rect 94200 2400 94400 2841
rect 95160 2159 95360 3452
rect 95160 2041 95201 2159
rect 95319 2041 95360 2159
rect 95160 1600 95360 2041
rect 96120 1359 96320 3452
rect 96120 1241 96161 1359
rect 96279 1241 96320 1359
rect 96120 800 96320 1241
rect 92080 41 92121 159
rect 92239 41 92280 159
rect 92080 0 92280 41
rect 97080 559 97280 3452
rect 99200 2559 99400 3452
rect 99200 2441 99241 2559
rect 99359 2441 99400 2559
rect 99200 2400 99400 2441
rect 100160 1759 100360 3452
rect 100160 1641 100201 1759
rect 100319 1641 100360 1759
rect 100160 1600 100360 1641
rect 101120 959 101320 3452
rect 101120 841 101161 959
rect 101279 841 101320 959
rect 101120 800 101320 841
rect 97080 441 97121 559
rect 97239 441 97280 559
rect 97080 0 97280 441
rect 102080 159 102280 3452
rect 104200 2959 104400 3452
rect 104200 2841 104241 2959
rect 104359 2841 104400 2959
rect 104200 2400 104400 2841
rect 105160 2159 105360 3452
rect 105160 2041 105201 2159
rect 105319 2041 105360 2159
rect 105160 1600 105360 2041
rect 106120 1359 106320 3452
rect 106120 1241 106161 1359
rect 106279 1241 106320 1359
rect 106120 800 106320 1241
rect 102080 41 102121 159
rect 102239 41 102280 159
rect 102080 0 102280 41
rect 107080 559 107280 3452
rect 109200 2559 109400 3452
rect 109200 2441 109241 2559
rect 109359 2441 109400 2559
rect 109200 2400 109400 2441
rect 110160 1759 110360 3452
rect 110160 1641 110201 1759
rect 110319 1641 110360 1759
rect 110160 1600 110360 1641
rect 111120 959 111320 3452
rect 111120 841 111161 959
rect 111279 841 111320 959
rect 111120 800 111320 841
rect 107080 441 107121 559
rect 107239 441 107280 559
rect 107080 0 107280 441
rect 112080 159 112280 3452
rect 114200 2959 114400 3452
rect 114200 2841 114241 2959
rect 114359 2841 114400 2959
rect 114200 2400 114400 2841
rect 115160 2159 115360 3452
rect 115160 2041 115201 2159
rect 115319 2041 115360 2159
rect 115160 1600 115360 2041
rect 116120 1359 116320 3452
rect 116120 1241 116161 1359
rect 116279 1241 116320 1359
rect 116120 800 116320 1241
rect 112080 41 112121 159
rect 112239 41 112280 159
rect 112080 0 112280 41
rect 117080 559 117280 3452
rect 119200 2559 119400 3452
rect 119200 2441 119241 2559
rect 119359 2441 119400 2559
rect 119200 2400 119400 2441
rect 120160 1759 120360 3452
rect 120160 1641 120201 1759
rect 120319 1641 120360 1759
rect 120160 1600 120360 1641
rect 121120 959 121320 3452
rect 121120 841 121161 959
rect 121279 841 121320 959
rect 121120 800 121320 841
rect 117080 441 117121 559
rect 117239 441 117280 559
rect 117080 0 117280 441
rect 122080 159 122280 3452
rect 124200 2959 124400 3452
rect 124200 2841 124241 2959
rect 124359 2841 124400 2959
rect 124200 2400 124400 2841
rect 125160 2159 125360 3452
rect 125160 2041 125201 2159
rect 125319 2041 125360 2159
rect 125160 1600 125360 2041
rect 126120 1359 126320 3452
rect 126120 1241 126161 1359
rect 126279 1241 126320 1359
rect 126120 800 126320 1241
rect 122080 41 122121 159
rect 122239 41 122280 159
rect 122080 0 122280 41
rect 127080 559 127280 3452
rect 129200 2559 129400 3452
rect 129200 2441 129241 2559
rect 129359 2441 129400 2559
rect 129200 2400 129400 2441
rect 130160 1759 130360 3452
rect 130160 1641 130201 1759
rect 130319 1641 130360 1759
rect 130160 1600 130360 1641
rect 131120 959 131320 3452
rect 131120 841 131161 959
rect 131279 841 131320 959
rect 131120 800 131320 841
rect 127080 441 127121 559
rect 127239 441 127280 559
rect 127080 0 127280 441
rect 132080 159 132280 3452
rect 134200 2959 134400 3452
rect 134200 2841 134241 2959
rect 134359 2841 134400 2959
rect 134200 2400 134400 2841
rect 135160 2159 135360 3452
rect 135160 2041 135201 2159
rect 135319 2041 135360 2159
rect 135160 1600 135360 2041
rect 136120 1359 136320 3452
rect 136120 1241 136161 1359
rect 136279 1241 136320 1359
rect 136120 800 136320 1241
rect 132080 41 132121 159
rect 132239 41 132280 159
rect 132080 0 132280 41
rect 137080 559 137280 3452
rect 139200 2559 139400 3452
rect 139200 2441 139241 2559
rect 139359 2441 139400 2559
rect 139200 2400 139400 2441
rect 140160 1759 140360 3452
rect 140160 1641 140201 1759
rect 140319 1641 140360 1759
rect 140160 1600 140360 1641
rect 141120 959 141320 3452
rect 141120 841 141161 959
rect 141279 841 141320 959
rect 141120 800 141320 841
rect 137080 441 137121 559
rect 137239 441 137280 559
rect 137080 0 137280 441
rect 142080 159 142280 3452
rect 144200 2959 144400 3452
rect 144200 2841 144241 2959
rect 144359 2841 144400 2959
rect 144200 2400 144400 2841
rect 145160 2159 145360 3452
rect 145160 2041 145201 2159
rect 145319 2041 145360 2159
rect 145160 1600 145360 2041
rect 146120 1359 146320 3452
rect 146120 1241 146161 1359
rect 146279 1241 146320 1359
rect 146120 800 146320 1241
rect 142080 41 142121 159
rect 142239 41 142280 159
rect 142080 0 142280 41
rect 147080 559 147280 3452
rect 149200 2559 149400 3452
rect 149200 2441 149241 2559
rect 149359 2441 149400 2559
rect 149200 2400 149400 2441
rect 150160 1759 150360 3452
rect 150160 1641 150201 1759
rect 150319 1641 150360 1759
rect 150160 1600 150360 1641
rect 151120 959 151320 3452
rect 151120 841 151161 959
rect 151279 841 151320 959
rect 151120 800 151320 841
rect 147080 441 147121 559
rect 147239 441 147280 559
rect 147080 0 147280 441
rect 152080 159 152280 3452
rect 154200 2959 154400 3452
rect 154200 2841 154241 2959
rect 154359 2841 154400 2959
rect 154200 2400 154400 2841
rect 155160 2159 155360 3452
rect 155160 2041 155201 2159
rect 155319 2041 155360 2159
rect 155160 1600 155360 2041
rect 156120 1359 156320 3452
rect 156120 1241 156161 1359
rect 156279 1241 156320 1359
rect 156120 800 156320 1241
rect 152080 41 152121 159
rect 152239 41 152280 159
rect 152080 0 152280 41
rect 157080 559 157280 3452
rect 159200 2559 159400 3452
rect 159200 2441 159241 2559
rect 159359 2441 159400 2559
rect 159200 2400 159400 2441
rect 160160 1759 160360 3452
rect 160160 1641 160201 1759
rect 160319 1641 160360 1759
rect 160160 1600 160360 1641
rect 161120 959 161320 3452
rect 161120 841 161161 959
rect 161279 841 161320 959
rect 161120 800 161320 841
rect 157080 441 157121 559
rect 157239 441 157280 559
rect 157080 0 157280 441
rect 162080 159 162280 3452
rect 164200 2959 164400 3452
rect 164200 2841 164241 2959
rect 164359 2841 164400 2959
rect 164200 2400 164400 2841
rect 165160 2159 165360 3452
rect 165160 2041 165201 2159
rect 165319 2041 165360 2159
rect 165160 1600 165360 2041
rect 166120 1359 166320 3452
rect 166120 1241 166161 1359
rect 166279 1241 166320 1359
rect 166120 800 166320 1241
rect 162080 41 162121 159
rect 162239 41 162280 159
rect 162080 0 162280 41
rect 167080 559 167280 3452
rect 169200 2559 169400 3452
rect 169200 2441 169241 2559
rect 169359 2441 169400 2559
rect 169200 2400 169400 2441
rect 170160 1759 170360 3452
rect 170160 1641 170201 1759
rect 170319 1641 170360 1759
rect 170160 1600 170360 1641
rect 171120 959 171320 3452
rect 171120 841 171161 959
rect 171279 841 171320 959
rect 171120 800 171320 841
rect 167080 441 167121 559
rect 167239 441 167280 559
rect 167080 0 167280 441
rect 172080 159 172280 3452
rect 174200 2959 174400 3452
rect 174200 2841 174241 2959
rect 174359 2841 174400 2959
rect 174200 2400 174400 2841
rect 175160 2159 175360 3452
rect 175160 2041 175201 2159
rect 175319 2041 175360 2159
rect 175160 1600 175360 2041
rect 176120 1359 176320 3452
rect 176120 1241 176161 1359
rect 176279 1241 176320 1359
rect 176120 800 176320 1241
rect 172080 41 172121 159
rect 172239 41 172280 159
rect 172080 0 172280 41
rect 177080 559 177280 3452
rect 179200 2559 179400 3452
rect 179200 2441 179241 2559
rect 179359 2441 179400 2559
rect 179200 2400 179400 2441
rect 180160 1759 180360 3452
rect 180160 1641 180201 1759
rect 180319 1641 180360 1759
rect 180160 1600 180360 1641
rect 181120 959 181320 3452
rect 181120 841 181161 959
rect 181279 841 181320 959
rect 181120 800 181320 841
rect 177080 441 177121 559
rect 177239 441 177280 559
rect 177080 0 177280 441
rect 182080 159 182280 3452
rect 184200 2959 184400 3452
rect 184200 2841 184241 2959
rect 184359 2841 184400 2959
rect 184200 2400 184400 2841
rect 185160 2159 185360 3452
rect 185160 2041 185201 2159
rect 185319 2041 185360 2159
rect 185160 1600 185360 2041
rect 186120 1359 186320 3452
rect 186120 1241 186161 1359
rect 186279 1241 186320 1359
rect 186120 800 186320 1241
rect 182080 41 182121 159
rect 182239 41 182280 159
rect 182080 0 182280 41
rect 187080 559 187280 3452
rect 189200 2559 189400 3452
rect 189200 2441 189241 2559
rect 189359 2441 189400 2559
rect 189200 2400 189400 2441
rect 190160 1759 190360 3452
rect 190160 1641 190201 1759
rect 190319 1641 190360 1759
rect 190160 1600 190360 1641
rect 191120 959 191320 3452
rect 191120 841 191161 959
rect 191279 841 191320 959
rect 191120 800 191320 841
rect 187080 441 187121 559
rect 187239 441 187280 559
rect 187080 0 187280 441
rect 192080 159 192280 3452
rect 194200 2959 194400 3452
rect 194200 2841 194241 2959
rect 194359 2841 194400 2959
rect 194200 2400 194400 2841
rect 195160 2159 195360 3452
rect 195160 2041 195201 2159
rect 195319 2041 195360 2159
rect 195160 1600 195360 2041
rect 196120 1359 196320 3452
rect 196120 1241 196161 1359
rect 196279 1241 196320 1359
rect 196120 800 196320 1241
rect 192080 41 192121 159
rect 192239 41 192280 159
rect 192080 0 192280 41
rect 197080 559 197280 3452
rect 199200 2559 199400 3452
rect 199200 2441 199241 2559
rect 199359 2441 199400 2559
rect 199200 2400 199400 2441
rect 200160 1759 200360 3452
rect 200160 1641 200201 1759
rect 200319 1641 200360 1759
rect 200160 1600 200360 1641
rect 201120 959 201320 3452
rect 201120 841 201161 959
rect 201279 841 201320 959
rect 201120 800 201320 841
rect 197080 441 197121 559
rect 197239 441 197280 559
rect 197080 0 197280 441
rect 202080 159 202280 3452
rect 204200 2959 204400 3452
rect 204200 2841 204241 2959
rect 204359 2841 204400 2959
rect 204200 2400 204400 2841
rect 205160 2159 205360 3452
rect 205160 2041 205201 2159
rect 205319 2041 205360 2159
rect 205160 1600 205360 2041
rect 206120 1359 206320 3452
rect 206120 1241 206161 1359
rect 206279 1241 206320 1359
rect 206120 800 206320 1241
rect 202080 41 202121 159
rect 202239 41 202280 159
rect 202080 0 202280 41
rect 207080 559 207280 3452
rect 209200 2559 209400 3452
rect 209200 2441 209241 2559
rect 209359 2441 209400 2559
rect 209200 2400 209400 2441
rect 210160 1759 210360 3452
rect 210160 1641 210201 1759
rect 210319 1641 210360 1759
rect 210160 1600 210360 1641
rect 211120 959 211320 3452
rect 211120 841 211161 959
rect 211279 841 211320 959
rect 211120 800 211320 841
rect 207080 441 207121 559
rect 207239 441 207280 559
rect 207080 0 207280 441
rect 212080 159 212280 3452
rect 214200 2959 214400 3452
rect 214200 2841 214241 2959
rect 214359 2841 214400 2959
rect 214200 2400 214400 2841
rect 215160 2159 215360 3452
rect 215160 2041 215201 2159
rect 215319 2041 215360 2159
rect 215160 1600 215360 2041
rect 216120 1359 216320 3452
rect 216120 1241 216161 1359
rect 216279 1241 216320 1359
rect 216120 800 216320 1241
rect 212080 41 212121 159
rect 212239 41 212280 159
rect 212080 0 212280 41
rect 217080 559 217280 3452
rect 219200 2559 219400 3452
rect 219200 2441 219241 2559
rect 219359 2441 219400 2559
rect 219200 2400 219400 2441
rect 220160 1759 220360 3452
rect 220160 1641 220201 1759
rect 220319 1641 220360 1759
rect 220160 1600 220360 1641
rect 221120 959 221320 3452
rect 221120 841 221161 959
rect 221279 841 221320 959
rect 221120 800 221320 841
rect 217080 441 217121 559
rect 217239 441 217280 559
rect 217080 0 217280 441
rect 222080 159 222280 3452
rect 224200 2959 224400 3452
rect 224200 2841 224241 2959
rect 224359 2841 224400 2959
rect 224200 2400 224400 2841
rect 225160 2159 225360 3452
rect 225160 2041 225201 2159
rect 225319 2041 225360 2159
rect 225160 1600 225360 2041
rect 226120 1359 226320 3452
rect 226120 1241 226161 1359
rect 226279 1241 226320 1359
rect 226120 800 226320 1241
rect 222080 41 222121 159
rect 222239 41 222280 159
rect 222080 0 222280 41
rect 227080 559 227280 3452
rect 229200 2559 229400 3452
rect 229200 2441 229241 2559
rect 229359 2441 229400 2559
rect 229200 2400 229400 2441
rect 230160 1759 230360 3452
rect 230160 1641 230201 1759
rect 230319 1641 230360 1759
rect 230160 1600 230360 1641
rect 231120 959 231320 3452
rect 231120 841 231161 959
rect 231279 841 231320 959
rect 231120 800 231320 841
rect 227080 441 227121 559
rect 227239 441 227280 559
rect 227080 0 227280 441
rect 232080 159 232280 3452
rect 234200 2959 234400 3452
rect 234200 2841 234241 2959
rect 234359 2841 234400 2959
rect 234200 2400 234400 2841
rect 235160 2159 235360 3452
rect 235160 2041 235201 2159
rect 235319 2041 235360 2159
rect 235160 1600 235360 2041
rect 236120 1359 236320 3452
rect 236120 1241 236161 1359
rect 236279 1241 236320 1359
rect 236120 800 236320 1241
rect 232080 41 232121 159
rect 232239 41 232280 159
rect 232080 0 232280 41
rect 237080 559 237280 3452
rect 239200 2559 239400 3452
rect 239200 2441 239241 2559
rect 239359 2441 239400 2559
rect 239200 2400 239400 2441
rect 240160 1759 240360 3452
rect 240160 1641 240201 1759
rect 240319 1641 240360 1759
rect 240160 1600 240360 1641
rect 241120 959 241320 3452
rect 241120 841 241161 959
rect 241279 841 241320 959
rect 241120 800 241320 841
rect 237080 441 237121 559
rect 237239 441 237280 559
rect 237080 0 237280 441
rect 242080 159 242280 3452
rect 244200 2959 244400 3452
rect 244200 2841 244241 2959
rect 244359 2841 244400 2959
rect 244200 2400 244400 2841
rect 245160 2159 245360 3452
rect 245160 2041 245201 2159
rect 245319 2041 245360 2159
rect 245160 1600 245360 2041
rect 246120 1359 246320 3452
rect 246120 1241 246161 1359
rect 246279 1241 246320 1359
rect 246120 800 246320 1241
rect 242080 41 242121 159
rect 242239 41 242280 159
rect 242080 0 242280 41
rect 247080 559 247280 3452
rect 249200 2559 249400 3452
rect 249200 2441 249241 2559
rect 249359 2441 249400 2559
rect 249200 2400 249400 2441
rect 250160 1759 250360 3452
rect 250160 1641 250201 1759
rect 250319 1641 250360 1759
rect 250160 1600 250360 1641
rect 251120 959 251320 3452
rect 251120 841 251161 959
rect 251279 841 251320 959
rect 251120 800 251320 841
rect 247080 441 247121 559
rect 247239 441 247280 559
rect 247080 0 247280 441
rect 252080 159 252280 3452
rect 254200 2959 254400 3452
rect 254200 2841 254241 2959
rect 254359 2841 254400 2959
rect 254200 2400 254400 2841
rect 255160 2159 255360 3452
rect 255160 2041 255201 2159
rect 255319 2041 255360 2159
rect 255160 1600 255360 2041
rect 256120 1359 256320 3452
rect 256120 1241 256161 1359
rect 256279 1241 256320 1359
rect 256120 800 256320 1241
rect 252080 41 252121 159
rect 252239 41 252280 159
rect 252080 0 252280 41
rect 257080 559 257280 3452
rect 259200 2559 259400 3452
rect 259200 2441 259241 2559
rect 259359 2441 259400 2559
rect 259200 2400 259400 2441
rect 260160 1759 260360 3452
rect 260160 1641 260201 1759
rect 260319 1641 260360 1759
rect 260160 1600 260360 1641
rect 261120 959 261320 3452
rect 261120 841 261161 959
rect 261279 841 261320 959
rect 261120 800 261320 841
rect 257080 441 257121 559
rect 257239 441 257280 559
rect 257080 0 257280 441
rect 262080 159 262280 3452
rect 264200 2959 264400 3452
rect 264200 2841 264241 2959
rect 264359 2841 264400 2959
rect 264200 2400 264400 2841
rect 265160 2159 265360 3452
rect 265160 2041 265201 2159
rect 265319 2041 265360 2159
rect 265160 1600 265360 2041
rect 266120 1359 266320 3452
rect 266120 1241 266161 1359
rect 266279 1241 266320 1359
rect 266120 800 266320 1241
rect 262080 41 262121 159
rect 262239 41 262280 159
rect 262080 0 262280 41
rect 267080 559 267280 3452
rect 269200 2559 269400 3452
rect 269200 2441 269241 2559
rect 269359 2441 269400 2559
rect 269200 2400 269400 2441
rect 270160 1759 270360 3452
rect 270160 1641 270201 1759
rect 270319 1641 270360 1759
rect 270160 1600 270360 1641
rect 271120 959 271320 3452
rect 271120 841 271161 959
rect 271279 841 271320 959
rect 271120 800 271320 841
rect 267080 441 267121 559
rect 267239 441 267280 559
rect 267080 0 267280 441
rect 272080 159 272280 3452
rect 274200 2959 274400 3452
rect 274200 2841 274241 2959
rect 274359 2841 274400 2959
rect 274200 2400 274400 2841
rect 275160 2159 275360 3452
rect 275160 2041 275201 2159
rect 275319 2041 275360 2159
rect 275160 1600 275360 2041
rect 276120 1359 276320 3452
rect 276120 1241 276161 1359
rect 276279 1241 276320 1359
rect 276120 800 276320 1241
rect 272080 41 272121 159
rect 272239 41 272280 159
rect 272080 0 272280 41
rect 277080 559 277280 3452
rect 279200 2559 279400 3452
rect 279200 2441 279241 2559
rect 279359 2441 279400 2559
rect 279200 2400 279400 2441
rect 280160 1759 280360 3452
rect 280160 1641 280201 1759
rect 280319 1641 280360 1759
rect 280160 1600 280360 1641
rect 281120 959 281320 3452
rect 281120 841 281161 959
rect 281279 841 281320 959
rect 281120 800 281320 841
rect 277080 441 277121 559
rect 277239 441 277280 559
rect 277080 0 277280 441
rect 282080 159 282280 3452
rect 284200 2959 284400 3452
rect 284200 2841 284241 2959
rect 284359 2841 284400 2959
rect 284200 2400 284400 2841
rect 285160 2159 285360 3452
rect 285160 2041 285201 2159
rect 285319 2041 285360 2159
rect 285160 1600 285360 2041
rect 286120 1359 286320 3452
rect 286120 1241 286161 1359
rect 286279 1241 286320 1359
rect 286120 800 286320 1241
rect 282080 41 282121 159
rect 282239 41 282280 159
rect 282080 0 282280 41
rect 287080 559 287280 3452
rect 289200 2559 289400 3452
rect 289200 2441 289241 2559
rect 289359 2441 289400 2559
rect 289200 2400 289400 2441
rect 290160 1759 290360 3452
rect 290160 1641 290201 1759
rect 290319 1641 290360 1759
rect 290160 1600 290360 1641
rect 291120 959 291320 3452
rect 291120 841 291161 959
rect 291279 841 291320 959
rect 291120 800 291320 841
rect 287080 441 287121 559
rect 287239 441 287280 559
rect 287080 0 287280 441
rect 292080 159 292280 3452
rect 294200 2959 294400 3452
rect 294200 2841 294241 2959
rect 294359 2841 294400 2959
rect 294200 2400 294400 2841
rect 296458 2959 296658 4241
rect 296458 2841 296499 2959
rect 296617 2841 296658 2959
rect 296458 2800 296658 2841
rect 296858 349359 297058 355833
rect 296858 349241 296899 349359
rect 297017 349241 297058 349359
rect 296858 339359 297058 349241
rect 296858 339241 296899 339359
rect 297017 339241 297058 339359
rect 296858 329359 297058 339241
rect 296858 329241 296899 329359
rect 297017 329241 297058 329359
rect 296858 319359 297058 329241
rect 296858 319241 296899 319359
rect 297017 319241 297058 319359
rect 296858 309359 297058 319241
rect 296858 309241 296899 309359
rect 297017 309241 297058 309359
rect 296858 299359 297058 309241
rect 296858 299241 296899 299359
rect 297017 299241 297058 299359
rect 296858 289359 297058 299241
rect 296858 289241 296899 289359
rect 297017 289241 297058 289359
rect 296858 279359 297058 289241
rect 296858 279241 296899 279359
rect 297017 279241 297058 279359
rect 296858 269359 297058 279241
rect 296858 269241 296899 269359
rect 297017 269241 297058 269359
rect 296858 259359 297058 269241
rect 296858 259241 296899 259359
rect 297017 259241 297058 259359
rect 296858 249359 297058 259241
rect 296858 249241 296899 249359
rect 297017 249241 297058 249359
rect 296858 239359 297058 249241
rect 296858 239241 296899 239359
rect 297017 239241 297058 239359
rect 296858 229359 297058 239241
rect 296858 229241 296899 229359
rect 297017 229241 297058 229359
rect 296858 219359 297058 229241
rect 296858 219241 296899 219359
rect 297017 219241 297058 219359
rect 296858 209359 297058 219241
rect 296858 209241 296899 209359
rect 297017 209241 297058 209359
rect 296858 199359 297058 209241
rect 296858 199241 296899 199359
rect 297017 199241 297058 199359
rect 296858 189359 297058 199241
rect 296858 189241 296899 189359
rect 297017 189241 297058 189359
rect 296858 179359 297058 189241
rect 296858 179241 296899 179359
rect 297017 179241 297058 179359
rect 296858 169359 297058 179241
rect 296858 169241 296899 169359
rect 297017 169241 297058 169359
rect 296858 159359 297058 169241
rect 296858 159241 296899 159359
rect 297017 159241 297058 159359
rect 296858 149359 297058 159241
rect 296858 149241 296899 149359
rect 297017 149241 297058 149359
rect 296858 139359 297058 149241
rect 296858 139241 296899 139359
rect 297017 139241 297058 139359
rect 296858 129359 297058 139241
rect 296858 129241 296899 129359
rect 297017 129241 297058 129359
rect 296858 119359 297058 129241
rect 296858 119241 296899 119359
rect 297017 119241 297058 119359
rect 296858 109359 297058 119241
rect 296858 109241 296899 109359
rect 297017 109241 297058 109359
rect 296858 99359 297058 109241
rect 296858 99241 296899 99359
rect 297017 99241 297058 99359
rect 296858 89359 297058 99241
rect 296858 89241 296899 89359
rect 297017 89241 297058 89359
rect 296858 79359 297058 89241
rect 296858 79241 296899 79359
rect 297017 79241 297058 79359
rect 296858 69359 297058 79241
rect 296858 69241 296899 69359
rect 297017 69241 297058 69359
rect 296858 59359 297058 69241
rect 296858 59241 296899 59359
rect 297017 59241 297058 59359
rect 296858 49359 297058 59241
rect 296858 49241 296899 49359
rect 297017 49241 297058 49359
rect 296858 39359 297058 49241
rect 296858 39241 296899 39359
rect 297017 39241 297058 39359
rect 296858 29359 297058 39241
rect 296858 29241 296899 29359
rect 297017 29241 297058 29359
rect 296858 19359 297058 29241
rect 296858 19241 296899 19359
rect 297017 19241 297058 19359
rect 296858 9359 297058 19241
rect 296858 9241 296899 9359
rect 297017 9241 297058 9359
rect 296858 2559 297058 9241
rect 296858 2441 296899 2559
rect 297017 2441 297058 2559
rect 296858 2400 297058 2441
rect 297258 345319 297458 356233
rect 297258 345201 297299 345319
rect 297417 345201 297458 345319
rect 297258 335319 297458 345201
rect 297258 335201 297299 335319
rect 297417 335201 297458 335319
rect 297258 325319 297458 335201
rect 297258 325201 297299 325319
rect 297417 325201 297458 325319
rect 297258 315319 297458 325201
rect 297258 315201 297299 315319
rect 297417 315201 297458 315319
rect 297258 305319 297458 315201
rect 297258 305201 297299 305319
rect 297417 305201 297458 305319
rect 297258 295319 297458 305201
rect 297258 295201 297299 295319
rect 297417 295201 297458 295319
rect 297258 285319 297458 295201
rect 297258 285201 297299 285319
rect 297417 285201 297458 285319
rect 297258 275319 297458 285201
rect 297258 275201 297299 275319
rect 297417 275201 297458 275319
rect 297258 265319 297458 275201
rect 297258 265201 297299 265319
rect 297417 265201 297458 265319
rect 297258 255319 297458 265201
rect 297258 255201 297299 255319
rect 297417 255201 297458 255319
rect 297258 245319 297458 255201
rect 297258 245201 297299 245319
rect 297417 245201 297458 245319
rect 297258 235319 297458 245201
rect 297258 235201 297299 235319
rect 297417 235201 297458 235319
rect 297258 225319 297458 235201
rect 297258 225201 297299 225319
rect 297417 225201 297458 225319
rect 297258 215319 297458 225201
rect 297258 215201 297299 215319
rect 297417 215201 297458 215319
rect 297258 205319 297458 215201
rect 297258 205201 297299 205319
rect 297417 205201 297458 205319
rect 297258 195319 297458 205201
rect 297258 195201 297299 195319
rect 297417 195201 297458 195319
rect 297258 185319 297458 195201
rect 297258 185201 297299 185319
rect 297417 185201 297458 185319
rect 297258 175319 297458 185201
rect 297258 175201 297299 175319
rect 297417 175201 297458 175319
rect 297258 165319 297458 175201
rect 297258 165201 297299 165319
rect 297417 165201 297458 165319
rect 297258 155319 297458 165201
rect 297258 155201 297299 155319
rect 297417 155201 297458 155319
rect 297258 145319 297458 155201
rect 297258 145201 297299 145319
rect 297417 145201 297458 145319
rect 297258 135319 297458 145201
rect 297258 135201 297299 135319
rect 297417 135201 297458 135319
rect 297258 125319 297458 135201
rect 297258 125201 297299 125319
rect 297417 125201 297458 125319
rect 297258 115319 297458 125201
rect 297258 115201 297299 115319
rect 297417 115201 297458 115319
rect 297258 105319 297458 115201
rect 297258 105201 297299 105319
rect 297417 105201 297458 105319
rect 297258 95319 297458 105201
rect 297258 95201 297299 95319
rect 297417 95201 297458 95319
rect 297258 85319 297458 95201
rect 297258 85201 297299 85319
rect 297417 85201 297458 85319
rect 297258 75319 297458 85201
rect 297258 75201 297299 75319
rect 297417 75201 297458 75319
rect 297258 65319 297458 75201
rect 297258 65201 297299 65319
rect 297417 65201 297458 65319
rect 297258 55319 297458 65201
rect 297258 55201 297299 55319
rect 297417 55201 297458 55319
rect 297258 45319 297458 55201
rect 297258 45201 297299 45319
rect 297417 45201 297458 45319
rect 297258 35319 297458 45201
rect 297258 35201 297299 35319
rect 297417 35201 297458 35319
rect 297258 25319 297458 35201
rect 297258 25201 297299 25319
rect 297417 25201 297458 25319
rect 297258 15319 297458 25201
rect 297258 15201 297299 15319
rect 297417 15201 297458 15319
rect 297258 5319 297458 15201
rect 297258 5201 297299 5319
rect 297417 5201 297458 5319
rect 297258 2159 297458 5201
rect 297258 2041 297299 2159
rect 297417 2041 297458 2159
rect 297258 2000 297458 2041
rect 297658 350319 297858 356633
rect 297658 350201 297699 350319
rect 297817 350201 297858 350319
rect 297658 340319 297858 350201
rect 297658 340201 297699 340319
rect 297817 340201 297858 340319
rect 297658 330319 297858 340201
rect 297658 330201 297699 330319
rect 297817 330201 297858 330319
rect 297658 320319 297858 330201
rect 297658 320201 297699 320319
rect 297817 320201 297858 320319
rect 297658 310319 297858 320201
rect 297658 310201 297699 310319
rect 297817 310201 297858 310319
rect 297658 300319 297858 310201
rect 297658 300201 297699 300319
rect 297817 300201 297858 300319
rect 297658 290319 297858 300201
rect 297658 290201 297699 290319
rect 297817 290201 297858 290319
rect 297658 280319 297858 290201
rect 297658 280201 297699 280319
rect 297817 280201 297858 280319
rect 297658 270319 297858 280201
rect 297658 270201 297699 270319
rect 297817 270201 297858 270319
rect 297658 260319 297858 270201
rect 297658 260201 297699 260319
rect 297817 260201 297858 260319
rect 297658 250319 297858 260201
rect 297658 250201 297699 250319
rect 297817 250201 297858 250319
rect 297658 240319 297858 250201
rect 297658 240201 297699 240319
rect 297817 240201 297858 240319
rect 297658 230319 297858 240201
rect 297658 230201 297699 230319
rect 297817 230201 297858 230319
rect 297658 220319 297858 230201
rect 297658 220201 297699 220319
rect 297817 220201 297858 220319
rect 297658 210319 297858 220201
rect 297658 210201 297699 210319
rect 297817 210201 297858 210319
rect 297658 200319 297858 210201
rect 297658 200201 297699 200319
rect 297817 200201 297858 200319
rect 297658 190319 297858 200201
rect 297658 190201 297699 190319
rect 297817 190201 297858 190319
rect 297658 180319 297858 190201
rect 297658 180201 297699 180319
rect 297817 180201 297858 180319
rect 297658 170319 297858 180201
rect 297658 170201 297699 170319
rect 297817 170201 297858 170319
rect 297658 160319 297858 170201
rect 297658 160201 297699 160319
rect 297817 160201 297858 160319
rect 297658 150319 297858 160201
rect 297658 150201 297699 150319
rect 297817 150201 297858 150319
rect 297658 140319 297858 150201
rect 297658 140201 297699 140319
rect 297817 140201 297858 140319
rect 297658 130319 297858 140201
rect 297658 130201 297699 130319
rect 297817 130201 297858 130319
rect 297658 120319 297858 130201
rect 297658 120201 297699 120319
rect 297817 120201 297858 120319
rect 297658 110319 297858 120201
rect 297658 110201 297699 110319
rect 297817 110201 297858 110319
rect 297658 100319 297858 110201
rect 297658 100201 297699 100319
rect 297817 100201 297858 100319
rect 297658 90319 297858 100201
rect 297658 90201 297699 90319
rect 297817 90201 297858 90319
rect 297658 80319 297858 90201
rect 297658 80201 297699 80319
rect 297817 80201 297858 80319
rect 297658 70319 297858 80201
rect 297658 70201 297699 70319
rect 297817 70201 297858 70319
rect 297658 60319 297858 70201
rect 297658 60201 297699 60319
rect 297817 60201 297858 60319
rect 297658 50319 297858 60201
rect 297658 50201 297699 50319
rect 297817 50201 297858 50319
rect 297658 40319 297858 50201
rect 297658 40201 297699 40319
rect 297817 40201 297858 40319
rect 297658 30319 297858 40201
rect 297658 30201 297699 30319
rect 297817 30201 297858 30319
rect 297658 20319 297858 30201
rect 297658 20201 297699 20319
rect 297817 20201 297858 20319
rect 297658 10319 297858 20201
rect 297658 10201 297699 10319
rect 297817 10201 297858 10319
rect 297658 1759 297858 10201
rect 297658 1641 297699 1759
rect 297817 1641 297858 1759
rect 297658 1600 297858 1641
rect 298058 346279 298258 357033
rect 298058 346161 298099 346279
rect 298217 346161 298258 346279
rect 298058 336279 298258 346161
rect 298058 336161 298099 336279
rect 298217 336161 298258 336279
rect 298058 326279 298258 336161
rect 298058 326161 298099 326279
rect 298217 326161 298258 326279
rect 298058 316279 298258 326161
rect 298058 316161 298099 316279
rect 298217 316161 298258 316279
rect 298058 306279 298258 316161
rect 298058 306161 298099 306279
rect 298217 306161 298258 306279
rect 298058 296279 298258 306161
rect 298058 296161 298099 296279
rect 298217 296161 298258 296279
rect 298058 286279 298258 296161
rect 298058 286161 298099 286279
rect 298217 286161 298258 286279
rect 298058 276279 298258 286161
rect 298058 276161 298099 276279
rect 298217 276161 298258 276279
rect 298058 266279 298258 276161
rect 298058 266161 298099 266279
rect 298217 266161 298258 266279
rect 298058 256279 298258 266161
rect 298058 256161 298099 256279
rect 298217 256161 298258 256279
rect 298058 246279 298258 256161
rect 298058 246161 298099 246279
rect 298217 246161 298258 246279
rect 298058 236279 298258 246161
rect 298058 236161 298099 236279
rect 298217 236161 298258 236279
rect 298058 226279 298258 236161
rect 298058 226161 298099 226279
rect 298217 226161 298258 226279
rect 298058 216279 298258 226161
rect 298058 216161 298099 216279
rect 298217 216161 298258 216279
rect 298058 206279 298258 216161
rect 298058 206161 298099 206279
rect 298217 206161 298258 206279
rect 298058 196279 298258 206161
rect 298058 196161 298099 196279
rect 298217 196161 298258 196279
rect 298058 186279 298258 196161
rect 298058 186161 298099 186279
rect 298217 186161 298258 186279
rect 298058 176279 298258 186161
rect 298058 176161 298099 176279
rect 298217 176161 298258 176279
rect 298058 166279 298258 176161
rect 298058 166161 298099 166279
rect 298217 166161 298258 166279
rect 298058 156279 298258 166161
rect 298058 156161 298099 156279
rect 298217 156161 298258 156279
rect 298058 146279 298258 156161
rect 298058 146161 298099 146279
rect 298217 146161 298258 146279
rect 298058 136279 298258 146161
rect 298058 136161 298099 136279
rect 298217 136161 298258 136279
rect 298058 126279 298258 136161
rect 298058 126161 298099 126279
rect 298217 126161 298258 126279
rect 298058 116279 298258 126161
rect 298058 116161 298099 116279
rect 298217 116161 298258 116279
rect 298058 106279 298258 116161
rect 298058 106161 298099 106279
rect 298217 106161 298258 106279
rect 298058 96279 298258 106161
rect 298058 96161 298099 96279
rect 298217 96161 298258 96279
rect 298058 86279 298258 96161
rect 298058 86161 298099 86279
rect 298217 86161 298258 86279
rect 298058 76279 298258 86161
rect 298058 76161 298099 76279
rect 298217 76161 298258 76279
rect 298058 66279 298258 76161
rect 298058 66161 298099 66279
rect 298217 66161 298258 66279
rect 298058 56279 298258 66161
rect 298058 56161 298099 56279
rect 298217 56161 298258 56279
rect 298058 46279 298258 56161
rect 298058 46161 298099 46279
rect 298217 46161 298258 46279
rect 298058 36279 298258 46161
rect 298058 36161 298099 36279
rect 298217 36161 298258 36279
rect 298058 26279 298258 36161
rect 298058 26161 298099 26279
rect 298217 26161 298258 26279
rect 298058 16279 298258 26161
rect 298058 16161 298099 16279
rect 298217 16161 298258 16279
rect 298058 6279 298258 16161
rect 298058 6161 298099 6279
rect 298217 6161 298258 6279
rect 298058 1359 298258 6161
rect 298058 1241 298099 1359
rect 298217 1241 298258 1359
rect 298058 1200 298258 1241
rect 298458 351279 298658 357433
rect 298458 351161 298499 351279
rect 298617 351161 298658 351279
rect 298458 341279 298658 351161
rect 298458 341161 298499 341279
rect 298617 341161 298658 341279
rect 298458 331279 298658 341161
rect 298458 331161 298499 331279
rect 298617 331161 298658 331279
rect 298458 321279 298658 331161
rect 298458 321161 298499 321279
rect 298617 321161 298658 321279
rect 298458 311279 298658 321161
rect 298458 311161 298499 311279
rect 298617 311161 298658 311279
rect 298458 301279 298658 311161
rect 298458 301161 298499 301279
rect 298617 301161 298658 301279
rect 298458 291279 298658 301161
rect 298458 291161 298499 291279
rect 298617 291161 298658 291279
rect 298458 281279 298658 291161
rect 298458 281161 298499 281279
rect 298617 281161 298658 281279
rect 298458 271279 298658 281161
rect 298458 271161 298499 271279
rect 298617 271161 298658 271279
rect 298458 261279 298658 271161
rect 298458 261161 298499 261279
rect 298617 261161 298658 261279
rect 298458 251279 298658 261161
rect 298458 251161 298499 251279
rect 298617 251161 298658 251279
rect 298458 241279 298658 251161
rect 298458 241161 298499 241279
rect 298617 241161 298658 241279
rect 298458 231279 298658 241161
rect 298458 231161 298499 231279
rect 298617 231161 298658 231279
rect 298458 221279 298658 231161
rect 298458 221161 298499 221279
rect 298617 221161 298658 221279
rect 298458 211279 298658 221161
rect 298458 211161 298499 211279
rect 298617 211161 298658 211279
rect 298458 201279 298658 211161
rect 298458 201161 298499 201279
rect 298617 201161 298658 201279
rect 298458 191279 298658 201161
rect 298458 191161 298499 191279
rect 298617 191161 298658 191279
rect 298458 181279 298658 191161
rect 298458 181161 298499 181279
rect 298617 181161 298658 181279
rect 298458 171279 298658 181161
rect 298458 171161 298499 171279
rect 298617 171161 298658 171279
rect 298458 161279 298658 171161
rect 298458 161161 298499 161279
rect 298617 161161 298658 161279
rect 298458 151279 298658 161161
rect 298458 151161 298499 151279
rect 298617 151161 298658 151279
rect 298458 141279 298658 151161
rect 298458 141161 298499 141279
rect 298617 141161 298658 141279
rect 298458 131279 298658 141161
rect 298458 131161 298499 131279
rect 298617 131161 298658 131279
rect 298458 121279 298658 131161
rect 298458 121161 298499 121279
rect 298617 121161 298658 121279
rect 298458 111279 298658 121161
rect 298458 111161 298499 111279
rect 298617 111161 298658 111279
rect 298458 101279 298658 111161
rect 298458 101161 298499 101279
rect 298617 101161 298658 101279
rect 298458 91279 298658 101161
rect 298458 91161 298499 91279
rect 298617 91161 298658 91279
rect 298458 81279 298658 91161
rect 298458 81161 298499 81279
rect 298617 81161 298658 81279
rect 298458 71279 298658 81161
rect 298458 71161 298499 71279
rect 298617 71161 298658 71279
rect 298458 61279 298658 71161
rect 298458 61161 298499 61279
rect 298617 61161 298658 61279
rect 298458 51279 298658 61161
rect 298458 51161 298499 51279
rect 298617 51161 298658 51279
rect 298458 41279 298658 51161
rect 298458 41161 298499 41279
rect 298617 41161 298658 41279
rect 298458 31279 298658 41161
rect 298458 31161 298499 31279
rect 298617 31161 298658 31279
rect 298458 21279 298658 31161
rect 298458 21161 298499 21279
rect 298617 21161 298658 21279
rect 298458 11279 298658 21161
rect 298458 11161 298499 11279
rect 298617 11161 298658 11279
rect 298458 959 298658 11161
rect 298458 841 298499 959
rect 298617 841 298658 959
rect 298458 800 298658 841
rect 298858 347239 299058 357833
rect 298858 347121 298899 347239
rect 299017 347121 299058 347239
rect 298858 337239 299058 347121
rect 298858 337121 298899 337239
rect 299017 337121 299058 337239
rect 298858 327239 299058 337121
rect 298858 327121 298899 327239
rect 299017 327121 299058 327239
rect 298858 317239 299058 327121
rect 298858 317121 298899 317239
rect 299017 317121 299058 317239
rect 298858 307239 299058 317121
rect 298858 307121 298899 307239
rect 299017 307121 299058 307239
rect 298858 297239 299058 307121
rect 298858 297121 298899 297239
rect 299017 297121 299058 297239
rect 298858 287239 299058 297121
rect 298858 287121 298899 287239
rect 299017 287121 299058 287239
rect 298858 277239 299058 287121
rect 298858 277121 298899 277239
rect 299017 277121 299058 277239
rect 298858 267239 299058 277121
rect 298858 267121 298899 267239
rect 299017 267121 299058 267239
rect 298858 257239 299058 267121
rect 298858 257121 298899 257239
rect 299017 257121 299058 257239
rect 298858 247239 299058 257121
rect 298858 247121 298899 247239
rect 299017 247121 299058 247239
rect 298858 237239 299058 247121
rect 298858 237121 298899 237239
rect 299017 237121 299058 237239
rect 298858 227239 299058 237121
rect 298858 227121 298899 227239
rect 299017 227121 299058 227239
rect 298858 217239 299058 227121
rect 298858 217121 298899 217239
rect 299017 217121 299058 217239
rect 298858 207239 299058 217121
rect 298858 207121 298899 207239
rect 299017 207121 299058 207239
rect 298858 197239 299058 207121
rect 298858 197121 298899 197239
rect 299017 197121 299058 197239
rect 298858 187239 299058 197121
rect 298858 187121 298899 187239
rect 299017 187121 299058 187239
rect 298858 177239 299058 187121
rect 298858 177121 298899 177239
rect 299017 177121 299058 177239
rect 298858 167239 299058 177121
rect 298858 167121 298899 167239
rect 299017 167121 299058 167239
rect 298858 157239 299058 167121
rect 298858 157121 298899 157239
rect 299017 157121 299058 157239
rect 298858 147239 299058 157121
rect 298858 147121 298899 147239
rect 299017 147121 299058 147239
rect 298858 137239 299058 147121
rect 298858 137121 298899 137239
rect 299017 137121 299058 137239
rect 298858 127239 299058 137121
rect 298858 127121 298899 127239
rect 299017 127121 299058 127239
rect 298858 117239 299058 127121
rect 298858 117121 298899 117239
rect 299017 117121 299058 117239
rect 298858 107239 299058 117121
rect 298858 107121 298899 107239
rect 299017 107121 299058 107239
rect 298858 97239 299058 107121
rect 298858 97121 298899 97239
rect 299017 97121 299058 97239
rect 298858 87239 299058 97121
rect 298858 87121 298899 87239
rect 299017 87121 299058 87239
rect 298858 77239 299058 87121
rect 298858 77121 298899 77239
rect 299017 77121 299058 77239
rect 298858 67239 299058 77121
rect 298858 67121 298899 67239
rect 299017 67121 299058 67239
rect 298858 57239 299058 67121
rect 298858 57121 298899 57239
rect 299017 57121 299058 57239
rect 298858 47239 299058 57121
rect 298858 47121 298899 47239
rect 299017 47121 299058 47239
rect 298858 37239 299058 47121
rect 298858 37121 298899 37239
rect 299017 37121 299058 37239
rect 298858 27239 299058 37121
rect 298858 27121 298899 27239
rect 299017 27121 299058 27239
rect 298858 17239 299058 27121
rect 298858 17121 298899 17239
rect 299017 17121 299058 17239
rect 298858 7239 299058 17121
rect 298858 7121 298899 7239
rect 299017 7121 299058 7239
rect 298858 559 299058 7121
rect 298858 441 298899 559
rect 299017 441 299058 559
rect 298858 400 299058 441
rect 299258 352239 299458 358233
rect 299258 352121 299299 352239
rect 299417 352121 299458 352239
rect 299258 342239 299458 352121
rect 299258 342121 299299 342239
rect 299417 342121 299458 342239
rect 299258 332239 299458 342121
rect 299258 332121 299299 332239
rect 299417 332121 299458 332239
rect 299258 322239 299458 332121
rect 299258 322121 299299 322239
rect 299417 322121 299458 322239
rect 299258 312239 299458 322121
rect 299258 312121 299299 312239
rect 299417 312121 299458 312239
rect 299258 302239 299458 312121
rect 299258 302121 299299 302239
rect 299417 302121 299458 302239
rect 299258 292239 299458 302121
rect 299258 292121 299299 292239
rect 299417 292121 299458 292239
rect 299258 282239 299458 292121
rect 299258 282121 299299 282239
rect 299417 282121 299458 282239
rect 299258 272239 299458 282121
rect 299258 272121 299299 272239
rect 299417 272121 299458 272239
rect 299258 262239 299458 272121
rect 299258 262121 299299 262239
rect 299417 262121 299458 262239
rect 299258 252239 299458 262121
rect 299258 252121 299299 252239
rect 299417 252121 299458 252239
rect 299258 242239 299458 252121
rect 299258 242121 299299 242239
rect 299417 242121 299458 242239
rect 299258 232239 299458 242121
rect 299258 232121 299299 232239
rect 299417 232121 299458 232239
rect 299258 222239 299458 232121
rect 299258 222121 299299 222239
rect 299417 222121 299458 222239
rect 299258 212239 299458 222121
rect 299258 212121 299299 212239
rect 299417 212121 299458 212239
rect 299258 202239 299458 212121
rect 299258 202121 299299 202239
rect 299417 202121 299458 202239
rect 299258 192239 299458 202121
rect 299258 192121 299299 192239
rect 299417 192121 299458 192239
rect 299258 182239 299458 192121
rect 299258 182121 299299 182239
rect 299417 182121 299458 182239
rect 299258 172239 299458 182121
rect 299258 172121 299299 172239
rect 299417 172121 299458 172239
rect 299258 162239 299458 172121
rect 299258 162121 299299 162239
rect 299417 162121 299458 162239
rect 299258 152239 299458 162121
rect 299258 152121 299299 152239
rect 299417 152121 299458 152239
rect 299258 142239 299458 152121
rect 299258 142121 299299 142239
rect 299417 142121 299458 142239
rect 299258 132239 299458 142121
rect 299258 132121 299299 132239
rect 299417 132121 299458 132239
rect 299258 122239 299458 132121
rect 299258 122121 299299 122239
rect 299417 122121 299458 122239
rect 299258 112239 299458 122121
rect 299258 112121 299299 112239
rect 299417 112121 299458 112239
rect 299258 102239 299458 112121
rect 299258 102121 299299 102239
rect 299417 102121 299458 102239
rect 299258 92239 299458 102121
rect 299258 92121 299299 92239
rect 299417 92121 299458 92239
rect 299258 82239 299458 92121
rect 299258 82121 299299 82239
rect 299417 82121 299458 82239
rect 299258 72239 299458 82121
rect 299258 72121 299299 72239
rect 299417 72121 299458 72239
rect 299258 62239 299458 72121
rect 299258 62121 299299 62239
rect 299417 62121 299458 62239
rect 299258 52239 299458 62121
rect 299258 52121 299299 52239
rect 299417 52121 299458 52239
rect 299258 42239 299458 52121
rect 299258 42121 299299 42239
rect 299417 42121 299458 42239
rect 299258 32239 299458 42121
rect 299258 32121 299299 32239
rect 299417 32121 299458 32239
rect 299258 22239 299458 32121
rect 299258 22121 299299 22239
rect 299417 22121 299458 22239
rect 299258 12239 299458 22121
rect 299258 12121 299299 12239
rect 299417 12121 299458 12239
rect 292080 41 292121 159
rect 292239 41 292280 159
rect 292080 0 292280 41
rect 299258 159 299458 12121
rect 299258 41 299299 159
rect 299417 41 299458 159
rect 299258 0 299458 41
<< via4 >>
rect 41 358233 159 358351
rect 41 352121 159 352239
rect 41 342121 159 342239
rect 41 332121 159 332239
rect 41 322121 159 322239
rect 41 312121 159 312239
rect 41 302121 159 302239
rect 41 292121 159 292239
rect 41 282121 159 282239
rect 41 272121 159 272239
rect 41 262121 159 262239
rect 41 252121 159 252239
rect 41 242121 159 242239
rect 41 232121 159 232239
rect 41 222121 159 222239
rect 41 212121 159 212239
rect 41 202121 159 202239
rect 41 192121 159 192239
rect 41 182121 159 182239
rect 41 172121 159 172239
rect 41 162121 159 162239
rect 41 152121 159 152239
rect 41 142121 159 142239
rect 41 132121 159 132239
rect 41 122121 159 122239
rect 41 112121 159 112239
rect 41 102121 159 102239
rect 41 92121 159 92239
rect 41 82121 159 82239
rect 41 72121 159 72239
rect 41 62121 159 62239
rect 41 52121 159 52239
rect 41 42121 159 42239
rect 41 32121 159 32239
rect 41 22121 159 22239
rect 41 12121 159 12239
rect 441 357833 559 357951
rect 7121 357833 7239 357951
rect 441 347121 559 347239
rect 441 337121 559 337239
rect 441 327121 559 327239
rect 441 317121 559 317239
rect 441 307121 559 307239
rect 441 297121 559 297239
rect 441 287121 559 287239
rect 441 277121 559 277239
rect 441 267121 559 267239
rect 441 257121 559 257239
rect 441 247121 559 247239
rect 441 237121 559 237239
rect 441 227121 559 227239
rect 441 217121 559 217239
rect 441 207121 559 207239
rect 441 197121 559 197239
rect 441 187121 559 187239
rect 441 177121 559 177239
rect 441 167121 559 167239
rect 441 157121 559 157239
rect 441 147121 559 147239
rect 441 137121 559 137239
rect 441 127121 559 127239
rect 441 117121 559 117239
rect 441 107121 559 107239
rect 441 97121 559 97239
rect 441 87121 559 87239
rect 441 77121 559 77239
rect 441 67121 559 67239
rect 441 57121 559 57239
rect 441 47121 559 47239
rect 441 37121 559 37239
rect 441 27121 559 27239
rect 441 17121 559 17239
rect 441 7121 559 7239
rect 841 357433 959 357551
rect 841 351161 959 351279
rect 841 341161 959 341279
rect 841 331161 959 331279
rect 841 321161 959 321279
rect 841 311161 959 311279
rect 841 301161 959 301279
rect 841 291161 959 291279
rect 841 281161 959 281279
rect 841 271161 959 271279
rect 841 261161 959 261279
rect 841 251161 959 251279
rect 841 241161 959 241279
rect 841 231161 959 231279
rect 841 221161 959 221279
rect 841 211161 959 211279
rect 841 201161 959 201279
rect 841 191161 959 191279
rect 841 181161 959 181279
rect 841 171161 959 171279
rect 841 161161 959 161279
rect 841 151161 959 151279
rect 841 141161 959 141279
rect 841 131161 959 131279
rect 841 121161 959 121279
rect 841 111161 959 111279
rect 841 101161 959 101279
rect 841 91161 959 91279
rect 841 81161 959 81279
rect 841 71161 959 71279
rect 841 61161 959 61279
rect 841 51161 959 51279
rect 841 41161 959 41279
rect 841 31161 959 31279
rect 841 21161 959 21279
rect 841 11161 959 11279
rect 1241 357033 1359 357151
rect 6161 357033 6279 357151
rect 1241 346161 1359 346279
rect 1241 336161 1359 336279
rect 1241 326161 1359 326279
rect 1241 316161 1359 316279
rect 1241 306161 1359 306279
rect 1241 296161 1359 296279
rect 1241 286161 1359 286279
rect 1241 276161 1359 276279
rect 1241 266161 1359 266279
rect 1241 256161 1359 256279
rect 1241 246161 1359 246279
rect 1241 236161 1359 236279
rect 1241 226161 1359 226279
rect 1241 216161 1359 216279
rect 1241 206161 1359 206279
rect 1241 196161 1359 196279
rect 1241 186161 1359 186279
rect 1241 176161 1359 176279
rect 1241 166161 1359 166279
rect 1241 156161 1359 156279
rect 1241 146161 1359 146279
rect 1241 136161 1359 136279
rect 1241 126161 1359 126279
rect 1241 116161 1359 116279
rect 1241 106161 1359 106279
rect 1241 96161 1359 96279
rect 1241 86161 1359 86279
rect 1241 76161 1359 76279
rect 1241 66161 1359 66279
rect 1241 56161 1359 56279
rect 1241 46161 1359 46279
rect 1241 36161 1359 36279
rect 1241 26161 1359 26279
rect 1241 16161 1359 16279
rect 1241 6161 1359 6279
rect 1641 356633 1759 356751
rect 1641 350201 1759 350319
rect 1641 340201 1759 340319
rect 1641 330201 1759 330319
rect 1641 320201 1759 320319
rect 1641 310201 1759 310319
rect 1641 300201 1759 300319
rect 1641 290201 1759 290319
rect 1641 280201 1759 280319
rect 1641 270201 1759 270319
rect 1641 260201 1759 260319
rect 1641 250201 1759 250319
rect 1641 240201 1759 240319
rect 1641 230201 1759 230319
rect 1641 220201 1759 220319
rect 1641 210201 1759 210319
rect 1641 200201 1759 200319
rect 1641 190201 1759 190319
rect 1641 180201 1759 180319
rect 1641 170201 1759 170319
rect 1641 160201 1759 160319
rect 1641 150201 1759 150319
rect 1641 140201 1759 140319
rect 1641 130201 1759 130319
rect 1641 120201 1759 120319
rect 1641 110201 1759 110319
rect 1641 100201 1759 100319
rect 1641 90201 1759 90319
rect 1641 80201 1759 80319
rect 1641 70201 1759 70319
rect 1641 60201 1759 60319
rect 1641 50201 1759 50319
rect 1641 40201 1759 40319
rect 1641 30201 1759 30319
rect 1641 20201 1759 20319
rect 1641 10201 1759 10319
rect 2041 356233 2159 356351
rect 5201 356233 5319 356351
rect 2041 345201 2159 345319
rect 2041 335201 2159 335319
rect 2041 325201 2159 325319
rect 2041 315201 2159 315319
rect 2041 305201 2159 305319
rect 2041 295201 2159 295319
rect 2041 285201 2159 285319
rect 2041 275201 2159 275319
rect 2041 265201 2159 265319
rect 2041 255201 2159 255319
rect 2041 245201 2159 245319
rect 2041 235201 2159 235319
rect 2041 225201 2159 225319
rect 2041 215201 2159 215319
rect 2041 205201 2159 205319
rect 2041 195201 2159 195319
rect 2041 185201 2159 185319
rect 2041 175201 2159 175319
rect 2041 165201 2159 165319
rect 2041 155201 2159 155319
rect 2041 145201 2159 145319
rect 2041 135201 2159 135319
rect 2041 125201 2159 125319
rect 2041 115201 2159 115319
rect 2041 105201 2159 105319
rect 2041 95201 2159 95319
rect 2041 85201 2159 85319
rect 2041 75201 2159 75319
rect 2041 65201 2159 65319
rect 2041 55201 2159 55319
rect 2041 45201 2159 45319
rect 2041 35201 2159 35319
rect 2041 25201 2159 25319
rect 2041 15201 2159 15319
rect 2041 5201 2159 5319
rect 2441 355833 2559 355951
rect 2441 349241 2559 349359
rect 2441 339241 2559 339359
rect 2441 329241 2559 329359
rect 2441 319241 2559 319359
rect 2441 309241 2559 309359
rect 2441 299241 2559 299359
rect 2441 289241 2559 289359
rect 2441 279241 2559 279359
rect 2441 269241 2559 269359
rect 2441 259241 2559 259359
rect 2441 249241 2559 249359
rect 2441 239241 2559 239359
rect 2441 229241 2559 229359
rect 2441 219241 2559 219359
rect 2441 209241 2559 209359
rect 2441 199241 2559 199359
rect 2441 189241 2559 189359
rect 2441 179241 2559 179359
rect 2441 169241 2559 169359
rect 2441 159241 2559 159359
rect 2441 149241 2559 149359
rect 2441 139241 2559 139359
rect 2441 129241 2559 129359
rect 2441 119241 2559 119359
rect 2441 109241 2559 109359
rect 2441 99241 2559 99359
rect 2441 89241 2559 89359
rect 2441 79241 2559 79359
rect 2441 69241 2559 69359
rect 2441 59241 2559 59359
rect 2441 49241 2559 49359
rect 2441 39241 2559 39359
rect 2441 29241 2559 29359
rect 2441 19241 2559 19359
rect 2441 9241 2559 9359
rect 2841 355433 2959 355551
rect 4241 355433 4359 355551
rect 12121 358233 12239 358351
rect 11161 357433 11279 357551
rect 10201 356633 10319 356751
rect 9241 355833 9359 355951
rect 17121 357833 17239 357951
rect 16161 357033 16279 357151
rect 15201 356233 15319 356351
rect 14241 355433 14359 355551
rect 22121 358233 22239 358351
rect 21161 357433 21279 357551
rect 20201 356633 20319 356751
rect 19241 355833 19359 355951
rect 27121 357833 27239 357951
rect 26161 357033 26279 357151
rect 25201 356233 25319 356351
rect 24241 355433 24359 355551
rect 32121 358233 32239 358351
rect 31161 357433 31279 357551
rect 30201 356633 30319 356751
rect 29241 355833 29359 355951
rect 37121 357833 37239 357951
rect 36161 357033 36279 357151
rect 35201 356233 35319 356351
rect 34241 355433 34359 355551
rect 42121 358233 42239 358351
rect 41161 357433 41279 357551
rect 40201 356633 40319 356751
rect 39241 355833 39359 355951
rect 47121 357833 47239 357951
rect 46161 357033 46279 357151
rect 45201 356233 45319 356351
rect 44241 355433 44359 355551
rect 52121 358233 52239 358351
rect 51161 357433 51279 357551
rect 50201 356633 50319 356751
rect 49241 355833 49359 355951
rect 57121 357833 57239 357951
rect 56161 357033 56279 357151
rect 55201 356233 55319 356351
rect 54241 355433 54359 355551
rect 62121 358233 62239 358351
rect 61161 357433 61279 357551
rect 60201 356633 60319 356751
rect 59241 355833 59359 355951
rect 67121 357833 67239 357951
rect 66161 357033 66279 357151
rect 65201 356233 65319 356351
rect 64241 355433 64359 355551
rect 72121 358233 72239 358351
rect 71161 357433 71279 357551
rect 70201 356633 70319 356751
rect 69241 355833 69359 355951
rect 77121 357833 77239 357951
rect 76161 357033 76279 357151
rect 75201 356233 75319 356351
rect 74241 355433 74359 355551
rect 82121 358233 82239 358351
rect 81161 357433 81279 357551
rect 80201 356633 80319 356751
rect 79241 355833 79359 355951
rect 87121 357833 87239 357951
rect 86161 357033 86279 357151
rect 85201 356233 85319 356351
rect 84241 355433 84359 355551
rect 92121 358233 92239 358351
rect 91161 357433 91279 357551
rect 90201 356633 90319 356751
rect 89241 355833 89359 355951
rect 97121 357833 97239 357951
rect 96161 357033 96279 357151
rect 95201 356233 95319 356351
rect 94241 355433 94359 355551
rect 102121 358233 102239 358351
rect 101161 357433 101279 357551
rect 100201 356633 100319 356751
rect 99241 355833 99359 355951
rect 107121 357833 107239 357951
rect 106161 357033 106279 357151
rect 105201 356233 105319 356351
rect 104241 355433 104359 355551
rect 112121 358233 112239 358351
rect 111161 357433 111279 357551
rect 110201 356633 110319 356751
rect 109241 355833 109359 355951
rect 117121 357833 117239 357951
rect 116161 357033 116279 357151
rect 115201 356233 115319 356351
rect 114241 355433 114359 355551
rect 122121 358233 122239 358351
rect 121161 357433 121279 357551
rect 120201 356633 120319 356751
rect 119241 355833 119359 355951
rect 127121 357833 127239 357951
rect 126161 357033 126279 357151
rect 125201 356233 125319 356351
rect 124241 355433 124359 355551
rect 132121 358233 132239 358351
rect 131161 357433 131279 357551
rect 130201 356633 130319 356751
rect 129241 355833 129359 355951
rect 137121 357833 137239 357951
rect 136161 357033 136279 357151
rect 135201 356233 135319 356351
rect 134241 355433 134359 355551
rect 142121 358233 142239 358351
rect 141161 357433 141279 357551
rect 140201 356633 140319 356751
rect 139241 355833 139359 355951
rect 147121 357833 147239 357951
rect 146161 357033 146279 357151
rect 145201 356233 145319 356351
rect 144241 355433 144359 355551
rect 152121 358233 152239 358351
rect 151161 357433 151279 357551
rect 150201 356633 150319 356751
rect 149241 355833 149359 355951
rect 157121 357833 157239 357951
rect 156161 357033 156279 357151
rect 155201 356233 155319 356351
rect 154241 355433 154359 355551
rect 162121 358233 162239 358351
rect 161161 357433 161279 357551
rect 160201 356633 160319 356751
rect 159241 355833 159359 355951
rect 167121 357833 167239 357951
rect 166161 357033 166279 357151
rect 165201 356233 165319 356351
rect 164241 355433 164359 355551
rect 172121 358233 172239 358351
rect 171161 357433 171279 357551
rect 170201 356633 170319 356751
rect 169241 355833 169359 355951
rect 177121 357833 177239 357951
rect 176161 357033 176279 357151
rect 175201 356233 175319 356351
rect 174241 355433 174359 355551
rect 182121 358233 182239 358351
rect 181161 357433 181279 357551
rect 180201 356633 180319 356751
rect 179241 355833 179359 355951
rect 187121 357833 187239 357951
rect 186161 357033 186279 357151
rect 185201 356233 185319 356351
rect 184241 355433 184359 355551
rect 192121 358233 192239 358351
rect 191161 357433 191279 357551
rect 190201 356633 190319 356751
rect 189241 355833 189359 355951
rect 197121 357833 197239 357951
rect 196161 357033 196279 357151
rect 195201 356233 195319 356351
rect 194241 355433 194359 355551
rect 202121 358233 202239 358351
rect 201161 357433 201279 357551
rect 200201 356633 200319 356751
rect 199241 355833 199359 355951
rect 207121 357833 207239 357951
rect 206161 357033 206279 357151
rect 205201 356233 205319 356351
rect 204241 355433 204359 355551
rect 212121 358233 212239 358351
rect 211161 357433 211279 357551
rect 210201 356633 210319 356751
rect 209241 355833 209359 355951
rect 217121 357833 217239 357951
rect 216161 357033 216279 357151
rect 215201 356233 215319 356351
rect 214241 355433 214359 355551
rect 222121 358233 222239 358351
rect 221161 357433 221279 357551
rect 220201 356633 220319 356751
rect 219241 355833 219359 355951
rect 227121 357833 227239 357951
rect 226161 357033 226279 357151
rect 225201 356233 225319 356351
rect 224241 355433 224359 355551
rect 232121 358233 232239 358351
rect 231161 357433 231279 357551
rect 230201 356633 230319 356751
rect 229241 355833 229359 355951
rect 237121 357833 237239 357951
rect 236161 357033 236279 357151
rect 235201 356233 235319 356351
rect 234241 355433 234359 355551
rect 242121 358233 242239 358351
rect 241161 357433 241279 357551
rect 240201 356633 240319 356751
rect 239241 355833 239359 355951
rect 247121 357833 247239 357951
rect 246161 357033 246279 357151
rect 245201 356233 245319 356351
rect 244241 355433 244359 355551
rect 252121 358233 252239 358351
rect 251161 357433 251279 357551
rect 250201 356633 250319 356751
rect 249241 355833 249359 355951
rect 257121 357833 257239 357951
rect 256161 357033 256279 357151
rect 255201 356233 255319 356351
rect 254241 355433 254359 355551
rect 262121 358233 262239 358351
rect 261161 357433 261279 357551
rect 260201 356633 260319 356751
rect 259241 355833 259359 355951
rect 267121 357833 267239 357951
rect 266161 357033 266279 357151
rect 265201 356233 265319 356351
rect 264241 355433 264359 355551
rect 272121 358233 272239 358351
rect 271161 357433 271279 357551
rect 270201 356633 270319 356751
rect 269241 355833 269359 355951
rect 277121 357833 277239 357951
rect 276161 357033 276279 357151
rect 275201 356233 275319 356351
rect 274241 355433 274359 355551
rect 282121 358233 282239 358351
rect 281161 357433 281279 357551
rect 280201 356633 280319 356751
rect 279241 355833 279359 355951
rect 287121 357833 287239 357951
rect 286161 357033 286279 357151
rect 285201 356233 285319 356351
rect 284241 355433 284359 355551
rect 292121 358233 292239 358351
rect 291161 357433 291279 357551
rect 290201 356633 290319 356751
rect 289241 355833 289359 355951
rect 299299 358233 299417 358351
rect 298899 357833 299017 357951
rect 298499 357433 298617 357551
rect 298099 357033 298217 357151
rect 297699 356633 297817 356751
rect 297299 356233 297417 356351
rect 296899 355833 297017 355951
rect 294241 355433 294359 355551
rect 296499 355433 296617 355551
rect 2841 344241 2959 344359
rect 2841 334241 2959 334359
rect 2841 324241 2959 324359
rect 2841 314241 2959 314359
rect 2841 304241 2959 304359
rect 2841 294241 2959 294359
rect 2841 284241 2959 284359
rect 2841 274241 2959 274359
rect 2841 264241 2959 264359
rect 2841 254241 2959 254359
rect 2841 244241 2959 244359
rect 2841 234241 2959 234359
rect 2841 224241 2959 224359
rect 2841 214241 2959 214359
rect 2841 204241 2959 204359
rect 2841 194241 2959 194359
rect 2841 184241 2959 184359
rect 2841 174241 2959 174359
rect 2841 164241 2959 164359
rect 2841 154241 2959 154359
rect 2841 144241 2959 144359
rect 2841 134241 2959 134359
rect 2841 124241 2959 124359
rect 2841 114241 2959 114359
rect 2841 104241 2959 104359
rect 2841 94241 2959 94359
rect 2841 84241 2959 84359
rect 2841 74241 2959 74359
rect 2841 64241 2959 64359
rect 2841 54241 2959 54359
rect 2841 44241 2959 44359
rect 2841 34241 2959 34359
rect 2841 24241 2959 24359
rect 2841 14241 2959 14359
rect 2841 4241 2959 4359
rect 296499 344241 296617 344359
rect 296499 334241 296617 334359
rect 296499 324241 296617 324359
rect 296499 314241 296617 314359
rect 296499 304241 296617 304359
rect 296499 294241 296617 294359
rect 296499 284241 296617 284359
rect 296499 274241 296617 274359
rect 296499 264241 296617 264359
rect 296499 254241 296617 254359
rect 296499 244241 296617 244359
rect 296499 234241 296617 234359
rect 296499 224241 296617 224359
rect 296499 214241 296617 214359
rect 296499 204241 296617 204359
rect 296499 194241 296617 194359
rect 296499 184241 296617 184359
rect 296499 174241 296617 174359
rect 296499 164241 296617 164359
rect 296499 154241 296617 154359
rect 296499 144241 296617 144359
rect 296499 134241 296617 134359
rect 296499 124241 296617 124359
rect 296499 114241 296617 114359
rect 296499 104241 296617 104359
rect 296499 94241 296617 94359
rect 296499 84241 296617 84359
rect 296499 74241 296617 74359
rect 296499 64241 296617 64359
rect 296499 54241 296617 54359
rect 296499 44241 296617 44359
rect 296499 34241 296617 34359
rect 296499 24241 296617 24359
rect 296499 14241 296617 14359
rect 296499 4241 296617 4359
rect 2841 2841 2959 2959
rect 4241 2841 4359 2959
rect 2441 2441 2559 2559
rect 2041 2041 2159 2159
rect 5201 2041 5319 2159
rect 1641 1641 1759 1759
rect 1241 1241 1359 1359
rect 6161 1241 6279 1359
rect 841 841 959 959
rect 441 441 559 559
rect 9241 2441 9359 2559
rect 10201 1641 10319 1759
rect 11161 841 11279 959
rect 7121 441 7239 559
rect 41 41 159 159
rect 14241 2841 14359 2959
rect 15201 2041 15319 2159
rect 16161 1241 16279 1359
rect 12121 41 12239 159
rect 19241 2441 19359 2559
rect 20201 1641 20319 1759
rect 21161 841 21279 959
rect 17121 441 17239 559
rect 24241 2841 24359 2959
rect 25201 2041 25319 2159
rect 26161 1241 26279 1359
rect 22121 41 22239 159
rect 29241 2441 29359 2559
rect 30201 1641 30319 1759
rect 31161 841 31279 959
rect 27121 441 27239 559
rect 34241 2841 34359 2959
rect 35201 2041 35319 2159
rect 36161 1241 36279 1359
rect 32121 41 32239 159
rect 39241 2441 39359 2559
rect 40201 1641 40319 1759
rect 41161 841 41279 959
rect 37121 441 37239 559
rect 44241 2841 44359 2959
rect 45201 2041 45319 2159
rect 46161 1241 46279 1359
rect 42121 41 42239 159
rect 49241 2441 49359 2559
rect 50201 1641 50319 1759
rect 51161 841 51279 959
rect 47121 441 47239 559
rect 54241 2841 54359 2959
rect 55201 2041 55319 2159
rect 56161 1241 56279 1359
rect 52121 41 52239 159
rect 59241 2441 59359 2559
rect 60201 1641 60319 1759
rect 61161 841 61279 959
rect 57121 441 57239 559
rect 64241 2841 64359 2959
rect 65201 2041 65319 2159
rect 66161 1241 66279 1359
rect 62121 41 62239 159
rect 69241 2441 69359 2559
rect 70201 1641 70319 1759
rect 71161 841 71279 959
rect 67121 441 67239 559
rect 74241 2841 74359 2959
rect 75201 2041 75319 2159
rect 76161 1241 76279 1359
rect 72121 41 72239 159
rect 79241 2441 79359 2559
rect 80201 1641 80319 1759
rect 81161 841 81279 959
rect 77121 441 77239 559
rect 84241 2841 84359 2959
rect 85201 2041 85319 2159
rect 86161 1241 86279 1359
rect 82121 41 82239 159
rect 89241 2441 89359 2559
rect 90201 1641 90319 1759
rect 91161 841 91279 959
rect 87121 441 87239 559
rect 94241 2841 94359 2959
rect 95201 2041 95319 2159
rect 96161 1241 96279 1359
rect 92121 41 92239 159
rect 99241 2441 99359 2559
rect 100201 1641 100319 1759
rect 101161 841 101279 959
rect 97121 441 97239 559
rect 104241 2841 104359 2959
rect 105201 2041 105319 2159
rect 106161 1241 106279 1359
rect 102121 41 102239 159
rect 109241 2441 109359 2559
rect 110201 1641 110319 1759
rect 111161 841 111279 959
rect 107121 441 107239 559
rect 114241 2841 114359 2959
rect 115201 2041 115319 2159
rect 116161 1241 116279 1359
rect 112121 41 112239 159
rect 119241 2441 119359 2559
rect 120201 1641 120319 1759
rect 121161 841 121279 959
rect 117121 441 117239 559
rect 124241 2841 124359 2959
rect 125201 2041 125319 2159
rect 126161 1241 126279 1359
rect 122121 41 122239 159
rect 129241 2441 129359 2559
rect 130201 1641 130319 1759
rect 131161 841 131279 959
rect 127121 441 127239 559
rect 134241 2841 134359 2959
rect 135201 2041 135319 2159
rect 136161 1241 136279 1359
rect 132121 41 132239 159
rect 139241 2441 139359 2559
rect 140201 1641 140319 1759
rect 141161 841 141279 959
rect 137121 441 137239 559
rect 144241 2841 144359 2959
rect 145201 2041 145319 2159
rect 146161 1241 146279 1359
rect 142121 41 142239 159
rect 149241 2441 149359 2559
rect 150201 1641 150319 1759
rect 151161 841 151279 959
rect 147121 441 147239 559
rect 154241 2841 154359 2959
rect 155201 2041 155319 2159
rect 156161 1241 156279 1359
rect 152121 41 152239 159
rect 159241 2441 159359 2559
rect 160201 1641 160319 1759
rect 161161 841 161279 959
rect 157121 441 157239 559
rect 164241 2841 164359 2959
rect 165201 2041 165319 2159
rect 166161 1241 166279 1359
rect 162121 41 162239 159
rect 169241 2441 169359 2559
rect 170201 1641 170319 1759
rect 171161 841 171279 959
rect 167121 441 167239 559
rect 174241 2841 174359 2959
rect 175201 2041 175319 2159
rect 176161 1241 176279 1359
rect 172121 41 172239 159
rect 179241 2441 179359 2559
rect 180201 1641 180319 1759
rect 181161 841 181279 959
rect 177121 441 177239 559
rect 184241 2841 184359 2959
rect 185201 2041 185319 2159
rect 186161 1241 186279 1359
rect 182121 41 182239 159
rect 189241 2441 189359 2559
rect 190201 1641 190319 1759
rect 191161 841 191279 959
rect 187121 441 187239 559
rect 194241 2841 194359 2959
rect 195201 2041 195319 2159
rect 196161 1241 196279 1359
rect 192121 41 192239 159
rect 199241 2441 199359 2559
rect 200201 1641 200319 1759
rect 201161 841 201279 959
rect 197121 441 197239 559
rect 204241 2841 204359 2959
rect 205201 2041 205319 2159
rect 206161 1241 206279 1359
rect 202121 41 202239 159
rect 209241 2441 209359 2559
rect 210201 1641 210319 1759
rect 211161 841 211279 959
rect 207121 441 207239 559
rect 214241 2841 214359 2959
rect 215201 2041 215319 2159
rect 216161 1241 216279 1359
rect 212121 41 212239 159
rect 219241 2441 219359 2559
rect 220201 1641 220319 1759
rect 221161 841 221279 959
rect 217121 441 217239 559
rect 224241 2841 224359 2959
rect 225201 2041 225319 2159
rect 226161 1241 226279 1359
rect 222121 41 222239 159
rect 229241 2441 229359 2559
rect 230201 1641 230319 1759
rect 231161 841 231279 959
rect 227121 441 227239 559
rect 234241 2841 234359 2959
rect 235201 2041 235319 2159
rect 236161 1241 236279 1359
rect 232121 41 232239 159
rect 239241 2441 239359 2559
rect 240201 1641 240319 1759
rect 241161 841 241279 959
rect 237121 441 237239 559
rect 244241 2841 244359 2959
rect 245201 2041 245319 2159
rect 246161 1241 246279 1359
rect 242121 41 242239 159
rect 249241 2441 249359 2559
rect 250201 1641 250319 1759
rect 251161 841 251279 959
rect 247121 441 247239 559
rect 254241 2841 254359 2959
rect 255201 2041 255319 2159
rect 256161 1241 256279 1359
rect 252121 41 252239 159
rect 259241 2441 259359 2559
rect 260201 1641 260319 1759
rect 261161 841 261279 959
rect 257121 441 257239 559
rect 264241 2841 264359 2959
rect 265201 2041 265319 2159
rect 266161 1241 266279 1359
rect 262121 41 262239 159
rect 269241 2441 269359 2559
rect 270201 1641 270319 1759
rect 271161 841 271279 959
rect 267121 441 267239 559
rect 274241 2841 274359 2959
rect 275201 2041 275319 2159
rect 276161 1241 276279 1359
rect 272121 41 272239 159
rect 279241 2441 279359 2559
rect 280201 1641 280319 1759
rect 281161 841 281279 959
rect 277121 441 277239 559
rect 284241 2841 284359 2959
rect 285201 2041 285319 2159
rect 286161 1241 286279 1359
rect 282121 41 282239 159
rect 289241 2441 289359 2559
rect 290201 1641 290319 1759
rect 291161 841 291279 959
rect 287121 441 287239 559
rect 294241 2841 294359 2959
rect 296499 2841 296617 2959
rect 296899 349241 297017 349359
rect 296899 339241 297017 339359
rect 296899 329241 297017 329359
rect 296899 319241 297017 319359
rect 296899 309241 297017 309359
rect 296899 299241 297017 299359
rect 296899 289241 297017 289359
rect 296899 279241 297017 279359
rect 296899 269241 297017 269359
rect 296899 259241 297017 259359
rect 296899 249241 297017 249359
rect 296899 239241 297017 239359
rect 296899 229241 297017 229359
rect 296899 219241 297017 219359
rect 296899 209241 297017 209359
rect 296899 199241 297017 199359
rect 296899 189241 297017 189359
rect 296899 179241 297017 179359
rect 296899 169241 297017 169359
rect 296899 159241 297017 159359
rect 296899 149241 297017 149359
rect 296899 139241 297017 139359
rect 296899 129241 297017 129359
rect 296899 119241 297017 119359
rect 296899 109241 297017 109359
rect 296899 99241 297017 99359
rect 296899 89241 297017 89359
rect 296899 79241 297017 79359
rect 296899 69241 297017 69359
rect 296899 59241 297017 59359
rect 296899 49241 297017 49359
rect 296899 39241 297017 39359
rect 296899 29241 297017 29359
rect 296899 19241 297017 19359
rect 296899 9241 297017 9359
rect 296899 2441 297017 2559
rect 297299 345201 297417 345319
rect 297299 335201 297417 335319
rect 297299 325201 297417 325319
rect 297299 315201 297417 315319
rect 297299 305201 297417 305319
rect 297299 295201 297417 295319
rect 297299 285201 297417 285319
rect 297299 275201 297417 275319
rect 297299 265201 297417 265319
rect 297299 255201 297417 255319
rect 297299 245201 297417 245319
rect 297299 235201 297417 235319
rect 297299 225201 297417 225319
rect 297299 215201 297417 215319
rect 297299 205201 297417 205319
rect 297299 195201 297417 195319
rect 297299 185201 297417 185319
rect 297299 175201 297417 175319
rect 297299 165201 297417 165319
rect 297299 155201 297417 155319
rect 297299 145201 297417 145319
rect 297299 135201 297417 135319
rect 297299 125201 297417 125319
rect 297299 115201 297417 115319
rect 297299 105201 297417 105319
rect 297299 95201 297417 95319
rect 297299 85201 297417 85319
rect 297299 75201 297417 75319
rect 297299 65201 297417 65319
rect 297299 55201 297417 55319
rect 297299 45201 297417 45319
rect 297299 35201 297417 35319
rect 297299 25201 297417 25319
rect 297299 15201 297417 15319
rect 297299 5201 297417 5319
rect 297299 2041 297417 2159
rect 297699 350201 297817 350319
rect 297699 340201 297817 340319
rect 297699 330201 297817 330319
rect 297699 320201 297817 320319
rect 297699 310201 297817 310319
rect 297699 300201 297817 300319
rect 297699 290201 297817 290319
rect 297699 280201 297817 280319
rect 297699 270201 297817 270319
rect 297699 260201 297817 260319
rect 297699 250201 297817 250319
rect 297699 240201 297817 240319
rect 297699 230201 297817 230319
rect 297699 220201 297817 220319
rect 297699 210201 297817 210319
rect 297699 200201 297817 200319
rect 297699 190201 297817 190319
rect 297699 180201 297817 180319
rect 297699 170201 297817 170319
rect 297699 160201 297817 160319
rect 297699 150201 297817 150319
rect 297699 140201 297817 140319
rect 297699 130201 297817 130319
rect 297699 120201 297817 120319
rect 297699 110201 297817 110319
rect 297699 100201 297817 100319
rect 297699 90201 297817 90319
rect 297699 80201 297817 80319
rect 297699 70201 297817 70319
rect 297699 60201 297817 60319
rect 297699 50201 297817 50319
rect 297699 40201 297817 40319
rect 297699 30201 297817 30319
rect 297699 20201 297817 20319
rect 297699 10201 297817 10319
rect 297699 1641 297817 1759
rect 298099 346161 298217 346279
rect 298099 336161 298217 336279
rect 298099 326161 298217 326279
rect 298099 316161 298217 316279
rect 298099 306161 298217 306279
rect 298099 296161 298217 296279
rect 298099 286161 298217 286279
rect 298099 276161 298217 276279
rect 298099 266161 298217 266279
rect 298099 256161 298217 256279
rect 298099 246161 298217 246279
rect 298099 236161 298217 236279
rect 298099 226161 298217 226279
rect 298099 216161 298217 216279
rect 298099 206161 298217 206279
rect 298099 196161 298217 196279
rect 298099 186161 298217 186279
rect 298099 176161 298217 176279
rect 298099 166161 298217 166279
rect 298099 156161 298217 156279
rect 298099 146161 298217 146279
rect 298099 136161 298217 136279
rect 298099 126161 298217 126279
rect 298099 116161 298217 116279
rect 298099 106161 298217 106279
rect 298099 96161 298217 96279
rect 298099 86161 298217 86279
rect 298099 76161 298217 76279
rect 298099 66161 298217 66279
rect 298099 56161 298217 56279
rect 298099 46161 298217 46279
rect 298099 36161 298217 36279
rect 298099 26161 298217 26279
rect 298099 16161 298217 16279
rect 298099 6161 298217 6279
rect 298099 1241 298217 1359
rect 298499 351161 298617 351279
rect 298499 341161 298617 341279
rect 298499 331161 298617 331279
rect 298499 321161 298617 321279
rect 298499 311161 298617 311279
rect 298499 301161 298617 301279
rect 298499 291161 298617 291279
rect 298499 281161 298617 281279
rect 298499 271161 298617 271279
rect 298499 261161 298617 261279
rect 298499 251161 298617 251279
rect 298499 241161 298617 241279
rect 298499 231161 298617 231279
rect 298499 221161 298617 221279
rect 298499 211161 298617 211279
rect 298499 201161 298617 201279
rect 298499 191161 298617 191279
rect 298499 181161 298617 181279
rect 298499 171161 298617 171279
rect 298499 161161 298617 161279
rect 298499 151161 298617 151279
rect 298499 141161 298617 141279
rect 298499 131161 298617 131279
rect 298499 121161 298617 121279
rect 298499 111161 298617 111279
rect 298499 101161 298617 101279
rect 298499 91161 298617 91279
rect 298499 81161 298617 81279
rect 298499 71161 298617 71279
rect 298499 61161 298617 61279
rect 298499 51161 298617 51279
rect 298499 41161 298617 41279
rect 298499 31161 298617 31279
rect 298499 21161 298617 21279
rect 298499 11161 298617 11279
rect 298499 841 298617 959
rect 298899 347121 299017 347239
rect 298899 337121 299017 337239
rect 298899 327121 299017 327239
rect 298899 317121 299017 317239
rect 298899 307121 299017 307239
rect 298899 297121 299017 297239
rect 298899 287121 299017 287239
rect 298899 277121 299017 277239
rect 298899 267121 299017 267239
rect 298899 257121 299017 257239
rect 298899 247121 299017 247239
rect 298899 237121 299017 237239
rect 298899 227121 299017 227239
rect 298899 217121 299017 217239
rect 298899 207121 299017 207239
rect 298899 197121 299017 197239
rect 298899 187121 299017 187239
rect 298899 177121 299017 177239
rect 298899 167121 299017 167239
rect 298899 157121 299017 157239
rect 298899 147121 299017 147239
rect 298899 137121 299017 137239
rect 298899 127121 299017 127239
rect 298899 117121 299017 117239
rect 298899 107121 299017 107239
rect 298899 97121 299017 97239
rect 298899 87121 299017 87239
rect 298899 77121 299017 77239
rect 298899 67121 299017 67239
rect 298899 57121 299017 57239
rect 298899 47121 299017 47239
rect 298899 37121 299017 37239
rect 298899 27121 299017 27239
rect 298899 17121 299017 17239
rect 298899 7121 299017 7239
rect 298899 441 299017 559
rect 299299 352121 299417 352239
rect 299299 342121 299417 342239
rect 299299 332121 299417 332239
rect 299299 322121 299417 322239
rect 299299 312121 299417 312239
rect 299299 302121 299417 302239
rect 299299 292121 299417 292239
rect 299299 282121 299417 282239
rect 299299 272121 299417 272239
rect 299299 262121 299417 262239
rect 299299 252121 299417 252239
rect 299299 242121 299417 242239
rect 299299 232121 299417 232239
rect 299299 222121 299417 222239
rect 299299 212121 299417 212239
rect 299299 202121 299417 202239
rect 299299 192121 299417 192239
rect 299299 182121 299417 182239
rect 299299 172121 299417 172239
rect 299299 162121 299417 162239
rect 299299 152121 299417 152239
rect 299299 142121 299417 142239
rect 299299 132121 299417 132239
rect 299299 122121 299417 122239
rect 299299 112121 299417 112239
rect 299299 102121 299417 102239
rect 299299 92121 299417 92239
rect 299299 82121 299417 82239
rect 299299 72121 299417 72239
rect 299299 62121 299417 62239
rect 299299 52121 299417 52239
rect 299299 42121 299417 42239
rect 299299 32121 299417 32239
rect 299299 22121 299417 22239
rect 299299 12121 299417 12239
rect 292121 41 292239 159
rect 299299 41 299417 159
<< metal5 >>
rect 0 358351 299458 358392
rect 0 358233 41 358351
rect 159 358233 12121 358351
rect 12239 358233 22121 358351
rect 22239 358233 32121 358351
rect 32239 358233 42121 358351
rect 42239 358233 52121 358351
rect 52239 358233 62121 358351
rect 62239 358233 72121 358351
rect 72239 358233 82121 358351
rect 82239 358233 92121 358351
rect 92239 358233 102121 358351
rect 102239 358233 112121 358351
rect 112239 358233 122121 358351
rect 122239 358233 132121 358351
rect 132239 358233 142121 358351
rect 142239 358233 152121 358351
rect 152239 358233 162121 358351
rect 162239 358233 172121 358351
rect 172239 358233 182121 358351
rect 182239 358233 192121 358351
rect 192239 358233 202121 358351
rect 202239 358233 212121 358351
rect 212239 358233 222121 358351
rect 222239 358233 232121 358351
rect 232239 358233 242121 358351
rect 242239 358233 252121 358351
rect 252239 358233 262121 358351
rect 262239 358233 272121 358351
rect 272239 358233 282121 358351
rect 282239 358233 292121 358351
rect 292239 358233 299299 358351
rect 299417 358233 299458 358351
rect 0 358192 299458 358233
rect 400 357951 299058 357992
rect 400 357833 441 357951
rect 559 357833 7121 357951
rect 7239 357833 17121 357951
rect 17239 357833 27121 357951
rect 27239 357833 37121 357951
rect 37239 357833 47121 357951
rect 47239 357833 57121 357951
rect 57239 357833 67121 357951
rect 67239 357833 77121 357951
rect 77239 357833 87121 357951
rect 87239 357833 97121 357951
rect 97239 357833 107121 357951
rect 107239 357833 117121 357951
rect 117239 357833 127121 357951
rect 127239 357833 137121 357951
rect 137239 357833 147121 357951
rect 147239 357833 157121 357951
rect 157239 357833 167121 357951
rect 167239 357833 177121 357951
rect 177239 357833 187121 357951
rect 187239 357833 197121 357951
rect 197239 357833 207121 357951
rect 207239 357833 217121 357951
rect 217239 357833 227121 357951
rect 227239 357833 237121 357951
rect 237239 357833 247121 357951
rect 247239 357833 257121 357951
rect 257239 357833 267121 357951
rect 267239 357833 277121 357951
rect 277239 357833 287121 357951
rect 287239 357833 298899 357951
rect 299017 357833 299058 357951
rect 400 357792 299058 357833
rect 800 357551 298658 357592
rect 800 357433 841 357551
rect 959 357433 11161 357551
rect 11279 357433 21161 357551
rect 21279 357433 31161 357551
rect 31279 357433 41161 357551
rect 41279 357433 51161 357551
rect 51279 357433 61161 357551
rect 61279 357433 71161 357551
rect 71279 357433 81161 357551
rect 81279 357433 91161 357551
rect 91279 357433 101161 357551
rect 101279 357433 111161 357551
rect 111279 357433 121161 357551
rect 121279 357433 131161 357551
rect 131279 357433 141161 357551
rect 141279 357433 151161 357551
rect 151279 357433 161161 357551
rect 161279 357433 171161 357551
rect 171279 357433 181161 357551
rect 181279 357433 191161 357551
rect 191279 357433 201161 357551
rect 201279 357433 211161 357551
rect 211279 357433 221161 357551
rect 221279 357433 231161 357551
rect 231279 357433 241161 357551
rect 241279 357433 251161 357551
rect 251279 357433 261161 357551
rect 261279 357433 271161 357551
rect 271279 357433 281161 357551
rect 281279 357433 291161 357551
rect 291279 357433 298499 357551
rect 298617 357433 298658 357551
rect 800 357392 298658 357433
rect 1200 357151 298258 357192
rect 1200 357033 1241 357151
rect 1359 357033 6161 357151
rect 6279 357033 16161 357151
rect 16279 357033 26161 357151
rect 26279 357033 36161 357151
rect 36279 357033 46161 357151
rect 46279 357033 56161 357151
rect 56279 357033 66161 357151
rect 66279 357033 76161 357151
rect 76279 357033 86161 357151
rect 86279 357033 96161 357151
rect 96279 357033 106161 357151
rect 106279 357033 116161 357151
rect 116279 357033 126161 357151
rect 126279 357033 136161 357151
rect 136279 357033 146161 357151
rect 146279 357033 156161 357151
rect 156279 357033 166161 357151
rect 166279 357033 176161 357151
rect 176279 357033 186161 357151
rect 186279 357033 196161 357151
rect 196279 357033 206161 357151
rect 206279 357033 216161 357151
rect 216279 357033 226161 357151
rect 226279 357033 236161 357151
rect 236279 357033 246161 357151
rect 246279 357033 256161 357151
rect 256279 357033 266161 357151
rect 266279 357033 276161 357151
rect 276279 357033 286161 357151
rect 286279 357033 298099 357151
rect 298217 357033 298258 357151
rect 1200 356992 298258 357033
rect 1600 356751 297858 356792
rect 1600 356633 1641 356751
rect 1759 356633 10201 356751
rect 10319 356633 20201 356751
rect 20319 356633 30201 356751
rect 30319 356633 40201 356751
rect 40319 356633 50201 356751
rect 50319 356633 60201 356751
rect 60319 356633 70201 356751
rect 70319 356633 80201 356751
rect 80319 356633 90201 356751
rect 90319 356633 100201 356751
rect 100319 356633 110201 356751
rect 110319 356633 120201 356751
rect 120319 356633 130201 356751
rect 130319 356633 140201 356751
rect 140319 356633 150201 356751
rect 150319 356633 160201 356751
rect 160319 356633 170201 356751
rect 170319 356633 180201 356751
rect 180319 356633 190201 356751
rect 190319 356633 200201 356751
rect 200319 356633 210201 356751
rect 210319 356633 220201 356751
rect 220319 356633 230201 356751
rect 230319 356633 240201 356751
rect 240319 356633 250201 356751
rect 250319 356633 260201 356751
rect 260319 356633 270201 356751
rect 270319 356633 280201 356751
rect 280319 356633 290201 356751
rect 290319 356633 297699 356751
rect 297817 356633 297858 356751
rect 1600 356592 297858 356633
rect 2000 356351 297458 356392
rect 2000 356233 2041 356351
rect 2159 356233 5201 356351
rect 5319 356233 15201 356351
rect 15319 356233 25201 356351
rect 25319 356233 35201 356351
rect 35319 356233 45201 356351
rect 45319 356233 55201 356351
rect 55319 356233 65201 356351
rect 65319 356233 75201 356351
rect 75319 356233 85201 356351
rect 85319 356233 95201 356351
rect 95319 356233 105201 356351
rect 105319 356233 115201 356351
rect 115319 356233 125201 356351
rect 125319 356233 135201 356351
rect 135319 356233 145201 356351
rect 145319 356233 155201 356351
rect 155319 356233 165201 356351
rect 165319 356233 175201 356351
rect 175319 356233 185201 356351
rect 185319 356233 195201 356351
rect 195319 356233 205201 356351
rect 205319 356233 215201 356351
rect 215319 356233 225201 356351
rect 225319 356233 235201 356351
rect 235319 356233 245201 356351
rect 245319 356233 255201 356351
rect 255319 356233 265201 356351
rect 265319 356233 275201 356351
rect 275319 356233 285201 356351
rect 285319 356233 297299 356351
rect 297417 356233 297458 356351
rect 2000 356192 297458 356233
rect 2400 355951 297058 355992
rect 2400 355833 2441 355951
rect 2559 355833 9241 355951
rect 9359 355833 19241 355951
rect 19359 355833 29241 355951
rect 29359 355833 39241 355951
rect 39359 355833 49241 355951
rect 49359 355833 59241 355951
rect 59359 355833 69241 355951
rect 69359 355833 79241 355951
rect 79359 355833 89241 355951
rect 89359 355833 99241 355951
rect 99359 355833 109241 355951
rect 109359 355833 119241 355951
rect 119359 355833 129241 355951
rect 129359 355833 139241 355951
rect 139359 355833 149241 355951
rect 149359 355833 159241 355951
rect 159359 355833 169241 355951
rect 169359 355833 179241 355951
rect 179359 355833 189241 355951
rect 189359 355833 199241 355951
rect 199359 355833 209241 355951
rect 209359 355833 219241 355951
rect 219359 355833 229241 355951
rect 229359 355833 239241 355951
rect 239359 355833 249241 355951
rect 249359 355833 259241 355951
rect 259359 355833 269241 355951
rect 269359 355833 279241 355951
rect 279359 355833 289241 355951
rect 289359 355833 296899 355951
rect 297017 355833 297058 355951
rect 2400 355792 297058 355833
rect 2800 355551 296658 355592
rect 2800 355433 2841 355551
rect 2959 355433 4241 355551
rect 4359 355433 14241 355551
rect 14359 355433 24241 355551
rect 24359 355433 34241 355551
rect 34359 355433 44241 355551
rect 44359 355433 54241 355551
rect 54359 355433 64241 355551
rect 64359 355433 74241 355551
rect 74359 355433 84241 355551
rect 84359 355433 94241 355551
rect 94359 355433 104241 355551
rect 104359 355433 114241 355551
rect 114359 355433 124241 355551
rect 124359 355433 134241 355551
rect 134359 355433 144241 355551
rect 144359 355433 154241 355551
rect 154359 355433 164241 355551
rect 164359 355433 174241 355551
rect 174359 355433 184241 355551
rect 184359 355433 194241 355551
rect 194359 355433 204241 355551
rect 204359 355433 214241 355551
rect 214359 355433 224241 355551
rect 224359 355433 234241 355551
rect 234359 355433 244241 355551
rect 244359 355433 254241 355551
rect 254359 355433 264241 355551
rect 264359 355433 274241 355551
rect 274359 355433 284241 355551
rect 284359 355433 294241 355551
rect 294359 355433 296499 355551
rect 296617 355433 296658 355551
rect 2800 355392 296658 355433
rect 0 352239 3988 352280
rect 0 352121 41 352239
rect 159 352121 3988 352239
rect 0 352080 3988 352121
rect 295508 352239 299458 352280
rect 295508 352121 299299 352239
rect 299417 352121 299458 352239
rect 295508 352080 299458 352121
rect 800 351279 3988 351320
rect 800 351161 841 351279
rect 959 351161 3988 351279
rect 800 351120 3988 351161
rect 295508 351279 298658 351320
rect 295508 351161 298499 351279
rect 298617 351161 298658 351279
rect 295508 351120 298658 351161
rect 1600 350319 3988 350360
rect 1600 350201 1641 350319
rect 1759 350201 3988 350319
rect 1600 350160 3988 350201
rect 295508 350319 297858 350360
rect 295508 350201 297699 350319
rect 297817 350201 297858 350319
rect 295508 350160 297858 350201
rect 2400 349359 3988 349400
rect 2400 349241 2441 349359
rect 2559 349241 3988 349359
rect 2400 349200 3988 349241
rect 295508 349359 297058 349400
rect 295508 349241 296899 349359
rect 297017 349241 297058 349359
rect 295508 349200 297058 349241
rect 0 347239 3988 347280
rect 0 347121 441 347239
rect 559 347121 3988 347239
rect 0 347080 3988 347121
rect 295508 347239 299458 347280
rect 295508 347121 298899 347239
rect 299017 347121 299458 347239
rect 295508 347080 299458 347121
rect 800 346279 3988 346320
rect 800 346161 1241 346279
rect 1359 346161 3988 346279
rect 800 346120 3988 346161
rect 295508 346279 298658 346320
rect 295508 346161 298099 346279
rect 298217 346161 298658 346279
rect 295508 346120 298658 346161
rect 1600 345319 3988 345360
rect 1600 345201 2041 345319
rect 2159 345201 3988 345319
rect 1600 345160 3988 345201
rect 295508 345319 297858 345360
rect 295508 345201 297299 345319
rect 297417 345201 297858 345319
rect 295508 345160 297858 345201
rect 2400 344359 3988 344400
rect 2400 344241 2841 344359
rect 2959 344241 3988 344359
rect 2400 344200 3988 344241
rect 295508 344359 297058 344400
rect 295508 344241 296499 344359
rect 296617 344241 297058 344359
rect 295508 344200 297058 344241
rect 0 342239 3988 342280
rect 0 342121 41 342239
rect 159 342121 3988 342239
rect 0 342080 3988 342121
rect 295508 342239 299458 342280
rect 295508 342121 299299 342239
rect 299417 342121 299458 342239
rect 295508 342080 299458 342121
rect 800 341279 3988 341320
rect 800 341161 841 341279
rect 959 341161 3988 341279
rect 800 341120 3988 341161
rect 295508 341279 298658 341320
rect 295508 341161 298499 341279
rect 298617 341161 298658 341279
rect 295508 341120 298658 341161
rect 1600 340319 3988 340360
rect 1600 340201 1641 340319
rect 1759 340201 3988 340319
rect 1600 340160 3988 340201
rect 295508 340319 297858 340360
rect 295508 340201 297699 340319
rect 297817 340201 297858 340319
rect 295508 340160 297858 340201
rect 2400 339359 3988 339400
rect 2400 339241 2441 339359
rect 2559 339241 3988 339359
rect 2400 339200 3988 339241
rect 295508 339359 297058 339400
rect 295508 339241 296899 339359
rect 297017 339241 297058 339359
rect 295508 339200 297058 339241
rect 0 337239 3988 337280
rect 0 337121 441 337239
rect 559 337121 3988 337239
rect 0 337080 3988 337121
rect 295508 337239 299458 337280
rect 295508 337121 298899 337239
rect 299017 337121 299458 337239
rect 295508 337080 299458 337121
rect 800 336279 3988 336320
rect 800 336161 1241 336279
rect 1359 336161 3988 336279
rect 800 336120 3988 336161
rect 295508 336279 298658 336320
rect 295508 336161 298099 336279
rect 298217 336161 298658 336279
rect 295508 336120 298658 336161
rect 1600 335319 3988 335360
rect 1600 335201 2041 335319
rect 2159 335201 3988 335319
rect 1600 335160 3988 335201
rect 295508 335319 297858 335360
rect 295508 335201 297299 335319
rect 297417 335201 297858 335319
rect 295508 335160 297858 335201
rect 2400 334359 3988 334400
rect 2400 334241 2841 334359
rect 2959 334241 3988 334359
rect 2400 334200 3988 334241
rect 295508 334359 297058 334400
rect 295508 334241 296499 334359
rect 296617 334241 297058 334359
rect 295508 334200 297058 334241
rect 0 332239 3988 332280
rect 0 332121 41 332239
rect 159 332121 3988 332239
rect 0 332080 3988 332121
rect 295508 332239 299458 332280
rect 295508 332121 299299 332239
rect 299417 332121 299458 332239
rect 295508 332080 299458 332121
rect 800 331279 3988 331320
rect 800 331161 841 331279
rect 959 331161 3988 331279
rect 800 331120 3988 331161
rect 295508 331279 298658 331320
rect 295508 331161 298499 331279
rect 298617 331161 298658 331279
rect 295508 331120 298658 331161
rect 1600 330319 3988 330360
rect 1600 330201 1641 330319
rect 1759 330201 3988 330319
rect 1600 330160 3988 330201
rect 295508 330319 297858 330360
rect 295508 330201 297699 330319
rect 297817 330201 297858 330319
rect 295508 330160 297858 330201
rect 2400 329359 3988 329400
rect 2400 329241 2441 329359
rect 2559 329241 3988 329359
rect 2400 329200 3988 329241
rect 295508 329359 297058 329400
rect 295508 329241 296899 329359
rect 297017 329241 297058 329359
rect 295508 329200 297058 329241
rect 0 327239 3988 327280
rect 0 327121 441 327239
rect 559 327121 3988 327239
rect 0 327080 3988 327121
rect 295508 327239 299458 327280
rect 295508 327121 298899 327239
rect 299017 327121 299458 327239
rect 295508 327080 299458 327121
rect 800 326279 3988 326320
rect 800 326161 1241 326279
rect 1359 326161 3988 326279
rect 800 326120 3988 326161
rect 295508 326279 298658 326320
rect 295508 326161 298099 326279
rect 298217 326161 298658 326279
rect 295508 326120 298658 326161
rect 1600 325319 3988 325360
rect 1600 325201 2041 325319
rect 2159 325201 3988 325319
rect 1600 325160 3988 325201
rect 295508 325319 297858 325360
rect 295508 325201 297299 325319
rect 297417 325201 297858 325319
rect 295508 325160 297858 325201
rect 2400 324359 3988 324400
rect 2400 324241 2841 324359
rect 2959 324241 3988 324359
rect 2400 324200 3988 324241
rect 295508 324359 297058 324400
rect 295508 324241 296499 324359
rect 296617 324241 297058 324359
rect 295508 324200 297058 324241
rect 0 322239 3988 322280
rect 0 322121 41 322239
rect 159 322121 3988 322239
rect 0 322080 3988 322121
rect 295508 322239 299458 322280
rect 295508 322121 299299 322239
rect 299417 322121 299458 322239
rect 295508 322080 299458 322121
rect 800 321279 3988 321320
rect 800 321161 841 321279
rect 959 321161 3988 321279
rect 800 321120 3988 321161
rect 295508 321279 298658 321320
rect 295508 321161 298499 321279
rect 298617 321161 298658 321279
rect 295508 321120 298658 321161
rect 1600 320319 3988 320360
rect 1600 320201 1641 320319
rect 1759 320201 3988 320319
rect 1600 320160 3988 320201
rect 295508 320319 297858 320360
rect 295508 320201 297699 320319
rect 297817 320201 297858 320319
rect 295508 320160 297858 320201
rect 2400 319359 3988 319400
rect 2400 319241 2441 319359
rect 2559 319241 3988 319359
rect 2400 319200 3988 319241
rect 295508 319359 297058 319400
rect 295508 319241 296899 319359
rect 297017 319241 297058 319359
rect 295508 319200 297058 319241
rect 0 317239 3988 317280
rect 0 317121 441 317239
rect 559 317121 3988 317239
rect 0 317080 3988 317121
rect 295508 317239 299458 317280
rect 295508 317121 298899 317239
rect 299017 317121 299458 317239
rect 295508 317080 299458 317121
rect 800 316279 3988 316320
rect 800 316161 1241 316279
rect 1359 316161 3988 316279
rect 800 316120 3988 316161
rect 295508 316279 298658 316320
rect 295508 316161 298099 316279
rect 298217 316161 298658 316279
rect 295508 316120 298658 316161
rect 1600 315319 3988 315360
rect 1600 315201 2041 315319
rect 2159 315201 3988 315319
rect 1600 315160 3988 315201
rect 295508 315319 297858 315360
rect 295508 315201 297299 315319
rect 297417 315201 297858 315319
rect 295508 315160 297858 315201
rect 2400 314359 3988 314400
rect 2400 314241 2841 314359
rect 2959 314241 3988 314359
rect 2400 314200 3988 314241
rect 295508 314359 297058 314400
rect 295508 314241 296499 314359
rect 296617 314241 297058 314359
rect 295508 314200 297058 314241
rect 0 312239 3988 312280
rect 0 312121 41 312239
rect 159 312121 3988 312239
rect 0 312080 3988 312121
rect 295508 312239 299458 312280
rect 295508 312121 299299 312239
rect 299417 312121 299458 312239
rect 295508 312080 299458 312121
rect 800 311279 3988 311320
rect 800 311161 841 311279
rect 959 311161 3988 311279
rect 800 311120 3988 311161
rect 295508 311279 298658 311320
rect 295508 311161 298499 311279
rect 298617 311161 298658 311279
rect 295508 311120 298658 311161
rect 1600 310319 3988 310360
rect 1600 310201 1641 310319
rect 1759 310201 3988 310319
rect 1600 310160 3988 310201
rect 295508 310319 297858 310360
rect 295508 310201 297699 310319
rect 297817 310201 297858 310319
rect 295508 310160 297858 310201
rect 2400 309359 3988 309400
rect 2400 309241 2441 309359
rect 2559 309241 3988 309359
rect 2400 309200 3988 309241
rect 295508 309359 297058 309400
rect 295508 309241 296899 309359
rect 297017 309241 297058 309359
rect 295508 309200 297058 309241
rect 0 307239 3988 307280
rect 0 307121 441 307239
rect 559 307121 3988 307239
rect 0 307080 3988 307121
rect 295508 307239 299458 307280
rect 295508 307121 298899 307239
rect 299017 307121 299458 307239
rect 295508 307080 299458 307121
rect 800 306279 3988 306320
rect 800 306161 1241 306279
rect 1359 306161 3988 306279
rect 800 306120 3988 306161
rect 295508 306279 298658 306320
rect 295508 306161 298099 306279
rect 298217 306161 298658 306279
rect 295508 306120 298658 306161
rect 1600 305319 3988 305360
rect 1600 305201 2041 305319
rect 2159 305201 3988 305319
rect 1600 305160 3988 305201
rect 295508 305319 297858 305360
rect 295508 305201 297299 305319
rect 297417 305201 297858 305319
rect 295508 305160 297858 305201
rect 2400 304359 3988 304400
rect 2400 304241 2841 304359
rect 2959 304241 3988 304359
rect 2400 304200 3988 304241
rect 295508 304359 297058 304400
rect 295508 304241 296499 304359
rect 296617 304241 297058 304359
rect 295508 304200 297058 304241
rect 0 302239 3988 302280
rect 0 302121 41 302239
rect 159 302121 3988 302239
rect 0 302080 3988 302121
rect 295508 302239 299458 302280
rect 295508 302121 299299 302239
rect 299417 302121 299458 302239
rect 295508 302080 299458 302121
rect 800 301279 3988 301320
rect 800 301161 841 301279
rect 959 301161 3988 301279
rect 800 301120 3988 301161
rect 295508 301279 298658 301320
rect 295508 301161 298499 301279
rect 298617 301161 298658 301279
rect 295508 301120 298658 301161
rect 1600 300319 3988 300360
rect 1600 300201 1641 300319
rect 1759 300201 3988 300319
rect 1600 300160 3988 300201
rect 295508 300319 297858 300360
rect 295508 300201 297699 300319
rect 297817 300201 297858 300319
rect 295508 300160 297858 300201
rect 2400 299359 3988 299400
rect 2400 299241 2441 299359
rect 2559 299241 3988 299359
rect 2400 299200 3988 299241
rect 295508 299359 297058 299400
rect 295508 299241 296899 299359
rect 297017 299241 297058 299359
rect 295508 299200 297058 299241
rect 0 297239 3988 297280
rect 0 297121 441 297239
rect 559 297121 3988 297239
rect 0 297080 3988 297121
rect 295508 297239 299458 297280
rect 295508 297121 298899 297239
rect 299017 297121 299458 297239
rect 295508 297080 299458 297121
rect 800 296279 3988 296320
rect 800 296161 1241 296279
rect 1359 296161 3988 296279
rect 800 296120 3988 296161
rect 295508 296279 298658 296320
rect 295508 296161 298099 296279
rect 298217 296161 298658 296279
rect 295508 296120 298658 296161
rect 1600 295319 3988 295360
rect 1600 295201 2041 295319
rect 2159 295201 3988 295319
rect 1600 295160 3988 295201
rect 295508 295319 297858 295360
rect 295508 295201 297299 295319
rect 297417 295201 297858 295319
rect 295508 295160 297858 295201
rect 2400 294359 3988 294400
rect 2400 294241 2841 294359
rect 2959 294241 3988 294359
rect 2400 294200 3988 294241
rect 295508 294359 297058 294400
rect 295508 294241 296499 294359
rect 296617 294241 297058 294359
rect 295508 294200 297058 294241
rect 0 292239 3988 292280
rect 0 292121 41 292239
rect 159 292121 3988 292239
rect 0 292080 3988 292121
rect 295508 292239 299458 292280
rect 295508 292121 299299 292239
rect 299417 292121 299458 292239
rect 295508 292080 299458 292121
rect 800 291279 3988 291320
rect 800 291161 841 291279
rect 959 291161 3988 291279
rect 800 291120 3988 291161
rect 295508 291279 298658 291320
rect 295508 291161 298499 291279
rect 298617 291161 298658 291279
rect 295508 291120 298658 291161
rect 1600 290319 3988 290360
rect 1600 290201 1641 290319
rect 1759 290201 3988 290319
rect 1600 290160 3988 290201
rect 295508 290319 297858 290360
rect 295508 290201 297699 290319
rect 297817 290201 297858 290319
rect 295508 290160 297858 290201
rect 2400 289359 3988 289400
rect 2400 289241 2441 289359
rect 2559 289241 3988 289359
rect 2400 289200 3988 289241
rect 295508 289359 297058 289400
rect 295508 289241 296899 289359
rect 297017 289241 297058 289359
rect 295508 289200 297058 289241
rect 0 287239 3988 287280
rect 0 287121 441 287239
rect 559 287121 3988 287239
rect 0 287080 3988 287121
rect 295508 287239 299458 287280
rect 295508 287121 298899 287239
rect 299017 287121 299458 287239
rect 295508 287080 299458 287121
rect 800 286279 3988 286320
rect 800 286161 1241 286279
rect 1359 286161 3988 286279
rect 800 286120 3988 286161
rect 295508 286279 298658 286320
rect 295508 286161 298099 286279
rect 298217 286161 298658 286279
rect 295508 286120 298658 286161
rect 1600 285319 3988 285360
rect 1600 285201 2041 285319
rect 2159 285201 3988 285319
rect 1600 285160 3988 285201
rect 295508 285319 297858 285360
rect 295508 285201 297299 285319
rect 297417 285201 297858 285319
rect 295508 285160 297858 285201
rect 2400 284359 3988 284400
rect 2400 284241 2841 284359
rect 2959 284241 3988 284359
rect 2400 284200 3988 284241
rect 295508 284359 297058 284400
rect 295508 284241 296499 284359
rect 296617 284241 297058 284359
rect 295508 284200 297058 284241
rect 0 282239 3988 282280
rect 0 282121 41 282239
rect 159 282121 3988 282239
rect 0 282080 3988 282121
rect 295508 282239 299458 282280
rect 295508 282121 299299 282239
rect 299417 282121 299458 282239
rect 295508 282080 299458 282121
rect 800 281279 3988 281320
rect 800 281161 841 281279
rect 959 281161 3988 281279
rect 800 281120 3988 281161
rect 295508 281279 298658 281320
rect 295508 281161 298499 281279
rect 298617 281161 298658 281279
rect 295508 281120 298658 281161
rect 1600 280319 3988 280360
rect 1600 280201 1641 280319
rect 1759 280201 3988 280319
rect 1600 280160 3988 280201
rect 295508 280319 297858 280360
rect 295508 280201 297699 280319
rect 297817 280201 297858 280319
rect 295508 280160 297858 280201
rect 2400 279359 3988 279400
rect 2400 279241 2441 279359
rect 2559 279241 3988 279359
rect 2400 279200 3988 279241
rect 295508 279359 297058 279400
rect 295508 279241 296899 279359
rect 297017 279241 297058 279359
rect 295508 279200 297058 279241
rect 0 277239 3988 277280
rect 0 277121 441 277239
rect 559 277121 3988 277239
rect 0 277080 3988 277121
rect 295508 277239 299458 277280
rect 295508 277121 298899 277239
rect 299017 277121 299458 277239
rect 295508 277080 299458 277121
rect 800 276279 3988 276320
rect 800 276161 1241 276279
rect 1359 276161 3988 276279
rect 800 276120 3988 276161
rect 295508 276279 298658 276320
rect 295508 276161 298099 276279
rect 298217 276161 298658 276279
rect 295508 276120 298658 276161
rect 1600 275319 3988 275360
rect 1600 275201 2041 275319
rect 2159 275201 3988 275319
rect 1600 275160 3988 275201
rect 295508 275319 297858 275360
rect 295508 275201 297299 275319
rect 297417 275201 297858 275319
rect 295508 275160 297858 275201
rect 2400 274359 3988 274400
rect 2400 274241 2841 274359
rect 2959 274241 3988 274359
rect 2400 274200 3988 274241
rect 295508 274359 297058 274400
rect 295508 274241 296499 274359
rect 296617 274241 297058 274359
rect 295508 274200 297058 274241
rect 0 272239 3988 272280
rect 0 272121 41 272239
rect 159 272121 3988 272239
rect 0 272080 3988 272121
rect 295508 272239 299458 272280
rect 295508 272121 299299 272239
rect 299417 272121 299458 272239
rect 295508 272080 299458 272121
rect 800 271279 3988 271320
rect 800 271161 841 271279
rect 959 271161 3988 271279
rect 800 271120 3988 271161
rect 295508 271279 298658 271320
rect 295508 271161 298499 271279
rect 298617 271161 298658 271279
rect 295508 271120 298658 271161
rect 1600 270319 3988 270360
rect 1600 270201 1641 270319
rect 1759 270201 3988 270319
rect 1600 270160 3988 270201
rect 295508 270319 297858 270360
rect 295508 270201 297699 270319
rect 297817 270201 297858 270319
rect 295508 270160 297858 270201
rect 2400 269359 3988 269400
rect 2400 269241 2441 269359
rect 2559 269241 3988 269359
rect 2400 269200 3988 269241
rect 295508 269359 297058 269400
rect 295508 269241 296899 269359
rect 297017 269241 297058 269359
rect 295508 269200 297058 269241
rect 0 267239 3988 267280
rect 0 267121 441 267239
rect 559 267121 3988 267239
rect 0 267080 3988 267121
rect 295508 267239 299458 267280
rect 295508 267121 298899 267239
rect 299017 267121 299458 267239
rect 295508 267080 299458 267121
rect 800 266279 3988 266320
rect 800 266161 1241 266279
rect 1359 266161 3988 266279
rect 800 266120 3988 266161
rect 295508 266279 298658 266320
rect 295508 266161 298099 266279
rect 298217 266161 298658 266279
rect 295508 266120 298658 266161
rect 1600 265319 3988 265360
rect 1600 265201 2041 265319
rect 2159 265201 3988 265319
rect 1600 265160 3988 265201
rect 295508 265319 297858 265360
rect 295508 265201 297299 265319
rect 297417 265201 297858 265319
rect 295508 265160 297858 265201
rect 2400 264359 3988 264400
rect 2400 264241 2841 264359
rect 2959 264241 3988 264359
rect 2400 264200 3988 264241
rect 295508 264359 297058 264400
rect 295508 264241 296499 264359
rect 296617 264241 297058 264359
rect 295508 264200 297058 264241
rect 0 262239 3988 262280
rect 0 262121 41 262239
rect 159 262121 3988 262239
rect 0 262080 3988 262121
rect 295508 262239 299458 262280
rect 295508 262121 299299 262239
rect 299417 262121 299458 262239
rect 295508 262080 299458 262121
rect 800 261279 3988 261320
rect 800 261161 841 261279
rect 959 261161 3988 261279
rect 800 261120 3988 261161
rect 295508 261279 298658 261320
rect 295508 261161 298499 261279
rect 298617 261161 298658 261279
rect 295508 261120 298658 261161
rect 1600 260319 3988 260360
rect 1600 260201 1641 260319
rect 1759 260201 3988 260319
rect 1600 260160 3988 260201
rect 295508 260319 297858 260360
rect 295508 260201 297699 260319
rect 297817 260201 297858 260319
rect 295508 260160 297858 260201
rect 2400 259359 3988 259400
rect 2400 259241 2441 259359
rect 2559 259241 3988 259359
rect 2400 259200 3988 259241
rect 295508 259359 297058 259400
rect 295508 259241 296899 259359
rect 297017 259241 297058 259359
rect 295508 259200 297058 259241
rect 0 257239 3988 257280
rect 0 257121 441 257239
rect 559 257121 3988 257239
rect 0 257080 3988 257121
rect 295508 257239 299458 257280
rect 295508 257121 298899 257239
rect 299017 257121 299458 257239
rect 295508 257080 299458 257121
rect 800 256279 3988 256320
rect 800 256161 1241 256279
rect 1359 256161 3988 256279
rect 800 256120 3988 256161
rect 295508 256279 298658 256320
rect 295508 256161 298099 256279
rect 298217 256161 298658 256279
rect 295508 256120 298658 256161
rect 1600 255319 3988 255360
rect 1600 255201 2041 255319
rect 2159 255201 3988 255319
rect 1600 255160 3988 255201
rect 295508 255319 297858 255360
rect 295508 255201 297299 255319
rect 297417 255201 297858 255319
rect 295508 255160 297858 255201
rect 2400 254359 3988 254400
rect 2400 254241 2841 254359
rect 2959 254241 3988 254359
rect 2400 254200 3988 254241
rect 295508 254359 297058 254400
rect 295508 254241 296499 254359
rect 296617 254241 297058 254359
rect 295508 254200 297058 254241
rect 0 252239 3988 252280
rect 0 252121 41 252239
rect 159 252121 3988 252239
rect 0 252080 3988 252121
rect 295508 252239 299458 252280
rect 295508 252121 299299 252239
rect 299417 252121 299458 252239
rect 295508 252080 299458 252121
rect 800 251279 3988 251320
rect 800 251161 841 251279
rect 959 251161 3988 251279
rect 800 251120 3988 251161
rect 295508 251279 298658 251320
rect 295508 251161 298499 251279
rect 298617 251161 298658 251279
rect 295508 251120 298658 251161
rect 1600 250319 3988 250360
rect 1600 250201 1641 250319
rect 1759 250201 3988 250319
rect 1600 250160 3988 250201
rect 295508 250319 297858 250360
rect 295508 250201 297699 250319
rect 297817 250201 297858 250319
rect 295508 250160 297858 250201
rect 2400 249359 3988 249400
rect 2400 249241 2441 249359
rect 2559 249241 3988 249359
rect 2400 249200 3988 249241
rect 295508 249359 297058 249400
rect 295508 249241 296899 249359
rect 297017 249241 297058 249359
rect 295508 249200 297058 249241
rect 0 247239 3988 247280
rect 0 247121 441 247239
rect 559 247121 3988 247239
rect 0 247080 3988 247121
rect 295508 247239 299458 247280
rect 295508 247121 298899 247239
rect 299017 247121 299458 247239
rect 295508 247080 299458 247121
rect 800 246279 3988 246320
rect 800 246161 1241 246279
rect 1359 246161 3988 246279
rect 800 246120 3988 246161
rect 295508 246279 298658 246320
rect 295508 246161 298099 246279
rect 298217 246161 298658 246279
rect 295508 246120 298658 246161
rect 1600 245319 3988 245360
rect 1600 245201 2041 245319
rect 2159 245201 3988 245319
rect 1600 245160 3988 245201
rect 295508 245319 297858 245360
rect 295508 245201 297299 245319
rect 297417 245201 297858 245319
rect 295508 245160 297858 245201
rect 2400 244359 3988 244400
rect 2400 244241 2841 244359
rect 2959 244241 3988 244359
rect 2400 244200 3988 244241
rect 295508 244359 297058 244400
rect 295508 244241 296499 244359
rect 296617 244241 297058 244359
rect 295508 244200 297058 244241
rect 0 242239 3988 242280
rect 0 242121 41 242239
rect 159 242121 3988 242239
rect 0 242080 3988 242121
rect 295508 242239 299458 242280
rect 295508 242121 299299 242239
rect 299417 242121 299458 242239
rect 295508 242080 299458 242121
rect 800 241279 3988 241320
rect 800 241161 841 241279
rect 959 241161 3988 241279
rect 800 241120 3988 241161
rect 295508 241279 298658 241320
rect 295508 241161 298499 241279
rect 298617 241161 298658 241279
rect 295508 241120 298658 241161
rect 1600 240319 3988 240360
rect 1600 240201 1641 240319
rect 1759 240201 3988 240319
rect 1600 240160 3988 240201
rect 295508 240319 297858 240360
rect 295508 240201 297699 240319
rect 297817 240201 297858 240319
rect 295508 240160 297858 240201
rect 2400 239359 3988 239400
rect 2400 239241 2441 239359
rect 2559 239241 3988 239359
rect 2400 239200 3988 239241
rect 295508 239359 297058 239400
rect 295508 239241 296899 239359
rect 297017 239241 297058 239359
rect 295508 239200 297058 239241
rect 0 237239 3988 237280
rect 0 237121 441 237239
rect 559 237121 3988 237239
rect 0 237080 3988 237121
rect 295508 237239 299458 237280
rect 295508 237121 298899 237239
rect 299017 237121 299458 237239
rect 295508 237080 299458 237121
rect 800 236279 3988 236320
rect 800 236161 1241 236279
rect 1359 236161 3988 236279
rect 800 236120 3988 236161
rect 295508 236279 298658 236320
rect 295508 236161 298099 236279
rect 298217 236161 298658 236279
rect 295508 236120 298658 236161
rect 1600 235319 3988 235360
rect 1600 235201 2041 235319
rect 2159 235201 3988 235319
rect 1600 235160 3988 235201
rect 295508 235319 297858 235360
rect 295508 235201 297299 235319
rect 297417 235201 297858 235319
rect 295508 235160 297858 235201
rect 2400 234359 3988 234400
rect 2400 234241 2841 234359
rect 2959 234241 3988 234359
rect 2400 234200 3988 234241
rect 295508 234359 297058 234400
rect 295508 234241 296499 234359
rect 296617 234241 297058 234359
rect 295508 234200 297058 234241
rect 0 232239 3988 232280
rect 0 232121 41 232239
rect 159 232121 3988 232239
rect 0 232080 3988 232121
rect 295508 232239 299458 232280
rect 295508 232121 299299 232239
rect 299417 232121 299458 232239
rect 295508 232080 299458 232121
rect 800 231279 3988 231320
rect 800 231161 841 231279
rect 959 231161 3988 231279
rect 800 231120 3988 231161
rect 295508 231279 298658 231320
rect 295508 231161 298499 231279
rect 298617 231161 298658 231279
rect 295508 231120 298658 231161
rect 1600 230319 3988 230360
rect 1600 230201 1641 230319
rect 1759 230201 3988 230319
rect 1600 230160 3988 230201
rect 295508 230319 297858 230360
rect 295508 230201 297699 230319
rect 297817 230201 297858 230319
rect 295508 230160 297858 230201
rect 2400 229359 3988 229400
rect 2400 229241 2441 229359
rect 2559 229241 3988 229359
rect 2400 229200 3988 229241
rect 295508 229359 297058 229400
rect 295508 229241 296899 229359
rect 297017 229241 297058 229359
rect 295508 229200 297058 229241
rect 0 227239 3988 227280
rect 0 227121 441 227239
rect 559 227121 3988 227239
rect 0 227080 3988 227121
rect 295508 227239 299458 227280
rect 295508 227121 298899 227239
rect 299017 227121 299458 227239
rect 295508 227080 299458 227121
rect 800 226279 3988 226320
rect 800 226161 1241 226279
rect 1359 226161 3988 226279
rect 800 226120 3988 226161
rect 295508 226279 298658 226320
rect 295508 226161 298099 226279
rect 298217 226161 298658 226279
rect 295508 226120 298658 226161
rect 1600 225319 3988 225360
rect 1600 225201 2041 225319
rect 2159 225201 3988 225319
rect 1600 225160 3988 225201
rect 295508 225319 297858 225360
rect 295508 225201 297299 225319
rect 297417 225201 297858 225319
rect 295508 225160 297858 225201
rect 2400 224359 3988 224400
rect 2400 224241 2841 224359
rect 2959 224241 3988 224359
rect 2400 224200 3988 224241
rect 295508 224359 297058 224400
rect 295508 224241 296499 224359
rect 296617 224241 297058 224359
rect 295508 224200 297058 224241
rect 0 222239 3988 222280
rect 0 222121 41 222239
rect 159 222121 3988 222239
rect 0 222080 3988 222121
rect 295508 222239 299458 222280
rect 295508 222121 299299 222239
rect 299417 222121 299458 222239
rect 295508 222080 299458 222121
rect 800 221279 3988 221320
rect 800 221161 841 221279
rect 959 221161 3988 221279
rect 800 221120 3988 221161
rect 295508 221279 298658 221320
rect 295508 221161 298499 221279
rect 298617 221161 298658 221279
rect 295508 221120 298658 221161
rect 1600 220319 3988 220360
rect 1600 220201 1641 220319
rect 1759 220201 3988 220319
rect 1600 220160 3988 220201
rect 295508 220319 297858 220360
rect 295508 220201 297699 220319
rect 297817 220201 297858 220319
rect 295508 220160 297858 220201
rect 2400 219359 3988 219400
rect 2400 219241 2441 219359
rect 2559 219241 3988 219359
rect 2400 219200 3988 219241
rect 295508 219359 297058 219400
rect 295508 219241 296899 219359
rect 297017 219241 297058 219359
rect 295508 219200 297058 219241
rect 0 217239 3988 217280
rect 0 217121 441 217239
rect 559 217121 3988 217239
rect 0 217080 3988 217121
rect 295508 217239 299458 217280
rect 295508 217121 298899 217239
rect 299017 217121 299458 217239
rect 295508 217080 299458 217121
rect 800 216279 3988 216320
rect 800 216161 1241 216279
rect 1359 216161 3988 216279
rect 800 216120 3988 216161
rect 295508 216279 298658 216320
rect 295508 216161 298099 216279
rect 298217 216161 298658 216279
rect 295508 216120 298658 216161
rect 1600 215319 3988 215360
rect 1600 215201 2041 215319
rect 2159 215201 3988 215319
rect 1600 215160 3988 215201
rect 295508 215319 297858 215360
rect 295508 215201 297299 215319
rect 297417 215201 297858 215319
rect 295508 215160 297858 215201
rect 2400 214359 3988 214400
rect 2400 214241 2841 214359
rect 2959 214241 3988 214359
rect 2400 214200 3988 214241
rect 295508 214359 297058 214400
rect 295508 214241 296499 214359
rect 296617 214241 297058 214359
rect 295508 214200 297058 214241
rect 0 212239 3988 212280
rect 0 212121 41 212239
rect 159 212121 3988 212239
rect 0 212080 3988 212121
rect 295508 212239 299458 212280
rect 295508 212121 299299 212239
rect 299417 212121 299458 212239
rect 295508 212080 299458 212121
rect 800 211279 3988 211320
rect 800 211161 841 211279
rect 959 211161 3988 211279
rect 800 211120 3988 211161
rect 295508 211279 298658 211320
rect 295508 211161 298499 211279
rect 298617 211161 298658 211279
rect 295508 211120 298658 211161
rect 1600 210319 3988 210360
rect 1600 210201 1641 210319
rect 1759 210201 3988 210319
rect 1600 210160 3988 210201
rect 295508 210319 297858 210360
rect 295508 210201 297699 210319
rect 297817 210201 297858 210319
rect 295508 210160 297858 210201
rect 2400 209359 3988 209400
rect 2400 209241 2441 209359
rect 2559 209241 3988 209359
rect 2400 209200 3988 209241
rect 295508 209359 297058 209400
rect 295508 209241 296899 209359
rect 297017 209241 297058 209359
rect 295508 209200 297058 209241
rect 0 207239 3988 207280
rect 0 207121 441 207239
rect 559 207121 3988 207239
rect 0 207080 3988 207121
rect 295508 207239 299458 207280
rect 295508 207121 298899 207239
rect 299017 207121 299458 207239
rect 295508 207080 299458 207121
rect 800 206279 3988 206320
rect 800 206161 1241 206279
rect 1359 206161 3988 206279
rect 800 206120 3988 206161
rect 295508 206279 298658 206320
rect 295508 206161 298099 206279
rect 298217 206161 298658 206279
rect 295508 206120 298658 206161
rect 1600 205319 3988 205360
rect 1600 205201 2041 205319
rect 2159 205201 3988 205319
rect 1600 205160 3988 205201
rect 295508 205319 297858 205360
rect 295508 205201 297299 205319
rect 297417 205201 297858 205319
rect 295508 205160 297858 205201
rect 2400 204359 3988 204400
rect 2400 204241 2841 204359
rect 2959 204241 3988 204359
rect 2400 204200 3988 204241
rect 295508 204359 297058 204400
rect 295508 204241 296499 204359
rect 296617 204241 297058 204359
rect 295508 204200 297058 204241
rect 0 202239 3988 202280
rect 0 202121 41 202239
rect 159 202121 3988 202239
rect 0 202080 3988 202121
rect 295508 202239 299458 202280
rect 295508 202121 299299 202239
rect 299417 202121 299458 202239
rect 295508 202080 299458 202121
rect 800 201279 3988 201320
rect 800 201161 841 201279
rect 959 201161 3988 201279
rect 800 201120 3988 201161
rect 295508 201279 298658 201320
rect 295508 201161 298499 201279
rect 298617 201161 298658 201279
rect 295508 201120 298658 201161
rect 1600 200319 3988 200360
rect 1600 200201 1641 200319
rect 1759 200201 3988 200319
rect 1600 200160 3988 200201
rect 295508 200319 297858 200360
rect 295508 200201 297699 200319
rect 297817 200201 297858 200319
rect 295508 200160 297858 200201
rect 2400 199359 3988 199400
rect 2400 199241 2441 199359
rect 2559 199241 3988 199359
rect 2400 199200 3988 199241
rect 295508 199359 297058 199400
rect 295508 199241 296899 199359
rect 297017 199241 297058 199359
rect 295508 199200 297058 199241
rect 0 197239 3988 197280
rect 0 197121 441 197239
rect 559 197121 3988 197239
rect 0 197080 3988 197121
rect 295508 197239 299458 197280
rect 295508 197121 298899 197239
rect 299017 197121 299458 197239
rect 295508 197080 299458 197121
rect 800 196279 3988 196320
rect 800 196161 1241 196279
rect 1359 196161 3988 196279
rect 800 196120 3988 196161
rect 295508 196279 298658 196320
rect 295508 196161 298099 196279
rect 298217 196161 298658 196279
rect 295508 196120 298658 196161
rect 1600 195319 3988 195360
rect 1600 195201 2041 195319
rect 2159 195201 3988 195319
rect 1600 195160 3988 195201
rect 295508 195319 297858 195360
rect 295508 195201 297299 195319
rect 297417 195201 297858 195319
rect 295508 195160 297858 195201
rect 2400 194359 3988 194400
rect 2400 194241 2841 194359
rect 2959 194241 3988 194359
rect 2400 194200 3988 194241
rect 295508 194359 297058 194400
rect 295508 194241 296499 194359
rect 296617 194241 297058 194359
rect 295508 194200 297058 194241
rect 0 192239 3988 192280
rect 0 192121 41 192239
rect 159 192121 3988 192239
rect 0 192080 3988 192121
rect 295508 192239 299458 192280
rect 295508 192121 299299 192239
rect 299417 192121 299458 192239
rect 295508 192080 299458 192121
rect 800 191279 3988 191320
rect 800 191161 841 191279
rect 959 191161 3988 191279
rect 800 191120 3988 191161
rect 295508 191279 298658 191320
rect 295508 191161 298499 191279
rect 298617 191161 298658 191279
rect 295508 191120 298658 191161
rect 1600 190319 3988 190360
rect 1600 190201 1641 190319
rect 1759 190201 3988 190319
rect 1600 190160 3988 190201
rect 295508 190319 297858 190360
rect 295508 190201 297699 190319
rect 297817 190201 297858 190319
rect 295508 190160 297858 190201
rect 2400 189359 3988 189400
rect 2400 189241 2441 189359
rect 2559 189241 3988 189359
rect 2400 189200 3988 189241
rect 295508 189359 297058 189400
rect 295508 189241 296899 189359
rect 297017 189241 297058 189359
rect 295508 189200 297058 189241
rect 0 187239 3988 187280
rect 0 187121 441 187239
rect 559 187121 3988 187239
rect 0 187080 3988 187121
rect 295508 187239 299458 187280
rect 295508 187121 298899 187239
rect 299017 187121 299458 187239
rect 295508 187080 299458 187121
rect 800 186279 3988 186320
rect 800 186161 1241 186279
rect 1359 186161 3988 186279
rect 800 186120 3988 186161
rect 295508 186279 298658 186320
rect 295508 186161 298099 186279
rect 298217 186161 298658 186279
rect 295508 186120 298658 186161
rect 1600 185319 3988 185360
rect 1600 185201 2041 185319
rect 2159 185201 3988 185319
rect 1600 185160 3988 185201
rect 295508 185319 297858 185360
rect 295508 185201 297299 185319
rect 297417 185201 297858 185319
rect 295508 185160 297858 185201
rect 2400 184359 3988 184400
rect 2400 184241 2841 184359
rect 2959 184241 3988 184359
rect 2400 184200 3988 184241
rect 295508 184359 297058 184400
rect 295508 184241 296499 184359
rect 296617 184241 297058 184359
rect 295508 184200 297058 184241
rect 0 182239 3988 182280
rect 0 182121 41 182239
rect 159 182121 3988 182239
rect 0 182080 3988 182121
rect 295508 182239 299458 182280
rect 295508 182121 299299 182239
rect 299417 182121 299458 182239
rect 295508 182080 299458 182121
rect 800 181279 3988 181320
rect 800 181161 841 181279
rect 959 181161 3988 181279
rect 800 181120 3988 181161
rect 295508 181279 298658 181320
rect 295508 181161 298499 181279
rect 298617 181161 298658 181279
rect 295508 181120 298658 181161
rect 1600 180319 3988 180360
rect 1600 180201 1641 180319
rect 1759 180201 3988 180319
rect 1600 180160 3988 180201
rect 295508 180319 297858 180360
rect 295508 180201 297699 180319
rect 297817 180201 297858 180319
rect 295508 180160 297858 180201
rect 2400 179359 3988 179400
rect 2400 179241 2441 179359
rect 2559 179241 3988 179359
rect 2400 179200 3988 179241
rect 295508 179359 297058 179400
rect 295508 179241 296899 179359
rect 297017 179241 297058 179359
rect 295508 179200 297058 179241
rect 0 177239 3988 177280
rect 0 177121 441 177239
rect 559 177121 3988 177239
rect 0 177080 3988 177121
rect 295508 177239 299458 177280
rect 295508 177121 298899 177239
rect 299017 177121 299458 177239
rect 295508 177080 299458 177121
rect 800 176279 3988 176320
rect 800 176161 1241 176279
rect 1359 176161 3988 176279
rect 800 176120 3988 176161
rect 295508 176279 298658 176320
rect 295508 176161 298099 176279
rect 298217 176161 298658 176279
rect 295508 176120 298658 176161
rect 1600 175319 3988 175360
rect 1600 175201 2041 175319
rect 2159 175201 3988 175319
rect 1600 175160 3988 175201
rect 295508 175319 297858 175360
rect 295508 175201 297299 175319
rect 297417 175201 297858 175319
rect 295508 175160 297858 175201
rect 2400 174359 3988 174400
rect 2400 174241 2841 174359
rect 2959 174241 3988 174359
rect 2400 174200 3988 174241
rect 295508 174359 297058 174400
rect 295508 174241 296499 174359
rect 296617 174241 297058 174359
rect 295508 174200 297058 174241
rect 0 172239 3988 172280
rect 0 172121 41 172239
rect 159 172121 3988 172239
rect 0 172080 3988 172121
rect 295508 172239 299458 172280
rect 295508 172121 299299 172239
rect 299417 172121 299458 172239
rect 295508 172080 299458 172121
rect 800 171279 3988 171320
rect 800 171161 841 171279
rect 959 171161 3988 171279
rect 800 171120 3988 171161
rect 295508 171279 298658 171320
rect 295508 171161 298499 171279
rect 298617 171161 298658 171279
rect 295508 171120 298658 171161
rect 1600 170319 3988 170360
rect 1600 170201 1641 170319
rect 1759 170201 3988 170319
rect 1600 170160 3988 170201
rect 295508 170319 297858 170360
rect 295508 170201 297699 170319
rect 297817 170201 297858 170319
rect 295508 170160 297858 170201
rect 2400 169359 3988 169400
rect 2400 169241 2441 169359
rect 2559 169241 3988 169359
rect 2400 169200 3988 169241
rect 295508 169359 297058 169400
rect 295508 169241 296899 169359
rect 297017 169241 297058 169359
rect 295508 169200 297058 169241
rect 0 167239 3988 167280
rect 0 167121 441 167239
rect 559 167121 3988 167239
rect 0 167080 3988 167121
rect 295508 167239 299458 167280
rect 295508 167121 298899 167239
rect 299017 167121 299458 167239
rect 295508 167080 299458 167121
rect 800 166279 3988 166320
rect 800 166161 1241 166279
rect 1359 166161 3988 166279
rect 800 166120 3988 166161
rect 295508 166279 298658 166320
rect 295508 166161 298099 166279
rect 298217 166161 298658 166279
rect 295508 166120 298658 166161
rect 1600 165319 3988 165360
rect 1600 165201 2041 165319
rect 2159 165201 3988 165319
rect 1600 165160 3988 165201
rect 295508 165319 297858 165360
rect 295508 165201 297299 165319
rect 297417 165201 297858 165319
rect 295508 165160 297858 165201
rect 2400 164359 3988 164400
rect 2400 164241 2841 164359
rect 2959 164241 3988 164359
rect 2400 164200 3988 164241
rect 295508 164359 297058 164400
rect 295508 164241 296499 164359
rect 296617 164241 297058 164359
rect 295508 164200 297058 164241
rect 0 162239 3988 162280
rect 0 162121 41 162239
rect 159 162121 3988 162239
rect 0 162080 3988 162121
rect 295508 162239 299458 162280
rect 295508 162121 299299 162239
rect 299417 162121 299458 162239
rect 295508 162080 299458 162121
rect 800 161279 3988 161320
rect 800 161161 841 161279
rect 959 161161 3988 161279
rect 800 161120 3988 161161
rect 295508 161279 298658 161320
rect 295508 161161 298499 161279
rect 298617 161161 298658 161279
rect 295508 161120 298658 161161
rect 1600 160319 3988 160360
rect 1600 160201 1641 160319
rect 1759 160201 3988 160319
rect 1600 160160 3988 160201
rect 295508 160319 297858 160360
rect 295508 160201 297699 160319
rect 297817 160201 297858 160319
rect 295508 160160 297858 160201
rect 2400 159359 3988 159400
rect 2400 159241 2441 159359
rect 2559 159241 3988 159359
rect 2400 159200 3988 159241
rect 295508 159359 297058 159400
rect 295508 159241 296899 159359
rect 297017 159241 297058 159359
rect 295508 159200 297058 159241
rect 0 157239 3988 157280
rect 0 157121 441 157239
rect 559 157121 3988 157239
rect 0 157080 3988 157121
rect 295508 157239 299458 157280
rect 295508 157121 298899 157239
rect 299017 157121 299458 157239
rect 295508 157080 299458 157121
rect 800 156279 3988 156320
rect 800 156161 1241 156279
rect 1359 156161 3988 156279
rect 800 156120 3988 156161
rect 295508 156279 298658 156320
rect 295508 156161 298099 156279
rect 298217 156161 298658 156279
rect 295508 156120 298658 156161
rect 1600 155319 3988 155360
rect 1600 155201 2041 155319
rect 2159 155201 3988 155319
rect 1600 155160 3988 155201
rect 295508 155319 297858 155360
rect 295508 155201 297299 155319
rect 297417 155201 297858 155319
rect 295508 155160 297858 155201
rect 2400 154359 3988 154400
rect 2400 154241 2841 154359
rect 2959 154241 3988 154359
rect 2400 154200 3988 154241
rect 295508 154359 297058 154400
rect 295508 154241 296499 154359
rect 296617 154241 297058 154359
rect 295508 154200 297058 154241
rect 0 152239 3988 152280
rect 0 152121 41 152239
rect 159 152121 3988 152239
rect 0 152080 3988 152121
rect 295508 152239 299458 152280
rect 295508 152121 299299 152239
rect 299417 152121 299458 152239
rect 295508 152080 299458 152121
rect 800 151279 3988 151320
rect 800 151161 841 151279
rect 959 151161 3988 151279
rect 800 151120 3988 151161
rect 295508 151279 298658 151320
rect 295508 151161 298499 151279
rect 298617 151161 298658 151279
rect 295508 151120 298658 151161
rect 1600 150319 3988 150360
rect 1600 150201 1641 150319
rect 1759 150201 3988 150319
rect 1600 150160 3988 150201
rect 295508 150319 297858 150360
rect 295508 150201 297699 150319
rect 297817 150201 297858 150319
rect 295508 150160 297858 150201
rect 2400 149359 3988 149400
rect 2400 149241 2441 149359
rect 2559 149241 3988 149359
rect 2400 149200 3988 149241
rect 295508 149359 297058 149400
rect 295508 149241 296899 149359
rect 297017 149241 297058 149359
rect 295508 149200 297058 149241
rect 0 147239 3988 147280
rect 0 147121 441 147239
rect 559 147121 3988 147239
rect 0 147080 3988 147121
rect 295508 147239 299458 147280
rect 295508 147121 298899 147239
rect 299017 147121 299458 147239
rect 295508 147080 299458 147121
rect 800 146279 3988 146320
rect 800 146161 1241 146279
rect 1359 146161 3988 146279
rect 800 146120 3988 146161
rect 295508 146279 298658 146320
rect 295508 146161 298099 146279
rect 298217 146161 298658 146279
rect 295508 146120 298658 146161
rect 1600 145319 3988 145360
rect 1600 145201 2041 145319
rect 2159 145201 3988 145319
rect 1600 145160 3988 145201
rect 295508 145319 297858 145360
rect 295508 145201 297299 145319
rect 297417 145201 297858 145319
rect 295508 145160 297858 145201
rect 2400 144359 3988 144400
rect 2400 144241 2841 144359
rect 2959 144241 3988 144359
rect 2400 144200 3988 144241
rect 295508 144359 297058 144400
rect 295508 144241 296499 144359
rect 296617 144241 297058 144359
rect 295508 144200 297058 144241
rect 0 142239 3988 142280
rect 0 142121 41 142239
rect 159 142121 3988 142239
rect 0 142080 3988 142121
rect 295508 142239 299458 142280
rect 295508 142121 299299 142239
rect 299417 142121 299458 142239
rect 295508 142080 299458 142121
rect 800 141279 3988 141320
rect 800 141161 841 141279
rect 959 141161 3988 141279
rect 800 141120 3988 141161
rect 295508 141279 298658 141320
rect 295508 141161 298499 141279
rect 298617 141161 298658 141279
rect 295508 141120 298658 141161
rect 1600 140319 3988 140360
rect 1600 140201 1641 140319
rect 1759 140201 3988 140319
rect 1600 140160 3988 140201
rect 295508 140319 297858 140360
rect 295508 140201 297699 140319
rect 297817 140201 297858 140319
rect 295508 140160 297858 140201
rect 2400 139359 3988 139400
rect 2400 139241 2441 139359
rect 2559 139241 3988 139359
rect 2400 139200 3988 139241
rect 295508 139359 297058 139400
rect 295508 139241 296899 139359
rect 297017 139241 297058 139359
rect 295508 139200 297058 139241
rect 0 137239 3988 137280
rect 0 137121 441 137239
rect 559 137121 3988 137239
rect 0 137080 3988 137121
rect 295508 137239 299458 137280
rect 295508 137121 298899 137239
rect 299017 137121 299458 137239
rect 295508 137080 299458 137121
rect 800 136279 3988 136320
rect 800 136161 1241 136279
rect 1359 136161 3988 136279
rect 800 136120 3988 136161
rect 295508 136279 298658 136320
rect 295508 136161 298099 136279
rect 298217 136161 298658 136279
rect 295508 136120 298658 136161
rect 1600 135319 3988 135360
rect 1600 135201 2041 135319
rect 2159 135201 3988 135319
rect 1600 135160 3988 135201
rect 295508 135319 297858 135360
rect 295508 135201 297299 135319
rect 297417 135201 297858 135319
rect 295508 135160 297858 135201
rect 2400 134359 3988 134400
rect 2400 134241 2841 134359
rect 2959 134241 3988 134359
rect 2400 134200 3988 134241
rect 295508 134359 297058 134400
rect 295508 134241 296499 134359
rect 296617 134241 297058 134359
rect 295508 134200 297058 134241
rect 0 132239 3988 132280
rect 0 132121 41 132239
rect 159 132121 3988 132239
rect 0 132080 3988 132121
rect 295508 132239 299458 132280
rect 295508 132121 299299 132239
rect 299417 132121 299458 132239
rect 295508 132080 299458 132121
rect 800 131279 3988 131320
rect 800 131161 841 131279
rect 959 131161 3988 131279
rect 800 131120 3988 131161
rect 295508 131279 298658 131320
rect 295508 131161 298499 131279
rect 298617 131161 298658 131279
rect 295508 131120 298658 131161
rect 1600 130319 3988 130360
rect 1600 130201 1641 130319
rect 1759 130201 3988 130319
rect 1600 130160 3988 130201
rect 295508 130319 297858 130360
rect 295508 130201 297699 130319
rect 297817 130201 297858 130319
rect 295508 130160 297858 130201
rect 2400 129359 3988 129400
rect 2400 129241 2441 129359
rect 2559 129241 3988 129359
rect 2400 129200 3988 129241
rect 295508 129359 297058 129400
rect 295508 129241 296899 129359
rect 297017 129241 297058 129359
rect 295508 129200 297058 129241
rect 0 127239 3988 127280
rect 0 127121 441 127239
rect 559 127121 3988 127239
rect 0 127080 3988 127121
rect 295508 127239 299458 127280
rect 295508 127121 298899 127239
rect 299017 127121 299458 127239
rect 295508 127080 299458 127121
rect 800 126279 3988 126320
rect 800 126161 1241 126279
rect 1359 126161 3988 126279
rect 800 126120 3988 126161
rect 295508 126279 298658 126320
rect 295508 126161 298099 126279
rect 298217 126161 298658 126279
rect 295508 126120 298658 126161
rect 1600 125319 3988 125360
rect 1600 125201 2041 125319
rect 2159 125201 3988 125319
rect 1600 125160 3988 125201
rect 295508 125319 297858 125360
rect 295508 125201 297299 125319
rect 297417 125201 297858 125319
rect 295508 125160 297858 125201
rect 2400 124359 3988 124400
rect 2400 124241 2841 124359
rect 2959 124241 3988 124359
rect 2400 124200 3988 124241
rect 295508 124359 297058 124400
rect 295508 124241 296499 124359
rect 296617 124241 297058 124359
rect 295508 124200 297058 124241
rect 0 122239 3988 122280
rect 0 122121 41 122239
rect 159 122121 3988 122239
rect 0 122080 3988 122121
rect 295508 122239 299458 122280
rect 295508 122121 299299 122239
rect 299417 122121 299458 122239
rect 295508 122080 299458 122121
rect 800 121279 3988 121320
rect 800 121161 841 121279
rect 959 121161 3988 121279
rect 800 121120 3988 121161
rect 295508 121279 298658 121320
rect 295508 121161 298499 121279
rect 298617 121161 298658 121279
rect 295508 121120 298658 121161
rect 1600 120319 3988 120360
rect 1600 120201 1641 120319
rect 1759 120201 3988 120319
rect 1600 120160 3988 120201
rect 295508 120319 297858 120360
rect 295508 120201 297699 120319
rect 297817 120201 297858 120319
rect 295508 120160 297858 120201
rect 2400 119359 3988 119400
rect 2400 119241 2441 119359
rect 2559 119241 3988 119359
rect 2400 119200 3988 119241
rect 295508 119359 297058 119400
rect 295508 119241 296899 119359
rect 297017 119241 297058 119359
rect 295508 119200 297058 119241
rect 0 117239 3988 117280
rect 0 117121 441 117239
rect 559 117121 3988 117239
rect 0 117080 3988 117121
rect 295508 117239 299458 117280
rect 295508 117121 298899 117239
rect 299017 117121 299458 117239
rect 295508 117080 299458 117121
rect 800 116279 3988 116320
rect 800 116161 1241 116279
rect 1359 116161 3988 116279
rect 800 116120 3988 116161
rect 295508 116279 298658 116320
rect 295508 116161 298099 116279
rect 298217 116161 298658 116279
rect 295508 116120 298658 116161
rect 1600 115319 3988 115360
rect 1600 115201 2041 115319
rect 2159 115201 3988 115319
rect 1600 115160 3988 115201
rect 295508 115319 297858 115360
rect 295508 115201 297299 115319
rect 297417 115201 297858 115319
rect 295508 115160 297858 115201
rect 2400 114359 3988 114400
rect 2400 114241 2841 114359
rect 2959 114241 3988 114359
rect 2400 114200 3988 114241
rect 295508 114359 297058 114400
rect 295508 114241 296499 114359
rect 296617 114241 297058 114359
rect 295508 114200 297058 114241
rect 0 112239 3988 112280
rect 0 112121 41 112239
rect 159 112121 3988 112239
rect 0 112080 3988 112121
rect 295508 112239 299458 112280
rect 295508 112121 299299 112239
rect 299417 112121 299458 112239
rect 295508 112080 299458 112121
rect 800 111279 3988 111320
rect 800 111161 841 111279
rect 959 111161 3988 111279
rect 800 111120 3988 111161
rect 295508 111279 298658 111320
rect 295508 111161 298499 111279
rect 298617 111161 298658 111279
rect 295508 111120 298658 111161
rect 1600 110319 3988 110360
rect 1600 110201 1641 110319
rect 1759 110201 3988 110319
rect 1600 110160 3988 110201
rect 295508 110319 297858 110360
rect 295508 110201 297699 110319
rect 297817 110201 297858 110319
rect 295508 110160 297858 110201
rect 2400 109359 3988 109400
rect 2400 109241 2441 109359
rect 2559 109241 3988 109359
rect 2400 109200 3988 109241
rect 295508 109359 297058 109400
rect 295508 109241 296899 109359
rect 297017 109241 297058 109359
rect 295508 109200 297058 109241
rect 0 107239 3988 107280
rect 0 107121 441 107239
rect 559 107121 3988 107239
rect 0 107080 3988 107121
rect 295508 107239 299458 107280
rect 295508 107121 298899 107239
rect 299017 107121 299458 107239
rect 295508 107080 299458 107121
rect 800 106279 3988 106320
rect 800 106161 1241 106279
rect 1359 106161 3988 106279
rect 800 106120 3988 106161
rect 295508 106279 298658 106320
rect 295508 106161 298099 106279
rect 298217 106161 298658 106279
rect 295508 106120 298658 106161
rect 1600 105319 3988 105360
rect 1600 105201 2041 105319
rect 2159 105201 3988 105319
rect 1600 105160 3988 105201
rect 295508 105319 297858 105360
rect 295508 105201 297299 105319
rect 297417 105201 297858 105319
rect 295508 105160 297858 105201
rect 2400 104359 3988 104400
rect 2400 104241 2841 104359
rect 2959 104241 3988 104359
rect 2400 104200 3988 104241
rect 295508 104359 297058 104400
rect 295508 104241 296499 104359
rect 296617 104241 297058 104359
rect 295508 104200 297058 104241
rect 0 102239 3988 102280
rect 0 102121 41 102239
rect 159 102121 3988 102239
rect 0 102080 3988 102121
rect 295508 102239 299458 102280
rect 295508 102121 299299 102239
rect 299417 102121 299458 102239
rect 295508 102080 299458 102121
rect 800 101279 3988 101320
rect 800 101161 841 101279
rect 959 101161 3988 101279
rect 800 101120 3988 101161
rect 295508 101279 298658 101320
rect 295508 101161 298499 101279
rect 298617 101161 298658 101279
rect 295508 101120 298658 101161
rect 1600 100319 3988 100360
rect 1600 100201 1641 100319
rect 1759 100201 3988 100319
rect 1600 100160 3988 100201
rect 295508 100319 297858 100360
rect 295508 100201 297699 100319
rect 297817 100201 297858 100319
rect 295508 100160 297858 100201
rect 2400 99359 3988 99400
rect 2400 99241 2441 99359
rect 2559 99241 3988 99359
rect 2400 99200 3988 99241
rect 295508 99359 297058 99400
rect 295508 99241 296899 99359
rect 297017 99241 297058 99359
rect 295508 99200 297058 99241
rect 0 97239 3988 97280
rect 0 97121 441 97239
rect 559 97121 3988 97239
rect 0 97080 3988 97121
rect 295508 97239 299458 97280
rect 295508 97121 298899 97239
rect 299017 97121 299458 97239
rect 295508 97080 299458 97121
rect 800 96279 3988 96320
rect 800 96161 1241 96279
rect 1359 96161 3988 96279
rect 800 96120 3988 96161
rect 295508 96279 298658 96320
rect 295508 96161 298099 96279
rect 298217 96161 298658 96279
rect 295508 96120 298658 96161
rect 1600 95319 3988 95360
rect 1600 95201 2041 95319
rect 2159 95201 3988 95319
rect 1600 95160 3988 95201
rect 295508 95319 297858 95360
rect 295508 95201 297299 95319
rect 297417 95201 297858 95319
rect 295508 95160 297858 95201
rect 2400 94359 3988 94400
rect 2400 94241 2841 94359
rect 2959 94241 3988 94359
rect 2400 94200 3988 94241
rect 295508 94359 297058 94400
rect 295508 94241 296499 94359
rect 296617 94241 297058 94359
rect 295508 94200 297058 94241
rect 0 92239 3988 92280
rect 0 92121 41 92239
rect 159 92121 3988 92239
rect 0 92080 3988 92121
rect 295508 92239 299458 92280
rect 295508 92121 299299 92239
rect 299417 92121 299458 92239
rect 295508 92080 299458 92121
rect 800 91279 3988 91320
rect 800 91161 841 91279
rect 959 91161 3988 91279
rect 800 91120 3988 91161
rect 295508 91279 298658 91320
rect 295508 91161 298499 91279
rect 298617 91161 298658 91279
rect 295508 91120 298658 91161
rect 1600 90319 3988 90360
rect 1600 90201 1641 90319
rect 1759 90201 3988 90319
rect 1600 90160 3988 90201
rect 295508 90319 297858 90360
rect 295508 90201 297699 90319
rect 297817 90201 297858 90319
rect 295508 90160 297858 90201
rect 2400 89359 3988 89400
rect 2400 89241 2441 89359
rect 2559 89241 3988 89359
rect 2400 89200 3988 89241
rect 295508 89359 297058 89400
rect 295508 89241 296899 89359
rect 297017 89241 297058 89359
rect 295508 89200 297058 89241
rect 0 87239 3988 87280
rect 0 87121 441 87239
rect 559 87121 3988 87239
rect 0 87080 3988 87121
rect 295508 87239 299458 87280
rect 295508 87121 298899 87239
rect 299017 87121 299458 87239
rect 295508 87080 299458 87121
rect 800 86279 3988 86320
rect 800 86161 1241 86279
rect 1359 86161 3988 86279
rect 800 86120 3988 86161
rect 295508 86279 298658 86320
rect 295508 86161 298099 86279
rect 298217 86161 298658 86279
rect 295508 86120 298658 86161
rect 1600 85319 3988 85360
rect 1600 85201 2041 85319
rect 2159 85201 3988 85319
rect 1600 85160 3988 85201
rect 295508 85319 297858 85360
rect 295508 85201 297299 85319
rect 297417 85201 297858 85319
rect 295508 85160 297858 85201
rect 2400 84359 3988 84400
rect 2400 84241 2841 84359
rect 2959 84241 3988 84359
rect 2400 84200 3988 84241
rect 295508 84359 297058 84400
rect 295508 84241 296499 84359
rect 296617 84241 297058 84359
rect 295508 84200 297058 84241
rect 0 82239 3988 82280
rect 0 82121 41 82239
rect 159 82121 3988 82239
rect 0 82080 3988 82121
rect 295508 82239 299458 82280
rect 295508 82121 299299 82239
rect 299417 82121 299458 82239
rect 295508 82080 299458 82121
rect 800 81279 3988 81320
rect 800 81161 841 81279
rect 959 81161 3988 81279
rect 800 81120 3988 81161
rect 295508 81279 298658 81320
rect 295508 81161 298499 81279
rect 298617 81161 298658 81279
rect 295508 81120 298658 81161
rect 1600 80319 3988 80360
rect 1600 80201 1641 80319
rect 1759 80201 3988 80319
rect 1600 80160 3988 80201
rect 295508 80319 297858 80360
rect 295508 80201 297699 80319
rect 297817 80201 297858 80319
rect 295508 80160 297858 80201
rect 2400 79359 3988 79400
rect 2400 79241 2441 79359
rect 2559 79241 3988 79359
rect 2400 79200 3988 79241
rect 295508 79359 297058 79400
rect 295508 79241 296899 79359
rect 297017 79241 297058 79359
rect 295508 79200 297058 79241
rect 0 77239 3988 77280
rect 0 77121 441 77239
rect 559 77121 3988 77239
rect 0 77080 3988 77121
rect 295508 77239 299458 77280
rect 295508 77121 298899 77239
rect 299017 77121 299458 77239
rect 295508 77080 299458 77121
rect 800 76279 3988 76320
rect 800 76161 1241 76279
rect 1359 76161 3988 76279
rect 800 76120 3988 76161
rect 295508 76279 298658 76320
rect 295508 76161 298099 76279
rect 298217 76161 298658 76279
rect 295508 76120 298658 76161
rect 1600 75319 3988 75360
rect 1600 75201 2041 75319
rect 2159 75201 3988 75319
rect 1600 75160 3988 75201
rect 295508 75319 297858 75360
rect 295508 75201 297299 75319
rect 297417 75201 297858 75319
rect 295508 75160 297858 75201
rect 2400 74359 3988 74400
rect 2400 74241 2841 74359
rect 2959 74241 3988 74359
rect 2400 74200 3988 74241
rect 295508 74359 297058 74400
rect 295508 74241 296499 74359
rect 296617 74241 297058 74359
rect 295508 74200 297058 74241
rect 0 72239 3988 72280
rect 0 72121 41 72239
rect 159 72121 3988 72239
rect 0 72080 3988 72121
rect 295508 72239 299458 72280
rect 295508 72121 299299 72239
rect 299417 72121 299458 72239
rect 295508 72080 299458 72121
rect 800 71279 3988 71320
rect 800 71161 841 71279
rect 959 71161 3988 71279
rect 800 71120 3988 71161
rect 295508 71279 298658 71320
rect 295508 71161 298499 71279
rect 298617 71161 298658 71279
rect 295508 71120 298658 71161
rect 1600 70319 3988 70360
rect 1600 70201 1641 70319
rect 1759 70201 3988 70319
rect 1600 70160 3988 70201
rect 295508 70319 297858 70360
rect 295508 70201 297699 70319
rect 297817 70201 297858 70319
rect 295508 70160 297858 70201
rect 2400 69359 3988 69400
rect 2400 69241 2441 69359
rect 2559 69241 3988 69359
rect 2400 69200 3988 69241
rect 295508 69359 297058 69400
rect 295508 69241 296899 69359
rect 297017 69241 297058 69359
rect 295508 69200 297058 69241
rect 0 67239 3988 67280
rect 0 67121 441 67239
rect 559 67121 3988 67239
rect 0 67080 3988 67121
rect 295508 67239 299458 67280
rect 295508 67121 298899 67239
rect 299017 67121 299458 67239
rect 295508 67080 299458 67121
rect 800 66279 3988 66320
rect 800 66161 1241 66279
rect 1359 66161 3988 66279
rect 800 66120 3988 66161
rect 295508 66279 298658 66320
rect 295508 66161 298099 66279
rect 298217 66161 298658 66279
rect 295508 66120 298658 66161
rect 1600 65319 3988 65360
rect 1600 65201 2041 65319
rect 2159 65201 3988 65319
rect 1600 65160 3988 65201
rect 295508 65319 297858 65360
rect 295508 65201 297299 65319
rect 297417 65201 297858 65319
rect 295508 65160 297858 65201
rect 2400 64359 3988 64400
rect 2400 64241 2841 64359
rect 2959 64241 3988 64359
rect 2400 64200 3988 64241
rect 295508 64359 297058 64400
rect 295508 64241 296499 64359
rect 296617 64241 297058 64359
rect 295508 64200 297058 64241
rect 0 62239 3988 62280
rect 0 62121 41 62239
rect 159 62121 3988 62239
rect 0 62080 3988 62121
rect 295508 62239 299458 62280
rect 295508 62121 299299 62239
rect 299417 62121 299458 62239
rect 295508 62080 299458 62121
rect 800 61279 3988 61320
rect 800 61161 841 61279
rect 959 61161 3988 61279
rect 800 61120 3988 61161
rect 295508 61279 298658 61320
rect 295508 61161 298499 61279
rect 298617 61161 298658 61279
rect 295508 61120 298658 61161
rect 1600 60319 3988 60360
rect 1600 60201 1641 60319
rect 1759 60201 3988 60319
rect 1600 60160 3988 60201
rect 295508 60319 297858 60360
rect 295508 60201 297699 60319
rect 297817 60201 297858 60319
rect 295508 60160 297858 60201
rect 2400 59359 3988 59400
rect 2400 59241 2441 59359
rect 2559 59241 3988 59359
rect 2400 59200 3988 59241
rect 295508 59359 297058 59400
rect 295508 59241 296899 59359
rect 297017 59241 297058 59359
rect 295508 59200 297058 59241
rect 0 57239 3988 57280
rect 0 57121 441 57239
rect 559 57121 3988 57239
rect 0 57080 3988 57121
rect 295508 57239 299458 57280
rect 295508 57121 298899 57239
rect 299017 57121 299458 57239
rect 295508 57080 299458 57121
rect 800 56279 3988 56320
rect 800 56161 1241 56279
rect 1359 56161 3988 56279
rect 800 56120 3988 56161
rect 295508 56279 298658 56320
rect 295508 56161 298099 56279
rect 298217 56161 298658 56279
rect 295508 56120 298658 56161
rect 1600 55319 3988 55360
rect 1600 55201 2041 55319
rect 2159 55201 3988 55319
rect 1600 55160 3988 55201
rect 295508 55319 297858 55360
rect 295508 55201 297299 55319
rect 297417 55201 297858 55319
rect 295508 55160 297858 55201
rect 2400 54359 3988 54400
rect 2400 54241 2841 54359
rect 2959 54241 3988 54359
rect 2400 54200 3988 54241
rect 295508 54359 297058 54400
rect 295508 54241 296499 54359
rect 296617 54241 297058 54359
rect 295508 54200 297058 54241
rect 0 52239 3988 52280
rect 0 52121 41 52239
rect 159 52121 3988 52239
rect 0 52080 3988 52121
rect 295508 52239 299458 52280
rect 295508 52121 299299 52239
rect 299417 52121 299458 52239
rect 295508 52080 299458 52121
rect 800 51279 3988 51320
rect 800 51161 841 51279
rect 959 51161 3988 51279
rect 800 51120 3988 51161
rect 295508 51279 298658 51320
rect 295508 51161 298499 51279
rect 298617 51161 298658 51279
rect 295508 51120 298658 51161
rect 1600 50319 3988 50360
rect 1600 50201 1641 50319
rect 1759 50201 3988 50319
rect 1600 50160 3988 50201
rect 295508 50319 297858 50360
rect 295508 50201 297699 50319
rect 297817 50201 297858 50319
rect 295508 50160 297858 50201
rect 2400 49359 3988 49400
rect 2400 49241 2441 49359
rect 2559 49241 3988 49359
rect 2400 49200 3988 49241
rect 295508 49359 297058 49400
rect 295508 49241 296899 49359
rect 297017 49241 297058 49359
rect 295508 49200 297058 49241
rect 0 47239 3988 47280
rect 0 47121 441 47239
rect 559 47121 3988 47239
rect 0 47080 3988 47121
rect 295508 47239 299458 47280
rect 295508 47121 298899 47239
rect 299017 47121 299458 47239
rect 295508 47080 299458 47121
rect 800 46279 3988 46320
rect 800 46161 1241 46279
rect 1359 46161 3988 46279
rect 800 46120 3988 46161
rect 295508 46279 298658 46320
rect 295508 46161 298099 46279
rect 298217 46161 298658 46279
rect 295508 46120 298658 46161
rect 1600 45319 3988 45360
rect 1600 45201 2041 45319
rect 2159 45201 3988 45319
rect 1600 45160 3988 45201
rect 295508 45319 297858 45360
rect 295508 45201 297299 45319
rect 297417 45201 297858 45319
rect 295508 45160 297858 45201
rect 2400 44359 3988 44400
rect 2400 44241 2841 44359
rect 2959 44241 3988 44359
rect 2400 44200 3988 44241
rect 295508 44359 297058 44400
rect 295508 44241 296499 44359
rect 296617 44241 297058 44359
rect 295508 44200 297058 44241
rect 0 42239 3988 42280
rect 0 42121 41 42239
rect 159 42121 3988 42239
rect 0 42080 3988 42121
rect 295508 42239 299458 42280
rect 295508 42121 299299 42239
rect 299417 42121 299458 42239
rect 295508 42080 299458 42121
rect 800 41279 3988 41320
rect 800 41161 841 41279
rect 959 41161 3988 41279
rect 800 41120 3988 41161
rect 295508 41279 298658 41320
rect 295508 41161 298499 41279
rect 298617 41161 298658 41279
rect 295508 41120 298658 41161
rect 1600 40319 3988 40360
rect 1600 40201 1641 40319
rect 1759 40201 3988 40319
rect 1600 40160 3988 40201
rect 295508 40319 297858 40360
rect 295508 40201 297699 40319
rect 297817 40201 297858 40319
rect 295508 40160 297858 40201
rect 2400 39359 3988 39400
rect 2400 39241 2441 39359
rect 2559 39241 3988 39359
rect 2400 39200 3988 39241
rect 295508 39359 297058 39400
rect 295508 39241 296899 39359
rect 297017 39241 297058 39359
rect 295508 39200 297058 39241
rect 0 37239 3988 37280
rect 0 37121 441 37239
rect 559 37121 3988 37239
rect 0 37080 3988 37121
rect 295508 37239 299458 37280
rect 295508 37121 298899 37239
rect 299017 37121 299458 37239
rect 295508 37080 299458 37121
rect 800 36279 3988 36320
rect 800 36161 1241 36279
rect 1359 36161 3988 36279
rect 800 36120 3988 36161
rect 295508 36279 298658 36320
rect 295508 36161 298099 36279
rect 298217 36161 298658 36279
rect 295508 36120 298658 36161
rect 1600 35319 3988 35360
rect 1600 35201 2041 35319
rect 2159 35201 3988 35319
rect 1600 35160 3988 35201
rect 295508 35319 297858 35360
rect 295508 35201 297299 35319
rect 297417 35201 297858 35319
rect 295508 35160 297858 35201
rect 2400 34359 3988 34400
rect 2400 34241 2841 34359
rect 2959 34241 3988 34359
rect 2400 34200 3988 34241
rect 295508 34359 297058 34400
rect 295508 34241 296499 34359
rect 296617 34241 297058 34359
rect 295508 34200 297058 34241
rect 0 32239 3988 32280
rect 0 32121 41 32239
rect 159 32121 3988 32239
rect 0 32080 3988 32121
rect 295508 32239 299458 32280
rect 295508 32121 299299 32239
rect 299417 32121 299458 32239
rect 295508 32080 299458 32121
rect 800 31279 3988 31320
rect 800 31161 841 31279
rect 959 31161 3988 31279
rect 800 31120 3988 31161
rect 295508 31279 298658 31320
rect 295508 31161 298499 31279
rect 298617 31161 298658 31279
rect 295508 31120 298658 31161
rect 1600 30319 3988 30360
rect 1600 30201 1641 30319
rect 1759 30201 3988 30319
rect 1600 30160 3988 30201
rect 295508 30319 297858 30360
rect 295508 30201 297699 30319
rect 297817 30201 297858 30319
rect 295508 30160 297858 30201
rect 2400 29359 3988 29400
rect 2400 29241 2441 29359
rect 2559 29241 3988 29359
rect 2400 29200 3988 29241
rect 295508 29359 297058 29400
rect 295508 29241 296899 29359
rect 297017 29241 297058 29359
rect 295508 29200 297058 29241
rect 0 27239 3988 27280
rect 0 27121 441 27239
rect 559 27121 3988 27239
rect 0 27080 3988 27121
rect 295508 27239 299458 27280
rect 295508 27121 298899 27239
rect 299017 27121 299458 27239
rect 295508 27080 299458 27121
rect 800 26279 3988 26320
rect 800 26161 1241 26279
rect 1359 26161 3988 26279
rect 800 26120 3988 26161
rect 295508 26279 298658 26320
rect 295508 26161 298099 26279
rect 298217 26161 298658 26279
rect 295508 26120 298658 26161
rect 1600 25319 3988 25360
rect 1600 25201 2041 25319
rect 2159 25201 3988 25319
rect 1600 25160 3988 25201
rect 295508 25319 297858 25360
rect 295508 25201 297299 25319
rect 297417 25201 297858 25319
rect 295508 25160 297858 25201
rect 2400 24359 3988 24400
rect 2400 24241 2841 24359
rect 2959 24241 3988 24359
rect 2400 24200 3988 24241
rect 295508 24359 297058 24400
rect 295508 24241 296499 24359
rect 296617 24241 297058 24359
rect 295508 24200 297058 24241
rect 0 22239 3988 22280
rect 0 22121 41 22239
rect 159 22121 3988 22239
rect 0 22080 3988 22121
rect 295508 22239 299458 22280
rect 295508 22121 299299 22239
rect 299417 22121 299458 22239
rect 295508 22080 299458 22121
rect 800 21279 3988 21320
rect 800 21161 841 21279
rect 959 21161 3988 21279
rect 800 21120 3988 21161
rect 295508 21279 298658 21320
rect 295508 21161 298499 21279
rect 298617 21161 298658 21279
rect 295508 21120 298658 21161
rect 1600 20319 3988 20360
rect 1600 20201 1641 20319
rect 1759 20201 3988 20319
rect 1600 20160 3988 20201
rect 295508 20319 297858 20360
rect 295508 20201 297699 20319
rect 297817 20201 297858 20319
rect 295508 20160 297858 20201
rect 2400 19359 3988 19400
rect 2400 19241 2441 19359
rect 2559 19241 3988 19359
rect 2400 19200 3988 19241
rect 295508 19359 297058 19400
rect 295508 19241 296899 19359
rect 297017 19241 297058 19359
rect 295508 19200 297058 19241
rect 0 17239 3988 17280
rect 0 17121 441 17239
rect 559 17121 3988 17239
rect 0 17080 3988 17121
rect 295508 17239 299458 17280
rect 295508 17121 298899 17239
rect 299017 17121 299458 17239
rect 295508 17080 299458 17121
rect 800 16279 3988 16320
rect 800 16161 1241 16279
rect 1359 16161 3988 16279
rect 800 16120 3988 16161
rect 295508 16279 298658 16320
rect 295508 16161 298099 16279
rect 298217 16161 298658 16279
rect 295508 16120 298658 16161
rect 1600 15319 3988 15360
rect 1600 15201 2041 15319
rect 2159 15201 3988 15319
rect 1600 15160 3988 15201
rect 295508 15319 297858 15360
rect 295508 15201 297299 15319
rect 297417 15201 297858 15319
rect 295508 15160 297858 15201
rect 2400 14359 3988 14400
rect 2400 14241 2841 14359
rect 2959 14241 3988 14359
rect 2400 14200 3988 14241
rect 295508 14359 297058 14400
rect 295508 14241 296499 14359
rect 296617 14241 297058 14359
rect 295508 14200 297058 14241
rect 0 12239 3988 12280
rect 0 12121 41 12239
rect 159 12121 3988 12239
rect 0 12080 3988 12121
rect 295508 12239 299458 12280
rect 295508 12121 299299 12239
rect 299417 12121 299458 12239
rect 295508 12080 299458 12121
rect 800 11279 3988 11320
rect 800 11161 841 11279
rect 959 11161 3988 11279
rect 800 11120 3988 11161
rect 295508 11279 298658 11320
rect 295508 11161 298499 11279
rect 298617 11161 298658 11279
rect 295508 11120 298658 11161
rect 1600 10319 3988 10360
rect 1600 10201 1641 10319
rect 1759 10201 3988 10319
rect 1600 10160 3988 10201
rect 295508 10319 297858 10360
rect 295508 10201 297699 10319
rect 297817 10201 297858 10319
rect 295508 10160 297858 10201
rect 2400 9359 3988 9400
rect 2400 9241 2441 9359
rect 2559 9241 3988 9359
rect 2400 9200 3988 9241
rect 295508 9359 297058 9400
rect 295508 9241 296899 9359
rect 297017 9241 297058 9359
rect 295508 9200 297058 9241
rect 0 7239 3988 7280
rect 0 7121 441 7239
rect 559 7121 3988 7239
rect 0 7080 3988 7121
rect 295508 7239 299458 7280
rect 295508 7121 298899 7239
rect 299017 7121 299458 7239
rect 295508 7080 299458 7121
rect 800 6279 3988 6320
rect 800 6161 1241 6279
rect 1359 6161 3988 6279
rect 800 6120 3988 6161
rect 295508 6279 298658 6320
rect 295508 6161 298099 6279
rect 298217 6161 298658 6279
rect 295508 6120 298658 6161
rect 1600 5319 3988 5360
rect 1600 5201 2041 5319
rect 2159 5201 3988 5319
rect 1600 5160 3988 5201
rect 295508 5319 297858 5360
rect 295508 5201 297299 5319
rect 297417 5201 297858 5319
rect 295508 5160 297858 5201
rect 2400 4359 3988 4400
rect 2400 4241 2841 4359
rect 2959 4241 3988 4359
rect 2400 4200 3988 4241
rect 295508 4359 297058 4400
rect 295508 4241 296499 4359
rect 296617 4241 297058 4359
rect 295508 4200 297058 4241
rect 2800 2959 296658 3000
rect 2800 2841 2841 2959
rect 2959 2841 4241 2959
rect 4359 2841 14241 2959
rect 14359 2841 24241 2959
rect 24359 2841 34241 2959
rect 34359 2841 44241 2959
rect 44359 2841 54241 2959
rect 54359 2841 64241 2959
rect 64359 2841 74241 2959
rect 74359 2841 84241 2959
rect 84359 2841 94241 2959
rect 94359 2841 104241 2959
rect 104359 2841 114241 2959
rect 114359 2841 124241 2959
rect 124359 2841 134241 2959
rect 134359 2841 144241 2959
rect 144359 2841 154241 2959
rect 154359 2841 164241 2959
rect 164359 2841 174241 2959
rect 174359 2841 184241 2959
rect 184359 2841 194241 2959
rect 194359 2841 204241 2959
rect 204359 2841 214241 2959
rect 214359 2841 224241 2959
rect 224359 2841 234241 2959
rect 234359 2841 244241 2959
rect 244359 2841 254241 2959
rect 254359 2841 264241 2959
rect 264359 2841 274241 2959
rect 274359 2841 284241 2959
rect 284359 2841 294241 2959
rect 294359 2841 296499 2959
rect 296617 2841 296658 2959
rect 2800 2800 296658 2841
rect 2400 2559 297058 2600
rect 2400 2441 2441 2559
rect 2559 2441 9241 2559
rect 9359 2441 19241 2559
rect 19359 2441 29241 2559
rect 29359 2441 39241 2559
rect 39359 2441 49241 2559
rect 49359 2441 59241 2559
rect 59359 2441 69241 2559
rect 69359 2441 79241 2559
rect 79359 2441 89241 2559
rect 89359 2441 99241 2559
rect 99359 2441 109241 2559
rect 109359 2441 119241 2559
rect 119359 2441 129241 2559
rect 129359 2441 139241 2559
rect 139359 2441 149241 2559
rect 149359 2441 159241 2559
rect 159359 2441 169241 2559
rect 169359 2441 179241 2559
rect 179359 2441 189241 2559
rect 189359 2441 199241 2559
rect 199359 2441 209241 2559
rect 209359 2441 219241 2559
rect 219359 2441 229241 2559
rect 229359 2441 239241 2559
rect 239359 2441 249241 2559
rect 249359 2441 259241 2559
rect 259359 2441 269241 2559
rect 269359 2441 279241 2559
rect 279359 2441 289241 2559
rect 289359 2441 296899 2559
rect 297017 2441 297058 2559
rect 2400 2400 297058 2441
rect 2000 2159 297458 2200
rect 2000 2041 2041 2159
rect 2159 2041 5201 2159
rect 5319 2041 15201 2159
rect 15319 2041 25201 2159
rect 25319 2041 35201 2159
rect 35319 2041 45201 2159
rect 45319 2041 55201 2159
rect 55319 2041 65201 2159
rect 65319 2041 75201 2159
rect 75319 2041 85201 2159
rect 85319 2041 95201 2159
rect 95319 2041 105201 2159
rect 105319 2041 115201 2159
rect 115319 2041 125201 2159
rect 125319 2041 135201 2159
rect 135319 2041 145201 2159
rect 145319 2041 155201 2159
rect 155319 2041 165201 2159
rect 165319 2041 175201 2159
rect 175319 2041 185201 2159
rect 185319 2041 195201 2159
rect 195319 2041 205201 2159
rect 205319 2041 215201 2159
rect 215319 2041 225201 2159
rect 225319 2041 235201 2159
rect 235319 2041 245201 2159
rect 245319 2041 255201 2159
rect 255319 2041 265201 2159
rect 265319 2041 275201 2159
rect 275319 2041 285201 2159
rect 285319 2041 297299 2159
rect 297417 2041 297458 2159
rect 2000 2000 297458 2041
rect 1600 1759 297858 1800
rect 1600 1641 1641 1759
rect 1759 1641 10201 1759
rect 10319 1641 20201 1759
rect 20319 1641 30201 1759
rect 30319 1641 40201 1759
rect 40319 1641 50201 1759
rect 50319 1641 60201 1759
rect 60319 1641 70201 1759
rect 70319 1641 80201 1759
rect 80319 1641 90201 1759
rect 90319 1641 100201 1759
rect 100319 1641 110201 1759
rect 110319 1641 120201 1759
rect 120319 1641 130201 1759
rect 130319 1641 140201 1759
rect 140319 1641 150201 1759
rect 150319 1641 160201 1759
rect 160319 1641 170201 1759
rect 170319 1641 180201 1759
rect 180319 1641 190201 1759
rect 190319 1641 200201 1759
rect 200319 1641 210201 1759
rect 210319 1641 220201 1759
rect 220319 1641 230201 1759
rect 230319 1641 240201 1759
rect 240319 1641 250201 1759
rect 250319 1641 260201 1759
rect 260319 1641 270201 1759
rect 270319 1641 280201 1759
rect 280319 1641 290201 1759
rect 290319 1641 297699 1759
rect 297817 1641 297858 1759
rect 1600 1600 297858 1641
rect 1200 1359 298258 1400
rect 1200 1241 1241 1359
rect 1359 1241 6161 1359
rect 6279 1241 16161 1359
rect 16279 1241 26161 1359
rect 26279 1241 36161 1359
rect 36279 1241 46161 1359
rect 46279 1241 56161 1359
rect 56279 1241 66161 1359
rect 66279 1241 76161 1359
rect 76279 1241 86161 1359
rect 86279 1241 96161 1359
rect 96279 1241 106161 1359
rect 106279 1241 116161 1359
rect 116279 1241 126161 1359
rect 126279 1241 136161 1359
rect 136279 1241 146161 1359
rect 146279 1241 156161 1359
rect 156279 1241 166161 1359
rect 166279 1241 176161 1359
rect 176279 1241 186161 1359
rect 186279 1241 196161 1359
rect 196279 1241 206161 1359
rect 206279 1241 216161 1359
rect 216279 1241 226161 1359
rect 226279 1241 236161 1359
rect 236279 1241 246161 1359
rect 246279 1241 256161 1359
rect 256279 1241 266161 1359
rect 266279 1241 276161 1359
rect 276279 1241 286161 1359
rect 286279 1241 298099 1359
rect 298217 1241 298258 1359
rect 1200 1200 298258 1241
rect 800 959 298658 1000
rect 800 841 841 959
rect 959 841 11161 959
rect 11279 841 21161 959
rect 21279 841 31161 959
rect 31279 841 41161 959
rect 41279 841 51161 959
rect 51279 841 61161 959
rect 61279 841 71161 959
rect 71279 841 81161 959
rect 81279 841 91161 959
rect 91279 841 101161 959
rect 101279 841 111161 959
rect 111279 841 121161 959
rect 121279 841 131161 959
rect 131279 841 141161 959
rect 141279 841 151161 959
rect 151279 841 161161 959
rect 161279 841 171161 959
rect 171279 841 181161 959
rect 181279 841 191161 959
rect 191279 841 201161 959
rect 201279 841 211161 959
rect 211279 841 221161 959
rect 221279 841 231161 959
rect 231279 841 241161 959
rect 241279 841 251161 959
rect 251279 841 261161 959
rect 261279 841 271161 959
rect 271279 841 281161 959
rect 281279 841 291161 959
rect 291279 841 298499 959
rect 298617 841 298658 959
rect 800 800 298658 841
rect 400 559 299058 600
rect 400 441 441 559
rect 559 441 7121 559
rect 7239 441 17121 559
rect 17239 441 27121 559
rect 27239 441 37121 559
rect 37239 441 47121 559
rect 47239 441 57121 559
rect 57239 441 67121 559
rect 67239 441 77121 559
rect 77239 441 87121 559
rect 87239 441 97121 559
rect 97239 441 107121 559
rect 107239 441 117121 559
rect 117239 441 127121 559
rect 127239 441 137121 559
rect 137239 441 147121 559
rect 147239 441 157121 559
rect 157239 441 167121 559
rect 167239 441 177121 559
rect 177239 441 187121 559
rect 187239 441 197121 559
rect 197239 441 207121 559
rect 207239 441 217121 559
rect 217239 441 227121 559
rect 227239 441 237121 559
rect 237239 441 247121 559
rect 247239 441 257121 559
rect 257239 441 267121 559
rect 267239 441 277121 559
rect 277239 441 287121 559
rect 287239 441 298899 559
rect 299017 441 299058 559
rect 400 400 299058 441
rect 0 159 299458 200
rect 0 41 41 159
rect 159 41 12121 159
rect 12239 41 22121 159
rect 22239 41 32121 159
rect 32239 41 42121 159
rect 42239 41 52121 159
rect 52239 41 62121 159
rect 62239 41 72121 159
rect 72239 41 82121 159
rect 82239 41 92121 159
rect 92239 41 102121 159
rect 102239 41 112121 159
rect 112239 41 122121 159
rect 122239 41 132121 159
rect 132239 41 142121 159
rect 142239 41 152121 159
rect 152239 41 162121 159
rect 162239 41 172121 159
rect 172239 41 182121 159
rect 182239 41 192121 159
rect 192239 41 202121 159
rect 202239 41 212121 159
rect 212239 41 222121 159
rect 222239 41 232121 159
rect 232239 41 242121 159
rect 242239 41 252121 159
rect 252239 41 262121 159
rect 262239 41 272121 159
rect 272239 41 282121 159
rect 282239 41 292121 159
rect 292239 41 299299 159
rect 299417 41 299458 159
rect 0 0 299458 41
use user_proj_example  mprj
timestamp 1606369131
transform 1 0 3748 0 1 3212
box 0 0 59876 60000
<< labels >>
rlabel metal3 s 295508 6140 295748 6200 4 analog_io[0]
port 1 nsew
rlabel metal3 s 295508 240740 295748 240800 4 analog_io[10]
port 2 nsew
rlabel metal3 s 295508 264200 295748 264260 4 analog_io[11]
port 3 nsew
rlabel metal3 s 295508 287660 295748 287720 4 analog_io[12]
port 4 nsew
rlabel metal3 s 295508 311120 295748 311180 4 analog_io[13]
port 5 nsew
rlabel metal3 s 295508 334580 295748 334640 4 analog_io[14]
port 6 nsew
rlabel metal2 s 291671 354972 291699 355212 4 analog_io[15]
port 7 nsew
rlabel metal2 s 259241 354972 259269 355212 4 analog_io[16]
port 8 nsew
rlabel metal2 s 226811 354972 226839 355212 4 analog_io[17]
port 9 nsew
rlabel metal2 s 194335 354972 194363 355212 4 analog_io[18]
port 10 nsew
rlabel metal2 s 161905 354972 161933 355212 4 analog_io[19]
port 11 nsew
rlabel metal3 s 295508 29600 295748 29660 4 analog_io[1]
port 12 nsew
rlabel metal2 s 129475 354972 129503 355212 4 analog_io[20]
port 13 nsew
rlabel metal2 s 96999 354972 97027 355212 4 analog_io[21]
port 14 nsew
rlabel metal2 s 64569 354972 64597 355212 4 analog_io[22]
port 15 nsew
rlabel metal2 s 32139 354972 32167 355212 4 analog_io[23]
port 16 nsew
rlabel metal3 s 3748 351512 3988 351572 4 analog_io[24]
port 17 nsew
rlabel metal3 s 3748 322748 3988 322808 4 analog_io[25]
port 18 nsew
rlabel metal3 s 3748 294052 3988 294112 4 analog_io[26]
port 19 nsew
rlabel metal3 s 3748 265288 3988 265348 4 analog_io[27]
port 20 nsew
rlabel metal3 s 3748 236592 3988 236652 4 analog_io[28]
port 21 nsew
rlabel metal3 s 3748 207828 3988 207888 4 analog_io[29]
port 22 nsew
rlabel metal3 s 295508 53060 295748 53120 4 analog_io[2]
port 23 nsew
rlabel metal3 s 3748 179132 3988 179192 4 analog_io[30]
port 24 nsew
rlabel metal3 s 295508 76520 295748 76580 4 analog_io[3]
port 25 nsew
rlabel metal3 s 295508 99980 295748 100040 4 analog_io[4]
port 26 nsew
rlabel metal3 s 295508 123440 295748 123500 4 analog_io[5]
port 27 nsew
rlabel metal3 s 295508 146900 295748 146960 4 analog_io[6]
port 28 nsew
rlabel metal3 s 295508 170360 295748 170420 4 analog_io[7]
port 29 nsew
rlabel metal3 s 295508 193820 295748 193880 4 analog_io[8]
port 30 nsew
rlabel metal3 s 295508 217280 295748 217340 4 analog_io[9]
port 31 nsew
rlabel metal3 s 295508 11988 295748 12048 4 io_in[0]
port 32 nsew
rlabel metal3 s 295508 246588 295748 246648 4 io_in[10]
port 33 nsew
rlabel metal3 s 295508 270116 295748 270176 4 io_in[11]
port 34 nsew
rlabel metal3 s 295508 293576 295748 293636 4 io_in[12]
port 35 nsew
rlabel metal3 s 295508 317036 295748 317096 4 io_in[13]
port 36 nsew
rlabel metal3 s 295508 340496 295748 340556 4 io_in[14]
port 37 nsew
rlabel metal2 s 283575 354972 283603 355212 4 io_in[15]
port 38 nsew
rlabel metal2 s 251145 354972 251173 355212 4 io_in[16]
port 39 nsew
rlabel metal2 s 218669 354972 218697 355212 4 io_in[17]
port 40 nsew
rlabel metal2 s 186239 354972 186267 355212 4 io_in[18]
port 41 nsew
rlabel metal2 s 153809 354972 153837 355212 4 io_in[19]
port 42 nsew
rlabel metal3 s 295508 35448 295748 35508 4 io_in[1]
port 43 nsew
rlabel metal2 s 121333 354972 121361 355212 4 io_in[20]
port 44 nsew
rlabel metal2 s 88903 354972 88931 355212 4 io_in[21]
port 45 nsew
rlabel metal2 s 56473 354972 56501 355212 4 io_in[22]
port 46 nsew
rlabel metal2 s 23997 354972 24025 355212 4 io_in[23]
port 47 nsew
rlabel metal3 s 3748 344304 3988 344364 4 io_in[24]
port 48 nsew
rlabel metal3 s 3748 315608 3988 315668 4 io_in[25]
port 49 nsew
rlabel metal3 s 3748 286844 3988 286904 4 io_in[26]
port 50 nsew
rlabel metal3 s 3748 258148 3988 258208 4 io_in[27]
port 51 nsew
rlabel metal3 s 3748 229384 3988 229444 4 io_in[28]
port 52 nsew
rlabel metal3 s 3748 200688 3988 200748 4 io_in[29]
port 53 nsew
rlabel metal3 s 295508 58908 295748 58968 4 io_in[2]
port 54 nsew
rlabel metal3 s 3748 171924 3988 171984 4 io_in[30]
port 55 nsew
rlabel metal3 s 3748 150368 3988 150428 4 io_in[31]
port 56 nsew
rlabel metal3 s 3748 128812 3988 128872 4 io_in[32]
port 57 nsew
rlabel metal3 s 3748 107256 3988 107316 4 io_in[33]
port 58 nsew
rlabel metal3 s 3748 85700 3988 85760 4 io_in[34]
port 59 nsew
rlabel metal3 s 3748 64212 3988 64272 4 io_in[35]
port 60 nsew
rlabel metal3 s 3748 42656 3988 42716 4 io_in[36]
port 61 nsew
rlabel metal3 s 3748 21100 3988 21160 4 io_in[37]
port 62 nsew
rlabel metal3 s 295508 82368 295748 82428 4 io_in[3]
port 63 nsew
rlabel metal3 s 295508 105828 295748 105888 4 io_in[4]
port 64 nsew
rlabel metal3 s 295508 129288 295748 129348 4 io_in[5]
port 65 nsew
rlabel metal3 s 295508 152748 295748 152808 4 io_in[6]
port 66 nsew
rlabel metal3 s 295508 176208 295748 176268 4 io_in[7]
port 67 nsew
rlabel metal3 s 295508 199668 295748 199728 4 io_in[8]
port 68 nsew
rlabel metal3 s 295508 223128 295748 223188 4 io_in[9]
port 69 nsew
rlabel metal3 s 295508 23684 295748 23744 4 io_oeb[0]
port 70 nsew
rlabel metal3 s 295508 258352 295748 258412 4 io_oeb[10]
port 71 nsew
rlabel metal3 s 295508 281812 295748 281872 4 io_oeb[11]
port 72 nsew
rlabel metal3 s 295508 305272 295748 305332 4 io_oeb[12]
port 73 nsew
rlabel metal3 s 295508 328732 295748 328792 4 io_oeb[13]
port 74 nsew
rlabel metal3 s 295508 352192 295748 352252 4 io_oeb[14]
port 75 nsew
rlabel metal2 s 267337 354972 267365 355212 4 io_oeb[15]
port 76 nsew
rlabel metal2 s 234907 354972 234935 355212 4 io_oeb[16]
port 77 nsew
rlabel metal2 s 202477 354972 202505 355212 4 io_oeb[17]
port 78 nsew
rlabel metal2 s 170001 354972 170029 355212 4 io_oeb[18]
port 79 nsew
rlabel metal2 s 137571 354972 137599 355212 4 io_oeb[19]
port 80 nsew
rlabel metal3 s 295508 47144 295748 47204 4 io_oeb[1]
port 81 nsew
rlabel metal2 s 105141 354972 105169 355212 4 io_oeb[20]
port 82 nsew
rlabel metal2 s 72665 354972 72693 355212 4 io_oeb[21]
port 83 nsew
rlabel metal2 s 40235 354972 40263 355212 4 io_oeb[22]
port 84 nsew
rlabel metal2 s 7805 354972 7833 355212 4 io_oeb[23]
port 85 nsew
rlabel metal3 s 3748 329956 3988 330016 4 io_oeb[24]
port 86 nsew
rlabel metal3 s 3748 301192 3988 301252 4 io_oeb[25]
port 87 nsew
rlabel metal3 s 3748 272496 3988 272556 4 io_oeb[26]
port 88 nsew
rlabel metal3 s 3748 243732 3988 243792 4 io_oeb[27]
port 89 nsew
rlabel metal3 s 3748 215036 3988 215096 4 io_oeb[28]
port 90 nsew
rlabel metal3 s 3748 186272 3988 186332 4 io_oeb[29]
port 91 nsew
rlabel metal3 s 295508 70604 295748 70664 4 io_oeb[2]
port 92 nsew
rlabel metal3 s 3748 157576 3988 157636 4 io_oeb[30]
port 93 nsew
rlabel metal3 s 3748 136020 3988 136080 4 io_oeb[31]
port 94 nsew
rlabel metal3 s 3748 114464 3988 114524 4 io_oeb[32]
port 95 nsew
rlabel metal3 s 3748 92908 3988 92968 4 io_oeb[33]
port 96 nsew
rlabel metal3 s 3748 71352 3988 71412 4 io_oeb[34]
port 97 nsew
rlabel metal3 s 3748 49796 3988 49856 4 io_oeb[35]
port 98 nsew
rlabel metal3 s 3748 28240 3988 28300 4 io_oeb[36]
port 99 nsew
rlabel metal3 s 3748 6752 3988 6812 4 io_oeb[37]
port 100 nsew
rlabel metal3 s 295508 94132 295748 94192 4 io_oeb[3]
port 101 nsew
rlabel metal3 s 295508 117592 295748 117652 4 io_oeb[4]
port 102 nsew
rlabel metal3 s 295508 141052 295748 141112 4 io_oeb[5]
port 103 nsew
rlabel metal3 s 295508 164512 295748 164572 4 io_oeb[6]
port 104 nsew
rlabel metal3 s 295508 187972 295748 188032 4 io_oeb[7]
port 105 nsew
rlabel metal3 s 295508 211432 295748 211492 4 io_oeb[8]
port 106 nsew
rlabel metal3 s 295508 234892 295748 234952 4 io_oeb[9]
port 107 nsew
rlabel metal3 s 295508 17836 295748 17896 4 io_out[0]
port 108 nsew
rlabel metal3 s 295508 252504 295748 252564 4 io_out[10]
port 109 nsew
rlabel metal3 s 295508 275964 295748 276024 4 io_out[11]
port 110 nsew
rlabel metal3 s 295508 299424 295748 299484 4 io_out[12]
port 111 nsew
rlabel metal3 s 295508 322884 295748 322944 4 io_out[13]
port 112 nsew
rlabel metal3 s 295508 346344 295748 346404 4 io_out[14]
port 113 nsew
rlabel metal2 s 275479 354972 275507 355212 4 io_out[15]
port 114 nsew
rlabel metal2 s 243003 354972 243031 355212 4 io_out[16]
port 115 nsew
rlabel metal2 s 210573 354972 210601 355212 4 io_out[17]
port 116 nsew
rlabel metal2 s 178143 354972 178171 355212 4 io_out[18]
port 117 nsew
rlabel metal2 s 145667 354972 145695 355212 4 io_out[19]
port 118 nsew
rlabel metal3 s 295508 41296 295748 41356 4 io_out[1]
port 119 nsew
rlabel metal2 s 113237 354972 113265 355212 4 io_out[20]
port 120 nsew
rlabel metal2 s 80807 354972 80835 355212 4 io_out[21]
port 121 nsew
rlabel metal2 s 48331 354972 48359 355212 4 io_out[22]
port 122 nsew
rlabel metal2 s 15901 354972 15929 355212 4 io_out[23]
port 123 nsew
rlabel metal3 s 3748 337164 3988 337224 4 io_out[24]
port 124 nsew
rlabel metal3 s 3748 308400 3988 308460 4 io_out[25]
port 125 nsew
rlabel metal3 s 3748 279704 3988 279764 4 io_out[26]
port 126 nsew
rlabel metal3 s 3748 250940 3988 251000 4 io_out[27]
port 127 nsew
rlabel metal3 s 3748 222176 3988 222236 4 io_out[28]
port 128 nsew
rlabel metal3 s 3748 193480 3988 193540 4 io_out[29]
port 129 nsew
rlabel metal3 s 295508 64756 295748 64816 4 io_out[2]
port 130 nsew
rlabel metal3 s 3748 164716 3988 164776 4 io_out[30]
port 131 nsew
rlabel metal3 s 3748 143228 3988 143288 4 io_out[31]
port 132 nsew
rlabel metal3 s 3748 121672 3988 121732 4 io_out[32]
port 133 nsew
rlabel metal3 s 3748 100116 3988 100176 4 io_out[33]
port 134 nsew
rlabel metal3 s 3748 78560 3988 78620 4 io_out[34]
port 135 nsew
rlabel metal3 s 3748 57004 3988 57064 4 io_out[35]
port 136 nsew
rlabel metal3 s 3748 35448 3988 35508 4 io_out[36]
port 137 nsew
rlabel metal3 s 3748 13892 3988 13952 4 io_out[37]
port 138 nsew
rlabel metal3 s 295508 88216 295748 88276 4 io_out[3]
port 139 nsew
rlabel metal3 s 295508 111676 295748 111736 4 io_out[4]
port 140 nsew
rlabel metal3 s 295508 135136 295748 135196 4 io_out[5]
port 141 nsew
rlabel metal3 s 295508 158596 295748 158656 4 io_out[6]
port 142 nsew
rlabel metal3 s 295508 182124 295748 182184 4 io_out[7]
port 143 nsew
rlabel metal3 s 295508 205584 295748 205644 4 io_out[8]
port 144 nsew
rlabel metal3 s 295508 229044 295748 229104 4 io_out[9]
port 145 nsew
rlabel metal2 s 67053 3212 67081 3452 4 la_data_in[0]
port 146 nsew
rlabel metal2 s 245487 3212 245515 3452 4 la_data_in[100]
port 147 nsew
rlabel metal2 s 247235 3212 247263 3452 4 la_data_in[101]
port 148 nsew
rlabel metal2 s 249029 3212 249057 3452 4 la_data_in[102]
port 149 nsew
rlabel metal2 s 250823 3212 250851 3452 4 la_data_in[103]
port 150 nsew
rlabel metal2 s 252617 3212 252645 3452 4 la_data_in[104]
port 151 nsew
rlabel metal2 s 254365 3212 254393 3452 4 la_data_in[105]
port 152 nsew
rlabel metal2 s 256159 3212 256187 3452 4 la_data_in[106]
port 153 nsew
rlabel metal2 s 257953 3212 257981 3452 4 la_data_in[107]
port 154 nsew
rlabel metal2 s 259747 3212 259775 3452 4 la_data_in[108]
port 155 nsew
rlabel metal2 s 261541 3212 261569 3452 4 la_data_in[109]
port 156 nsew
rlabel metal2 s 84901 3212 84929 3452 4 la_data_in[10]
port 157 nsew
rlabel metal2 s 263289 3212 263317 3452 4 la_data_in[110]
port 158 nsew
rlabel metal2 s 265083 3212 265111 3452 4 la_data_in[111]
port 159 nsew
rlabel metal2 s 266877 3212 266905 3452 4 la_data_in[112]
port 160 nsew
rlabel metal2 s 268671 3212 268699 3452 4 la_data_in[113]
port 161 nsew
rlabel metal2 s 270465 3212 270493 3452 4 la_data_in[114]
port 162 nsew
rlabel metal2 s 272213 3212 272241 3452 4 la_data_in[115]
port 163 nsew
rlabel metal2 s 274007 3212 274035 3452 4 la_data_in[116]
port 164 nsew
rlabel metal2 s 275801 3212 275829 3452 4 la_data_in[117]
port 165 nsew
rlabel metal2 s 277595 3212 277623 3452 4 la_data_in[118]
port 166 nsew
rlabel metal2 s 279343 3212 279371 3452 4 la_data_in[119]
port 167 nsew
rlabel metal2 s 86695 3212 86723 3452 4 la_data_in[11]
port 168 nsew
rlabel metal2 s 281137 3212 281165 3452 4 la_data_in[120]
port 169 nsew
rlabel metal2 s 282931 3212 282959 3452 4 la_data_in[121]
port 170 nsew
rlabel metal2 s 284725 3212 284753 3452 4 la_data_in[122]
port 171 nsew
rlabel metal2 s 286519 3212 286547 3452 4 la_data_in[123]
port 172 nsew
rlabel metal2 s 288267 3212 288295 3452 4 la_data_in[124]
port 173 nsew
rlabel metal2 s 290061 3212 290089 3452 4 la_data_in[125]
port 174 nsew
rlabel metal2 s 291855 3212 291883 3452 4 la_data_in[126]
port 175 nsew
rlabel metal2 s 293649 3212 293677 3452 4 la_data_in[127]
port 176 nsew
rlabel metal2 s 88443 3212 88471 3452 4 la_data_in[12]
port 177 nsew
rlabel metal2 s 90237 3212 90265 3452 4 la_data_in[13]
port 178 nsew
rlabel metal2 s 92031 3212 92059 3452 4 la_data_in[14]
port 179 nsew
rlabel metal2 s 93825 3212 93853 3452 4 la_data_in[15]
port 180 nsew
rlabel metal2 s 95619 3212 95647 3452 4 la_data_in[16]
port 181 nsew
rlabel metal2 s 97367 3212 97395 3452 4 la_data_in[17]
port 182 nsew
rlabel metal2 s 99161 3212 99189 3452 4 la_data_in[18]
port 183 nsew
rlabel metal2 s 100955 3212 100983 3452 4 la_data_in[19]
port 184 nsew
rlabel metal2 s 68847 3212 68875 3452 4 la_data_in[1]
port 185 nsew
rlabel metal2 s 102749 3212 102777 3452 4 la_data_in[20]
port 186 nsew
rlabel metal2 s 104497 3212 104525 3452 4 la_data_in[21]
port 187 nsew
rlabel metal2 s 106291 3212 106319 3452 4 la_data_in[22]
port 188 nsew
rlabel metal2 s 108085 3212 108113 3452 4 la_data_in[23]
port 189 nsew
rlabel metal2 s 109879 3212 109907 3452 4 la_data_in[24]
port 190 nsew
rlabel metal2 s 111673 3212 111701 3452 4 la_data_in[25]
port 191 nsew
rlabel metal2 s 113421 3212 113449 3452 4 la_data_in[26]
port 192 nsew
rlabel metal2 s 115215 3212 115243 3452 4 la_data_in[27]
port 193 nsew
rlabel metal2 s 117009 3212 117037 3452 4 la_data_in[28]
port 194 nsew
rlabel metal2 s 118803 3212 118831 3452 4 la_data_in[29]
port 195 nsew
rlabel metal2 s 70641 3212 70669 3452 4 la_data_in[2]
port 196 nsew
rlabel metal2 s 120597 3212 120625 3452 4 la_data_in[30]
port 197 nsew
rlabel metal2 s 122345 3212 122373 3452 4 la_data_in[31]
port 198 nsew
rlabel metal2 s 124139 3212 124167 3452 4 la_data_in[32]
port 199 nsew
rlabel metal2 s 125933 3212 125961 3452 4 la_data_in[33]
port 200 nsew
rlabel metal2 s 127727 3212 127755 3452 4 la_data_in[34]
port 201 nsew
rlabel metal2 s 129475 3212 129503 3452 4 la_data_in[35]
port 202 nsew
rlabel metal2 s 131269 3212 131297 3452 4 la_data_in[36]
port 203 nsew
rlabel metal2 s 133063 3212 133091 3452 4 la_data_in[37]
port 204 nsew
rlabel metal2 s 134857 3212 134885 3452 4 la_data_in[38]
port 205 nsew
rlabel metal2 s 136651 3212 136679 3452 4 la_data_in[39]
port 206 nsew
rlabel metal2 s 72389 3212 72417 3452 4 la_data_in[3]
port 207 nsew
rlabel metal2 s 138399 3212 138427 3452 4 la_data_in[40]
port 208 nsew
rlabel metal2 s 140193 3212 140221 3452 4 la_data_in[41]
port 209 nsew
rlabel metal2 s 141987 3212 142015 3452 4 la_data_in[42]
port 210 nsew
rlabel metal2 s 143781 3212 143809 3452 4 la_data_in[43]
port 211 nsew
rlabel metal2 s 145575 3212 145603 3452 4 la_data_in[44]
port 212 nsew
rlabel metal2 s 147323 3212 147351 3452 4 la_data_in[45]
port 213 nsew
rlabel metal2 s 149117 3212 149145 3452 4 la_data_in[46]
port 214 nsew
rlabel metal2 s 150911 3212 150939 3452 4 la_data_in[47]
port 215 nsew
rlabel metal2 s 152705 3212 152733 3452 4 la_data_in[48]
port 216 nsew
rlabel metal2 s 154453 3212 154481 3452 4 la_data_in[49]
port 217 nsew
rlabel metal2 s 74183 3212 74211 3452 4 la_data_in[4]
port 218 nsew
rlabel metal2 s 156247 3212 156275 3452 4 la_data_in[50]
port 219 nsew
rlabel metal2 s 158041 3212 158069 3452 4 la_data_in[51]
port 220 nsew
rlabel metal2 s 159835 3212 159863 3452 4 la_data_in[52]
port 221 nsew
rlabel metal2 s 161629 3212 161657 3452 4 la_data_in[53]
port 222 nsew
rlabel metal2 s 163377 3212 163405 3452 4 la_data_in[54]
port 223 nsew
rlabel metal2 s 165171 3212 165199 3452 4 la_data_in[55]
port 224 nsew
rlabel metal2 s 166965 3212 166993 3452 4 la_data_in[56]
port 225 nsew
rlabel metal2 s 168759 3212 168787 3452 4 la_data_in[57]
port 226 nsew
rlabel metal2 s 170553 3212 170581 3452 4 la_data_in[58]
port 227 nsew
rlabel metal2 s 172301 3212 172329 3452 4 la_data_in[59]
port 228 nsew
rlabel metal2 s 75977 3212 76005 3452 4 la_data_in[5]
port 229 nsew
rlabel metal2 s 174095 3212 174123 3452 4 la_data_in[60]
port 230 nsew
rlabel metal2 s 175889 3212 175917 3452 4 la_data_in[61]
port 231 nsew
rlabel metal2 s 177683 3212 177711 3452 4 la_data_in[62]
port 232 nsew
rlabel metal2 s 179431 3212 179459 3452 4 la_data_in[63]
port 233 nsew
rlabel metal2 s 181225 3212 181253 3452 4 la_data_in[64]
port 234 nsew
rlabel metal2 s 183019 3212 183047 3452 4 la_data_in[65]
port 235 nsew
rlabel metal2 s 184813 3212 184841 3452 4 la_data_in[66]
port 236 nsew
rlabel metal2 s 186607 3212 186635 3452 4 la_data_in[67]
port 237 nsew
rlabel metal2 s 188355 3212 188383 3452 4 la_data_in[68]
port 238 nsew
rlabel metal2 s 190149 3212 190177 3452 4 la_data_in[69]
port 239 nsew
rlabel metal2 s 77771 3212 77799 3452 4 la_data_in[6]
port 240 nsew
rlabel metal2 s 191943 3212 191971 3452 4 la_data_in[70]
port 241 nsew
rlabel metal2 s 193737 3212 193765 3452 4 la_data_in[71]
port 242 nsew
rlabel metal2 s 195531 3212 195559 3452 4 la_data_in[72]
port 243 nsew
rlabel metal2 s 197279 3212 197307 3452 4 la_data_in[73]
port 244 nsew
rlabel metal2 s 199073 3212 199101 3452 4 la_data_in[74]
port 245 nsew
rlabel metal2 s 200867 3212 200895 3452 4 la_data_in[75]
port 246 nsew
rlabel metal2 s 202661 3212 202689 3452 4 la_data_in[76]
port 247 nsew
rlabel metal2 s 204409 3212 204437 3452 4 la_data_in[77]
port 248 nsew
rlabel metal2 s 206203 3212 206231 3452 4 la_data_in[78]
port 249 nsew
rlabel metal2 s 207997 3212 208025 3452 4 la_data_in[79]
port 250 nsew
rlabel metal2 s 79519 3212 79547 3452 4 la_data_in[7]
port 251 nsew
rlabel metal2 s 209791 3212 209819 3452 4 la_data_in[80]
port 252 nsew
rlabel metal2 s 211585 3212 211613 3452 4 la_data_in[81]
port 253 nsew
rlabel metal2 s 213333 3212 213361 3452 4 la_data_in[82]
port 254 nsew
rlabel metal2 s 215127 3212 215155 3452 4 la_data_in[83]
port 255 nsew
rlabel metal2 s 216921 3212 216949 3452 4 la_data_in[84]
port 256 nsew
rlabel metal2 s 218715 3212 218743 3452 4 la_data_in[85]
port 257 nsew
rlabel metal2 s 220509 3212 220537 3452 4 la_data_in[86]
port 258 nsew
rlabel metal2 s 222257 3212 222285 3452 4 la_data_in[87]
port 259 nsew
rlabel metal2 s 224051 3212 224079 3452 4 la_data_in[88]
port 260 nsew
rlabel metal2 s 225845 3212 225873 3452 4 la_data_in[89]
port 261 nsew
rlabel metal2 s 81313 3212 81341 3452 4 la_data_in[8]
port 262 nsew
rlabel metal2 s 227639 3212 227667 3452 4 la_data_in[90]
port 263 nsew
rlabel metal2 s 229387 3212 229415 3452 4 la_data_in[91]
port 264 nsew
rlabel metal2 s 231181 3212 231209 3452 4 la_data_in[92]
port 265 nsew
rlabel metal2 s 232975 3212 233003 3452 4 la_data_in[93]
port 266 nsew
rlabel metal2 s 234769 3212 234797 3452 4 la_data_in[94]
port 267 nsew
rlabel metal2 s 236563 3212 236591 3452 4 la_data_in[95]
port 268 nsew
rlabel metal2 s 238311 3212 238339 3452 4 la_data_in[96]
port 269 nsew
rlabel metal2 s 240105 3212 240133 3452 4 la_data_in[97]
port 270 nsew
rlabel metal2 s 241899 3212 241927 3452 4 la_data_in[98]
port 271 nsew
rlabel metal2 s 243693 3212 243721 3452 4 la_data_in[99]
port 272 nsew
rlabel metal2 s 83107 3212 83135 3452 4 la_data_in[9]
port 273 nsew
rlabel metal2 s 67651 3212 67679 3452 4 la_data_out[0]
port 274 nsew
rlabel metal2 s 246039 3212 246067 3452 4 la_data_out[100]
port 275 nsew
rlabel metal2 s 247833 3212 247861 3452 4 la_data_out[101]
port 276 nsew
rlabel metal2 s 249627 3212 249655 3452 4 la_data_out[102]
port 277 nsew
rlabel metal2 s 251421 3212 251449 3452 4 la_data_out[103]
port 278 nsew
rlabel metal2 s 253215 3212 253243 3452 4 la_data_out[104]
port 279 nsew
rlabel metal2 s 254963 3212 254991 3452 4 la_data_out[105]
port 280 nsew
rlabel metal2 s 256757 3212 256785 3452 4 la_data_out[106]
port 281 nsew
rlabel metal2 s 258551 3212 258579 3452 4 la_data_out[107]
port 282 nsew
rlabel metal2 s 260345 3212 260373 3452 4 la_data_out[108]
port 283 nsew
rlabel metal2 s 262139 3212 262167 3452 4 la_data_out[109]
port 284 nsew
rlabel metal2 s 85499 3212 85527 3452 4 la_data_out[10]
port 285 nsew
rlabel metal2 s 263887 3212 263915 3452 4 la_data_out[110]
port 286 nsew
rlabel metal2 s 265681 3212 265709 3452 4 la_data_out[111]
port 287 nsew
rlabel metal2 s 267475 3212 267503 3452 4 la_data_out[112]
port 288 nsew
rlabel metal2 s 269269 3212 269297 3452 4 la_data_out[113]
port 289 nsew
rlabel metal2 s 271017 3212 271045 3452 4 la_data_out[114]
port 290 nsew
rlabel metal2 s 272811 3212 272839 3452 4 la_data_out[115]
port 291 nsew
rlabel metal2 s 274605 3212 274633 3452 4 la_data_out[116]
port 292 nsew
rlabel metal2 s 276399 3212 276427 3452 4 la_data_out[117]
port 293 nsew
rlabel metal2 s 278193 3212 278221 3452 4 la_data_out[118]
port 294 nsew
rlabel metal2 s 279941 3212 279969 3452 4 la_data_out[119]
port 295 nsew
rlabel metal2 s 87293 3212 87321 3452 4 la_data_out[11]
port 296 nsew
rlabel metal2 s 281735 3212 281763 3452 4 la_data_out[120]
port 297 nsew
rlabel metal2 s 283529 3212 283557 3452 4 la_data_out[121]
port 298 nsew
rlabel metal2 s 285323 3212 285351 3452 4 la_data_out[122]
port 299 nsew
rlabel metal2 s 287117 3212 287145 3452 4 la_data_out[123]
port 300 nsew
rlabel metal2 s 288865 3212 288893 3452 4 la_data_out[124]
port 301 nsew
rlabel metal2 s 290659 3212 290687 3452 4 la_data_out[125]
port 302 nsew
rlabel metal2 s 292453 3212 292481 3452 4 la_data_out[126]
port 303 nsew
rlabel metal2 s 294247 3212 294275 3452 4 la_data_out[127]
port 304 nsew
rlabel metal2 s 89041 3212 89069 3452 4 la_data_out[12]
port 305 nsew
rlabel metal2 s 90835 3212 90863 3452 4 la_data_out[13]
port 306 nsew
rlabel metal2 s 92629 3212 92657 3452 4 la_data_out[14]
port 307 nsew
rlabel metal2 s 94423 3212 94451 3452 4 la_data_out[15]
port 308 nsew
rlabel metal2 s 96171 3212 96199 3452 4 la_data_out[16]
port 309 nsew
rlabel metal2 s 97965 3212 97993 3452 4 la_data_out[17]
port 310 nsew
rlabel metal2 s 99759 3212 99787 3452 4 la_data_out[18]
port 311 nsew
rlabel metal2 s 101553 3212 101581 3452 4 la_data_out[19]
port 312 nsew
rlabel metal2 s 69445 3212 69473 3452 4 la_data_out[1]
port 313 nsew
rlabel metal2 s 103347 3212 103375 3452 4 la_data_out[20]
port 314 nsew
rlabel metal2 s 105095 3212 105123 3452 4 la_data_out[21]
port 315 nsew
rlabel metal2 s 106889 3212 106917 3452 4 la_data_out[22]
port 316 nsew
rlabel metal2 s 108683 3212 108711 3452 4 la_data_out[23]
port 317 nsew
rlabel metal2 s 110477 3212 110505 3452 4 la_data_out[24]
port 318 nsew
rlabel metal2 s 112271 3212 112299 3452 4 la_data_out[25]
port 319 nsew
rlabel metal2 s 114019 3212 114047 3452 4 la_data_out[26]
port 320 nsew
rlabel metal2 s 115813 3212 115841 3452 4 la_data_out[27]
port 321 nsew
rlabel metal2 s 117607 3212 117635 3452 4 la_data_out[28]
port 322 nsew
rlabel metal2 s 119401 3212 119429 3452 4 la_data_out[29]
port 323 nsew
rlabel metal2 s 71193 3212 71221 3452 4 la_data_out[2]
port 324 nsew
rlabel metal2 s 121149 3212 121177 3452 4 la_data_out[30]
port 325 nsew
rlabel metal2 s 122943 3212 122971 3452 4 la_data_out[31]
port 326 nsew
rlabel metal2 s 124737 3212 124765 3452 4 la_data_out[32]
port 327 nsew
rlabel metal2 s 126531 3212 126559 3452 4 la_data_out[33]
port 328 nsew
rlabel metal2 s 128325 3212 128353 3452 4 la_data_out[34]
port 329 nsew
rlabel metal2 s 130073 3212 130101 3452 4 la_data_out[35]
port 330 nsew
rlabel metal2 s 131867 3212 131895 3452 4 la_data_out[36]
port 331 nsew
rlabel metal2 s 133661 3212 133689 3452 4 la_data_out[37]
port 332 nsew
rlabel metal2 s 135455 3212 135483 3452 4 la_data_out[38]
port 333 nsew
rlabel metal2 s 137249 3212 137277 3452 4 la_data_out[39]
port 334 nsew
rlabel metal2 s 72987 3212 73015 3452 4 la_data_out[3]
port 335 nsew
rlabel metal2 s 138997 3212 139025 3452 4 la_data_out[40]
port 336 nsew
rlabel metal2 s 140791 3212 140819 3452 4 la_data_out[41]
port 337 nsew
rlabel metal2 s 142585 3212 142613 3452 4 la_data_out[42]
port 338 nsew
rlabel metal2 s 144379 3212 144407 3452 4 la_data_out[43]
port 339 nsew
rlabel metal2 s 146127 3212 146155 3452 4 la_data_out[44]
port 340 nsew
rlabel metal2 s 147921 3212 147949 3452 4 la_data_out[45]
port 341 nsew
rlabel metal2 s 149715 3212 149743 3452 4 la_data_out[46]
port 342 nsew
rlabel metal2 s 151509 3212 151537 3452 4 la_data_out[47]
port 343 nsew
rlabel metal2 s 153303 3212 153331 3452 4 la_data_out[48]
port 344 nsew
rlabel metal2 s 155051 3212 155079 3452 4 la_data_out[49]
port 345 nsew
rlabel metal2 s 74781 3212 74809 3452 4 la_data_out[4]
port 346 nsew
rlabel metal2 s 156845 3212 156873 3452 4 la_data_out[50]
port 347 nsew
rlabel metal2 s 158639 3212 158667 3452 4 la_data_out[51]
port 348 nsew
rlabel metal2 s 160433 3212 160461 3452 4 la_data_out[52]
port 349 nsew
rlabel metal2 s 162227 3212 162255 3452 4 la_data_out[53]
port 350 nsew
rlabel metal2 s 163975 3212 164003 3452 4 la_data_out[54]
port 351 nsew
rlabel metal2 s 165769 3212 165797 3452 4 la_data_out[55]
port 352 nsew
rlabel metal2 s 167563 3212 167591 3452 4 la_data_out[56]
port 353 nsew
rlabel metal2 s 169357 3212 169385 3452 4 la_data_out[57]
port 354 nsew
rlabel metal2 s 171105 3212 171133 3452 4 la_data_out[58]
port 355 nsew
rlabel metal2 s 172899 3212 172927 3452 4 la_data_out[59]
port 356 nsew
rlabel metal2 s 76575 3212 76603 3452 4 la_data_out[5]
port 357 nsew
rlabel metal2 s 174693 3212 174721 3452 4 la_data_out[60]
port 358 nsew
rlabel metal2 s 176487 3212 176515 3452 4 la_data_out[61]
port 359 nsew
rlabel metal2 s 178281 3212 178309 3452 4 la_data_out[62]
port 360 nsew
rlabel metal2 s 180029 3212 180057 3452 4 la_data_out[63]
port 361 nsew
rlabel metal2 s 181823 3212 181851 3452 4 la_data_out[64]
port 362 nsew
rlabel metal2 s 183617 3212 183645 3452 4 la_data_out[65]
port 363 nsew
rlabel metal2 s 185411 3212 185439 3452 4 la_data_out[66]
port 364 nsew
rlabel metal2 s 187205 3212 187233 3452 4 la_data_out[67]
port 365 nsew
rlabel metal2 s 188953 3212 188981 3452 4 la_data_out[68]
port 366 nsew
rlabel metal2 s 190747 3212 190775 3452 4 la_data_out[69]
port 367 nsew
rlabel metal2 s 78369 3212 78397 3452 4 la_data_out[6]
port 368 nsew
rlabel metal2 s 192541 3212 192569 3452 4 la_data_out[70]
port 369 nsew
rlabel metal2 s 194335 3212 194363 3452 4 la_data_out[71]
port 370 nsew
rlabel metal2 s 196083 3212 196111 3452 4 la_data_out[72]
port 371 nsew
rlabel metal2 s 197877 3212 197905 3452 4 la_data_out[73]
port 372 nsew
rlabel metal2 s 199671 3212 199699 3452 4 la_data_out[74]
port 373 nsew
rlabel metal2 s 201465 3212 201493 3452 4 la_data_out[75]
port 374 nsew
rlabel metal2 s 203259 3212 203287 3452 4 la_data_out[76]
port 375 nsew
rlabel metal2 s 205007 3212 205035 3452 4 la_data_out[77]
port 376 nsew
rlabel metal2 s 206801 3212 206829 3452 4 la_data_out[78]
port 377 nsew
rlabel metal2 s 208595 3212 208623 3452 4 la_data_out[79]
port 378 nsew
rlabel metal2 s 80117 3212 80145 3452 4 la_data_out[7]
port 379 nsew
rlabel metal2 s 210389 3212 210417 3452 4 la_data_out[80]
port 380 nsew
rlabel metal2 s 212183 3212 212211 3452 4 la_data_out[81]
port 381 nsew
rlabel metal2 s 213931 3212 213959 3452 4 la_data_out[82]
port 382 nsew
rlabel metal2 s 215725 3212 215753 3452 4 la_data_out[83]
port 383 nsew
rlabel metal2 s 217519 3212 217547 3452 4 la_data_out[84]
port 384 nsew
rlabel metal2 s 219313 3212 219341 3452 4 la_data_out[85]
port 385 nsew
rlabel metal2 s 221061 3212 221089 3452 4 la_data_out[86]
port 386 nsew
rlabel metal2 s 222855 3212 222883 3452 4 la_data_out[87]
port 387 nsew
rlabel metal2 s 224649 3212 224677 3452 4 la_data_out[88]
port 388 nsew
rlabel metal2 s 226443 3212 226471 3452 4 la_data_out[89]
port 389 nsew
rlabel metal2 s 81911 3212 81939 3452 4 la_data_out[8]
port 390 nsew
rlabel metal2 s 228237 3212 228265 3452 4 la_data_out[90]
port 391 nsew
rlabel metal2 s 229985 3212 230013 3452 4 la_data_out[91]
port 392 nsew
rlabel metal2 s 231779 3212 231807 3452 4 la_data_out[92]
port 393 nsew
rlabel metal2 s 233573 3212 233601 3452 4 la_data_out[93]
port 394 nsew
rlabel metal2 s 235367 3212 235395 3452 4 la_data_out[94]
port 395 nsew
rlabel metal2 s 237161 3212 237189 3452 4 la_data_out[95]
port 396 nsew
rlabel metal2 s 238909 3212 238937 3452 4 la_data_out[96]
port 397 nsew
rlabel metal2 s 240703 3212 240731 3452 4 la_data_out[97]
port 398 nsew
rlabel metal2 s 242497 3212 242525 3452 4 la_data_out[98]
port 399 nsew
rlabel metal2 s 244291 3212 244319 3452 4 la_data_out[99]
port 400 nsew
rlabel metal2 s 83705 3212 83733 3452 4 la_data_out[9]
port 401 nsew
rlabel metal2 s 68249 3212 68277 3452 4 la_oen[0]
port 402 nsew
rlabel metal2 s 246637 3212 246665 3452 4 la_oen[100]
port 403 nsew
rlabel metal2 s 248431 3212 248459 3452 4 la_oen[101]
port 404 nsew
rlabel metal2 s 250225 3212 250253 3452 4 la_oen[102]
port 405 nsew
rlabel metal2 s 252019 3212 252047 3452 4 la_oen[103]
port 406 nsew
rlabel metal2 s 253813 3212 253841 3452 4 la_oen[104]
port 407 nsew
rlabel metal2 s 255561 3212 255589 3452 4 la_oen[105]
port 408 nsew
rlabel metal2 s 257355 3212 257383 3452 4 la_oen[106]
port 409 nsew
rlabel metal2 s 259149 3212 259177 3452 4 la_oen[107]
port 410 nsew
rlabel metal2 s 260943 3212 260971 3452 4 la_oen[108]
port 411 nsew
rlabel metal2 s 262691 3212 262719 3452 4 la_oen[109]
port 412 nsew
rlabel metal2 s 86097 3212 86125 3452 4 la_oen[10]
port 413 nsew
rlabel metal2 s 264485 3212 264513 3452 4 la_oen[110]
port 414 nsew
rlabel metal2 s 266279 3212 266307 3452 4 la_oen[111]
port 415 nsew
rlabel metal2 s 268073 3212 268101 3452 4 la_oen[112]
port 416 nsew
rlabel metal2 s 269867 3212 269895 3452 4 la_oen[113]
port 417 nsew
rlabel metal2 s 271615 3212 271643 3452 4 la_oen[114]
port 418 nsew
rlabel metal2 s 273409 3212 273437 3452 4 la_oen[115]
port 419 nsew
rlabel metal2 s 275203 3212 275231 3452 4 la_oen[116]
port 420 nsew
rlabel metal2 s 276997 3212 277025 3452 4 la_oen[117]
port 421 nsew
rlabel metal2 s 278791 3212 278819 3452 4 la_oen[118]
port 422 nsew
rlabel metal2 s 280539 3212 280567 3452 4 la_oen[119]
port 423 nsew
rlabel metal2 s 87845 3212 87873 3452 4 la_oen[11]
port 424 nsew
rlabel metal2 s 282333 3212 282361 3452 4 la_oen[120]
port 425 nsew
rlabel metal2 s 284127 3212 284155 3452 4 la_oen[121]
port 426 nsew
rlabel metal2 s 285921 3212 285949 3452 4 la_oen[122]
port 427 nsew
rlabel metal2 s 287669 3212 287697 3452 4 la_oen[123]
port 428 nsew
rlabel metal2 s 289463 3212 289491 3452 4 la_oen[124]
port 429 nsew
rlabel metal2 s 291257 3212 291285 3452 4 la_oen[125]
port 430 nsew
rlabel metal2 s 293051 3212 293079 3452 4 la_oen[126]
port 431 nsew
rlabel metal2 s 294845 3212 294873 3452 4 la_oen[127]
port 432 nsew
rlabel metal2 s 89639 3212 89667 3452 4 la_oen[12]
port 433 nsew
rlabel metal2 s 91433 3212 91461 3452 4 la_oen[13]
port 434 nsew
rlabel metal2 s 93227 3212 93255 3452 4 la_oen[14]
port 435 nsew
rlabel metal2 s 95021 3212 95049 3452 4 la_oen[15]
port 436 nsew
rlabel metal2 s 96769 3212 96797 3452 4 la_oen[16]
port 437 nsew
rlabel metal2 s 98563 3212 98591 3452 4 la_oen[17]
port 438 nsew
rlabel metal2 s 100357 3212 100385 3452 4 la_oen[18]
port 439 nsew
rlabel metal2 s 102151 3212 102179 3452 4 la_oen[19]
port 440 nsew
rlabel metal2 s 70043 3212 70071 3452 4 la_oen[1]
port 441 nsew
rlabel metal2 s 103945 3212 103973 3452 4 la_oen[20]
port 442 nsew
rlabel metal2 s 105693 3212 105721 3452 4 la_oen[21]
port 443 nsew
rlabel metal2 s 107487 3212 107515 3452 4 la_oen[22]
port 444 nsew
rlabel metal2 s 109281 3212 109309 3452 4 la_oen[23]
port 445 nsew
rlabel metal2 s 111075 3212 111103 3452 4 la_oen[24]
port 446 nsew
rlabel metal2 s 112823 3212 112851 3452 4 la_oen[25]
port 447 nsew
rlabel metal2 s 114617 3212 114645 3452 4 la_oen[26]
port 448 nsew
rlabel metal2 s 116411 3212 116439 3452 4 la_oen[27]
port 449 nsew
rlabel metal2 s 118205 3212 118233 3452 4 la_oen[28]
port 450 nsew
rlabel metal2 s 119999 3212 120027 3452 4 la_oen[29]
port 451 nsew
rlabel metal2 s 71791 3212 71819 3452 4 la_oen[2]
port 452 nsew
rlabel metal2 s 121747 3212 121775 3452 4 la_oen[30]
port 453 nsew
rlabel metal2 s 123541 3212 123569 3452 4 la_oen[31]
port 454 nsew
rlabel metal2 s 125335 3212 125363 3452 4 la_oen[32]
port 455 nsew
rlabel metal2 s 127129 3212 127157 3452 4 la_oen[33]
port 456 nsew
rlabel metal2 s 128923 3212 128951 3452 4 la_oen[34]
port 457 nsew
rlabel metal2 s 130671 3212 130699 3452 4 la_oen[35]
port 458 nsew
rlabel metal2 s 132465 3212 132493 3452 4 la_oen[36]
port 459 nsew
rlabel metal2 s 134259 3212 134287 3452 4 la_oen[37]
port 460 nsew
rlabel metal2 s 136053 3212 136081 3452 4 la_oen[38]
port 461 nsew
rlabel metal2 s 137801 3212 137829 3452 4 la_oen[39]
port 462 nsew
rlabel metal2 s 73585 3212 73613 3452 4 la_oen[3]
port 463 nsew
rlabel metal2 s 139595 3212 139623 3452 4 la_oen[40]
port 464 nsew
rlabel metal2 s 141389 3212 141417 3452 4 la_oen[41]
port 465 nsew
rlabel metal2 s 143183 3212 143211 3452 4 la_oen[42]
port 466 nsew
rlabel metal2 s 144977 3212 145005 3452 4 la_oen[43]
port 467 nsew
rlabel metal2 s 146725 3212 146753 3452 4 la_oen[44]
port 468 nsew
rlabel metal2 s 148519 3212 148547 3452 4 la_oen[45]
port 469 nsew
rlabel metal2 s 150313 3212 150341 3452 4 la_oen[46]
port 470 nsew
rlabel metal2 s 152107 3212 152135 3452 4 la_oen[47]
port 471 nsew
rlabel metal2 s 153901 3212 153929 3452 4 la_oen[48]
port 472 nsew
rlabel metal2 s 155649 3212 155677 3452 4 la_oen[49]
port 473 nsew
rlabel metal2 s 75379 3212 75407 3452 4 la_oen[4]
port 474 nsew
rlabel metal2 s 157443 3212 157471 3452 4 la_oen[50]
port 475 nsew
rlabel metal2 s 159237 3212 159265 3452 4 la_oen[51]
port 476 nsew
rlabel metal2 s 161031 3212 161059 3452 4 la_oen[52]
port 477 nsew
rlabel metal2 s 162779 3212 162807 3452 4 la_oen[53]
port 478 nsew
rlabel metal2 s 164573 3212 164601 3452 4 la_oen[54]
port 479 nsew
rlabel metal2 s 166367 3212 166395 3452 4 la_oen[55]
port 480 nsew
rlabel metal2 s 168161 3212 168189 3452 4 la_oen[56]
port 481 nsew
rlabel metal2 s 169955 3212 169983 3452 4 la_oen[57]
port 482 nsew
rlabel metal2 s 171703 3212 171731 3452 4 la_oen[58]
port 483 nsew
rlabel metal2 s 173497 3212 173525 3452 4 la_oen[59]
port 484 nsew
rlabel metal2 s 77173 3212 77201 3452 4 la_oen[5]
port 485 nsew
rlabel metal2 s 175291 3212 175319 3452 4 la_oen[60]
port 486 nsew
rlabel metal2 s 177085 3212 177113 3452 4 la_oen[61]
port 487 nsew
rlabel metal2 s 178879 3212 178907 3452 4 la_oen[62]
port 488 nsew
rlabel metal2 s 180627 3212 180655 3452 4 la_oen[63]
port 489 nsew
rlabel metal2 s 182421 3212 182449 3452 4 la_oen[64]
port 490 nsew
rlabel metal2 s 184215 3212 184243 3452 4 la_oen[65]
port 491 nsew
rlabel metal2 s 186009 3212 186037 3452 4 la_oen[66]
port 492 nsew
rlabel metal2 s 187757 3212 187785 3452 4 la_oen[67]
port 493 nsew
rlabel metal2 s 189551 3212 189579 3452 4 la_oen[68]
port 494 nsew
rlabel metal2 s 191345 3212 191373 3452 4 la_oen[69]
port 495 nsew
rlabel metal2 s 78967 3212 78995 3452 4 la_oen[6]
port 496 nsew
rlabel metal2 s 193139 3212 193167 3452 4 la_oen[70]
port 497 nsew
rlabel metal2 s 194933 3212 194961 3452 4 la_oen[71]
port 498 nsew
rlabel metal2 s 196681 3212 196709 3452 4 la_oen[72]
port 499 nsew
rlabel metal2 s 198475 3212 198503 3452 4 la_oen[73]
port 500 nsew
rlabel metal2 s 200269 3212 200297 3452 4 la_oen[74]
port 501 nsew
rlabel metal2 s 202063 3212 202091 3452 4 la_oen[75]
port 502 nsew
rlabel metal2 s 203857 3212 203885 3452 4 la_oen[76]
port 503 nsew
rlabel metal2 s 205605 3212 205633 3452 4 la_oen[77]
port 504 nsew
rlabel metal2 s 207399 3212 207427 3452 4 la_oen[78]
port 505 nsew
rlabel metal2 s 209193 3212 209221 3452 4 la_oen[79]
port 506 nsew
rlabel metal2 s 80715 3212 80743 3452 4 la_oen[7]
port 507 nsew
rlabel metal2 s 210987 3212 211015 3452 4 la_oen[80]
port 508 nsew
rlabel metal2 s 212735 3212 212763 3452 4 la_oen[81]
port 509 nsew
rlabel metal2 s 214529 3212 214557 3452 4 la_oen[82]
port 510 nsew
rlabel metal2 s 216323 3212 216351 3452 4 la_oen[83]
port 511 nsew
rlabel metal2 s 218117 3212 218145 3452 4 la_oen[84]
port 512 nsew
rlabel metal2 s 219911 3212 219939 3452 4 la_oen[85]
port 513 nsew
rlabel metal2 s 221659 3212 221687 3452 4 la_oen[86]
port 514 nsew
rlabel metal2 s 223453 3212 223481 3452 4 la_oen[87]
port 515 nsew
rlabel metal2 s 225247 3212 225275 3452 4 la_oen[88]
port 516 nsew
rlabel metal2 s 227041 3212 227069 3452 4 la_oen[89]
port 517 nsew
rlabel metal2 s 82509 3212 82537 3452 4 la_oen[8]
port 518 nsew
rlabel metal2 s 228835 3212 228863 3452 4 la_oen[90]
port 519 nsew
rlabel metal2 s 230583 3212 230611 3452 4 la_oen[91]
port 520 nsew
rlabel metal2 s 232377 3212 232405 3452 4 la_oen[92]
port 521 nsew
rlabel metal2 s 234171 3212 234199 3452 4 la_oen[93]
port 522 nsew
rlabel metal2 s 235965 3212 235993 3452 4 la_oen[94]
port 523 nsew
rlabel metal2 s 237713 3212 237741 3452 4 la_oen[95]
port 524 nsew
rlabel metal2 s 239507 3212 239535 3452 4 la_oen[96]
port 525 nsew
rlabel metal2 s 241301 3212 241329 3452 4 la_oen[97]
port 526 nsew
rlabel metal2 s 243095 3212 243123 3452 4 la_oen[98]
port 527 nsew
rlabel metal2 s 244889 3212 244917 3452 4 la_oen[99]
port 528 nsew
rlabel metal2 s 84303 3212 84331 3452 4 la_oen[9]
port 529 nsew
rlabel metal2 s 295443 3212 295471 3452 4 user_clock2
port 530 nsew
rlabel metal2 s 4033 3212 4061 3452 4 wb_clk_i
port 531 nsew
rlabel metal2 s 4585 3212 4613 3452 4 wb_rst_i
port 532 nsew
rlabel metal2 s 5183 3212 5211 3452 4 wbs_ack_o
port 533 nsew
rlabel metal2 s 7575 3212 7603 3452 4 wbs_adr_i[0]
port 534 nsew
rlabel metal2 s 27815 3212 27843 3452 4 wbs_adr_i[10]
port 535 nsew
rlabel metal2 s 29563 3212 29591 3452 4 wbs_adr_i[11]
port 536 nsew
rlabel metal2 s 31357 3212 31385 3452 4 wbs_adr_i[12]
port 537 nsew
rlabel metal2 s 33151 3212 33179 3452 4 wbs_adr_i[13]
port 538 nsew
rlabel metal2 s 34945 3212 34973 3452 4 wbs_adr_i[14]
port 539 nsew
rlabel metal2 s 36739 3212 36767 3452 4 wbs_adr_i[15]
port 540 nsew
rlabel metal2 s 38487 3212 38515 3452 4 wbs_adr_i[16]
port 541 nsew
rlabel metal2 s 40281 3212 40309 3452 4 wbs_adr_i[17]
port 542 nsew
rlabel metal2 s 42075 3212 42103 3452 4 wbs_adr_i[18]
port 543 nsew
rlabel metal2 s 43869 3212 43897 3452 4 wbs_adr_i[19]
port 544 nsew
rlabel metal2 s 9967 3212 9995 3452 4 wbs_adr_i[1]
port 545 nsew
rlabel metal2 s 45663 3212 45691 3452 4 wbs_adr_i[20]
port 546 nsew
rlabel metal2 s 47411 3212 47439 3452 4 wbs_adr_i[21]
port 547 nsew
rlabel metal2 s 49205 3212 49233 3452 4 wbs_adr_i[22]
port 548 nsew
rlabel metal2 s 50999 3212 51027 3452 4 wbs_adr_i[23]
port 549 nsew
rlabel metal2 s 52793 3212 52821 3452 4 wbs_adr_i[24]
port 550 nsew
rlabel metal2 s 54541 3212 54569 3452 4 wbs_adr_i[25]
port 551 nsew
rlabel metal2 s 56335 3212 56363 3452 4 wbs_adr_i[26]
port 552 nsew
rlabel metal2 s 58129 3212 58157 3452 4 wbs_adr_i[27]
port 553 nsew
rlabel metal2 s 59923 3212 59951 3452 4 wbs_adr_i[28]
port 554 nsew
rlabel metal2 s 61717 3212 61745 3452 4 wbs_adr_i[29]
port 555 nsew
rlabel metal2 s 12359 3212 12387 3452 4 wbs_adr_i[2]
port 556 nsew
rlabel metal2 s 63465 3212 63493 3452 4 wbs_adr_i[30]
port 557 nsew
rlabel metal2 s 65259 3212 65287 3452 4 wbs_adr_i[31]
port 558 nsew
rlabel metal2 s 14705 3212 14733 3452 4 wbs_adr_i[3]
port 559 nsew
rlabel metal2 s 17097 3212 17125 3452 4 wbs_adr_i[4]
port 560 nsew
rlabel metal2 s 18891 3212 18919 3452 4 wbs_adr_i[5]
port 561 nsew
rlabel metal2 s 20685 3212 20713 3452 4 wbs_adr_i[6]
port 562 nsew
rlabel metal2 s 22433 3212 22461 3452 4 wbs_adr_i[7]
port 563 nsew
rlabel metal2 s 24227 3212 24255 3452 4 wbs_adr_i[8]
port 564 nsew
rlabel metal2 s 26021 3212 26049 3452 4 wbs_adr_i[9]
port 565 nsew
rlabel metal2 s 5781 3212 5809 3452 4 wbs_cyc_i
port 566 nsew
rlabel metal2 s 8173 3212 8201 3452 4 wbs_dat_i[0]
port 567 nsew
rlabel metal2 s 28413 3212 28441 3452 4 wbs_dat_i[10]
port 568 nsew
rlabel metal2 s 30161 3212 30189 3452 4 wbs_dat_i[11]
port 569 nsew
rlabel metal2 s 31955 3212 31983 3452 4 wbs_dat_i[12]
port 570 nsew
rlabel metal2 s 33749 3212 33777 3452 4 wbs_dat_i[13]
port 571 nsew
rlabel metal2 s 35543 3212 35571 3452 4 wbs_dat_i[14]
port 572 nsew
rlabel metal2 s 37337 3212 37365 3452 4 wbs_dat_i[15]
port 573 nsew
rlabel metal2 s 39085 3212 39113 3452 4 wbs_dat_i[16]
port 574 nsew
rlabel metal2 s 40879 3212 40907 3452 4 wbs_dat_i[17]
port 575 nsew
rlabel metal2 s 42673 3212 42701 3452 4 wbs_dat_i[18]
port 576 nsew
rlabel metal2 s 44467 3212 44495 3452 4 wbs_dat_i[19]
port 577 nsew
rlabel metal2 s 10565 3212 10593 3452 4 wbs_dat_i[1]
port 578 nsew
rlabel metal2 s 46215 3212 46243 3452 4 wbs_dat_i[20]
port 579 nsew
rlabel metal2 s 48009 3212 48037 3452 4 wbs_dat_i[21]
port 580 nsew
rlabel metal2 s 49803 3212 49831 3452 4 wbs_dat_i[22]
port 581 nsew
rlabel metal2 s 51597 3212 51625 3452 4 wbs_dat_i[23]
port 582 nsew
rlabel metal2 s 53391 3212 53419 3452 4 wbs_dat_i[24]
port 583 nsew
rlabel metal2 s 55139 3212 55167 3452 4 wbs_dat_i[25]
port 584 nsew
rlabel metal2 s 56933 3212 56961 3452 4 wbs_dat_i[26]
port 585 nsew
rlabel metal2 s 58727 3212 58755 3452 4 wbs_dat_i[27]
port 586 nsew
rlabel metal2 s 60521 3212 60549 3452 4 wbs_dat_i[28]
port 587 nsew
rlabel metal2 s 62315 3212 62343 3452 4 wbs_dat_i[29]
port 588 nsew
rlabel metal2 s 12911 3212 12939 3452 4 wbs_dat_i[2]
port 589 nsew
rlabel metal2 s 64063 3212 64091 3452 4 wbs_dat_i[30]
port 590 nsew
rlabel metal2 s 65857 3212 65885 3452 4 wbs_dat_i[31]
port 591 nsew
rlabel metal2 s 15303 3212 15331 3452 4 wbs_dat_i[3]
port 592 nsew
rlabel metal2 s 17695 3212 17723 3452 4 wbs_dat_i[4]
port 593 nsew
rlabel metal2 s 19489 3212 19517 3452 4 wbs_dat_i[5]
port 594 nsew
rlabel metal2 s 21237 3212 21265 3452 4 wbs_dat_i[6]
port 595 nsew
rlabel metal2 s 23031 3212 23059 3452 4 wbs_dat_i[7]
port 596 nsew
rlabel metal2 s 24825 3212 24853 3452 4 wbs_dat_i[8]
port 597 nsew
rlabel metal2 s 26619 3212 26647 3452 4 wbs_dat_i[9]
port 598 nsew
rlabel metal2 s 8771 3212 8799 3452 4 wbs_dat_o[0]
port 599 nsew
rlabel metal2 s 29011 3212 29039 3452 4 wbs_dat_o[10]
port 600 nsew
rlabel metal2 s 30759 3212 30787 3452 4 wbs_dat_o[11]
port 601 nsew
rlabel metal2 s 32553 3212 32581 3452 4 wbs_dat_o[12]
port 602 nsew
rlabel metal2 s 34347 3212 34375 3452 4 wbs_dat_o[13]
port 603 nsew
rlabel metal2 s 36141 3212 36169 3452 4 wbs_dat_o[14]
port 604 nsew
rlabel metal2 s 37889 3212 37917 3452 4 wbs_dat_o[15]
port 605 nsew
rlabel metal2 s 39683 3212 39711 3452 4 wbs_dat_o[16]
port 606 nsew
rlabel metal2 s 41477 3212 41505 3452 4 wbs_dat_o[17]
port 607 nsew
rlabel metal2 s 43271 3212 43299 3452 4 wbs_dat_o[18]
port 608 nsew
rlabel metal2 s 45065 3212 45093 3452 4 wbs_dat_o[19]
port 609 nsew
rlabel metal2 s 11163 3212 11191 3452 4 wbs_dat_o[1]
port 610 nsew
rlabel metal2 s 46813 3212 46841 3452 4 wbs_dat_o[20]
port 611 nsew
rlabel metal2 s 48607 3212 48635 3452 4 wbs_dat_o[21]
port 612 nsew
rlabel metal2 s 50401 3212 50429 3452 4 wbs_dat_o[22]
port 613 nsew
rlabel metal2 s 52195 3212 52223 3452 4 wbs_dat_o[23]
port 614 nsew
rlabel metal2 s 53989 3212 54017 3452 4 wbs_dat_o[24]
port 615 nsew
rlabel metal2 s 55737 3212 55765 3452 4 wbs_dat_o[25]
port 616 nsew
rlabel metal2 s 57531 3212 57559 3452 4 wbs_dat_o[26]
port 617 nsew
rlabel metal2 s 59325 3212 59353 3452 4 wbs_dat_o[27]
port 618 nsew
rlabel metal2 s 61119 3212 61147 3452 4 wbs_dat_o[28]
port 619 nsew
rlabel metal2 s 62867 3212 62895 3452 4 wbs_dat_o[29]
port 620 nsew
rlabel metal2 s 13509 3212 13537 3452 4 wbs_dat_o[2]
port 621 nsew
rlabel metal2 s 64661 3212 64689 3452 4 wbs_dat_o[30]
port 622 nsew
rlabel metal2 s 66455 3212 66483 3452 4 wbs_dat_o[31]
port 623 nsew
rlabel metal2 s 15901 3212 15929 3452 4 wbs_dat_o[3]
port 624 nsew
rlabel metal2 s 18293 3212 18321 3452 4 wbs_dat_o[4]
port 625 nsew
rlabel metal2 s 20087 3212 20115 3452 4 wbs_dat_o[5]
port 626 nsew
rlabel metal2 s 21835 3212 21863 3452 4 wbs_dat_o[6]
port 627 nsew
rlabel metal2 s 23629 3212 23657 3452 4 wbs_dat_o[7]
port 628 nsew
rlabel metal2 s 25423 3212 25451 3452 4 wbs_dat_o[8]
port 629 nsew
rlabel metal2 s 27217 3212 27245 3452 4 wbs_dat_o[9]
port 630 nsew
rlabel metal2 s 9369 3212 9397 3452 4 wbs_sel_i[0]
port 631 nsew
rlabel metal2 s 11761 3212 11789 3452 4 wbs_sel_i[1]
port 632 nsew
rlabel metal2 s 14107 3212 14135 3452 4 wbs_sel_i[2]
port 633 nsew
rlabel metal2 s 16499 3212 16527 3452 4 wbs_sel_i[3]
port 634 nsew
rlabel metal2 s 6379 3212 6407 3452 4 wbs_stb_i
port 635 nsew
rlabel metal2 s 6977 3212 7005 3452 4 wbs_we_i
port 636 nsew
rlabel metal5 s 2800 2800 296658 3000 4 vccd1
port 637 nsew
rlabel metal5 s 2400 2400 297058 2600 4 vssd1
port 638 nsew
rlabel metal5 s 2000 2000 297458 2200 4 vccd2
port 639 nsew
rlabel metal5 s 1600 1600 297858 1800 4 vssd2
port 640 nsew
rlabel metal5 s 1200 1200 298258 1400 4 vdda1
port 641 nsew
rlabel metal5 s 800 800 298658 1000 4 vssa1
port 642 nsew
rlabel metal5 s 400 400 299058 600 4 vdda2
port 643 nsew
rlabel metal5 s 0 0 299458 200 4 vssa2
port 644 nsew
<< properties >>
string FIXED_BBOX 0 0 299458 358392
string GDS_FILE /project/openlane/user_project_wrapper_empty/runs/user_project_wrapper/results/magic/user_project_wrapper.gds
string GDS_END 5390882
string GDS_START 5141968
<< end >>
