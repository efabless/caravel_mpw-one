magic
tech sky130A
magscale 1 2
timestamp 1606497726
<< checkpaint >>
rect -1260 -1259 6384 6344
<< viali >>
rect 1633 2694 1667 2728
rect 2113 1880 2147 1914
<< metal1 >>
rect 66 4994 5058 5019
rect 66 4942 1610 4994
rect 1662 4942 1674 4994
rect 1726 4942 1738 4994
rect 1790 4942 1802 4994
rect 1854 4942 3277 4994
rect 3329 4942 3341 4994
rect 3393 4942 3405 4994
rect 3457 4942 3469 4994
rect 3521 4942 5058 4994
rect 66 4917 5058 4942
rect 66 3366 5058 3391
rect 66 3314 777 3366
rect 829 3314 841 3366
rect 893 3314 905 3366
rect 957 3314 969 3366
rect 1021 3314 2444 3366
rect 2496 3314 2508 3366
rect 2560 3314 2572 3366
rect 2624 3314 2636 3366
rect 2688 3314 4110 3366
rect 4162 3314 4174 3366
rect 4226 3314 4238 3366
rect 4290 3314 4302 3366
rect 4354 3314 5058 3366
rect 66 3289 5058 3314
rect 1621 2728 1679 2734
rect 1621 2694 1633 2728
rect 1667 2725 1679 2728
rect 4402 2725 4408 2737
rect 1667 2697 4408 2725
rect 1667 2694 1679 2697
rect 1621 2688 1679 2694
rect 4402 2685 4408 2697
rect 4460 2685 4466 2737
rect 658 1871 664 1923
rect 716 1911 722 1923
rect 2101 1914 2159 1920
rect 2101 1911 2113 1914
rect 716 1883 2113 1911
rect 716 1871 722 1883
rect 2101 1880 2113 1883
rect 2147 1880 2159 1914
rect 2101 1874 2159 1880
rect 66 1738 5058 1763
rect 66 1686 1610 1738
rect 1662 1686 1674 1738
rect 1726 1686 1738 1738
rect 1790 1686 1802 1738
rect 1854 1686 3277 1738
rect 3329 1686 3341 1738
rect 3393 1686 3405 1738
rect 3457 1686 3469 1738
rect 3521 1686 5058 1738
rect 66 1661 5058 1686
rect 66 110 5058 135
rect 66 58 777 110
rect 829 58 841 110
rect 893 58 905 110
rect 957 58 969 110
rect 1021 58 2444 110
rect 2496 58 2508 110
rect 2560 58 2572 110
rect 2624 58 2636 110
rect 2688 58 4110 110
rect 4162 58 4174 110
rect 4226 58 4238 110
rect 4290 58 4302 110
rect 4354 58 5058 110
rect 66 33 5058 58
<< via1 >>
rect 1610 4942 1662 4994
rect 1674 4942 1726 4994
rect 1738 4942 1790 4994
rect 1802 4942 1854 4994
rect 3277 4942 3329 4994
rect 3341 4942 3393 4994
rect 3405 4942 3457 4994
rect 3469 4942 3521 4994
rect 777 3314 829 3366
rect 841 3314 893 3366
rect 905 3314 957 3366
rect 969 3314 1021 3366
rect 2444 3314 2496 3366
rect 2508 3314 2560 3366
rect 2572 3314 2624 3366
rect 2636 3314 2688 3366
rect 4110 3314 4162 3366
rect 4174 3314 4226 3366
rect 4238 3314 4290 3366
rect 4302 3314 4354 3366
rect 4408 2685 4460 2737
rect 664 1871 716 1923
rect 1610 1686 1662 1738
rect 1674 1686 1726 1738
rect 1738 1686 1790 1738
rect 1802 1686 1854 1738
rect 3277 1686 3329 1738
rect 3341 1686 3393 1738
rect 3405 1686 3457 1738
rect 3469 1686 3521 1738
rect 777 58 829 110
rect 841 58 893 110
rect 905 58 957 110
rect 969 58 1021 110
rect 2444 58 2496 110
rect 2508 58 2560 110
rect 2572 58 2624 110
rect 2636 58 2688 110
rect 4110 58 4162 110
rect 4174 58 4226 110
rect 4238 58 4290 110
rect 4302 58 4354 110
<< metal2 >>
rect 1584 4996 1880 5019
rect 1640 4994 1664 4996
rect 1720 4994 1744 4996
rect 1800 4994 1824 4996
rect 1662 4942 1664 4994
rect 1726 4942 1738 4994
rect 1800 4942 1802 4994
rect 1640 4940 1664 4942
rect 1720 4940 1744 4942
rect 1800 4940 1824 4942
rect 1584 4917 1880 4940
rect 3251 4996 3547 5019
rect 3307 4994 3331 4996
rect 3387 4994 3411 4996
rect 3467 4994 3491 4996
rect 3329 4942 3331 4994
rect 3393 4942 3405 4994
rect 3467 4942 3469 4994
rect 3307 4940 3331 4942
rect 3387 4940 3411 4942
rect 3467 4940 3491 4942
rect 3251 4917 3547 4940
rect 4310 4284 4366 5084
rect 4324 3576 4352 4284
rect 4324 3548 4448 3576
rect 751 3368 1047 3391
rect 807 3366 831 3368
rect 887 3366 911 3368
rect 967 3366 991 3368
rect 829 3314 831 3366
rect 893 3314 905 3366
rect 967 3314 969 3366
rect 807 3312 831 3314
rect 887 3312 911 3314
rect 967 3312 991 3314
rect 751 3289 1047 3312
rect 2418 3368 2714 3391
rect 2474 3366 2498 3368
rect 2554 3366 2578 3368
rect 2634 3366 2658 3368
rect 2496 3314 2498 3366
rect 2560 3314 2572 3366
rect 2634 3314 2636 3366
rect 2474 3312 2498 3314
rect 2554 3312 2578 3314
rect 2634 3312 2658 3314
rect 2418 3289 2714 3312
rect 4084 3368 4380 3391
rect 4140 3366 4164 3368
rect 4220 3366 4244 3368
rect 4300 3366 4324 3368
rect 4162 3314 4164 3366
rect 4226 3314 4238 3366
rect 4300 3314 4302 3366
rect 4140 3312 4164 3314
rect 4220 3312 4244 3314
rect 4300 3312 4324 3314
rect 4084 3289 4380 3312
rect 4420 2743 4448 3548
rect 4408 2737 4460 2743
rect 4408 2679 4460 2685
rect 664 1923 716 1929
rect 664 1865 716 1871
rect 676 884 704 1865
rect 1584 1740 1880 1763
rect 1640 1738 1664 1740
rect 1720 1738 1744 1740
rect 1800 1738 1824 1740
rect 1662 1686 1664 1738
rect 1726 1686 1738 1738
rect 1800 1686 1802 1738
rect 1640 1684 1664 1686
rect 1720 1684 1744 1686
rect 1800 1684 1824 1686
rect 1584 1661 1880 1684
rect 3251 1740 3547 1763
rect 3307 1738 3331 1740
rect 3387 1738 3411 1740
rect 3467 1738 3491 1740
rect 3329 1686 3331 1738
rect 3393 1686 3405 1738
rect 3467 1686 3469 1738
rect 3307 1684 3331 1686
rect 3387 1684 3411 1686
rect 3467 1684 3491 1686
rect 3251 1661 3547 1684
rect 662 84 718 884
rect 751 112 1047 135
rect 807 110 831 112
rect 887 110 911 112
rect 967 110 991 112
rect 829 58 831 110
rect 893 58 905 110
rect 967 58 969 110
rect 807 56 831 58
rect 887 56 911 58
rect 967 56 991 58
rect 751 33 1047 56
rect 2418 112 2714 135
rect 2474 110 2498 112
rect 2554 110 2578 112
rect 2634 110 2658 112
rect 2496 58 2498 110
rect 2560 58 2572 110
rect 2634 58 2636 110
rect 2474 56 2498 58
rect 2554 56 2578 58
rect 2634 56 2658 58
rect 2418 33 2714 56
rect 4084 112 4380 135
rect 4140 110 4164 112
rect 4220 110 4244 112
rect 4300 110 4324 112
rect 4162 58 4164 110
rect 4226 58 4238 110
rect 4300 58 4302 110
rect 4140 56 4164 58
rect 4220 56 4244 58
rect 4300 56 4324 58
rect 4084 33 4380 56
<< via2 >>
rect 1584 4994 1640 4996
rect 1664 4994 1720 4996
rect 1744 4994 1800 4996
rect 1824 4994 1880 4996
rect 1584 4942 1610 4994
rect 1610 4942 1640 4994
rect 1664 4942 1674 4994
rect 1674 4942 1720 4994
rect 1744 4942 1790 4994
rect 1790 4942 1800 4994
rect 1824 4942 1854 4994
rect 1854 4942 1880 4994
rect 1584 4940 1640 4942
rect 1664 4940 1720 4942
rect 1744 4940 1800 4942
rect 1824 4940 1880 4942
rect 3251 4994 3307 4996
rect 3331 4994 3387 4996
rect 3411 4994 3467 4996
rect 3491 4994 3547 4996
rect 3251 4942 3277 4994
rect 3277 4942 3307 4994
rect 3331 4942 3341 4994
rect 3341 4942 3387 4994
rect 3411 4942 3457 4994
rect 3457 4942 3467 4994
rect 3491 4942 3521 4994
rect 3521 4942 3547 4994
rect 3251 4940 3307 4942
rect 3331 4940 3387 4942
rect 3411 4940 3467 4942
rect 3491 4940 3547 4942
rect 751 3366 807 3368
rect 831 3366 887 3368
rect 911 3366 967 3368
rect 991 3366 1047 3368
rect 751 3314 777 3366
rect 777 3314 807 3366
rect 831 3314 841 3366
rect 841 3314 887 3366
rect 911 3314 957 3366
rect 957 3314 967 3366
rect 991 3314 1021 3366
rect 1021 3314 1047 3366
rect 751 3312 807 3314
rect 831 3312 887 3314
rect 911 3312 967 3314
rect 991 3312 1047 3314
rect 2418 3366 2474 3368
rect 2498 3366 2554 3368
rect 2578 3366 2634 3368
rect 2658 3366 2714 3368
rect 2418 3314 2444 3366
rect 2444 3314 2474 3366
rect 2498 3314 2508 3366
rect 2508 3314 2554 3366
rect 2578 3314 2624 3366
rect 2624 3314 2634 3366
rect 2658 3314 2688 3366
rect 2688 3314 2714 3366
rect 2418 3312 2474 3314
rect 2498 3312 2554 3314
rect 2578 3312 2634 3314
rect 2658 3312 2714 3314
rect 4084 3366 4140 3368
rect 4164 3366 4220 3368
rect 4244 3366 4300 3368
rect 4324 3366 4380 3368
rect 4084 3314 4110 3366
rect 4110 3314 4140 3366
rect 4164 3314 4174 3366
rect 4174 3314 4220 3366
rect 4244 3314 4290 3366
rect 4290 3314 4300 3366
rect 4324 3314 4354 3366
rect 4354 3314 4380 3366
rect 4084 3312 4140 3314
rect 4164 3312 4220 3314
rect 4244 3312 4300 3314
rect 4324 3312 4380 3314
rect 1584 1738 1640 1740
rect 1664 1738 1720 1740
rect 1744 1738 1800 1740
rect 1824 1738 1880 1740
rect 1584 1686 1610 1738
rect 1610 1686 1640 1738
rect 1664 1686 1674 1738
rect 1674 1686 1720 1738
rect 1744 1686 1790 1738
rect 1790 1686 1800 1738
rect 1824 1686 1854 1738
rect 1854 1686 1880 1738
rect 1584 1684 1640 1686
rect 1664 1684 1720 1686
rect 1744 1684 1800 1686
rect 1824 1684 1880 1686
rect 3251 1738 3307 1740
rect 3331 1738 3387 1740
rect 3411 1738 3467 1740
rect 3491 1738 3547 1740
rect 3251 1686 3277 1738
rect 3277 1686 3307 1738
rect 3331 1686 3341 1738
rect 3341 1686 3387 1738
rect 3411 1686 3457 1738
rect 3457 1686 3467 1738
rect 3491 1686 3521 1738
rect 3521 1686 3547 1738
rect 3251 1684 3307 1686
rect 3331 1684 3387 1686
rect 3411 1684 3467 1686
rect 3491 1684 3547 1686
rect 751 110 807 112
rect 831 110 887 112
rect 911 110 967 112
rect 991 110 1047 112
rect 751 58 777 110
rect 777 58 807 110
rect 831 58 841 110
rect 841 58 887 110
rect 911 58 957 110
rect 957 58 967 110
rect 991 58 1021 110
rect 1021 58 1047 110
rect 751 56 807 58
rect 831 56 887 58
rect 911 56 967 58
rect 991 56 1047 58
rect 2418 110 2474 112
rect 2498 110 2554 112
rect 2578 110 2634 112
rect 2658 110 2714 112
rect 2418 58 2444 110
rect 2444 58 2474 110
rect 2498 58 2508 110
rect 2508 58 2554 110
rect 2578 58 2624 110
rect 2624 58 2634 110
rect 2658 58 2688 110
rect 2688 58 2714 110
rect 2418 56 2474 58
rect 2498 56 2554 58
rect 2578 56 2634 58
rect 2658 56 2714 58
rect 4084 110 4140 112
rect 4164 110 4220 112
rect 4244 110 4300 112
rect 4324 110 4380 112
rect 4084 58 4110 110
rect 4110 58 4140 110
rect 4164 58 4174 110
rect 4174 58 4220 110
rect 4244 58 4290 110
rect 4290 58 4300 110
rect 4324 58 4354 110
rect 4354 58 4380 110
rect 4084 56 4140 58
rect 4164 56 4220 58
rect 4244 56 4300 58
rect 4324 56 4380 58
<< metal3 >>
rect 1572 5000 1892 5001
rect 1572 4936 1580 5000
rect 1644 4936 1660 5000
rect 1724 4936 1740 5000
rect 1804 4936 1820 5000
rect 1884 4936 1892 5000
rect 1572 4935 1892 4936
rect 3239 5000 3559 5001
rect 3239 4936 3247 5000
rect 3311 4936 3327 5000
rect 3391 4936 3407 5000
rect 3471 4936 3487 5000
rect 3551 4936 3559 5000
rect 3239 4935 3559 4936
rect 739 3372 1059 3373
rect 739 3308 747 3372
rect 811 3308 827 3372
rect 891 3308 907 3372
rect 971 3308 987 3372
rect 1051 3308 1059 3372
rect 739 3307 1059 3308
rect 2406 3372 2726 3373
rect 2406 3308 2414 3372
rect 2478 3308 2494 3372
rect 2558 3308 2574 3372
rect 2638 3308 2654 3372
rect 2718 3308 2726 3372
rect 2406 3307 2726 3308
rect 4072 3372 4392 3373
rect 4072 3308 4080 3372
rect 4144 3308 4160 3372
rect 4224 3308 4240 3372
rect 4304 3308 4320 3372
rect 4384 3308 4392 3372
rect 4072 3307 4392 3308
rect 1572 1744 1892 1745
rect 1572 1680 1580 1744
rect 1644 1680 1660 1744
rect 1724 1680 1740 1744
rect 1804 1680 1820 1744
rect 1884 1680 1892 1744
rect 1572 1679 1892 1680
rect 3239 1744 3559 1745
rect 3239 1680 3247 1744
rect 3311 1680 3327 1744
rect 3391 1680 3407 1744
rect 3471 1680 3487 1744
rect 3551 1680 3559 1744
rect 3239 1679 3559 1680
rect 739 116 1059 117
rect 739 52 747 116
rect 811 52 827 116
rect 891 52 907 116
rect 971 52 987 116
rect 1051 52 1059 116
rect 739 51 1059 52
rect 2406 116 2726 117
rect 2406 52 2414 116
rect 2478 52 2494 116
rect 2558 52 2574 116
rect 2638 52 2654 116
rect 2718 52 2726 116
rect 2406 51 2726 52
rect 4072 116 4392 117
rect 4072 52 4080 116
rect 4144 52 4160 116
rect 4224 52 4240 116
rect 4304 52 4320 116
rect 4384 52 4392 116
rect 4072 51 4392 52
<< via3 >>
rect 1580 4996 1644 5000
rect 1580 4940 1584 4996
rect 1584 4940 1640 4996
rect 1640 4940 1644 4996
rect 1580 4936 1644 4940
rect 1660 4996 1724 5000
rect 1660 4940 1664 4996
rect 1664 4940 1720 4996
rect 1720 4940 1724 4996
rect 1660 4936 1724 4940
rect 1740 4996 1804 5000
rect 1740 4940 1744 4996
rect 1744 4940 1800 4996
rect 1800 4940 1804 4996
rect 1740 4936 1804 4940
rect 1820 4996 1884 5000
rect 1820 4940 1824 4996
rect 1824 4940 1880 4996
rect 1880 4940 1884 4996
rect 1820 4936 1884 4940
rect 3247 4996 3311 5000
rect 3247 4940 3251 4996
rect 3251 4940 3307 4996
rect 3307 4940 3311 4996
rect 3247 4936 3311 4940
rect 3327 4996 3391 5000
rect 3327 4940 3331 4996
rect 3331 4940 3387 4996
rect 3387 4940 3391 4996
rect 3327 4936 3391 4940
rect 3407 4996 3471 5000
rect 3407 4940 3411 4996
rect 3411 4940 3467 4996
rect 3467 4940 3471 4996
rect 3407 4936 3471 4940
rect 3487 4996 3551 5000
rect 3487 4940 3491 4996
rect 3491 4940 3547 4996
rect 3547 4940 3551 4996
rect 3487 4936 3551 4940
rect 747 3368 811 3372
rect 747 3312 751 3368
rect 751 3312 807 3368
rect 807 3312 811 3368
rect 747 3308 811 3312
rect 827 3368 891 3372
rect 827 3312 831 3368
rect 831 3312 887 3368
rect 887 3312 891 3368
rect 827 3308 891 3312
rect 907 3368 971 3372
rect 907 3312 911 3368
rect 911 3312 967 3368
rect 967 3312 971 3368
rect 907 3308 971 3312
rect 987 3368 1051 3372
rect 987 3312 991 3368
rect 991 3312 1047 3368
rect 1047 3312 1051 3368
rect 987 3308 1051 3312
rect 2414 3368 2478 3372
rect 2414 3312 2418 3368
rect 2418 3312 2474 3368
rect 2474 3312 2478 3368
rect 2414 3308 2478 3312
rect 2494 3368 2558 3372
rect 2494 3312 2498 3368
rect 2498 3312 2554 3368
rect 2554 3312 2558 3368
rect 2494 3308 2558 3312
rect 2574 3368 2638 3372
rect 2574 3312 2578 3368
rect 2578 3312 2634 3368
rect 2634 3312 2638 3368
rect 2574 3308 2638 3312
rect 2654 3368 2718 3372
rect 2654 3312 2658 3368
rect 2658 3312 2714 3368
rect 2714 3312 2718 3368
rect 2654 3308 2718 3312
rect 4080 3368 4144 3372
rect 4080 3312 4084 3368
rect 4084 3312 4140 3368
rect 4140 3312 4144 3368
rect 4080 3308 4144 3312
rect 4160 3368 4224 3372
rect 4160 3312 4164 3368
rect 4164 3312 4220 3368
rect 4220 3312 4224 3368
rect 4160 3308 4224 3312
rect 4240 3368 4304 3372
rect 4240 3312 4244 3368
rect 4244 3312 4300 3368
rect 4300 3312 4304 3368
rect 4240 3308 4304 3312
rect 4320 3368 4384 3372
rect 4320 3312 4324 3368
rect 4324 3312 4380 3368
rect 4380 3312 4384 3368
rect 4320 3308 4384 3312
rect 1580 1740 1644 1744
rect 1580 1684 1584 1740
rect 1584 1684 1640 1740
rect 1640 1684 1644 1740
rect 1580 1680 1644 1684
rect 1660 1740 1724 1744
rect 1660 1684 1664 1740
rect 1664 1684 1720 1740
rect 1720 1684 1724 1740
rect 1660 1680 1724 1684
rect 1740 1740 1804 1744
rect 1740 1684 1744 1740
rect 1744 1684 1800 1740
rect 1800 1684 1804 1740
rect 1740 1680 1804 1684
rect 1820 1740 1884 1744
rect 1820 1684 1824 1740
rect 1824 1684 1880 1740
rect 1880 1684 1884 1740
rect 1820 1680 1884 1684
rect 3247 1740 3311 1744
rect 3247 1684 3251 1740
rect 3251 1684 3307 1740
rect 3307 1684 3311 1740
rect 3247 1680 3311 1684
rect 3327 1740 3391 1744
rect 3327 1684 3331 1740
rect 3331 1684 3387 1740
rect 3387 1684 3391 1740
rect 3327 1680 3391 1684
rect 3407 1740 3471 1744
rect 3407 1684 3411 1740
rect 3411 1684 3467 1740
rect 3467 1684 3471 1740
rect 3407 1680 3471 1684
rect 3487 1740 3551 1744
rect 3487 1684 3491 1740
rect 3491 1684 3547 1740
rect 3547 1684 3551 1740
rect 3487 1680 3551 1684
rect 747 112 811 116
rect 747 56 751 112
rect 751 56 807 112
rect 807 56 811 112
rect 747 52 811 56
rect 827 112 891 116
rect 827 56 831 112
rect 831 56 887 112
rect 887 56 891 112
rect 827 52 891 56
rect 907 112 971 116
rect 907 56 911 112
rect 911 56 967 112
rect 967 56 971 112
rect 907 52 971 56
rect 987 112 1051 116
rect 987 56 991 112
rect 991 56 1047 112
rect 1047 56 1051 112
rect 987 52 1051 56
rect 2414 112 2478 116
rect 2414 56 2418 112
rect 2418 56 2474 112
rect 2474 56 2478 112
rect 2414 52 2478 56
rect 2494 112 2558 116
rect 2494 56 2498 112
rect 2498 56 2554 112
rect 2554 56 2558 112
rect 2494 52 2558 56
rect 2574 112 2638 116
rect 2574 56 2578 112
rect 2578 56 2634 112
rect 2634 56 2638 112
rect 2574 52 2638 56
rect 2654 112 2718 116
rect 2654 56 2658 112
rect 2658 56 2714 112
rect 2714 56 2718 112
rect 2654 52 2718 56
rect 4080 112 4144 116
rect 4080 56 4084 112
rect 4084 56 4140 112
rect 4140 56 4144 112
rect 4080 52 4144 56
rect 4160 112 4224 116
rect 4160 56 4164 112
rect 4164 56 4220 112
rect 4220 56 4224 112
rect 4160 52 4224 56
rect 4240 112 4304 116
rect 4240 56 4244 112
rect 4244 56 4300 112
rect 4300 56 4304 112
rect 4240 52 4304 56
rect 4320 112 4384 116
rect 4320 56 4324 112
rect 4324 56 4380 112
rect 4380 56 4384 112
rect 4320 52 4384 56
<< metal4 >>
rect 739 4317 1059 5019
rect 739 4081 781 4317
rect 1017 4081 1059 4317
rect 739 3372 1059 4081
rect 739 3308 747 3372
rect 811 3308 827 3372
rect 891 3308 907 3372
rect 971 3308 987 3372
rect 1051 3308 1059 3372
rect 739 2651 1059 3308
rect 739 2415 781 2651
rect 1017 2415 1059 2651
rect 739 984 1059 2415
rect 739 748 781 984
rect 1017 748 1059 984
rect 739 116 1059 748
rect 739 52 747 116
rect 811 52 827 116
rect 891 52 907 116
rect 971 52 987 116
rect 1051 52 1059 116
rect 739 33 1059 52
rect 1572 5000 1892 5019
rect 1572 4936 1580 5000
rect 1644 4936 1660 5000
rect 1724 4936 1740 5000
rect 1804 4936 1820 5000
rect 1884 4936 1892 5000
rect 1572 3484 1892 4936
rect 1572 3248 1614 3484
rect 1850 3248 1892 3484
rect 1572 1817 1892 3248
rect 1572 1744 1614 1817
rect 1850 1744 1892 1817
rect 1572 1680 1580 1744
rect 1884 1680 1892 1744
rect 1572 1581 1614 1680
rect 1850 1581 1892 1680
rect 1572 33 1892 1581
rect 2406 4317 2726 5019
rect 2406 4081 2448 4317
rect 2684 4081 2726 4317
rect 2406 3372 2726 4081
rect 2406 3308 2414 3372
rect 2478 3308 2494 3372
rect 2558 3308 2574 3372
rect 2638 3308 2654 3372
rect 2718 3308 2726 3372
rect 2406 2651 2726 3308
rect 2406 2415 2448 2651
rect 2684 2415 2726 2651
rect 2406 984 2726 2415
rect 2406 748 2448 984
rect 2684 748 2726 984
rect 2406 116 2726 748
rect 2406 52 2414 116
rect 2478 52 2494 116
rect 2558 52 2574 116
rect 2638 52 2654 116
rect 2718 52 2726 116
rect 2406 33 2726 52
rect 3239 5000 3559 5019
rect 3239 4936 3247 5000
rect 3311 4936 3327 5000
rect 3391 4936 3407 5000
rect 3471 4936 3487 5000
rect 3551 4936 3559 5000
rect 3239 3484 3559 4936
rect 3239 3248 3281 3484
rect 3517 3248 3559 3484
rect 3239 1817 3559 3248
rect 3239 1744 3281 1817
rect 3517 1744 3559 1817
rect 3239 1680 3247 1744
rect 3551 1680 3559 1744
rect 3239 1581 3281 1680
rect 3517 1581 3559 1680
rect 3239 33 3559 1581
rect 4072 4317 4392 5019
rect 4072 4081 4114 4317
rect 4350 4081 4392 4317
rect 4072 3372 4392 4081
rect 4072 3308 4080 3372
rect 4144 3308 4160 3372
rect 4224 3308 4240 3372
rect 4304 3308 4320 3372
rect 4384 3308 4392 3372
rect 4072 2651 4392 3308
rect 4072 2415 4114 2651
rect 4350 2415 4392 2651
rect 4072 984 4392 2415
rect 4072 748 4114 984
rect 4350 748 4392 984
rect 4072 116 4392 748
rect 4072 52 4080 116
rect 4144 52 4160 116
rect 4224 52 4240 116
rect 4304 52 4320 116
rect 4384 52 4392 116
rect 4072 33 4392 52
<< via4 >>
rect 781 4081 1017 4317
rect 781 2415 1017 2651
rect 781 748 1017 984
rect 1614 3248 1850 3484
rect 1614 1744 1850 1817
rect 1614 1680 1644 1744
rect 1644 1680 1660 1744
rect 1660 1680 1724 1744
rect 1724 1680 1740 1744
rect 1740 1680 1804 1744
rect 1804 1680 1820 1744
rect 1820 1680 1850 1744
rect 1614 1581 1850 1680
rect 2448 4081 2684 4317
rect 2448 2415 2684 2651
rect 2448 748 2684 984
rect 3281 3248 3517 3484
rect 3281 1744 3517 1817
rect 3281 1680 3311 1744
rect 3311 1680 3327 1744
rect 3327 1680 3391 1744
rect 3391 1680 3407 1744
rect 3407 1680 3471 1744
rect 3471 1680 3487 1744
rect 3487 1680 3517 1744
rect 3281 1581 3517 1680
rect 4114 4081 4350 4317
rect 4114 2415 4350 2651
rect 4114 748 4350 984
<< metal5 >>
rect 66 4317 5058 4359
rect 66 4081 781 4317
rect 1017 4081 2448 4317
rect 2684 4081 4114 4317
rect 4350 4081 5058 4317
rect 66 4039 5058 4081
rect 66 3484 5058 3526
rect 66 3248 1614 3484
rect 1850 3248 3281 3484
rect 3517 3248 5058 3484
rect 66 3206 5058 3248
rect 66 2651 5058 2693
rect 66 2415 781 2651
rect 1017 2415 2448 2651
rect 2684 2415 4114 2651
rect 4350 2415 5058 2651
rect 66 2373 5058 2415
rect 66 1817 5058 1859
rect 66 1581 1614 1817
rect 1850 1581 3281 1817
rect 3517 1581 5058 1817
rect 66 1539 5058 1581
rect 66 984 5058 1026
rect 66 748 781 984
rect 1017 748 2448 984
rect 2684 748 4114 984
rect 4350 748 5058 984
rect 66 706 5058 748
use sky130_fd_sc_hvl__decap_8  FILLER_1_39
timestamp 1606497726
transform 1 0 3810 0 1 1712
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_1_47
timestamp 1606497726
transform 1 0 4578 0 1 1712
box -66 -23 450 897
use sky130_fd_sc_hvl__fill_1  FILLER_1_51
timestamp 1606497726
transform 1 0 4962 0 1 1712
box -66 -23 162 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_40
timestamp 1606497726
transform 1 0 3906 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_2_48
timestamp 1606497726
transform 1 0 4674 0 -1 4154
box -66 -23 450 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_31
timestamp 1606497726
transform 1 0 3042 0 1 1712
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_24
timestamp 1606497726
transform 1 0 2370 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_32
timestamp 1606497726
transform 1 0 3138 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__lsbufhv2lv_1  lvlshiftdown
timestamp 1606497726
transform 1 0 1410 0 1 1712
box -66 -23 1698 1651
use sky130_fd_sc_hvl__decap_8  FILLER_1_0
timestamp 1606497726
transform 1 0 66 0 1 1712
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_1_8
timestamp 1606497726
transform 1 0 834 0 1 1712
box -66 -23 450 897
use sky130_fd_sc_hvl__fill_2  FILLER_1_12
timestamp 1606497726
transform 1 0 1218 0 1 1712
box -66 -23 258 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_0
timestamp 1606497726
transform 1 0 66 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_8
timestamp 1606497726
transform 1 0 834 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_16
timestamp 1606497726
transform 1 0 1602 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_40
timestamp 1606497726
transform 1 0 3906 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_0_48
timestamp 1606497726
transform 1 0 4674 0 -1 898
box -66 -23 450 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_24
timestamp 1606497726
transform 1 0 2370 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_32
timestamp 1606497726
transform 1 0 3138 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_0
timestamp 1606497726
transform 1 0 66 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_8
timestamp 1606497726
transform 1 0 834 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_16
timestamp 1606497726
transform 1 0 1602 0 -1 898
box -66 -23 834 897
<< labels >>
rlabel metal2 s 4310 4284 4366 5084 4 A
port 1 nsew
rlabel metal2 s 662 84 718 884 4 X
port 2 nsew
rlabel metal1 s 66 3289 5058 3391 4 VPWR
port 3 nsew
rlabel metal1 s 66 4917 5058 5019 4 VGND
port 4 nsew
<< properties >>
string FIXED_BBOX 0 1 5124 5084
<< end >>
