magic
tech sky130A
magscale 12 1
timestamp 1598777472
<< metal5 >>
rect 0 30 15 75
rect 30 30 45 75
rect 0 15 45 30
rect 5 10 40 15
rect 15 0 30 10
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
