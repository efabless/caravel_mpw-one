* NGSPICE file created from decred_controller.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

.subckt decred_controller CLK_LED DATA_AVAILABLE[0] DATA_AVAILABLE[1] DATA_AVAILABLE[2]
+ DATA_AVAILABLE[3] DATA_FROM_HASH[0] DATA_FROM_HASH[1] DATA_FROM_HASH[2] DATA_FROM_HASH[3]
+ DATA_FROM_HASH[4] DATA_FROM_HASH[5] DATA_FROM_HASH[6] DATA_FROM_HASH[7] DATA_TO_HASH[0]
+ DATA_TO_HASH[1] DATA_TO_HASH[2] DATA_TO_HASH[3] DATA_TO_HASH[4] DATA_TO_HASH[5]
+ DATA_TO_HASH[6] DATA_TO_HASH[7] EXT_RESET_N_fromHost EXT_RESET_N_toClient HASH_ADDR[0]
+ HASH_ADDR[1] HASH_ADDR[2] HASH_ADDR[3] HASH_ADDR[4] HASH_ADDR[5] HASH_EN HASH_LED
+ ID_fromClient ID_toHost IRQ_OUT_fromClient IRQ_OUT_toHost M1_CLK_IN M1_CLK_SELECT
+ MACRO_RD_SELECT[0] MACRO_RD_SELECT[1] MACRO_RD_SELECT[2] MACRO_RD_SELECT[3] MACRO_WR_SELECT[0]
+ MACRO_WR_SELECT[1] MACRO_WR_SELECT[2] MACRO_WR_SELECT[3] MISO_fromClient MISO_toHost
+ MOSI_fromHost MOSI_toClient PLL_INPUT S1_CLK_IN S1_CLK_SELECT SCLK_fromHost SCLK_toClient
+ SCSN_fromHost SCSN_toClient THREAD_COUNT[0] THREAD_COUNT[1] THREAD_COUNT[2] THREAD_COUNT[3]
+ m1_clk_local one zero VPWR VGND
X_2037_ _2043_/C _2047_/A _2043_/D _2037_/D VGND VGND VPWR VPWR _2038_/B sky130_fd_sc_hd__nand4_4
XFILLER_39_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2106_ _1222_/A SCSN_fromHost VGND VGND VPWR VPWR _2106_/X sky130_fd_sc_hd__or2_4
XFILLER_26_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1270_ _1270_/A VGND VGND VPWR VPWR _2010_/B sky130_fd_sc_hd__buf_2
XFILLER_3_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1606_ _1426_/A _1428_/D VGND VGND VPWR VPWR _1609_/B sky130_fd_sc_hd__nor2_4
XFILLER_8_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1399_ _2618_/Q _1397_/Y _1398_/Y VGND VGND VPWR VPWR _1400_/A sky130_fd_sc_hd__a21o_4
XFILLER_47_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1537_ _1424_/Y VGND VGND VPWR VPWR _1537_/X sky130_fd_sc_hd__buf_2
X_1468_ _1428_/Y VGND VGND VPWR VPWR _1548_/D sky130_fd_sc_hd__buf_2
X_2586_ _2606_/CLK _2586_/D VGND VGND VPWR VPWR _1459_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_27_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2440_ _2598_/CLK _2143_/Y VGND VGND VPWR VPWR _1964_/A sky130_fd_sc_hd__dfxtp_4
X_2371_ _2370_/CLK _2371_/D VGND VGND VPWR VPWR _2371_/Q sky130_fd_sc_hd__dfxtp_4
X_1253_ _2363_/Q VGND VGND VPWR VPWR _1374_/A sky130_fd_sc_hd__inv_2
X_1322_ _1239_/Y _1321_/X _1316_/D VGND VGND VPWR VPWR _1323_/A sky130_fd_sc_hd__nand3_4
Xclkbuf_1_0_0_m1_clk_local clkbuf_0_m1_clk_local/X VGND VGND VPWR VPWR clkbuf_2_1_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1184_ _1528_/A VGND VGND VPWR VPWR _1185_/A sky130_fd_sc_hd__buf_2
XFILLER_24_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2569_ _2570_/CLK _2569_/D VGND VGND VPWR VPWR _1735_/D sky130_fd_sc_hd__dfxtp_4
X_2638_ _2638_/CLK _2638_/D VGND VGND VPWR VPWR _1295_/A sky130_fd_sc_hd__dfxtp_4
XINSDIODE2_4 _1955_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1871_ _1870_/X DATA_FROM_HASH[7] VGND VGND VPWR VPWR _2566_/D sky130_fd_sc_hd__and2_4
X_1940_ _1938_/A _1746_/Y VGND VGND VPWR VPWR _1940_/Y sky130_fd_sc_hd__nor2_4
XFILLER_14_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2423_ _2408_/CLK _2271_/Y VGND VGND VPWR VPWR _1746_/A sky130_fd_sc_hd__dfxtp_4
X_1236_ _1236_/A _2623_/Q VGND VGND VPWR VPWR _1237_/A sky130_fd_sc_hd__nand2_4
X_2354_ _2097_/B _1179_/A _2353_/X VGND VGND VPWR VPWR _2354_/Y sky130_fd_sc_hd__o21ai_4
X_1305_ _1318_/B _1308_/C _1243_/X _1246_/D VGND VGND VPWR VPWR _1305_/X sky130_fd_sc_hd__and4_4
Xclkbuf_0_m1_clk_local m1_clk_local VGND VGND VPWR VPWR clkbuf_0_m1_clk_local/X sky130_fd_sc_hd__clkbuf_16
X_2285_ _2276_/X _2253_/Y _2278_/X _1923_/Y _2280_/X VGND VGND VPWR VPWR _2285_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_64_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_3_0_m1_clk_local clkbuf_3_3_0_m1_clk_local/A VGND VGND VPWR VPWR clkbuf_4_7_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
X_2070_ _2070_/A VGND VGND VPWR VPWR _2070_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1785_ _1783_/Y _1784_/Y _1781_/X VGND VGND VPWR VPWR _2588_/D sky130_fd_sc_hd__a21oi_4
X_1854_ _1854_/A _1640_/X VGND VGND VPWR VPWR _1854_/X sky130_fd_sc_hd__or2_4
X_1923_ _2151_/B VGND VGND VPWR VPWR _1923_/Y sky130_fd_sc_hd__inv_2
X_2406_ _2408_/CLK _2303_/Y VGND VGND VPWR VPWR HASH_LED sky130_fd_sc_hd__dfxtp_4
X_1219_ _2384_/Q VGND VGND VPWR VPWR _1219_/X sky130_fd_sc_hd__buf_2
X_2337_ _2337_/A _1575_/Y _1683_/Y VGND VGND VPWR VPWR _2338_/A sky130_fd_sc_hd__nand3_4
XFILLER_25_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2199_ _1623_/Y _2428_/Q VGND VGND VPWR VPWR _2199_/Y sky130_fd_sc_hd__nand2_4
X_2268_ _2268_/A VGND VGND VPWR VPWR _2268_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1570_ _1570_/A VGND VGND VPWR VPWR _1571_/A sky130_fd_sc_hd__buf_2
X_2053_ _1992_/A _2060_/A _1992_/D VGND VGND VPWR VPWR _2053_/Y sky130_fd_sc_hd__nor3_4
X_2122_ _1874_/A _2121_/X _1420_/A VGND VGND VPWR VPWR _2122_/Y sky130_fd_sc_hd__nand3_4
XFILLER_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1837_ _1836_/X VGND VGND VPWR VPWR _2570_/D sky130_fd_sc_hd__inv_2
X_1906_ _2154_/B VGND VGND VPWR VPWR _1906_/Y sky130_fd_sc_hd__inv_2
X_1768_ _1438_/B _1768_/B VGND VGND VPWR VPWR _1768_/X sky130_fd_sc_hd__xor2_4
XFILLER_57_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1699_ _1693_/Y _1698_/Y _1454_/X VGND VGND VPWR VPWR _2594_/D sky130_fd_sc_hd__a21oi_4
XFILLER_57_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1622_ _2426_/Q VGND VGND VPWR VPWR _1622_/Y sky130_fd_sc_hd__inv_2
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1553_ _1490_/A _1527_/Y _1530_/Y _1552_/Y VGND VGND VPWR VPWR _1557_/A sky130_fd_sc_hd__a211o_4
X_1484_ _1484_/A VGND VGND VPWR VPWR _1505_/B sky130_fd_sc_hd__buf_2
X_2036_ _2037_/D _2035_/X _1374_/X VGND VGND VPWR VPWR _2038_/A sky130_fd_sc_hd__o21a_4
XFILLER_54_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2105_ _1222_/A _2105_/B VGND VGND VPWR VPWR _2105_/X sky130_fd_sc_hd__or2_4
XFILLER_22_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1605_ _1605_/A VGND VGND VPWR VPWR _1651_/A sky130_fd_sc_hd__buf_2
X_2585_ _2581_/CLK _1796_/X VGND VGND VPWR VPWR _1477_/A sky130_fd_sc_hd__dfxtp_4
X_1536_ _1525_/Y _1532_/Y _1535_/X VGND VGND VPWR VPWR _2604_/D sky130_fd_sc_hd__a21oi_4
X_1398_ _2618_/Q _1397_/Y _1374_/X VGND VGND VPWR VPWR _1398_/Y sky130_fd_sc_hd__o21ai_4
X_1467_ _2602_/Q VGND VGND VPWR VPWR _1467_/Y sky130_fd_sc_hd__inv_2
X_2019_ _1395_/A _2019_/B _2019_/C VGND VGND VPWR VPWR _2019_/Y sky130_fd_sc_hd__nor3_4
XFILLER_35_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2370_ _2370_/CLK _2369_/Q VGND VGND VPWR VPWR _2371_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_49_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1321_ _1241_/Y VGND VGND VPWR VPWR _1321_/X sky130_fd_sc_hd__buf_2
X_1252_ _1271_/C _1251_/Y VGND VGND VPWR VPWR _1263_/A sky130_fd_sc_hd__nand2_4
XFILLER_64_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1183_ _2353_/A _1179_/X _1182_/X VGND VGND VPWR VPWR _1183_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_32_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_4_0_addressalyzerBlock.SPI_CLK clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_4_9_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_20_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE2_5 _1920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2499_ _2470_/CLK _1971_/X VGND VGND VPWR VPWR MACRO_WR_SELECT[0] sky130_fd_sc_hd__dfxtp_4
X_2568_ _2550_/CLK _2568_/D VGND VGND VPWR VPWR _1862_/B sky130_fd_sc_hd__dfxtp_4
X_2637_ _2477_/CLK _2637_/D VGND VGND VPWR VPWR _1299_/A sky130_fd_sc_hd__dfxtp_4
X_1519_ _1473_/B _1440_/B _1518_/Y VGND VGND VPWR VPWR _1519_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_59_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1870_ _1840_/B VGND VGND VPWR VPWR _1870_/X sky130_fd_sc_hd__buf_2
X_2353_ _2353_/A _1180_/Y VGND VGND VPWR VPWR _2353_/X sky130_fd_sc_hd__or2_4
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2422_ _2408_/CLK _2422_/D VGND VGND VPWR VPWR _1941_/A sky130_fd_sc_hd__dfxtp_4
X_1235_ _1235_/A VGND VGND VPWR VPWR _1365_/D sky130_fd_sc_hd__inv_2
XFILLER_37_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1304_ _2635_/Q VGND VGND VPWR VPWR _1308_/C sky130_fd_sc_hd__buf_2
X_2284_ _2276_/X _2133_/Y _2278_/X _1744_/B _2280_/X VGND VGND VPWR VPWR _2415_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_20_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1999_ _1999_/A _1999_/B _2011_/A _2492_/Q VGND VGND VPWR VPWR _2010_/C sky130_fd_sc_hd__nand4_4
XFILLER_20_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1922_ _1932_/A _2537_/Q VGND VGND VPWR VPWR _2531_/D sky130_fd_sc_hd__and2_4
X_1784_ _1678_/Y _2349_/A VGND VGND VPWR VPWR _1784_/Y sky130_fd_sc_hd__nand2_4
X_1853_ _1850_/X _1852_/X _1471_/X VGND VGND VPWR VPWR _1853_/Y sky130_fd_sc_hd__a21oi_4
X_2336_ _1575_/Y _2328_/X _2335_/Y VGND VGND VPWR VPWR _2388_/D sky130_fd_sc_hd__o21ai_4
XFILLER_29_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2405_ _2557_/CLK _2305_/Y VGND VGND VPWR VPWR _1232_/A sky130_fd_sc_hd__dfxtp_4
X_1218_ _1218_/A _1218_/B VGND VGND VPWR VPWR _1218_/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2267_ _2266_/Y _2262_/X _2258_/X _1937_/Y _2264_/X VGND VGND VPWR VPWR _2425_/D
+ sky130_fd_sc_hd__o32ai_4
X_2198_ _2196_/Y _1708_/X _2198_/C VGND VGND VPWR VPWR _2198_/Y sky130_fd_sc_hd__nand3_4
XFILLER_52_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2052_ _2014_/X _2040_/X _2051_/Y VGND VGND VPWR VPWR _2052_/Y sky130_fd_sc_hd__a21oi_4
X_2121_ _1696_/A VGND VGND VPWR VPWR _2121_/X sky130_fd_sc_hd__buf_2
XFILLER_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1905_ _1901_/X _1905_/B VGND VGND VPWR VPWR _1905_/Y sky130_fd_sc_hd__nor2_4
X_1836_ _1735_/C _1834_/Y _1835_/Y VGND VGND VPWR VPWR _1836_/X sky130_fd_sc_hd__a21o_4
X_1698_ _1698_/A _1697_/Y _1689_/Y _2340_/B VGND VGND VPWR VPWR _1698_/Y sky130_fd_sc_hd__nand4_4
XFILLER_30_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1767_ _1483_/B _1767_/B VGND VGND VPWR VPWR _1767_/X sky130_fd_sc_hd__xor2_4
X_2319_ _1771_/Y _2310_/X _1503_/A _2312_/X VGND VGND VPWR VPWR _2319_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1552_ _1537_/X _1548_/D _1544_/Y VGND VGND VPWR VPWR _1552_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_8_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1621_ _2410_/Q _2181_/A _1617_/Y _1620_/Y VGND VGND VPWR VPWR _1621_/X sky130_fd_sc_hd__a211o_4
X_2104_ _2104_/A _2091_/Y _2103_/Y _2468_/Q VGND VGND VPWR VPWR _2104_/X sky130_fd_sc_hd__and4_4
X_1483_ _1482_/Y _1483_/B _2604_/Q _2603_/Q VGND VGND VPWR VPWR _1484_/A sky130_fd_sc_hd__and4_4
X_2035_ _2029_/Y _2030_/X _2017_/B _2043_/D VGND VGND VPWR VPWR _2035_/X sky130_fd_sc_hd__and4_4
XFILLER_22_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1819_ _2575_/Q _1809_/X _1818_/X VGND VGND VPWR VPWR _2576_/D sky130_fd_sc_hd__o21a_4
XFILLER_53_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1604_ _1559_/B _2600_/Q VGND VGND VPWR VPWR _1605_/A sky130_fd_sc_hd__and2_4
X_1535_ _1556_/A _1534_/X _1500_/X VGND VGND VPWR VPWR _1535_/X sky130_fd_sc_hd__a21o_4
X_2584_ _2606_/CLK _1798_/X VGND VGND VPWR VPWR _1490_/A sky130_fd_sc_hd__dfxtp_4
X_1397_ _1397_/A _1397_/B _1397_/C VGND VGND VPWR VPWR _1397_/Y sky130_fd_sc_hd__nor3_4
X_1466_ _1466_/A VGND VGND VPWR VPWR _1466_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2018_ _2488_/Q _2017_/X _1984_/A _1999_/A _2011_/A VGND VGND VPWR VPWR _2019_/C
+ sky130_fd_sc_hd__a41oi_4
XFILLER_42_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1320_ _1319_/Y VGND VGND VPWR VPWR _2634_/D sky130_fd_sc_hd__inv_2
XFILLER_64_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1182_ _1182_/A _1194_/B VGND VGND VPWR VPWR _1182_/X sky130_fd_sc_hd__or2_4
X_1251_ _1251_/A VGND VGND VPWR VPWR _1251_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2636_ _2477_/CLK _2636_/D VGND VGND VPWR VPWR _2636_/Q sky130_fd_sc_hd__dfxtp_4
X_2498_ _2498_/CLK _2498_/D VGND VGND VPWR VPWR _1973_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_59_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2567_ _2498_/CLK _1869_/Y VGND VGND VPWR VPWR _2567_/Q sky130_fd_sc_hd__dfxtp_4
X_1518_ _1473_/B _1482_/Y _1473_/C _1466_/A _2340_/C VGND VGND VPWR VPWR _1518_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1449_ _1441_/Y _1449_/B VGND VGND VPWR VPWR _1449_/Y sky130_fd_sc_hd__nand2_4
XFILLER_15_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2352_ _2543_/Q _2544_/Q _2352_/C VGND VGND VPWR VPWR IRQ_OUT_toHost sky130_fd_sc_hd__or3_4
X_1303_ _1258_/Y VGND VGND VPWR VPWR _1318_/B sky130_fd_sc_hd__buf_2
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2283_ _2276_/X _2130_/Y _2278_/X _1845_/B _2280_/X VGND VGND VPWR VPWR _2416_/D
+ sky130_fd_sc_hd__o32ai_4
X_2421_ _2408_/CLK _2421_/D VGND VGND VPWR VPWR _1944_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_52_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1234_ _1385_/A _2621_/Q VGND VGND VPWR VPWR _1235_/A sky130_fd_sc_hd__nand2_4
XFILLER_37_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1998_ _1998_/A _2008_/A VGND VGND VPWR VPWR _1999_/B sky130_fd_sc_hd__nor2_4
X_2619_ _2370_/CLK _1395_/Y VGND VGND VPWR VPWR _2619_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_18_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1921_ _1254_/X VGND VGND VPWR VPWR _1932_/A sky130_fd_sc_hd__buf_2
X_1852_ _2444_/Q _1751_/A _1633_/X _1851_/Y VGND VGND VPWR VPWR _1852_/X sky130_fd_sc_hd__a211o_4
X_1783_ _1678_/A _1783_/B _1779_/C _1783_/D VGND VGND VPWR VPWR _1783_/Y sky130_fd_sc_hd__nand4_4
X_2335_ _2335_/A _2335_/B _1218_/B _1577_/X VGND VGND VPWR VPWR _2335_/Y sky130_fd_sc_hd__nand4_4
X_2266_ _2266_/A VGND VGND VPWR VPWR _2266_/Y sky130_fd_sc_hd__inv_2
X_2404_ _2408_/CLK _2307_/Y VGND VGND VPWR VPWR _2404_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_25_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1217_ _1185_/A VGND VGND VPWR VPWR _1218_/B sky130_fd_sc_hd__buf_2
X_2197_ _2404_/Q _2175_/B VGND VGND VPWR VPWR _2198_/C sky130_fd_sc_hd__nand2_4
XFILLER_4_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2120_ _2123_/A VGND VGND VPWR VPWR _2120_/X sky130_fd_sc_hd__buf_2
X_2051_ _2014_/X _2040_/X _1346_/X VGND VGND VPWR VPWR _2051_/Y sky130_fd_sc_hd__o21ai_4
X_1835_ _1735_/C _1834_/Y _1831_/B VGND VGND VPWR VPWR _1835_/Y sky130_fd_sc_hd__o21ai_4
X_1904_ _2431_/Q VGND VGND VPWR VPWR _1905_/B sky130_fd_sc_hd__inv_2
XFILLER_15_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1697_ _1697_/A VGND VGND VPWR VPWR _1697_/Y sky130_fd_sc_hd__inv_2
X_1766_ _1438_/C _1766_/B VGND VGND VPWR VPWR _1766_/Y sky130_fd_sc_hd__nor2_4
XFILLER_57_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2249_ _2248_/X VGND VGND VPWR VPWR _2249_/X sky130_fd_sc_hd__buf_2
X_2318_ _2158_/B _2311_/X _2253_/C _2313_/X VGND VGND VPWR VPWR _2318_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_40_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1551_ _1546_/X _1550_/Y _1454_/X VGND VGND VPWR VPWR _1551_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_8_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1620_ _2175_/B _1620_/B VGND VGND VPWR VPWR _1620_/Y sky130_fd_sc_hd__nor2_4
X_1482_ _1467_/Y _1424_/Y _1428_/Y VGND VGND VPWR VPWR _1482_/Y sky130_fd_sc_hd__nor3_4
X_2103_ _2103_/A VGND VGND VPWR VPWR _2103_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2034_ _2017_/C _2032_/X _2033_/Y VGND VGND VPWR VPWR _2034_/X sky130_fd_sc_hd__o21a_4
X_1818_ _2576_/Q _1810_/X _1813_/X VGND VGND VPWR VPWR _1818_/X sky130_fd_sc_hd__o21a_4
X_1749_ _1745_/X _1748_/Y _1628_/X VGND VGND VPWR VPWR _1749_/X sky130_fd_sc_hd__a21o_4
XFILLER_45_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_4_0_addressalyzerBlock.SPI_CLK clkbuf_4_5_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2557_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_9_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2652_ _2570_/CLK _2652_/D VGND VGND VPWR VPWR _2097_/B sky130_fd_sc_hd__dfxtp_4
X_1534_ _1534_/A VGND VGND VPWR VPWR _1534_/X sky130_fd_sc_hd__buf_2
X_1603_ _1602_/Y VGND VGND VPWR VPWR _1603_/Y sky130_fd_sc_hd__inv_2
X_2583_ _2606_/CLK _2583_/D VGND VGND VPWR VPWR _1497_/A sky130_fd_sc_hd__dfxtp_4
X_1465_ _1458_/Y _1463_/Y _1464_/Y VGND VGND VPWR VPWR _2611_/D sky130_fd_sc_hd__a21oi_4
X_2017_ _2047_/A _2017_/B _2017_/C _2017_/D VGND VGND VPWR VPWR _2017_/X sky130_fd_sc_hd__and4_4
X_1396_ _1231_/B VGND VGND VPWR VPWR _1397_/A sky130_fd_sc_hd__inv_2
XFILLER_50_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1181_ _1180_/Y VGND VGND VPWR VPWR _1194_/B sky130_fd_sc_hd__buf_2
X_1250_ _1262_/C _1277_/B _1277_/D _1249_/Y VGND VGND VPWR VPWR _1271_/C sky130_fd_sc_hd__nand4_4
XFILLER_32_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2635_ _2477_/CLK _2635_/D VGND VGND VPWR VPWR _2635_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_4_8_0_m1_clk_local clkbuf_4_9_0_m1_clk_local/A VGND VGND VPWR VPWR _2618_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_2497_ _2496_/CLK _1978_/X VGND VGND VPWR VPWR _2497_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_55_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2566_ _2557_/CLK _2566_/D VGND VGND VPWR VPWR _2566_/Q sky130_fd_sc_hd__dfxtp_4
X_1517_ _1513_/X _1515_/Y _1516_/X VGND VGND VPWR VPWR _2606_/D sky130_fd_sc_hd__a21oi_4
X_1448_ _1448_/A VGND VGND VPWR VPWR _1449_/B sky130_fd_sc_hd__buf_2
X_1379_ _1379_/A VGND VGND VPWR VPWR _1379_/X sky130_fd_sc_hd__buf_2
XFILLER_55_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2420_ _2408_/CLK _2420_/D VGND VGND VPWR VPWR _2420_/Q sky130_fd_sc_hd__dfxtp_4
X_2351_ _2351_/A _2546_/Q _2351_/C VGND VGND VPWR VPWR _2352_/C sky130_fd_sc_hd__or3_4
X_1233_ _1233_/A _1397_/B _1233_/C _1397_/C VGND VGND VPWR VPWR _1379_/A sky130_fd_sc_hd__nor4_4
X_1302_ _1301_/Y VGND VGND VPWR VPWR _2637_/D sky130_fd_sc_hd__inv_2
X_2282_ _2276_/X _2127_/Y _2278_/X _1705_/Y _2280_/X VGND VGND VPWR VPWR _2417_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_64_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1997_ _2017_/C _1994_/Y _2488_/Q _2017_/D VGND VGND VPWR VPWR _2008_/A sky130_fd_sc_hd__nand4_4
XFILLER_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2549_ _2550_/CLK _2549_/D VGND VGND VPWR VPWR _1897_/B sky130_fd_sc_hd__dfxtp_4
X_2618_ _2618_/CLK _1400_/Y VGND VGND VPWR VPWR _2618_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_55_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0_addressalyzerBlock.SPI_CLK clkbuf_0_addressalyzerBlock.SPI_CLK/X VGND
+ VGND VPWR VPWR clkbuf_2_1_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_46_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1851_ _1635_/X _1766_/B VGND VGND VPWR VPWR _1851_/Y sky130_fd_sc_hd__nor2_4
X_1920_ _1918_/A _2538_/Q VGND VGND VPWR VPWR _1920_/X sky130_fd_sc_hd__and2_4
X_1782_ _1779_/Y _1780_/Y _1781_/X VGND VGND VPWR VPWR _1782_/Y sky130_fd_sc_hd__a21oi_4
X_2403_ _2408_/CLK _2403_/D VGND VGND VPWR VPWR _2089_/A sky130_fd_sc_hd__dfxtp_4
X_1216_ _1194_/B _1216_/B _2645_/Q VGND VGND VPWR VPWR _1216_/Y sky130_fd_sc_hd__nand3_4
X_2334_ _1529_/Y _2333_/Y _1781_/X VGND VGND VPWR VPWR _2389_/D sky130_fd_sc_hd__a21oi_4
X_2265_ _1420_/Y _2262_/X _2258_/X _1622_/Y _2264_/X VGND VGND VPWR VPWR _2426_/D
+ sky130_fd_sc_hd__o32ai_4
X_2196_ _2151_/A _1927_/A VGND VGND VPWR VPWR _2196_/Y sky130_fd_sc_hd__nand2_4
XFILLER_52_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2050_ _2049_/Y VGND VGND VPWR VPWR _2050_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1834_ _1834_/A VGND VGND VPWR VPWR _1834_/Y sky130_fd_sc_hd__inv_2
X_1903_ _1901_/X _1902_/Y VGND VGND VPWR VPWR _1903_/Y sky130_fd_sc_hd__nor2_4
X_1765_ _1765_/A VGND VGND VPWR VPWR _1766_/B sky130_fd_sc_hd__inv_2
X_1696_ _1696_/A VGND VGND VPWR VPWR _1698_/A sky130_fd_sc_hd__buf_2
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2317_ _1751_/B _2311_/X _1490_/A _2313_/X VGND VGND VPWR VPWR _2399_/D sky130_fd_sc_hd__a2bb2o_4
X_2179_ _2177_/Y _2179_/B _2179_/C VGND VGND VPWR VPWR _2179_/Y sky130_fd_sc_hd__nand3_4
X_2248_ _1583_/X _1594_/X _1600_/B _1696_/A _1736_/A VGND VGND VPWR VPWR _2248_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_25_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1550_ _1547_/X _1548_/Y _1549_/Y VGND VGND VPWR VPWR _1550_/Y sky130_fd_sc_hd__o21ai_4
X_1481_ _1436_/B VGND VGND VPWR VPWR _1487_/A sky130_fd_sc_hd__buf_2
X_2033_ _2043_/C _2047_/A _2017_/C _2017_/D _1275_/X VGND VGND VPWR VPWR _2033_/Y
+ sky130_fd_sc_hd__a41oi_4
X_2102_ _2102_/A _2103_/A _2468_/Q _2091_/Y VGND VGND VPWR VPWR _2461_/D sky130_fd_sc_hd__nor4_4
XFILLER_39_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1817_ _2576_/Q _1809_/X _1816_/X VGND VGND VPWR VPWR _1817_/X sky130_fd_sc_hd__o21a_4
X_1748_ _1746_/Y _1624_/X _1747_/Y VGND VGND VPWR VPWR _1748_/Y sky130_fd_sc_hd__o21ai_4
X_1679_ _1566_/X _1683_/A VGND VGND VPWR VPWR _1679_/Y sky130_fd_sc_hd__nor2_4
XFILLER_53_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2651_ _2457_/CLK _1193_/Y VGND VGND VPWR VPWR _2353_/A sky130_fd_sc_hd__dfxtp_4
X_1602_ _1602_/A _1600_/Y _1602_/C VGND VGND VPWR VPWR _1602_/Y sky130_fd_sc_hd__nand3_4
X_2582_ _2581_/CLK _2582_/D VGND VGND VPWR VPWR _1503_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_8_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1395_ _1395_/A _1379_/X _1394_/Y VGND VGND VPWR VPWR _1395_/Y sky130_fd_sc_hd__nor3_4
X_1464_ _1438_/B _1449_/B _1213_/X VGND VGND VPWR VPWR _1464_/Y sky130_fd_sc_hd__o21ai_4
X_1533_ _2604_/Q VGND VGND VPWR VPWR _1534_/A sky130_fd_sc_hd__inv_2
X_2016_ _1987_/A VGND VGND VPWR VPWR _2017_/B sky130_fd_sc_hd__buf_2
XFILLER_50_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1180_ _1178_/A VGND VGND VPWR VPWR _1180_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2634_ _2626_/CLK _2634_/D VGND VGND VPWR VPWR _1318_/A sky130_fd_sc_hd__dfxtp_4
X_2565_ _2562_/CLK _2565_/D VGND VGND VPWR VPWR _2565_/Q sky130_fd_sc_hd__dfxtp_4
X_1516_ _1450_/X _1512_/Y _1500_/X VGND VGND VPWR VPWR _1516_/X sky130_fd_sc_hd__a21o_4
X_2496_ _2496_/CLK _2496_/D VGND VGND VPWR VPWR _2496_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_59_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1378_ _1378_/A VGND VGND VPWR VPWR _2624_/D sky130_fd_sc_hd__inv_2
X_1447_ _1446_/Y VGND VGND VPWR VPWR _1448_/A sky130_fd_sc_hd__inv_2
XFILLER_55_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2350_ _2349_/A _2348_/Y _2349_/Y VGND VGND VPWR VPWR MISO_toHost sky130_fd_sc_hd__a21oi_4
XFILLER_49_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1232_ _1232_/A _2615_/Q _1409_/B _1232_/D VGND VGND VPWR VPWR _1397_/C sky130_fd_sc_hd__nand4_4
X_1301_ _1301_/A _2006_/B _1300_/Y VGND VGND VPWR VPWR _1301_/Y sky130_fd_sc_hd__nand3_4
X_2281_ _2276_/X _2122_/Y _2278_/X _1620_/B _2280_/X VGND VGND VPWR VPWR _2281_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_64_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1996_ _1995_/Y VGND VGND VPWR VPWR _2017_/D sky130_fd_sc_hd__inv_2
XFILLER_20_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2548_ _2550_/CLK _1894_/X VGND VGND VPWR VPWR _1899_/B sky130_fd_sc_hd__dfxtp_4
X_2617_ _2618_/CLK _1404_/Y VGND VGND VPWR VPWR _1231_/B sky130_fd_sc_hd__dfxtp_4
X_2479_ _2483_/CLK _2065_/X VGND VGND VPWR VPWR _1993_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_55_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1781_ _1781_/A VGND VGND VPWR VPWR _1781_/X sky130_fd_sc_hd__buf_2
X_1850_ _1846_/X _1849_/Y _1628_/X VGND VGND VPWR VPWR _1850_/X sky130_fd_sc_hd__a21o_4
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2333_ _1218_/B _2333_/B VGND VGND VPWR VPWR _2333_/Y sky130_fd_sc_hd__nand2_4
X_2402_ _2445_/CLK _2402_/D VGND VGND VPWR VPWR _1636_/A sky130_fd_sc_hd__dfxtp_4
X_1215_ _1211_/Y _2322_/A _1214_/Y VGND VGND VPWR VPWR _1215_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_37_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2195_ _1534_/A _2552_/Q _2148_/X VGND VGND VPWR VPWR _2195_/Y sky130_fd_sc_hd__o21ai_4
X_2264_ _2263_/X VGND VGND VPWR VPWR _2264_/X sky130_fd_sc_hd__buf_2
XFILLER_52_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1979_ _1979_/A _2496_/Q VGND VGND VPWR VPWR _1979_/X sky130_fd_sc_hd__or2_4
XFILLER_20_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1902_ _1902_/A VGND VGND VPWR VPWR _1902_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1833_ _1178_/A _1735_/D VGND VGND VPWR VPWR _1834_/A sky130_fd_sc_hd__nand2_4
XFILLER_30_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1764_ _1764_/A VGND VGND VPWR VPWR _1764_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2316_ _1766_/B _2311_/X _2268_/A _2313_/X VGND VGND VPWR VPWR _2316_/X sky130_fd_sc_hd__a2bb2o_4
X_1695_ _1694_/X VGND VGND VPWR VPWR _1696_/A sky130_fd_sc_hd__buf_2
X_2247_ _2246_/Y VGND VGND VPWR VPWR _2247_/X sky130_fd_sc_hd__buf_2
X_2178_ _1944_/A _1703_/A VGND VGND VPWR VPWR _2179_/C sky130_fd_sc_hd__nand2_4
XFILLER_40_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_9_0_addressalyzerBlock.SPI_CLK clkbuf_4_9_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2388_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1480_ _1476_/Y _1478_/Y _1479_/Y VGND VGND VPWR VPWR _1480_/Y sky130_fd_sc_hd__a21oi_4
X_2032_ _2029_/Y _2030_/X _2043_/C _2017_/D VGND VGND VPWR VPWR _2032_/X sky130_fd_sc_hd__and4_4
X_2101_ _1221_/A VGND VGND VPWR VPWR _2102_/A sky130_fd_sc_hd__buf_2
X_1678_ _1678_/A VGND VGND VPWR VPWR _1678_/Y sky130_fd_sc_hd__inv_2
X_1816_ _2577_/Q _1810_/X _1813_/X VGND VGND VPWR VPWR _1816_/X sky130_fd_sc_hd__o21a_4
X_1747_ _1625_/X _2431_/Q _1708_/X VGND VGND VPWR VPWR _1747_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2650_ _2457_/CLK _1197_/Y VGND VGND VPWR VPWR _1182_/A sky130_fd_sc_hd__dfxtp_4
X_2581_ _2581_/CLK _1805_/X VGND VGND VPWR VPWR _1514_/A sky130_fd_sc_hd__dfxtp_4
X_1601_ _1555_/A VGND VGND VPWR VPWR _1602_/C sky130_fd_sc_hd__buf_2
X_1532_ _1420_/A _1527_/Y _1556_/A VGND VGND VPWR VPWR _1532_/Y sky130_fd_sc_hd__a21oi_4
X_1394_ _2619_/Q _1383_/A VGND VGND VPWR VPWR _1394_/Y sky130_fd_sc_hd__nor2_4
XFILLER_4_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1463_ _2266_/A _2333_/B _1462_/X VGND VGND VPWR VPWR _1463_/Y sky130_fd_sc_hd__a21oi_4
X_2015_ _2014_/X _1986_/Y _1994_/D VGND VGND VPWR VPWR _2047_/A sky130_fd_sc_hd__nor3_4
XFILLER_35_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_1_0_m1_clk_local clkbuf_2_1_0_m1_clk_local/A VGND VGND VPWR VPWR clkbuf_3_3_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_0_0_addressalyzerBlock.SPI_CLK clkbuf_2_1_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_2_0_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2495_ _2496_/CLK _2495_/D VGND VGND VPWR VPWR _1979_/A sky130_fd_sc_hd__dfxtp_4
X_2633_ _2626_/CLK _2633_/D VGND VGND VPWR VPWR _1244_/B sky130_fd_sc_hd__dfxtp_4
X_2564_ _2557_/CLK _2564_/D VGND VGND VPWR VPWR _2564_/Q sky130_fd_sc_hd__dfxtp_4
X_1515_ _1514_/X _1460_/X _1462_/X VGND VGND VPWR VPWR _1515_/Y sky130_fd_sc_hd__a21oi_4
X_1377_ _1375_/X _1376_/Y VGND VGND VPWR VPWR _1378_/A sky130_fd_sc_hd__nand2_4
X_1446_ _1442_/X _1445_/A _1545_/A VGND VGND VPWR VPWR _1446_/Y sky130_fd_sc_hd__nand3_4
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1231_ _2618_/Q _1231_/B VGND VGND VPWR VPWR _1233_/C sky130_fd_sc_hd__nand2_4
X_1300_ _1260_/Y _1300_/B VGND VGND VPWR VPWR _1300_/Y sky130_fd_sc_hd__nand2_4
X_2280_ _2279_/X VGND VGND VPWR VPWR _2280_/X sky130_fd_sc_hd__buf_2
XFILLER_64_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1995_ _2043_/D _2037_/D VGND VGND VPWR VPWR _1995_/Y sky130_fd_sc_hd__nand2_4
X_2616_ _2618_/CLK _1408_/Y VGND VGND VPWR VPWR _2616_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_9_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2547_ _2550_/CLK _2547_/D VGND VGND VPWR VPWR _2547_/Q sky130_fd_sc_hd__dfxtp_4
X_2478_ _2483_/CLK _2478_/D VGND VGND VPWR VPWR _2478_/Q sky130_fd_sc_hd__dfxtp_4
X_1429_ _1424_/Y _1428_/Y VGND VGND VPWR VPWR _1429_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_4_4_0_m1_clk_local clkbuf_4_5_0_m1_clk_local/A VGND VGND VPWR VPWR _2477_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1780_ _1678_/Y _1780_/B VGND VGND VPWR VPWR _1780_/Y sky130_fd_sc_hd__nand2_4
X_2332_ _1218_/B _2392_/Q _2102_/A _1729_/Y VGND VGND VPWR VPWR _2391_/D sky130_fd_sc_hd__a211o_4
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2401_ _2410_/CLK _2401_/D VGND VGND VPWR VPWR _1768_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_52_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1214_ _2436_/Q _1187_/A _1213_/X VGND VGND VPWR VPWR _1214_/Y sky130_fd_sc_hd__o21ai_4
X_2194_ _1409_/B _1571_/A _1568_/A _1660_/A _2146_/Y VGND VGND VPWR VPWR _2194_/Y
+ sky130_fd_sc_hd__o41ai_4
XFILLER_37_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2263_ _1583_/X _1594_/X _1669_/B _1694_/X _1736_/A VGND VGND VPWR VPWR _2263_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_1_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1978_ _1980_/A _1978_/B _1978_/C VGND VGND VPWR VPWR _1978_/X sky130_fd_sc_hd__and3_4
XFILLER_45_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1832_ _1829_/Y _1830_/Y _1831_/Y VGND VGND VPWR VPWR _2571_/D sky130_fd_sc_hd__a21oi_4
XFILLER_34_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1901_ _2063_/A VGND VGND VPWR VPWR _1901_/X sky130_fd_sc_hd__buf_2
X_1763_ _1740_/Y _1760_/Y _1762_/Y VGND VGND VPWR VPWR _2590_/D sky130_fd_sc_hd__o21ai_4
X_1694_ _2594_/Q VGND VGND VPWR VPWR _1694_/X sky130_fd_sc_hd__buf_2
X_2315_ _1713_/Y _2311_/X _2266_/A _2313_/X VGND VGND VPWR VPWR _2401_/D sky130_fd_sc_hd__a2bb2o_4
X_2246_ _2246_/A VGND VGND VPWR VPWR _2246_/Y sky130_fd_sc_hd__inv_2
X_2177_ _2151_/A _2177_/B VGND VGND VPWR VPWR _2177_/Y sky130_fd_sc_hd__nand2_4
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_14_0_addressalyzerBlock.SPI_CLK clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR _2570_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_21_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2100_ _1781_/X _2099_/C _2098_/Y VGND VGND VPWR VPWR _2462_/D sky130_fd_sc_hd__nor3_4
X_2031_ _2017_/B VGND VGND VPWR VPWR _2043_/C sky130_fd_sc_hd__buf_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1815_ _2577_/Q _1809_/X _1814_/X VGND VGND VPWR VPWR _2578_/D sky130_fd_sc_hd__o21a_4
X_1677_ _1674_/Y _1676_/Y VGND VGND VPWR VPWR _2596_/D sky130_fd_sc_hd__nand2_4
X_1746_ _1746_/A VGND VGND VPWR VPWR _1746_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2229_ _1645_/A _1333_/A _1612_/A VGND VGND VPWR VPWR _2229_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_29_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1531_ _1530_/Y VGND VGND VPWR VPWR _1556_/A sky130_fd_sc_hd__buf_2
X_1600_ _1549_/A _1600_/B VGND VGND VPWR VPWR _1600_/Y sky130_fd_sc_hd__nand2_4
X_1462_ _1450_/X VGND VGND VPWR VPWR _1462_/X sky130_fd_sc_hd__buf_2
X_2580_ _2581_/CLK _1807_/X VGND VGND VPWR VPWR _1520_/A sky130_fd_sc_hd__dfxtp_4
X_1393_ _1385_/D _1379_/X _1392_/Y VGND VGND VPWR VPWR _2620_/D sky130_fd_sc_hd__o21a_4
X_2014_ _1985_/Y VGND VGND VPWR VPWR _2014_/X sky130_fd_sc_hd__buf_2
XFILLER_35_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1729_ _2386_/Q _1566_/A _1689_/Y VGND VGND VPWR VPWR _1729_/Y sky130_fd_sc_hd__nor3_4
XFILLER_64_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2632_ _2626_/CLK _1337_/Y VGND VGND VPWR VPWR _1335_/A sky130_fd_sc_hd__dfxtp_4
X_2563_ _2562_/CLK _1876_/X VGND VGND VPWR VPWR _2563_/Q sky130_fd_sc_hd__dfxtp_4
X_1445_ _1445_/A _1434_/Y _1444_/Y _1445_/D VGND VGND VPWR VPWR _1545_/A sky130_fd_sc_hd__nand4_4
X_2494_ _2388_/CLK _1983_/Y VGND VGND VPWR VPWR _1528_/A sky130_fd_sc_hd__dfxtp_4
X_1514_ _1514_/A VGND VGND VPWR VPWR _1514_/X sky130_fd_sc_hd__buf_2
X_1376_ _1366_/X _1236_/A _1373_/B VGND VGND VPWR VPWR _1376_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_4_12_0_m1_clk_local clkbuf_3_6_0_m1_clk_local/X VGND VGND VPWR VPWR _2367_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1230_ _2616_/Q VGND VGND VPWR VPWR _1397_/B sky130_fd_sc_hd__inv_2
X_1994_ _1985_/Y _1986_/Y _1994_/C _1994_/D VGND VGND VPWR VPWR _1994_/Y sky130_fd_sc_hd__nor4_4
XFILLER_60_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2615_ _2618_/CLK _1412_/X VGND VGND VPWR VPWR _2615_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_9_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2546_ _2550_/CLK _2546_/D VGND VGND VPWR VPWR _2546_/Q sky130_fd_sc_hd__dfxtp_4
X_2477_ _2477_/CLK _2070_/Y VGND VGND VPWR VPWR _2477_/Q sky130_fd_sc_hd__dfxtp_4
X_1428_ _1570_/A _1428_/B _1428_/C _1428_/D VGND VGND VPWR VPWR _1428_/Y sky130_fd_sc_hd__nand4_4
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1359_ _1358_/Y VGND VGND VPWR VPWR _2627_/D sky130_fd_sc_hd__inv_2
XFILLER_34_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2400_ _2606_/CLK _2316_/X VGND VGND VPWR VPWR _1765_/A sky130_fd_sc_hd__dfxtp_4
X_1213_ _2096_/A VGND VGND VPWR VPWR _1213_/X sky130_fd_sc_hd__buf_2
X_2331_ _1222_/X _2330_/Y VGND VGND VPWR VPWR _2390_/D sky130_fd_sc_hd__nor2_4
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2262_ _1649_/B VGND VGND VPWR VPWR _2262_/X sky130_fd_sc_hd__buf_2
X_2193_ _1726_/A _2191_/Y _2192_/Y VGND VGND VPWR VPWR _2193_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_37_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1977_ _1979_/A _2496_/Q _2497_/Q VGND VGND VPWR VPWR _1978_/C sky130_fd_sc_hd__a21o_4
XFILLER_33_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2529_ _2528_/CLK _2529_/D VGND VGND VPWR VPWR _2529_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1900_ _1900_/A _2547_/Q VGND VGND VPWR VPWR _2543_/D sky130_fd_sc_hd__and2_4
X_1831_ _1831_/A _1831_/B VGND VGND VPWR VPWR _1831_/Y sky130_fd_sc_hd__nand2_4
XFILLER_30_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1762_ _1762_/A _1762_/B VGND VGND VPWR VPWR _1762_/Y sky130_fd_sc_hd__nand2_4
X_1693_ _1688_/Y _1690_/Y _1692_/X VGND VGND VPWR VPWR _1693_/Y sky130_fd_sc_hd__o21ai_4
X_2245_ _1219_/X _2245_/B _1691_/Y VGND VGND VPWR VPWR _2246_/A sky130_fd_sc_hd__nor3_4
X_2314_ _1637_/B _2311_/X _1420_/A _2313_/X VGND VGND VPWR VPWR _2402_/D sky130_fd_sc_hd__a2bb2o_4
X_2176_ _2174_/Y _1708_/X _2176_/C VGND VGND VPWR VPWR _2176_/Y sky130_fd_sc_hd__nand3_4
XFILLER_56_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2030_ _2030_/A VGND VGND VPWR VPWR _2030_/X sky130_fd_sc_hd__buf_2
XFILLER_47_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1814_ _2578_/Q _1810_/X _1813_/X VGND VGND VPWR VPWR _1814_/X sky130_fd_sc_hd__o21a_4
X_1745_ _2300_/C _1703_/X _2179_/B _1744_/Y VGND VGND VPWR VPWR _1745_/X sky130_fd_sc_hd__a211o_4
X_1676_ _1726_/A _1676_/B VGND VGND VPWR VPWR _1676_/Y sky130_fd_sc_hd__nand2_4
XFILLER_7_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2228_ _2217_/Y _2226_/Y _2227_/Y VGND VGND VPWR VPWR _2228_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_26_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2159_ _1960_/A _1635_/X _1632_/Y _2158_/Y VGND VGND VPWR VPWR _2159_/X sky130_fd_sc_hd__a211o_4
XFILLER_42_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_0_0_addressalyzerBlock.SPI_CLK clkbuf_2_0_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR clkbuf_4_1_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_13_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1392_ _1379_/X _1385_/D _2063_/A VGND VGND VPWR VPWR _1392_/Y sky130_fd_sc_hd__a21oi_4
X_1530_ _1442_/X _1545_/A _1529_/Y VGND VGND VPWR VPWR _1530_/Y sky130_fd_sc_hd__nand3_4
X_1461_ _1460_/X VGND VGND VPWR VPWR _2333_/B sky130_fd_sc_hd__buf_2
X_2013_ _2002_/X _2003_/Y _2013_/C _2013_/D VGND VGND VPWR VPWR _2019_/B sky130_fd_sc_hd__nor4_4
XFILLER_35_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1728_ _1697_/A _1689_/A _1728_/C VGND VGND VPWR VPWR _1728_/Y sky130_fd_sc_hd__nor3_4
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1659_ _1659_/A VGND VGND VPWR VPWR _1660_/A sky130_fd_sc_hd__buf_2
XFILLER_26_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2562_ _2562_/CLK _2562_/D VGND VGND VPWR VPWR _2562_/Q sky130_fd_sc_hd__dfxtp_4
X_2631_ _2626_/CLK _1341_/X VGND VGND VPWR VPWR _1242_/B sky130_fd_sc_hd__dfxtp_4
X_2493_ _2470_/CLK _2493_/D VGND VGND VPWR VPWR CLK_LED sky130_fd_sc_hd__dfxtp_4
X_1375_ _1236_/A _1373_/X _1374_/X VGND VGND VPWR VPWR _1375_/X sky130_fd_sc_hd__o21a_4
X_1444_ _2385_/Q VGND VGND VPWR VPWR _1444_/Y sky130_fd_sc_hd__inv_2
X_1513_ _1511_/Y _1512_/Y _1508_/X VGND VGND VPWR VPWR _1513_/X sky130_fd_sc_hd__a21o_4
XFILLER_23_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1993_ _1993_/A _1993_/B _1993_/C _1993_/D VGND VGND VPWR VPWR _1994_/D sky130_fd_sc_hd__nand4_4
XFILLER_9_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2545_ _2550_/CLK _2545_/D VGND VGND VPWR VPWR _2351_/A sky130_fd_sc_hd__dfxtp_4
X_2614_ _2618_/CLK _2614_/D VGND VGND VPWR VPWR _1409_/B sky130_fd_sc_hd__dfxtp_4
X_2476_ _2483_/CLK _2075_/Y VGND VGND VPWR VPWR _1990_/B sky130_fd_sc_hd__dfxtp_4
X_1358_ _1358_/A _2006_/B _1358_/C VGND VGND VPWR VPWR _1358_/Y sky130_fd_sc_hd__nand3_4
X_1427_ _1427_/A VGND VGND VPWR VPWR _1428_/D sky130_fd_sc_hd__buf_2
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1289_ _1289_/A _1971_/A _1289_/C VGND VGND VPWR VPWR _1290_/A sky130_fd_sc_hd__nand3_4
XFILLER_11_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2192_ _1762_/A _2437_/Q VGND VGND VPWR VPWR _2192_/Y sky130_fd_sc_hd__nand2_4
X_1212_ _1188_/A VGND VGND VPWR VPWR _2322_/A sky130_fd_sc_hd__buf_2
X_2330_ _2463_/Q _2385_/Q _2322_/A _2333_/B VGND VGND VPWR VPWR _2330_/Y sky130_fd_sc_hd__a22oi_4
X_2261_ _2243_/Y _2260_/Y _2258_/X _1914_/B _2248_/X VGND VGND VPWR VPWR _2427_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_52_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1976_ _1976_/A _1976_/B VGND VGND VPWR VPWR _1980_/A sky130_fd_sc_hd__nor2_4
X_2528_ _2528_/CLK _2528_/D VGND VGND VPWR VPWR _1933_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_45_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2459_ _2570_/CLK _2105_/X VGND VGND VPWR VPWR _2103_/A sky130_fd_sc_hd__dfxtp_4
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_0_0_m1_clk_local clkbuf_4_1_0_m1_clk_local/A VGND VGND VPWR VPWR _2519_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1830_ _1179_/X _1735_/C _1735_/D VGND VGND VPWR VPWR _1830_/Y sky130_fd_sc_hd__nand3_4
X_1761_ _1739_/A VGND VGND VPWR VPWR _1762_/A sky130_fd_sc_hd__buf_2
X_1692_ _1691_/Y _1488_/X _1780_/B _1731_/B VGND VGND VPWR VPWR _1692_/X sky130_fd_sc_hd__a2bb2o_4
X_2313_ _2312_/X VGND VGND VPWR VPWR _2313_/X sky130_fd_sc_hd__buf_2
XFILLER_53_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2244_ _2243_/Y VGND VGND VPWR VPWR _2244_/X sky130_fd_sc_hd__buf_2
X_2175_ _1232_/A _2175_/B VGND VGND VPWR VPWR _2176_/C sky130_fd_sc_hd__nand2_4
XFILLER_15_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1959_ _1969_/A _2515_/Q VGND VGND VPWR VPWR _1959_/X sky130_fd_sc_hd__and2_4
XFILLER_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_6_0_m1_clk_local clkbuf_3_7_0_m1_clk_local/A VGND VGND VPWR VPWR clkbuf_3_6_0_m1_clk_local/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1813_ _1838_/A VGND VGND VPWR VPWR _1813_/X sky130_fd_sc_hd__buf_2
XFILLER_7_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1744_ _1630_/X _1744_/B VGND VGND VPWR VPWR _1744_/Y sky130_fd_sc_hd__nor2_4
X_1675_ _1739_/A VGND VGND VPWR VPWR _1726_/A sky130_fd_sc_hd__buf_2
X_2227_ _1300_/B _1640_/X _1651_/X _1856_/A VGND VGND VPWR VPWR _2227_/Y sky130_fd_sc_hd__a2bb2oi_4
X_2089_ _2089_/A VGND VGND VPWR VPWR _2089_/Y sky130_fd_sc_hd__inv_2
X_2158_ _1703_/X _2158_/B VGND VGND VPWR VPWR _2158_/Y sky130_fd_sc_hd__nor2_4
XFILLER_17_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1391_ _1274_/X VGND VGND VPWR VPWR _2063_/A sky130_fd_sc_hd__buf_2
X_1460_ _2390_/Q VGND VGND VPWR VPWR _1460_/X sky130_fd_sc_hd__buf_2
X_2012_ _2008_/A VGND VGND VPWR VPWR _2013_/D sky130_fd_sc_hd__buf_2
XFILLER_50_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1727_ _1725_/X _1726_/Y VGND VGND VPWR VPWR _2593_/D sky130_fd_sc_hd__nand2_4
X_1658_ _1612_/X _1653_/Y _1657_/Y VGND VGND VPWR VPWR _1658_/Y sky130_fd_sc_hd__o21ai_4
X_1589_ _1426_/A VGND VGND VPWR VPWR _1590_/B sky130_fd_sc_hd__inv_2
XFILLER_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2492_ _2372_/CLK _2492_/D VGND VGND VPWR VPWR _2492_/Q sky130_fd_sc_hd__dfxtp_4
X_2561_ _2550_/CLK _2561_/D VGND VGND VPWR VPWR _2561_/Q sky130_fd_sc_hd__dfxtp_4
X_2630_ _2477_/CLK _1343_/X VGND VGND VPWR VPWR _1242_/C sky130_fd_sc_hd__dfxtp_4
X_1512_ _1486_/A VGND VGND VPWR VPWR _1512_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1374_ _1374_/A VGND VGND VPWR VPWR _1374_/X sky130_fd_sc_hd__buf_2
X_1443_ _1443_/A VGND VGND VPWR VPWR _1445_/A sky130_fd_sc_hd__inv_2
XFILLER_4_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1992_ _1992_/A _1992_/B _2060_/A _1992_/D VGND VGND VPWR VPWR _1993_/B sky130_fd_sc_hd__nor4_4
X_2544_ _2550_/CLK _1899_/X VGND VGND VPWR VPWR _2544_/Q sky130_fd_sc_hd__dfxtp_4
X_2475_ _2477_/CLK _2475_/D VGND VGND VPWR VPWR _2071_/A sky130_fd_sc_hd__dfxtp_4
X_2613_ _2370_/CLK _1419_/X VGND VGND VPWR VPWR _1232_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_55_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1357_ _1228_/Y _1350_/X _1349_/Y VGND VGND VPWR VPWR _1358_/C sky130_fd_sc_hd__o21ai_4
X_1426_ _1426_/A VGND VGND VPWR VPWR _1428_/C sky130_fd_sc_hd__buf_2
X_1288_ _1257_/X _1260_/Y _1225_/X VGND VGND VPWR VPWR _1289_/C sky130_fd_sc_hd__o21ai_4
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2191_ _2351_/A _1739_/B _2190_/Y _2168_/Y VGND VGND VPWR VPWR _2191_/Y sky130_fd_sc_hd__a22oi_4
X_1211_ _2645_/Q _1194_/B _1210_/X VGND VGND VPWR VPWR _1211_/Y sky130_fd_sc_hd__o21ai_4
X_2260_ _1840_/B _1698_/A _1520_/X VGND VGND VPWR VPWR _2260_/Y sky130_fd_sc_hd__nand3_4
XFILLER_52_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1975_ _1976_/A _1976_/B _1975_/C VGND VGND VPWR VPWR _2498_/D sky130_fd_sc_hd__nor3_4
XFILLER_60_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1409_ _1409_/A _1409_/B _1409_/C VGND VGND VPWR VPWR _1409_/Y sky130_fd_sc_hd__nand3_4
X_2458_ _2570_/CLK _2106_/X VGND VGND VPWR VPWR _2105_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_29_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2527_ _2506_/CLK _2527_/D VGND VGND VPWR VPWR _2527_/Q sky130_fd_sc_hd__dfxtp_4
X_2389_ _2390_/CLK _2389_/D VGND VGND VPWR VPWR _1443_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_0_0_addressalyzerBlock.SPI_CLK clkbuf_4_1_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2428_/CLK sky130_fd_sc_hd__clkbuf_1
X_1760_ _1758_/Y _1759_/Y _1673_/C VGND VGND VPWR VPWR _1760_/Y sky130_fd_sc_hd__a21oi_4
X_1691_ _2594_/Q VGND VGND VPWR VPWR _1691_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2312_ _1609_/B _1189_/Y _2245_/B _1694_/X VGND VGND VPWR VPWR _2312_/X sky130_fd_sc_hd__and4_4
XFILLER_38_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2174_ _2151_/A _2174_/B VGND VGND VPWR VPWR _2174_/Y sky130_fd_sc_hd__nand2_4
X_2243_ _1609_/B VGND VGND VPWR VPWR _2243_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1889_ _1891_/A _2560_/Q VGND VGND VPWR VPWR _1889_/X sky130_fd_sc_hd__and2_4
X_1958_ _1969_/A _1958_/B VGND VGND VPWR VPWR _1958_/X sky130_fd_sc_hd__and2_4
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_5_0_addressalyzerBlock.SPI_CLK clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1674_ _1658_/Y _1661_/X _1673_/Y VGND VGND VPWR VPWR _1674_/Y sky130_fd_sc_hd__nand3_4
X_1743_ _2415_/Q VGND VGND VPWR VPWR _1744_/B sky130_fd_sc_hd__inv_2
X_1812_ _2578_/Q _1809_/X _1811_/X VGND VGND VPWR VPWR _2579_/D sky130_fd_sc_hd__o21a_4
X_2226_ _2222_/X _2225_/X _1471_/X VGND VGND VPWR VPWR _2226_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_53_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2088_ _1971_/A _2088_/B VGND VGND VPWR VPWR _2088_/X sky130_fd_sc_hd__and2_4
XFILLER_26_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2157_ _2153_/Y _2156_/Y _1628_/X VGND VGND VPWR VPWR _2157_/X sky130_fd_sc_hd__a21o_4
XFILLER_21_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1390_ _1395_/A _1390_/B _1390_/C VGND VGND VPWR VPWR _1390_/Y sky130_fd_sc_hd__nor3_4
X_2011_ _2011_/A VGND VGND VPWR VPWR _2013_/C sky130_fd_sc_hd__inv_2
XFILLER_50_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1726_ _1726_/A _2593_/Q VGND VGND VPWR VPWR _1726_/Y sky130_fd_sc_hd__nand2_4
X_1657_ _1612_/X _2628_/Q _1656_/X VGND VGND VPWR VPWR _1657_/Y sky130_fd_sc_hd__a21oi_4
X_1588_ _1577_/X _1460_/X _1514_/X VGND VGND VPWR VPWR _1588_/Y sky130_fd_sc_hd__o21ai_4
X_2209_ _1611_/A _1385_/A _1654_/Y VGND VGND VPWR VPWR _2209_/X sky130_fd_sc_hd__a21o_4
XFILLER_26_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2491_ _2470_/CLK _2019_/Y VGND VGND VPWR VPWR _2011_/A sky130_fd_sc_hd__dfxtp_4
X_2560_ _2554_/CLK _2560_/D VGND VGND VPWR VPWR _2560_/Q sky130_fd_sc_hd__dfxtp_4
X_1442_ _1434_/Y _1422_/A _1528_/A VGND VGND VPWR VPWR _1442_/X sky130_fd_sc_hd__a21o_4
XFILLER_4_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1511_ _1505_/B VGND VGND VPWR VPWR _1511_/Y sky130_fd_sc_hd__inv_2
X_1373_ _1379_/A _1373_/B _1383_/C _1365_/D VGND VGND VPWR VPWR _1373_/X sky130_fd_sc_hd__and4_4
XFILLER_63_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1709_ _1709_/A VGND VGND VPWR VPWR _1710_/B sky130_fd_sc_hd__inv_2
XFILLER_64_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1991_ _1991_/A _1991_/B _1991_/C _1991_/D VGND VGND VPWR VPWR _1992_/D sky130_fd_sc_hd__nand4_4
X_2612_ _2390_/CLK _1455_/Y VGND VGND VPWR VPWR _2335_/B sky130_fd_sc_hd__dfxtp_4
X_2543_ _2550_/CLK _2543_/D VGND VGND VPWR VPWR _2543_/Q sky130_fd_sc_hd__dfxtp_4
X_2474_ _2477_/CLK _2474_/D VGND VGND VPWR VPWR _1991_/D sky130_fd_sc_hd__dfxtp_4
X_1425_ _2600_/Q VGND VGND VPWR VPWR _1570_/A sky130_fd_sc_hd__buf_2
XFILLER_55_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1356_ _1356_/A VGND VGND VPWR VPWR _1358_/A sky130_fd_sc_hd__inv_2
X_1287_ _1277_/B VGND VGND VPWR VPWR _1289_/A sky130_fd_sc_hd__inv_2
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1210_ _1206_/A _1178_/A VGND VGND VPWR VPWR _1210_/X sky130_fd_sc_hd__or2_4
X_2190_ _2172_/Y _2188_/Y _2189_/Y VGND VGND VPWR VPWR _2190_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_37_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1974_ _1978_/B _1973_/A _1973_/Y VGND VGND VPWR VPWR _1975_/C sky130_fd_sc_hd__a21oi_4
XFILLER_33_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2457_ _2457_/CLK _2107_/X VGND VGND VPWR VPWR _2093_/B sky130_fd_sc_hd__dfxtp_4
X_1408_ _1395_/A _1408_/B _1407_/Y VGND VGND VPWR VPWR _1408_/Y sky130_fd_sc_hd__nor3_4
X_2388_ _2388_/CLK _2388_/D VGND VGND VPWR VPWR _1566_/A sky130_fd_sc_hd__dfxtp_4
X_2526_ _2528_/CLK _2526_/D VGND VGND VPWR VPWR MACRO_RD_SELECT[3] sky130_fd_sc_hd__dfxtp_4
X_1339_ _1274_/X VGND VGND VPWR VPWR _1339_/X sky130_fd_sc_hd__buf_2
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1690_ _1697_/A _1728_/C _1689_/Y VGND VGND VPWR VPWR _1690_/Y sky130_fd_sc_hd__nor3_4
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2311_ _2310_/X VGND VGND VPWR VPWR _2311_/X sky130_fd_sc_hd__buf_2
X_2242_ _2122_/Y _2239_/Y _2241_/Y VGND VGND VPWR VPWR _2434_/D sky130_fd_sc_hd__o21ai_4
X_2173_ _1534_/A _2553_/Q _2148_/X VGND VGND VPWR VPWR _2173_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_25_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1957_ _1969_/A _1957_/B VGND VGND VPWR VPWR _2509_/D sky130_fd_sc_hd__and2_4
XFILLER_21_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1888_ _1891_/A _2561_/Q VGND VGND VPWR VPWR _2553_/D sky130_fd_sc_hd__and2_4
X_2509_ _2519_/CLK _2509_/D VGND VGND VPWR VPWR DATA_TO_HASH[2] sky130_fd_sc_hd__dfxtp_4
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1811_ _2579_/Q _1810_/X _1799_/X VGND VGND VPWR VPWR _1811_/X sky130_fd_sc_hd__o21a_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1673_ _1739_/A _2166_/A _1673_/C _1739_/B VGND VGND VPWR VPWR _1673_/Y sky130_fd_sc_hd__nor4_4
X_1742_ _1316_/B _1646_/X _1741_/Y VGND VGND VPWR VPWR _1742_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_38_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2225_ _1966_/A _1751_/A _1633_/X _2224_/Y VGND VGND VPWR VPWR _2225_/X sky130_fd_sc_hd__a211o_4
X_2087_ _1284_/X _2078_/X VGND VGND VPWR VPWR _2087_/Y sky130_fd_sc_hd__nor2_4
XFILLER_38_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2156_ _2154_/Y _2179_/B _2156_/C VGND VGND VPWR VPWR _2156_/Y sky130_fd_sc_hd__nand3_4
XFILLER_21_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2010_ _2009_/X _2010_/B _2010_/C VGND VGND VPWR VPWR _2492_/D sky130_fd_sc_hd__and3_4
Xclkbuf_3_2_0_m1_clk_local clkbuf_3_3_0_m1_clk_local/A VGND VGND VPWR VPWR clkbuf_4_5_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
X_1725_ _1722_/Y _1723_/Y _1724_/X VGND VGND VPWR VPWR _1725_/X sky130_fd_sc_hd__a21o_4
X_1656_ _1656_/A VGND VGND VPWR VPWR _1656_/X sky130_fd_sc_hd__buf_2
X_1587_ _1545_/X _1576_/X _1578_/Y _1582_/Y _1586_/X VGND VGND VPWR VPWR _1587_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_7_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2208_ _1242_/C _1646_/A _1741_/Y VGND VGND VPWR VPWR _2208_/X sky130_fd_sc_hd__o21a_4
X_2139_ _1594_/X _2245_/B _1669_/B _2121_/X _1221_/A VGND VGND VPWR VPWR _2139_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_41_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2490_ _2470_/CLK _2490_/D VGND VGND VPWR VPWR _1999_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1510_ _1507_/Y _1509_/X _1454_/X VGND VGND VPWR VPWR _2607_/D sky130_fd_sc_hd__a21oi_4
X_1441_ _1420_/Y _1445_/D _1440_/Y VGND VGND VPWR VPWR _1441_/Y sky130_fd_sc_hd__o21ai_4
X_1372_ _2623_/Q VGND VGND VPWR VPWR _1373_/B sky130_fd_sc_hd__buf_2
XFILLER_48_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1708_ _2448_/Q VGND VGND VPWR VPWR _1708_/X sky130_fd_sc_hd__buf_2
XFILLER_58_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1639_ _1629_/X _1638_/X _1471_/X VGND VGND VPWR VPWR _1639_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_64_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1990_ _2071_/A _1990_/B VGND VGND VPWR VPWR _2060_/A sky130_fd_sc_hd__nand2_4
XFILLER_20_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2542_ _2519_/CLK _1903_/Y VGND VGND VPWR VPWR _2542_/Q sky130_fd_sc_hd__dfxtp_4
X_2611_ _2581_/CLK _2611_/D VGND VGND VPWR VPWR _1438_/B sky130_fd_sc_hd__dfxtp_4
X_1355_ _1354_/Y VGND VGND VPWR VPWR _2628_/D sky130_fd_sc_hd__inv_2
X_2473_ _2477_/CLK _2473_/D VGND VGND VPWR VPWR _1991_/C sky130_fd_sc_hd__dfxtp_4
X_1424_ _1608_/B VGND VGND VPWR VPWR _1424_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1286_ _1284_/X _1261_/Y _1286_/C VGND VGND VPWR VPWR _2640_/D sky130_fd_sc_hd__nor3_4
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_5_0_addressalyzerBlock.SPI_CLK clkbuf_4_5_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2562_/CLK sky130_fd_sc_hd__clkbuf_1
X_1973_ _1973_/A _1980_/B VGND VGND VPWR VPWR _1973_/Y sky130_fd_sc_hd__nor2_4
XFILLER_60_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2525_ _2528_/CLK _2525_/D VGND VGND VPWR VPWR MACRO_RD_SELECT[2] sky130_fd_sc_hd__dfxtp_4
X_2456_ _2457_/CLK _2456_/D VGND VGND VPWR VPWR _2456_/Q sky130_fd_sc_hd__dfxtp_4
X_1407_ _1409_/A _2615_/Q _1409_/B _1409_/C _2616_/Q VGND VGND VPWR VPWR _1407_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1338_ _1324_/X _1335_/D _1329_/X _1321_/X VGND VGND VPWR VPWR _1338_/X sky130_fd_sc_hd__and4_4
X_2387_ _2390_/CLK _2387_/D VGND VGND VPWR VPWR _1683_/A sky130_fd_sc_hd__dfxtp_4
X_1269_ _1374_/A VGND VGND VPWR VPWR _1270_/A sky130_fd_sc_hd__buf_2
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2172_ _2615_/Q _1571_/A _1568_/A _1660_/A _2146_/Y VGND VGND VPWR VPWR _2172_/Y
+ sky130_fd_sc_hd__o41ai_4
X_2241_ _2239_/Y _2298_/B _2434_/Q VGND VGND VPWR VPWR _2241_/Y sky130_fd_sc_hd__nand3_4
X_2310_ _1594_/X _1600_/B _2245_/B _1696_/A _1736_/A VGND VGND VPWR VPWR _2310_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_33_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1887_ _1891_/A _2562_/Q VGND VGND VPWR VPWR _1887_/X sky130_fd_sc_hd__and2_4
X_1956_ _1254_/X VGND VGND VPWR VPWR _1969_/A sky130_fd_sc_hd__buf_2
X_2508_ _2496_/CLK _1958_/X VGND VGND VPWR VPWR DATA_TO_HASH[1] sky130_fd_sc_hd__dfxtp_4
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2439_ _2557_/CLK _2439_/D VGND VGND VPWR VPWR _1966_/A sky130_fd_sc_hd__dfxtp_4
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1741_ _1611_/A VGND VGND VPWR VPWR _1741_/Y sky130_fd_sc_hd__inv_2
X_1810_ _2461_/Q VGND VGND VPWR VPWR _1810_/X sky130_fd_sc_hd__buf_2
XFILLER_11_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1672_ _1672_/A VGND VGND VPWR VPWR _1739_/B sky130_fd_sc_hd__buf_2
XFILLER_7_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2155_ _1941_/A _1703_/A VGND VGND VPWR VPWR _2156_/C sky130_fd_sc_hd__nand2_4
X_2224_ _1703_/X _2223_/Y VGND VGND VPWR VPWR _2224_/Y sky130_fd_sc_hd__nor2_4
XFILLER_53_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2086_ _2078_/X _1991_/B _2085_/Y VGND VGND VPWR VPWR _2086_/X sky130_fd_sc_hd__o21a_4
X_1939_ _1938_/A _1847_/Y VGND VGND VPWR VPWR _2520_/D sky130_fd_sc_hd__nor2_4
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_addressalyzerBlock.SPI_CLK clkbuf_0_addressalyzerBlock.SPI_CLK/X VGND
+ VGND VPWR VPWR clkbuf_2_3_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1724_ _1667_/A _1856_/A _1662_/Y _1672_/A VGND VGND VPWR VPWR _1724_/X sky130_fd_sc_hd__a211o_4
X_1655_ _1654_/Y VGND VGND VPWR VPWR _1656_/A sky130_fd_sc_hd__buf_2
X_1586_ _1549_/A _1583_/X _1781_/A VGND VGND VPWR VPWR _1586_/X sky130_fd_sc_hd__a21o_4
X_2069_ _2058_/X _2060_/Y _2068_/Y VGND VGND VPWR VPWR _2070_/A sky130_fd_sc_hd__o21ai_4
X_2207_ _2195_/Y _2205_/Y _2206_/Y VGND VGND VPWR VPWR _2207_/Y sky130_fd_sc_hd__o21ai_4
X_2138_ _2138_/A VGND VGND VPWR VPWR _2138_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1371_ _1360_/Y _1350_/X _1370_/Y VGND VGND VPWR VPWR _2625_/D sky130_fd_sc_hd__a21oi_4
XFILLER_4_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1440_ _1423_/Y _1440_/B _1435_/Y _1440_/D VGND VGND VPWR VPWR _1440_/Y sky130_fd_sc_hd__nand4_4
XFILLER_48_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1638_ _2125_/C _1751_/A _1633_/X _1637_/Y VGND VGND VPWR VPWR _1638_/X sky130_fd_sc_hd__a211o_4
X_1707_ _2295_/C _1703_/X _2179_/B _1706_/Y VGND VGND VPWR VPWR _1712_/A sky130_fd_sc_hd__a211o_4
X_1569_ _1731_/B _1566_/X _1661_/C VGND VGND VPWR VPWR _1569_/X sky130_fd_sc_hd__o21a_4
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2472_ _2477_/CLK _2086_/X VGND VGND VPWR VPWR _1991_/B sky130_fd_sc_hd__dfxtp_4
X_2541_ _2519_/CLK _1905_/Y VGND VGND VPWR VPWR _2541_/Q sky130_fd_sc_hd__dfxtp_4
X_2610_ _2581_/CLK _1480_/Y VGND VGND VPWR VPWR _1438_/C sky130_fd_sc_hd__dfxtp_4
X_1354_ _1352_/X _1353_/Y VGND VGND VPWR VPWR _1354_/Y sky130_fd_sc_hd__nand2_4
X_1285_ _1225_/X _1226_/Y _1257_/X _1246_/Y _1256_/Y VGND VGND VPWR VPWR _1286_/C
+ sky130_fd_sc_hd__o41a_4
X_1423_ _2335_/B VGND VGND VPWR VPWR _1423_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_10_0_addressalyzerBlock.SPI_CLK clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR _2581_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_6_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1972_ _1979_/A _2496_/Q _2497_/Q VGND VGND VPWR VPWR _1978_/B sky130_fd_sc_hd__nand3_4
XFILLER_33_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2455_ _2457_/CLK _2109_/X VGND VGND VPWR VPWR _2455_/Q sky130_fd_sc_hd__dfxtp_4
X_2524_ _2506_/CLK _2524_/D VGND VGND VPWR VPWR MACRO_RD_SELECT[1] sky130_fd_sc_hd__dfxtp_4
X_1337_ _1336_/Y VGND VGND VPWR VPWR _1337_/Y sky130_fd_sc_hd__inv_2
X_1406_ _1232_/D VGND VGND VPWR VPWR _1409_/C sky130_fd_sc_hd__buf_2
X_2386_ _2570_/CLK _2329_/Y VGND VGND VPWR VPWR _2386_/Q sky130_fd_sc_hd__dfxtp_4
X_1268_ _1268_/A _1719_/A VGND VGND VPWR VPWR _1268_/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1199_ _1194_/A _1179_/X _1198_/X VGND VGND VPWR VPWR _1199_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_51_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2171_ _1726_/A _2169_/Y _2170_/Y VGND VGND VPWR VPWR _2438_/D sky130_fd_sc_hd__o21ai_4
XFILLER_2_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2240_ _1555_/A VGND VGND VPWR VPWR _2298_/B sky130_fd_sc_hd__buf_2
XFILLER_33_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1886_ _1874_/A VGND VGND VPWR VPWR _1891_/A sky130_fd_sc_hd__buf_2
X_1955_ _1952_/A _2518_/Q VGND VGND VPWR VPWR _1955_/X sky130_fd_sc_hd__and2_4
X_2438_ _2550_/CLK _2438_/D VGND VGND VPWR VPWR _2170_/B sky130_fd_sc_hd__dfxtp_4
X_2507_ _2638_/CLK _1959_/X VGND VGND VPWR VPWR DATA_TO_HASH[0] sky130_fd_sc_hd__dfxtp_4
X_2369_ _2370_/CLK _2369_/D VGND VGND VPWR VPWR _2369_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1740_ _1739_/Y VGND VGND VPWR VPWR _1740_/Y sky130_fd_sc_hd__inv_2
X_1671_ _1571_/A _1660_/A _2234_/D VGND VGND VPWR VPWR _1672_/A sky130_fd_sc_hd__nor3_4
XFILLER_30_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2085_ _2078_/X _1991_/B _2063_/A VGND VGND VPWR VPWR _2085_/Y sky130_fd_sc_hd__a21oi_4
X_2223_ _1767_/B VGND VGND VPWR VPWR _2223_/Y sky130_fd_sc_hd__inv_2
X_2154_ _2151_/A _2154_/B VGND VGND VPWR VPWR _2154_/Y sky130_fd_sc_hd__nand2_4
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1869_ _1976_/A _1869_/B VGND VGND VPWR VPWR _1869_/Y sky130_fd_sc_hd__nor2_4
X_1938_ _1938_/A _1937_/Y VGND VGND VPWR VPWR _1938_/Y sky130_fd_sc_hd__nor2_4
XFILLER_29_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1723_ _1656_/X _2619_/Q _2166_/A VGND VGND VPWR VPWR _1723_/Y sky130_fd_sc_hd__a21oi_4
X_1654_ _1570_/A _1568_/A _1659_/A VGND VGND VPWR VPWR _1654_/Y sky130_fd_sc_hd__nor3_4
X_2206_ _1293_/Y _1613_/Y _1651_/A _1649_/Y VGND VGND VPWR VPWR _2206_/Y sky130_fd_sc_hd__a2bb2oi_4
X_1585_ _1736_/A VGND VGND VPWR VPWR _1781_/A sky130_fd_sc_hd__buf_2
X_2068_ _2060_/Y _2058_/X _1283_/X VGND VGND VPWR VPWR _2068_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2137_ _1221_/A _1691_/Y VGND VGND VPWR VPWR _2138_/A sky130_fd_sc_hd__nor2_4
XFILLER_43_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1370_ _1360_/Y _1350_/X _1346_/X VGND VGND VPWR VPWR _1370_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_63_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1706_ _1630_/X _1705_/Y VGND VGND VPWR VPWR _1706_/Y sky130_fd_sc_hd__nor2_4
X_1637_ _1635_/X _1637_/B VGND VGND VPWR VPWR _1637_/Y sky130_fd_sc_hd__nor2_4
XFILLER_58_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1568_ _1568_/A VGND VGND VPWR VPWR _1661_/C sky130_fd_sc_hd__buf_2
X_1499_ _1487_/A VGND VGND VPWR VPWR _1499_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2471_ _2477_/CLK _2087_/Y VGND VGND VPWR VPWR _1991_/A sky130_fd_sc_hd__dfxtp_4
X_2540_ _2519_/CLK _2540_/D VGND VGND VPWR VPWR _2540_/Q sky130_fd_sc_hd__dfxtp_4
X_1422_ _1422_/A VGND VGND VPWR VPWR _1445_/D sky130_fd_sc_hd__buf_2
X_1353_ _1324_/X _2628_/Q _1349_/A VGND VGND VPWR VPWR _1353_/Y sky130_fd_sc_hd__nand3_4
X_1284_ _1283_/X VGND VGND VPWR VPWR _1284_/X sky130_fd_sc_hd__buf_2
XFILLER_51_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1971_ _1971_/A _2503_/Q VGND VGND VPWR VPWR _1971_/X sky130_fd_sc_hd__and2_4
X_2454_ _2457_/CLK _2454_/D VGND VGND VPWR VPWR _2109_/B sky130_fd_sc_hd__dfxtp_4
X_1405_ _1232_/A VGND VGND VPWR VPWR _1409_/A sky130_fd_sc_hd__buf_2
X_2385_ _2570_/CLK _2385_/D VGND VGND VPWR VPWR _2385_/Q sky130_fd_sc_hd__dfxtp_4
X_2523_ _2506_/CLK _2523_/D VGND VGND VPWR VPWR MACRO_RD_SELECT[0] sky130_fd_sc_hd__dfxtp_4
X_1198_ _2648_/Q _1180_/Y VGND VGND VPWR VPWR _1198_/X sky130_fd_sc_hd__or2_4
X_1336_ _1331_/X _1335_/Y VGND VGND VPWR VPWR _1336_/Y sky130_fd_sc_hd__nand2_4
X_1267_ _1262_/C VGND VGND VPWR VPWR _1719_/A sky130_fd_sc_hd__inv_2
XFILLER_51_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0_addressalyzerBlock.SPI_CLK _2347_/X VGND VGND VPWR VPWR clkbuf_0_addressalyzerBlock.SPI_CLK/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_19_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2170_ _1762_/A _2170_/B VGND VGND VPWR VPWR _2170_/Y sky130_fd_sc_hd__nand2_4
XFILLER_18_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1954_ _1952_/A _2519_/Q VGND VGND VPWR VPWR _1954_/X sky130_fd_sc_hd__and2_4
XFILLER_21_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_1_0_addressalyzerBlock.SPI_CLK clkbuf_2_1_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_2_1_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
X_1885_ _1885_/A _2563_/Q VGND VGND VPWR VPWR _1885_/X sky130_fd_sc_hd__and2_4
X_2368_ _2372_/CLK _2367_/Q VGND VGND VPWR VPWR _2369_/D sky130_fd_sc_hd__dfxtp_4
Xclkbuf_4_7_0_m1_clk_local clkbuf_4_7_0_m1_clk_local/A VGND VGND VPWR VPWR _2470_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_2437_ _2590_/CLK _2193_/Y VGND VGND VPWR VPWR _2437_/Q sky130_fd_sc_hd__dfxtp_4
X_2506_ _2506_/CLK _2506_/D VGND VGND VPWR VPWR _1968_/B sky130_fd_sc_hd__dfxtp_4
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1319_ _1319_/A _1318_/Y VGND VGND VPWR VPWR _1319_/Y sky130_fd_sc_hd__nand2_4
XFILLER_24_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2299_ _2268_/Y _2291_/X _2298_/Y VGND VGND VPWR VPWR _2299_/Y sky130_fd_sc_hd__o21ai_4
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1670_ _1669_/Y VGND VGND VPWR VPWR _2234_/D sky130_fd_sc_hd__inv_2
XFILLER_7_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2222_ _2219_/Y _2221_/Y _1628_/X VGND VGND VPWR VPWR _2222_/X sky130_fd_sc_hd__a21o_4
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2084_ _2084_/A _2044_/B _2084_/C VGND VGND VPWR VPWR _2473_/D sky130_fd_sc_hd__and3_4
XFILLER_38_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2153_ _2151_/Y _1708_/X _2153_/C VGND VGND VPWR VPWR _2153_/Y sky130_fd_sc_hd__nand3_4
X_1937_ _1937_/A VGND VGND VPWR VPWR _1937_/Y sky130_fd_sc_hd__inv_2
X_1868_ _2567_/Q _1976_/B VGND VGND VPWR VPWR _1869_/B sky130_fd_sc_hd__xnor2_4
X_1799_ _1555_/A VGND VGND VPWR VPWR _1799_/X sky130_fd_sc_hd__buf_2
XFILLER_29_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1722_ _1700_/X _1720_/Y _1721_/Y VGND VGND VPWR VPWR _1722_/Y sky130_fd_sc_hd__o21ai_4
X_1653_ _1642_/Y _1646_/X _1652_/X VGND VGND VPWR VPWR _1653_/Y sky130_fd_sc_hd__a21oi_4
X_1584_ _1219_/X VGND VGND VPWR VPWR _1736_/A sky130_fd_sc_hd__buf_2
X_2205_ _2202_/X _2204_/X _1701_/A VGND VGND VPWR VPWR _2205_/Y sky130_fd_sc_hd__a21oi_4
X_2067_ _2063_/A _1993_/B _2066_/Y VGND VGND VPWR VPWR _2478_/D sky130_fd_sc_hd__nor3_4
XFILLER_41_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2136_ _2253_/C VGND VGND VPWR VPWR _2136_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1705_ _2417_/Q VGND VGND VPWR VPWR _1705_/Y sky130_fd_sc_hd__inv_2
X_1567_ _1428_/B _1428_/C _1428_/D VGND VGND VPWR VPWR _1568_/A sky130_fd_sc_hd__nand3_4
X_1636_ _1636_/A VGND VGND VPWR VPWR _1637_/B sky130_fd_sc_hd__inv_2
XFILLER_39_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2119_ _2119_/A VGND VGND VPWR VPWR _2123_/A sky130_fd_sc_hd__inv_2
X_1498_ _2253_/C _2333_/B _1462_/X VGND VGND VPWR VPWR _1498_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_13_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_15_0_addressalyzerBlock.SPI_CLK clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR _2457_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_54_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2470_ _2470_/CLK _2088_/X VGND VGND VPWR VPWR HASH_EN sky130_fd_sc_hd__dfxtp_4
X_1421_ _2390_/Q VGND VGND VPWR VPWR _1422_/A sky130_fd_sc_hd__inv_2
X_1283_ _2363_/Q VGND VGND VPWR VPWR _1283_/X sky130_fd_sc_hd__buf_2
XFILLER_48_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1352_ _2628_/Q _1356_/A _1306_/X VGND VGND VPWR VPWR _1352_/X sky130_fd_sc_hd__o21a_4
X_2599_ _2590_/CLK _1587_/Y VGND VGND VPWR VPWR _1428_/B sky130_fd_sc_hd__dfxtp_4
X_1619_ _1619_/A VGND VGND VPWR VPWR _1620_/B sky130_fd_sc_hd__inv_2
XFILLER_39_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1970_ _1971_/A _2504_/Q VGND VGND VPWR VPWR _2500_/D sky130_fd_sc_hd__and2_4
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2522_ _2528_/CLK _2522_/D VGND VGND VPWR VPWR _1951_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_4_15_0_m1_clk_local clkbuf_3_7_0_m1_clk_local/X VGND VGND VPWR VPWR _2496_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_2384_ _2550_/CLK _2384_/D VGND VGND VPWR VPWR _2384_/Q sky130_fd_sc_hd__dfxtp_4
X_1404_ _1404_/A VGND VGND VPWR VPWR _1404_/Y sky130_fd_sc_hd__inv_2
X_1335_ _1335_/A _1333_/Y _1335_/C _1335_/D VGND VGND VPWR VPWR _1335_/Y sky130_fd_sc_hd__nand4_4
X_2453_ _2390_/CLK _2111_/Y VGND VGND VPWR VPWR _2099_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_56_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1197_ _1195_/Y _1187_/X _1196_/Y VGND VGND VPWR VPWR _1197_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_36_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1266_ _1277_/D _1265_/Y _1224_/A _1249_/Y VGND VGND VPWR VPWR _1268_/A sky130_fd_sc_hd__nand4_4
XFILLER_51_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1884_ _1885_/A _2564_/Q VGND VGND VPWR VPWR _2556_/D sky130_fd_sc_hd__and2_4
X_1953_ _1952_/A _1953_/B VGND VGND VPWR VPWR _1953_/X sky130_fd_sc_hd__and2_4
X_2505_ _2641_/CLK _1963_/Y VGND VGND VPWR VPWR _2505_/Q sky130_fd_sc_hd__dfxtp_4
X_2367_ _2367_/CLK _1864_/A VGND VGND VPWR VPWR _2367_/Q sky130_fd_sc_hd__dfxtp_4
X_2436_ _2590_/CLK _2215_/Y VGND VGND VPWR VPWR _2436_/Q sky130_fd_sc_hd__dfxtp_4
X_1318_ _1318_/A _1318_/B _1316_/B _1316_/D VGND VGND VPWR VPWR _1318_/Y sky130_fd_sc_hd__nand4_4
X_2298_ _2304_/A _2298_/B ID_toHost VGND VGND VPWR VPWR _2298_/Y sky130_fd_sc_hd__nand3_4
XFILLER_64_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1249_ _1249_/A VGND VGND VPWR VPWR _1249_/Y sky130_fd_sc_hd__inv_2
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2221_ _1948_/Y _1624_/X _2220_/Y VGND VGND VPWR VPWR _2221_/Y sky130_fd_sc_hd__o21ai_4
X_2152_ HASH_LED _2175_/B VGND VGND VPWR VPWR _2153_/C sky130_fd_sc_hd__nand2_4
XFILLER_46_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2083_ _2078_/X _1991_/B _1991_/C VGND VGND VPWR VPWR _2084_/A sky130_fd_sc_hd__a21o_4
X_1867_ _1973_/A _2497_/Q _1980_/B VGND VGND VPWR VPWR _1976_/B sky130_fd_sc_hd__nor3_4
X_1936_ _1938_/A _1622_/Y VGND VGND VPWR VPWR _2522_/D sky130_fd_sc_hd__nor2_4
XFILLER_21_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1798_ _1983_/B _2576_/Q _1797_/X VGND VGND VPWR VPWR _1798_/X sky130_fd_sc_hd__o21a_4
XFILLER_16_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2419_ _2408_/CLK _2419_/D VGND VGND VPWR VPWR _1948_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_40_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1721_ _1612_/X _1349_/Y _1656_/X VGND VGND VPWR VPWR _1721_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_43_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1652_ _1856_/A _2636_/Q _1651_/X VGND VGND VPWR VPWR _1652_/X sky130_fd_sc_hd__and3_4
X_1583_ _1559_/B VGND VGND VPWR VPWR _1583_/X sky130_fd_sc_hd__buf_2
X_2135_ _2120_/X _2133_/Y _2134_/Y VGND VGND VPWR VPWR _2135_/Y sky130_fd_sc_hd__o21ai_4
X_2204_ _1964_/A _1635_/X _1632_/Y _2203_/Y VGND VGND VPWR VPWR _2204_/X sky130_fd_sc_hd__a211o_4
X_2066_ _2060_/Y _2058_/X _2062_/B VGND VGND VPWR VPWR _2066_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_22_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1919_ _1918_/A _2539_/Q VGND VGND VPWR VPWR _2533_/D sky130_fd_sc_hd__and2_4
XFILLER_57_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1704_ _1617_/Y VGND VGND VPWR VPWR _2179_/B sky130_fd_sc_hd__buf_2
X_1566_ _1566_/A VGND VGND VPWR VPWR _1566_/X sky130_fd_sc_hd__buf_2
X_1497_ _1497_/A VGND VGND VPWR VPWR _2253_/C sky130_fd_sc_hd__buf_2
X_1635_ _1703_/A VGND VGND VPWR VPWR _1635_/X sky130_fd_sc_hd__buf_2
X_2049_ _2049_/A _2006_/B _2048_/Y VGND VGND VPWR VPWR _2049_/Y sky130_fd_sc_hd__nand3_4
XFILLER_54_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2118_ _1590_/B _1579_/X _1669_/B _1694_/X VGND VGND VPWR VPWR _2119_/A sky130_fd_sc_hd__and4_4
XFILLER_14_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1351_ _1349_/Y _1228_/Y _1350_/X VGND VGND VPWR VPWR _1356_/A sky130_fd_sc_hd__nor3_4
X_1420_ _1420_/A VGND VGND VPWR VPWR _1420_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1282_ _1281_/Y _2010_/B _1282_/C VGND VGND VPWR VPWR _1282_/X sky130_fd_sc_hd__and3_4
XFILLER_0_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1618_ _2447_/Q VGND VGND VPWR VPWR _2175_/B sky130_fd_sc_hd__buf_2
XFILLER_59_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1549_ _1549_/A VGND VGND VPWR VPWR _1549_/Y sky130_fd_sc_hd__inv_2
X_2598_ _2598_/CLK _2598_/D VGND VGND VPWR VPWR _1426_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_54_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_1_0_addressalyzerBlock.SPI_CLK clkbuf_2_0_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR clkbuf_4_3_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_45_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2521_ _2641_/CLK _1938_/Y VGND VGND VPWR VPWR _2521_/Q sky130_fd_sc_hd__dfxtp_4
X_2383_ _2550_/CLK _2383_/D VGND VGND VPWR VPWR _2384_/D sky130_fd_sc_hd__dfxtp_4
X_1403_ _1231_/B _1408_/B _1402_/Y VGND VGND VPWR VPWR _1404_/A sky130_fd_sc_hd__o21ai_4
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1334_ _1242_/C VGND VGND VPWR VPWR _1335_/D sky130_fd_sc_hd__buf_2
X_2452_ _2570_/CLK _2112_/Y VGND VGND VPWR VPWR _2452_/Q sky130_fd_sc_hd__dfxtp_4
X_1265_ _1257_/X _1260_/Y VGND VGND VPWR VPWR _1265_/Y sky130_fd_sc_hd__nor2_4
X_1196_ _1862_/B _1216_/B _1191_/X VGND VGND VPWR VPWR _1196_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_24_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_0_0_m1_clk_local clkbuf_2_1_0_m1_clk_local/A VGND VGND VPWR VPWR clkbuf_3_1_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1883_ _1885_/A _2565_/Q VGND VGND VPWR VPWR _2557_/D sky130_fd_sc_hd__and2_4
X_1952_ _1952_/A _2521_/Q VGND VGND VPWR VPWR _1952_/X sky130_fd_sc_hd__and2_4
XFILLER_14_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2435_ _2590_/CLK _2237_/Y VGND VGND VPWR VPWR _1218_/A sky130_fd_sc_hd__dfxtp_4
X_2504_ _2638_/CLK _1965_/Y VGND VGND VPWR VPWR _2504_/Q sky130_fd_sc_hd__dfxtp_4
X_2366_ _2367_/CLK _2365_/Q VGND VGND VPWR VPWR _1864_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_56_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1317_ _1318_/A _1316_/X _1306_/X VGND VGND VPWR VPWR _1319_/A sky130_fd_sc_hd__o21a_4
X_1248_ _1277_/A _2641_/Q VGND VGND VPWR VPWR _1249_/A sky130_fd_sc_hd__nand2_4
X_2297_ _2290_/Y VGND VGND VPWR VPWR _2304_/A sky130_fd_sc_hd__buf_2
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1179_ _1179_/A VGND VGND VPWR VPWR _1179_/X sky130_fd_sc_hd__buf_2
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2082_ _2081_/X _2044_/B _2060_/B VGND VGND VPWR VPWR _2474_/D sky130_fd_sc_hd__and3_4
X_2220_ _1625_/X _1913_/A _2448_/Q VGND VGND VPWR VPWR _2220_/Y sky130_fd_sc_hd__a21oi_4
X_2151_ _2151_/A _2151_/B VGND VGND VPWR VPWR _2151_/Y sky130_fd_sc_hd__nand2_4
XFILLER_21_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1866_ _1979_/A _2496_/Q VGND VGND VPWR VPWR _1980_/B sky130_fd_sc_hd__nand2_4
X_1797_ _1788_/X _1490_/A _2326_/A VGND VGND VPWR VPWR _1797_/X sky130_fd_sc_hd__o21a_4
X_1935_ _1339_/X VGND VGND VPWR VPWR _1938_/A sky130_fd_sc_hd__buf_2
XFILLER_21_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2418_ _2445_/CLK _2281_/Y VGND VGND VPWR VPWR _1619_/A sky130_fd_sc_hd__dfxtp_4
X_2349_ _2349_/A MISO_fromClient VGND VGND VPWR VPWR _2349_/Y sky130_fd_sc_hd__nor2_4
XFILLER_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_3_0_m1_clk_local clkbuf_4_3_0_m1_clk_local/A VGND VGND VPWR VPWR _2641_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1651_ _1651_/A VGND VGND VPWR VPWR _1651_/X sky130_fd_sc_hd__buf_2
X_1720_ _1718_/Y _1719_/X _1645_/A VGND VGND VPWR VPWR _1720_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_7_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1582_ _1581_/X _1562_/Y _1569_/X VGND VGND VPWR VPWR _1582_/Y sky130_fd_sc_hd__o21ai_4
X_2065_ _2055_/X _1993_/B _2064_/Y VGND VGND VPWR VPWR _2065_/X sky130_fd_sc_hd__o21a_4
X_2134_ _2123_/A _2335_/A _2134_/C VGND VGND VPWR VPWR _2134_/Y sky130_fd_sc_hd__nand3_4
X_2203_ _2181_/A _1764_/Y VGND VGND VPWR VPWR _2203_/Y sky130_fd_sc_hd__nor2_4
XFILLER_34_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1849_ _1847_/Y _1624_/X _1848_/Y VGND VGND VPWR VPWR _1849_/Y sky130_fd_sc_hd__o21ai_4
X_1918_ _1918_/A _2540_/Q VGND VGND VPWR VPWR _1918_/X sky130_fd_sc_hd__and2_4
XFILLER_40_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1634_ _2447_/Q VGND VGND VPWR VPWR _1703_/A sky130_fd_sc_hd__buf_2
X_1703_ _1703_/A VGND VGND VPWR VPWR _1703_/X sky130_fd_sc_hd__buf_2
X_1565_ _2386_/Q VGND VGND VPWR VPWR _1731_/B sky130_fd_sc_hd__buf_2
X_1496_ _1487_/A _1494_/X _1495_/Y VGND VGND VPWR VPWR _1496_/Y sky130_fd_sc_hd__o21ai_4
X_2048_ _2014_/X _2040_/X _1986_/Y VGND VGND VPWR VPWR _2048_/Y sky130_fd_sc_hd__o21ai_4
X_2117_ _1602_/Y VGND VGND VPWR VPWR _2117_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1350_ _1238_/Y VGND VGND VPWR VPWR _1350_/X sky130_fd_sc_hd__buf_2
X_1281_ _1256_/Y _1225_/X _1257_/X _1260_/Y _1280_/Y VGND VGND VPWR VPWR _1281_/Y
+ sky130_fd_sc_hd__o41ai_4
X_2597_ _2598_/CLK _1603_/Y VGND VGND VPWR VPWR _1427_/A sky130_fd_sc_hd__dfxtp_4
X_1617_ _2448_/Q VGND VGND VPWR VPWR _1617_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1548_ _2602_/Q _1537_/X _1451_/X _1548_/D VGND VGND VPWR VPWR _1548_/Y sky130_fd_sc_hd__nor4_4
X_1479_ _1456_/X _1449_/B _1213_/X VGND VGND VPWR VPWR _1479_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_42_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1402_ _1408_/B _1231_/B _1283_/X VGND VGND VPWR VPWR _1402_/Y sky130_fd_sc_hd__a21oi_4
X_2451_ _2390_/CLK _2113_/X VGND VGND VPWR VPWR _1779_/C sky130_fd_sc_hd__dfxtp_4
X_2520_ _2528_/CLK _2520_/D VGND VGND VPWR VPWR _1953_/B sky130_fd_sc_hd__dfxtp_4
X_2382_ _2372_/CLK _2341_/Y VGND VGND VPWR VPWR _2363_/D sky130_fd_sc_hd__dfxtp_4
X_1333_ _1333_/A _1228_/Y _1240_/Y _1238_/Y VGND VGND VPWR VPWR _1333_/Y sky130_fd_sc_hd__nor4_4
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1264_ _1263_/Y VGND VGND VPWR VPWR _1264_/Y sky130_fd_sc_hd__inv_2
X_1195_ _1182_/A _1179_/X _1194_/X VGND VGND VPWR VPWR _1195_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_51_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2649_ _2457_/CLK _1201_/Y VGND VGND VPWR VPWR _1194_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_42_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1882_ _1885_/A _2566_/Q VGND VGND VPWR VPWR _2558_/D sky130_fd_sc_hd__and2_4
X_1951_ _1952_/A _1951_/B VGND VGND VPWR VPWR _1951_/X sky130_fd_sc_hd__and2_4
X_2365_ _2372_/CLK _2365_/D VGND VGND VPWR VPWR _2365_/Q sky130_fd_sc_hd__dfxtp_4
X_2503_ _2641_/CLK _2503_/D VGND VGND VPWR VPWR _2503_/Q sky130_fd_sc_hd__dfxtp_4
X_2434_ _2557_/CLK _2434_/D VGND VGND VPWR VPWR _2434_/Q sky130_fd_sc_hd__dfxtp_4
X_1178_ _1178_/A VGND VGND VPWR VPWR _1179_/A sky130_fd_sc_hd__buf_2
X_1316_ _1239_/Y _1316_/B _1241_/Y _1316_/D VGND VGND VPWR VPWR _1316_/X sky130_fd_sc_hd__and4_4
X_1247_ _1225_/X _1226_/Y _1257_/A _1246_/Y VGND VGND VPWR VPWR _1277_/B sky130_fd_sc_hd__nor4_4
X_2296_ _2266_/Y _2291_/X _2295_/Y VGND VGND VPWR VPWR _2296_/Y sky130_fd_sc_hd__o21ai_4
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_11_0_m1_clk_local clkbuf_3_5_0_m1_clk_local/X VGND VGND VPWR VPWR _2506_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2081_ _1991_/D _2080_/Y VGND VGND VPWR VPWR _2081_/X sky130_fd_sc_hd__or2_4
X_2150_ _1623_/Y VGND VGND VPWR VPWR _2151_/A sky130_fd_sc_hd__buf_2
XFILLER_46_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1934_ _1932_/A _2527_/Q VGND VGND VPWR VPWR _2523_/D sky130_fd_sc_hd__and2_4
X_1865_ _2365_/Q _2365_/D _1865_/C VGND VGND VPWR VPWR _1976_/A sky130_fd_sc_hd__nor3_4
X_1796_ _1983_/B _2577_/Q _1795_/X VGND VGND VPWR VPWR _1796_/X sky130_fd_sc_hd__o21a_4
X_2348_ _2464_/Q VGND VGND VPWR VPWR _2348_/Y sky130_fd_sc_hd__inv_2
X_2417_ _2428_/CLK _2417_/D VGND VGND VPWR VPWR _2417_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_29_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2279_ _1583_/X _1600_/B _1428_/C _1694_/X _1219_/X VGND VGND VPWR VPWR _2279_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_52_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1650_ _1649_/Y VGND VGND VPWR VPWR _1856_/A sky130_fd_sc_hd__buf_2
X_1581_ _2245_/B VGND VGND VPWR VPWR _1581_/X sky130_fd_sc_hd__buf_2
X_2202_ _2198_/Y _2201_/Y _2449_/Q VGND VGND VPWR VPWR _2202_/X sky130_fd_sc_hd__a21o_4
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2064_ _2058_/X _2060_/Y _2062_/B _2055_/X _1275_/X VGND VGND VPWR VPWR _2064_/Y
+ sky130_fd_sc_hd__a41oi_4
X_2133_ _1874_/A _2121_/X _1490_/A VGND VGND VPWR VPWR _2133_/Y sky130_fd_sc_hd__nand3_4
X_1917_ _1918_/A _2541_/Q VGND VGND VPWR VPWR _1917_/X sky130_fd_sc_hd__and2_4
X_1779_ _1778_/X _1678_/A _1779_/C VGND VGND VPWR VPWR _1779_/Y sky130_fd_sc_hd__nand3_4
XFILLER_1_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1848_ _1625_/X _1902_/A _2448_/Q VGND VGND VPWR VPWR _1848_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_17_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_1_0_addressalyzerBlock.SPI_CLK clkbuf_4_1_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2408_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_16_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1564_ _1530_/Y _1563_/Y VGND VGND VPWR VPWR _1564_/X sky130_fd_sc_hd__or2_4
X_1702_ _1701_/Y VGND VGND VPWR VPWR _1702_/Y sky130_fd_sc_hd__inv_2
X_1633_ _1632_/Y VGND VGND VPWR VPWR _1633_/X sky130_fd_sc_hd__buf_2
X_1495_ _1487_/A _1505_/B _1494_/B _1505_/C _2340_/C VGND VGND VPWR VPWR _1495_/Y
+ sky130_fd_sc_hd__a41oi_4
X_2047_ _2047_/A VGND VGND VPWR VPWR _2049_/A sky130_fd_sc_hd__inv_2
XFILLER_62_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2116_ _1545_/X _1576_/X _1588_/Y _1593_/Y _1595_/X VGND VGND VPWR VPWR _2448_/D
+ sky130_fd_sc_hd__a41oi_4
XFILLER_10_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_addressalyzerBlock.SPI_CLK clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_3_6_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1280_ _2641_/Q VGND VGND VPWR VPWR _1280_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2596_ _2590_/CLK _2596_/D VGND VGND VPWR VPWR _1676_/B sky130_fd_sc_hd__dfxtp_4
X_1547_ _1443_/A _2390_/Q _1477_/A VGND VGND VPWR VPWR _1547_/X sky130_fd_sc_hd__o21a_4
X_1616_ _2447_/Q VGND VGND VPWR VPWR _2181_/A sky130_fd_sc_hd__buf_2
XFILLER_27_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1478_ _2268_/A _2333_/B _1462_/X VGND VGND VPWR VPWR _1478_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_2_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2381_ _2498_/CLK _2381_/D VGND VGND VPWR VPWR _2383_/D sky130_fd_sc_hd__dfxtp_4
X_1401_ _1397_/B _1397_/C VGND VGND VPWR VPWR _1408_/B sky130_fd_sc_hd__nor2_4
XFILLER_5_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2450_ _2390_/CLK _2114_/X VGND VGND VPWR VPWR _2113_/B sky130_fd_sc_hd__dfxtp_4
X_1194_ _1194_/A _1194_/B VGND VGND VPWR VPWR _1194_/X sky130_fd_sc_hd__or2_4
X_1332_ _2629_/Q VGND VGND VPWR VPWR _1333_/A sky130_fd_sc_hd__inv_2
X_1263_ _1263_/A _1971_/A _1263_/C VGND VGND VPWR VPWR _1263_/Y sky130_fd_sc_hd__nand3_4
XFILLER_17_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2648_ _2457_/CLK _1205_/Y VGND VGND VPWR VPWR _2648_/Q sky130_fd_sc_hd__dfxtp_4
X_2579_ _2606_/CLK _2579_/D VGND VGND VPWR VPWR _2579_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_35_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1950_ _1254_/X VGND VGND VPWR VPWR _1952_/A sky130_fd_sc_hd__buf_2
X_1881_ _1885_/A DATA_FROM_HASH[0] VGND VGND VPWR VPWR _2559_/D sky130_fd_sc_hd__and2_4
X_2502_ _2513_/CLK _2502_/D VGND VGND VPWR VPWR MACRO_WR_SELECT[3] sky130_fd_sc_hd__dfxtp_4
X_2364_ _2372_/CLK _2363_/Q VGND VGND VPWR VPWR _2365_/D sky130_fd_sc_hd__dfxtp_4
X_1315_ _1244_/B VGND VGND VPWR VPWR _1316_/B sky130_fd_sc_hd__buf_2
X_2433_ _2428_/CLK _2433_/D VGND VGND VPWR VPWR _1709_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_52_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1246_ _1239_/Y _1241_/Y _1243_/X _1246_/D VGND VGND VPWR VPWR _1246_/Y sky130_fd_sc_hd__nand4_4
X_2295_ _2292_/X _2298_/B _2295_/C VGND VGND VPWR VPWR _2295_/Y sky130_fd_sc_hd__nand3_4
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2080_ _2084_/C VGND VGND VPWR VPWR _2080_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1933_ _1932_/A _1933_/B VGND VGND VPWR VPWR _2524_/D sky130_fd_sc_hd__and2_4
X_1864_ _1864_/A VGND VGND VPWR VPWR _1865_/C sky130_fd_sc_hd__inv_2
X_1795_ _1788_/X _2268_/A _2326_/A VGND VGND VPWR VPWR _1795_/X sky130_fd_sc_hd__o21a_4
X_2347_ _2567_/Q S1_CLK_SELECT _2346_/Y VGND VGND VPWR VPWR _2347_/X sky130_fd_sc_hd__o21a_4
XFILLER_29_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2416_ _2445_/CLK _2416_/D VGND VGND VPWR VPWR _1844_/A sky130_fd_sc_hd__dfxtp_4
X_2278_ _2278_/A VGND VGND VPWR VPWR _2278_/X sky130_fd_sc_hd__buf_2
X_1229_ _2619_/Q VGND VGND VPWR VPWR _1233_/A sky130_fd_sc_hd__inv_2
XFILLER_37_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1580_ _1579_/X VGND VGND VPWR VPWR _2245_/B sky130_fd_sc_hd__buf_2
XFILLER_7_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2132_ _2120_/X _2130_/Y _2131_/Y VGND VGND VPWR VPWR _2444_/D sky130_fd_sc_hd__o21ai_4
XFILLER_3_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2201_ _2199_/Y _2179_/B _2201_/C VGND VGND VPWR VPWR _2201_/Y sky130_fd_sc_hd__nand3_4
X_2063_ _2063_/A _2061_/Y _2062_/X VGND VGND VPWR VPWR _2480_/D sky130_fd_sc_hd__nor3_4
XFILLER_19_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1847_ _1847_/A VGND VGND VPWR VPWR _1847_/Y sky130_fd_sc_hd__inv_2
X_1916_ _1918_/A _2542_/Q VGND VGND VPWR VPWR _1916_/X sky130_fd_sc_hd__and2_4
X_1778_ _1783_/B _1783_/D _1440_/D VGND VGND VPWR VPWR _1778_/X sky130_fd_sc_hd__a21o_4
XFILLER_57_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1701_ _1701_/A _1701_/B VGND VGND VPWR VPWR _1701_/Y sky130_fd_sc_hd__nand2_4
XPHY_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1563_ _1435_/Y _1667_/A _1562_/Y _1497_/A _1527_/Y VGND VGND VPWR VPWR _1563_/Y
+ sky130_fd_sc_hd__a32oi_4
X_1494_ _1433_/A _1494_/B _1505_/C _1438_/D VGND VGND VPWR VPWR _1494_/X sky130_fd_sc_hd__and4_4
X_1632_ _2449_/Q VGND VGND VPWR VPWR _1632_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2115_ _1545_/X _1576_/X _1578_/Y _1582_/Y _1586_/X VGND VGND VPWR VPWR _2449_/D
+ sky130_fd_sc_hd__a41oi_4
X_2046_ _1395_/A _1994_/Y _2046_/C VGND VGND VPWR VPWR _2046_/Y sky130_fd_sc_hd__nor3_4
XFILLER_60_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_5_0_m1_clk_local clkbuf_3_4_0_m1_clk_local/A VGND VGND VPWR VPWR clkbuf_3_5_0_m1_clk_local/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2595_ _2390_/CLK _1686_/Y VGND VGND VPWR VPWR _1678_/A sky130_fd_sc_hd__dfxtp_4
X_1546_ _1544_/Y _1442_/X _1545_/X _1529_/Y _1467_/Y VGND VGND VPWR VPWR _1546_/X
+ sky130_fd_sc_hd__a41o_4
X_1615_ _1534_/X _2558_/Q _1614_/X VGND VGND VPWR VPWR _1615_/Y sky130_fd_sc_hd__o21ai_4
X_1477_ _1477_/A VGND VGND VPWR VPWR _2268_/A sky130_fd_sc_hd__buf_2
XFILLER_54_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2029_ _2014_/X _1994_/D VGND VGND VPWR VPWR _2029_/Y sky130_fd_sc_hd__nor2_4
XFILLER_24_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2380_ _2498_/CLK _2379_/Q VGND VGND VPWR VPWR _2381_/D sky130_fd_sc_hd__dfxtp_4
X_1400_ _1400_/A VGND VGND VPWR VPWR _1400_/Y sky130_fd_sc_hd__inv_2
X_1331_ _1335_/A _1330_/X _1306_/X VGND VGND VPWR VPWR _1331_/X sky130_fd_sc_hd__o21a_4
X_1193_ _1183_/Y _1187_/X _1192_/Y VGND VGND VPWR VPWR _1193_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_36_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1262_ _1251_/A _1261_/Y _1262_/C _1249_/Y VGND VGND VPWR VPWR _1263_/C sky130_fd_sc_hd__nand4_4
XFILLER_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2647_ _2457_/CLK _2647_/D VGND VGND VPWR VPWR _2647_/Q sky130_fd_sc_hd__dfxtp_4
X_1529_ _1528_/Y VGND VGND VPWR VPWR _1529_/Y sky130_fd_sc_hd__inv_2
X_2578_ _2606_/CLK _2578_/D VGND VGND VPWR VPWR _2578_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_19_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1880_ _1874_/A VGND VGND VPWR VPWR _1885_/A sky130_fd_sc_hd__buf_2
X_2501_ _2496_/CLK _1969_/X VGND VGND VPWR VPWR MACRO_WR_SELECT[2] sky130_fd_sc_hd__dfxtp_4
X_2363_ _2372_/CLK _2363_/D VGND VGND VPWR VPWR _2363_/Q sky130_fd_sc_hd__dfxtp_4
X_1314_ _1314_/A VGND VGND VPWR VPWR _2635_/D sky130_fd_sc_hd__inv_2
X_2432_ _2428_/CLK _2432_/D VGND VGND VPWR VPWR _1902_/A sky130_fd_sc_hd__dfxtp_4
X_2294_ _1420_/Y _2291_/X _2293_/Y VGND VGND VPWR VPWR _2410_/D sky130_fd_sc_hd__o21ai_4
X_1245_ _1245_/A VGND VGND VPWR VPWR _1246_/D sky130_fd_sc_hd__inv_2
XFILLER_32_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1863_ _1861_/Y _1862_/Y VGND VGND VPWR VPWR _2568_/D sky130_fd_sc_hd__nand2_4
X_1932_ _1932_/A _2529_/Q VGND VGND VPWR VPWR _2525_/D sky130_fd_sc_hd__and2_4
X_2415_ _2428_/CLK _2415_/D VGND VGND VPWR VPWR _2415_/Q sky130_fd_sc_hd__dfxtp_4
X_1794_ _1983_/B _2578_/Q _1793_/X VGND VGND VPWR VPWR _2586_/D sky130_fd_sc_hd__o21a_4
X_2346_ _2345_/Y S1_CLK_SELECT VGND VGND VPWR VPWR _2346_/Y sky130_fd_sc_hd__nand2_4
X_1228_ _1367_/A _1360_/A VGND VGND VPWR VPWR _1228_/Y sky130_fd_sc_hd__nand2_4
X_2277_ _1613_/A VGND VGND VPWR VPWR _2278_/A sky130_fd_sc_hd__inv_2
XFILLER_52_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2062_ _2053_/Y _2062_/B _2055_/X _1993_/C VGND VGND VPWR VPWR _2062_/X sky130_fd_sc_hd__and4_4
X_2131_ _2123_/A _2335_/A _2444_/Q VGND VGND VPWR VPWR _2131_/Y sky130_fd_sc_hd__nand3_4
X_2200_ _2420_/Q _1703_/A VGND VGND VPWR VPWR _2201_/C sky130_fd_sc_hd__nand2_4
XFILLER_19_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_6_0_addressalyzerBlock.SPI_CLK clkbuf_4_7_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2598_/CLK sky130_fd_sc_hd__clkbuf_1
X_1915_ _1254_/X VGND VGND VPWR VPWR _1918_/A sky130_fd_sc_hd__buf_2
X_1777_ _1777_/A _1777_/B _1777_/C _1777_/D VGND VGND VPWR VPWR _1783_/D sky130_fd_sc_hd__and4_4
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1846_ ID_toHost _2181_/A _1617_/Y _1845_/Y VGND VGND VPWR VPWR _1846_/X sky130_fd_sc_hd__a211o_4
X_2329_ _2102_/A _2322_/A _1683_/Y _2337_/A _2328_/X VGND VGND VPWR VPWR _2329_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_25_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1700_ _1645_/A _1308_/C _1612_/A VGND VGND VPWR VPWR _1700_/X sky130_fd_sc_hd__a21o_4
XPHY_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1631_ _1630_/X VGND VGND VPWR VPWR _1751_/A sky130_fd_sc_hd__buf_2
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1562_ _1562_/A VGND VGND VPWR VPWR _1562_/Y sky130_fd_sc_hd__inv_2
X_1493_ _1222_/X _1492_/Y VGND VGND VPWR VPWR _1493_/Y sky130_fd_sc_hd__nor2_4
X_2045_ _2029_/Y _2030_/X _2043_/C VGND VGND VPWR VPWR _2046_/C sky130_fd_sc_hd__a21oi_4
XFILLER_54_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2114_ _2104_/A ID_fromClient VGND VGND VPWR VPWR _2114_/X sky130_fd_sc_hd__and2_4
XFILLER_62_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1829_ _1829_/A VGND VGND VPWR VPWR _1829_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2594_ _2388_/CLK _2594_/D VGND VGND VPWR VPWR _2594_/Q sky130_fd_sc_hd__dfxtp_4
X_1614_ _1613_/Y VGND VGND VPWR VPWR _1614_/X sky130_fd_sc_hd__buf_2
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1545_ _1545_/A VGND VGND VPWR VPWR _1545_/X sky130_fd_sc_hd__buf_2
X_1476_ _1456_/X _1473_/X _1475_/Y VGND VGND VPWR VPWR _1476_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_54_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2028_ _2028_/A _2044_/B _2013_/D VGND VGND VPWR VPWR _2028_/X sky130_fd_sc_hd__and3_4
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1330_ _1318_/B _1335_/C _1242_/C _1329_/X VGND VGND VPWR VPWR _1330_/X sky130_fd_sc_hd__and4_4
X_1261_ _1256_/Y _1225_/X _1257_/X _1260_/Y VGND VGND VPWR VPWR _1261_/Y sky130_fd_sc_hd__nor4_4
X_1192_ _2593_/Q _1216_/B _1191_/X VGND VGND VPWR VPWR _1192_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_51_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2646_ _2570_/CLK _1215_/Y VGND VGND VPWR VPWR _1206_/A sky130_fd_sc_hd__dfxtp_4
X_2577_ _2581_/CLK _1817_/X VGND VGND VPWR VPWR _2577_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_59_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1528_ _1528_/A _1445_/A VGND VGND VPWR VPWR _1528_/Y sky130_fd_sc_hd__nor2_4
X_1459_ _1459_/A VGND VGND VPWR VPWR _2266_/A sky130_fd_sc_hd__buf_2
XFILLER_27_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2431_ _2428_/CLK _2431_/D VGND VGND VPWR VPWR _2431_/Q sky130_fd_sc_hd__dfxtp_4
X_2500_ _2519_/CLK _2500_/D VGND VGND VPWR VPWR MACRO_WR_SELECT[1] sky130_fd_sc_hd__dfxtp_4
XFILLER_56_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2362_ SCSN_fromHost VGND VGND VPWR VPWR SCSN_toClient sky130_fd_sc_hd__buf_2
X_1313_ _1308_/C _1308_/A _1312_/Y VGND VGND VPWR VPWR _1314_/A sky130_fd_sc_hd__o21ai_4
X_1244_ _1318_/A _1244_/B VGND VGND VPWR VPWR _1245_/A sky130_fd_sc_hd__nand2_4
XFILLER_2_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2293_ _2292_/X _2298_/B _2410_/Q VGND VGND VPWR VPWR _2293_/Y sky130_fd_sc_hd__nand3_4
XFILLER_64_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2629_ _2626_/CLK _2629_/D VGND VGND VPWR VPWR _2629_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_55_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1862_ _1762_/A _1862_/B VGND VGND VPWR VPWR _1862_/Y sky130_fd_sc_hd__nand2_4
X_1793_ _1788_/X _2266_/A _2326_/A VGND VGND VPWR VPWR _1793_/X sky130_fd_sc_hd__o21a_4
X_1931_ _1932_/A _1931_/B VGND VGND VPWR VPWR _2526_/D sky130_fd_sc_hd__and2_4
X_2414_ _2428_/CLK _2285_/Y VGND VGND VPWR VPWR _2151_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_6_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2345_ S1_CLK_IN VGND VGND VPWR VPWR _2345_/Y sky130_fd_sc_hd__inv_2
X_1227_ _1295_/A _1299_/A VGND VGND VPWR VPWR _1257_/A sky130_fd_sc_hd__nand2_4
X_2276_ _1581_/X VGND VGND VPWR VPWR _2276_/X sky130_fd_sc_hd__buf_2
XFILLER_20_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_11_0_addressalyzerBlock.SPI_CLK clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR _2390_/CLK sky130_fd_sc_hd__clkbuf_1
X_2061_ _2058_/X _2060_/Y _2062_/B _2055_/X _1993_/C VGND VGND VPWR VPWR _2061_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_34_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2130_ _1840_/B _2121_/X _2268_/A VGND VGND VPWR VPWR _2130_/Y sky130_fd_sc_hd__nand3_4
X_1914_ _1930_/A _1914_/B VGND VGND VPWR VPWR _2537_/D sky130_fd_sc_hd__nor2_4
XFILLER_19_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1776_ _1512_/Y _1764_/A _1494_/B _1771_/Y VGND VGND VPWR VPWR _1777_/D sky130_fd_sc_hd__a22oi_4
X_1845_ _2175_/B _1845_/B VGND VGND VPWR VPWR _1845_/Y sky130_fd_sc_hd__nor2_4
XFILLER_57_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2328_ _1187_/A _1680_/B _1781_/A VGND VGND VPWR VPWR _2328_/X sky130_fd_sc_hd__a21o_4
XFILLER_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2259_ _2243_/Y _2257_/Y _2258_/X _1911_/B _2248_/X VGND VGND VPWR VPWR _2428_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_63_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1630_ _2447_/Q VGND VGND VPWR VPWR _1630_/X sky130_fd_sc_hd__buf_2
XPHY_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1561_ _1428_/C _1669_/B VGND VGND VPWR VPWR _1562_/A sky130_fd_sc_hd__nand2_4
X_1492_ _2609_/Q _1489_/X _1491_/Y _1449_/B VGND VGND VPWR VPWR _1492_/Y sky130_fd_sc_hd__a22oi_4
X_2044_ _2044_/A _2044_/B _2044_/C VGND VGND VPWR VPWR _2044_/X sky130_fd_sc_hd__and3_4
X_2113_ _2104_/A _2113_/B VGND VGND VPWR VPWR _2113_/X sky130_fd_sc_hd__and2_4
X_1759_ _1656_/X _1397_/A _2166_/A VGND VGND VPWR VPWR _1759_/Y sky130_fd_sc_hd__a21oi_4
X_1828_ _1808_/Y _2455_/Q _1827_/X VGND VGND VPWR VPWR _2572_/D sky130_fd_sc_hd__o21a_4
XFILLER_53_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2593_ _2590_/CLK _2593_/D VGND VGND VPWR VPWR _2593_/Q sky130_fd_sc_hd__dfxtp_4
X_1613_ _1613_/A _1651_/A _1667_/C _1667_/D VGND VGND VPWR VPWR _1613_/Y sky130_fd_sc_hd__nand4_4
X_1544_ _1537_/X _1548_/D _1435_/Y VGND VGND VPWR VPWR _1544_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_39_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1475_ _1456_/X _1440_/B _1473_/B _1438_/A _2340_/C VGND VGND VPWR VPWR _1475_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_54_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2027_ _1270_/A VGND VGND VPWR VPWR _2044_/B sky130_fd_sc_hd__buf_2
XFILLER_50_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1191_ _2096_/A VGND VGND VPWR VPWR _1191_/X sky130_fd_sc_hd__buf_2
XFILLER_39_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1260_ _1258_/Y _1243_/X _1246_/D _1292_/C VGND VGND VPWR VPWR _1260_/Y sky130_fd_sc_hd__nand4_4
XFILLER_36_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_1_0_m1_clk_local clkbuf_3_1_0_m1_clk_local/A VGND VGND VPWR VPWR clkbuf_4_3_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2645_ _2570_/CLK _2645_/D VGND VGND VPWR VPWR _2645_/Q sky130_fd_sc_hd__dfxtp_4
X_1527_ _1526_/Y VGND VGND VPWR VPWR _1527_/Y sky130_fd_sc_hd__inv_2
X_2576_ _2581_/CLK _2576_/D VGND VGND VPWR VPWR _2576_/Q sky130_fd_sc_hd__dfxtp_4
X_1389_ _1379_/X _1385_/D _2621_/Q VGND VGND VPWR VPWR _1390_/C sky130_fd_sc_hd__a21oi_4
XFILLER_27_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1458_ _1438_/B _1457_/X _1452_/Y VGND VGND VPWR VPWR _1458_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_50_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2361_ SCLK_fromHost VGND VGND VPWR VPWR SCLK_toClient sky130_fd_sc_hd__buf_2
X_2430_ _2428_/CLK _2254_/Y VGND VGND VPWR VPWR _2154_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_64_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1243_ _1243_/A VGND VGND VPWR VPWR _1243_/X sky130_fd_sc_hd__buf_2
X_1312_ _1308_/C _1318_/B _1316_/D _1246_/D _1274_/X VGND VGND VPWR VPWR _1312_/Y
+ sky130_fd_sc_hd__a41oi_4
X_2292_ _2290_/Y VGND VGND VPWR VPWR _2292_/X sky130_fd_sc_hd__buf_2
XFILLER_2_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2628_ _2626_/CLK _2628_/D VGND VGND VPWR VPWR _2628_/Q sky130_fd_sc_hd__dfxtp_4
X_2559_ _2554_/CLK _2559_/D VGND VGND VPWR VPWR _2559_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_55_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1930_ _1930_/A _1929_/Y VGND VGND VPWR VPWR _2527_/D sky130_fd_sc_hd__nor2_4
X_1861_ _1859_/Y _1673_/Y _1860_/X VGND VGND VPWR VPWR _1861_/Y sky130_fd_sc_hd__nand3_4
X_1792_ _1983_/B _2579_/Q _1791_/X VGND VGND VPWR VPWR _1792_/X sky130_fd_sc_hd__o21a_4
XFILLER_14_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2413_ _2445_/CLK _2413_/D VGND VGND VPWR VPWR _2174_/B sky130_fd_sc_hd__dfxtp_4
X_2344_ _2342_/Y M1_CLK_SELECT _2343_/Y VGND VGND VPWR VPWR m1_clk_local sky130_fd_sc_hd__a21oi_4
XFILLER_37_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1226_ _2636_/Q _2635_/Q VGND VGND VPWR VPWR _1226_/Y sky130_fd_sc_hd__nand2_4
XFILLER_16_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2275_ _2144_/Y _1649_/B _2270_/X _1948_/Y _2263_/X VGND VGND VPWR VPWR _2419_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_52_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2060_ _2060_/A _2060_/B VGND VGND VPWR VPWR _2060_/Y sky130_fd_sc_hd__nor2_4
XFILLER_34_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1913_ _1913_/A VGND VGND VPWR VPWR _1914_/B sky130_fd_sc_hd__inv_2
X_1844_ _1844_/A VGND VGND VPWR VPWR _1845_/B sky130_fd_sc_hd__inv_2
X_1775_ _1499_/Y _1773_/A _1456_/X _1766_/B VGND VGND VPWR VPWR _1777_/C sky130_fd_sc_hd__a22oi_4
X_2327_ _1222_/A _1218_/B _1680_/B _1683_/Y _2326_/Y VGND VGND VPWR VPWR _2387_/D
+ sky130_fd_sc_hd__o41ai_4
X_2258_ _2246_/Y VGND VGND VPWR VPWR _2258_/X sky130_fd_sc_hd__buf_2
X_1209_ _1207_/Y _1187_/X _1208_/Y VGND VGND VPWR VPWR _2647_/D sky130_fd_sc_hd__a21oi_4
X_2189_ _2146_/A THREAD_COUNT[2] VGND VGND VPWR VPWR _2189_/Y sky130_fd_sc_hd__nand2_4
XFILLER_25_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1560_ _1428_/D VGND VGND VPWR VPWR _1669_/B sky130_fd_sc_hd__buf_2
X_2112_ _1870_/X _2103_/Y VGND VGND VPWR VPWR _2112_/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1491_ _2609_/Q _1451_/X _1487_/Y _1490_/Y _1445_/D VGND VGND VPWR VPWR _1491_/Y
+ sky130_fd_sc_hd__o32ai_4
X_2043_ _2030_/X _2029_/Y _2043_/C _2043_/D VGND VGND VPWR VPWR _2044_/C sky130_fd_sc_hd__nand4_4
XFILLER_54_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1827_ _2572_/Q _2461_/Q _2257_/A VGND VGND VPWR VPWR _1827_/X sky130_fd_sc_hd__o21a_4
X_1758_ _1742_/Y _1756_/Y _1757_/Y VGND VGND VPWR VPWR _1758_/Y sky130_fd_sc_hd__o21ai_4
X_1689_ _1689_/A VGND VGND VPWR VPWR _1689_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_2_0_addressalyzerBlock.SPI_CLK clkbuf_2_3_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1612_ _1612_/A VGND VGND VPWR VPWR _1612_/X sky130_fd_sc_hd__buf_2
X_2592_ _2590_/CLK _2592_/D VGND VGND VPWR VPWR _1662_/A sky130_fd_sc_hd__dfxtp_4
X_1474_ _1451_/X VGND VGND VPWR VPWR _2340_/C sky130_fd_sc_hd__buf_2
XFILLER_5_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1543_ _1539_/Y _1540_/Y _1542_/X VGND VGND VPWR VPWR _2603_/D sky130_fd_sc_hd__a21oi_4
XFILLER_39_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2026_ _2047_/A _2017_/B _2017_/C _2017_/D _2488_/Q VGND VGND VPWR VPWR _2028_/A
+ sky130_fd_sc_hd__a41o_4
XFILLER_2_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1190_ _1189_/Y VGND VGND VPWR VPWR _2096_/A sky130_fd_sc_hd__buf_2
XFILLER_39_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2644_ _2638_/CLK _1264_/Y VGND VGND VPWR VPWR _1251_/A sky130_fd_sc_hd__dfxtp_4
X_1526_ _1443_/A _2390_/Q VGND VGND VPWR VPWR _1526_/Y sky130_fd_sc_hd__nor2_4
X_2575_ _2581_/CLK _2575_/D VGND VGND VPWR VPWR _2575_/Q sky130_fd_sc_hd__dfxtp_4
X_1457_ _1440_/B _1456_/X _1438_/D _1438_/A VGND VGND VPWR VPWR _1457_/X sky130_fd_sc_hd__and4_4
X_1388_ _1283_/X VGND VGND VPWR VPWR _1395_/A sky130_fd_sc_hd__buf_2
X_2009_ _2008_/Y _1984_/A _1999_/A _2011_/A _2492_/Q VGND VGND VPWR VPWR _2009_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_18_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1311_ _1243_/X VGND VGND VPWR VPWR _1316_/D sky130_fd_sc_hd__buf_2
X_2360_ MOSI_fromHost VGND VGND VPWR VPWR MOSI_toClient sky130_fd_sc_hd__buf_2
X_2291_ _2290_/Y VGND VGND VPWR VPWR _2291_/X sky130_fd_sc_hd__buf_2
X_1242_ _1335_/A _1242_/B _1242_/C _2629_/Q VGND VGND VPWR VPWR _1243_/A sky130_fd_sc_hd__and4_4
XFILLER_2_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2627_ _2626_/CLK _2627_/D VGND VGND VPWR VPWR _1349_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_9_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2489_ _2470_/CLK _2025_/Y VGND VGND VPWR VPWR _1984_/A sky130_fd_sc_hd__dfxtp_4
X_2558_ _2562_/CLK _2558_/D VGND VGND VPWR VPWR _2558_/Q sky130_fd_sc_hd__dfxtp_4
X_1509_ _1508_/X _1448_/A _1505_/A VGND VGND VPWR VPWR _1509_/X sky130_fd_sc_hd__a21o_4
XFILLER_62_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1860_ _2618_/Q _1860_/B _1661_/C _1661_/D VGND VGND VPWR VPWR _1860_/X sky130_fd_sc_hd__or4_4
XFILLER_14_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1791_ _1788_/X _1420_/A _2326_/A VGND VGND VPWR VPWR _1791_/X sky130_fd_sc_hd__o21a_4
X_2343_ PLL_INPUT M1_CLK_SELECT VGND VGND VPWR VPWR _2343_/Y sky130_fd_sc_hd__nor2_4
X_2412_ _2410_/CLK _2412_/D VGND VGND VPWR VPWR _1927_/A sky130_fd_sc_hd__dfxtp_4
X_2274_ _2142_/Y _1649_/B _2270_/X _1947_/B _2263_/X VGND VGND VPWR VPWR _2420_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_52_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1225_ _1225_/A VGND VGND VPWR VPWR _1225_/X sky130_fd_sc_hd__buf_2
X_1989_ _2478_/Q VGND VGND VPWR VPWR _1992_/B sky130_fd_sc_hd__inv_2
XFILLER_57_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1843_ _1534_/X _2556_/Q _1614_/X VGND VGND VPWR VPWR _1843_/Y sky130_fd_sc_hd__o21ai_4
X_1912_ _1339_/X VGND VGND VPWR VPWR _1930_/A sky130_fd_sc_hd__buf_2
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1774_ _1751_/B _2609_/Q _1487_/A _2158_/B VGND VGND VPWR VPWR _1777_/B sky130_fd_sc_hd__a22oi_4
X_1208_ _2437_/Q _1187_/A _1191_/X VGND VGND VPWR VPWR _1208_/Y sky130_fd_sc_hd__o21ai_4
X_2326_ _2326_/A _1423_/Y _1185_/A _1577_/X VGND VGND VPWR VPWR _2326_/Y sky130_fd_sc_hd__nand4_4
X_2257_ _2257_/A _1698_/A _1514_/X VGND VGND VPWR VPWR _2257_/Y sky130_fd_sc_hd__nand3_4
XFILLER_40_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2188_ _2185_/Y _2186_/X _2187_/X VGND VGND VPWR VPWR _2188_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1490_ _1490_/A VGND VGND VPWR VPWR _1490_/Y sky130_fd_sc_hd__inv_2
X_2042_ _2041_/Y _1985_/A _2030_/X _2017_/B _2043_/D VGND VGND VPWR VPWR _2044_/A
+ sky130_fd_sc_hd__a41o_4
X_2111_ _1870_/X _2098_/Y VGND VGND VPWR VPWR _2111_/Y sky130_fd_sc_hd__nand2_4
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1826_ _2572_/Q _1808_/Y _1825_/X VGND VGND VPWR VPWR _2573_/D sky130_fd_sc_hd__o21a_4
X_1757_ _1612_/A _1360_/A _1656_/A VGND VGND VPWR VPWR _1757_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1688_ _1731_/B _1566_/X _2340_/B VGND VGND VPWR VPWR _1688_/Y sky130_fd_sc_hd__nor3_4
XFILLER_57_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2309_ _2144_/Y _2292_/X _2308_/Y VGND VGND VPWR VPWR _2403_/D sky130_fd_sc_hd__o21ai_4
XFILLER_48_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1611_ _1611_/A VGND VGND VPWR VPWR _1612_/A sky130_fd_sc_hd__buf_2
XFILLER_12_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1542_ _1549_/A _1466_/Y _1500_/X VGND VGND VPWR VPWR _1542_/X sky130_fd_sc_hd__a21o_4
X_2591_ _2581_/CLK _2591_/D VGND VGND VPWR VPWR _2591_/Q sky130_fd_sc_hd__dfxtp_4
X_1473_ _1469_/Y _1473_/B _1473_/C _1438_/A VGND VGND VPWR VPWR _1473_/X sky130_fd_sc_hd__and4_4
X_2025_ _2002_/X _2013_/D _2024_/Y VGND VGND VPWR VPWR _2025_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_54_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1809_ _1808_/Y VGND VGND VPWR VPWR _1809_/X sky130_fd_sc_hd__buf_2
XFILLER_18_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2643_ _2638_/CLK _2643_/D VGND VGND VPWR VPWR _1262_/C sky130_fd_sc_hd__dfxtp_4
X_2574_ _2581_/CLK _2574_/D VGND VGND VPWR VPWR _2574_/Q sky130_fd_sc_hd__dfxtp_4
X_1387_ _1387_/A VGND VGND VPWR VPWR _2622_/D sky130_fd_sc_hd__inv_2
X_1456_ _1438_/C VGND VGND VPWR VPWR _1456_/X sky130_fd_sc_hd__buf_2
X_1525_ _1473_/C _1469_/Y _1524_/Y VGND VGND VPWR VPWR _1525_/Y sky130_fd_sc_hd__o21ai_4
X_2008_ _2008_/A VGND VGND VPWR VPWR _2008_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1241_ _1240_/Y VGND VGND VPWR VPWR _1241_/Y sky130_fd_sc_hd__inv_2
X_1310_ _1309_/Y VGND VGND VPWR VPWR _2636_/D sky130_fd_sc_hd__inv_2
X_2290_ _2290_/A VGND VGND VPWR VPWR _2290_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2626_ _2626_/CLK _2626_/D VGND VGND VPWR VPWR _1367_/A sky130_fd_sc_hd__dfxtp_4
X_2557_ _2557_/CLK _2557_/D VGND VGND VPWR VPWR _1701_/B sky130_fd_sc_hd__dfxtp_4
X_2488_ _2470_/CLK _2028_/X VGND VGND VPWR VPWR _2488_/Q sky130_fd_sc_hd__dfxtp_4
X_1439_ _1439_/A VGND VGND VPWR VPWR _1440_/D sky130_fd_sc_hd__buf_2
X_1508_ _1469_/Y _1505_/C _1438_/D _1473_/C _1451_/X VGND VGND VPWR VPWR _1508_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_55_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1790_ _1838_/A VGND VGND VPWR VPWR _2326_/A sky130_fd_sc_hd__buf_2
X_2411_ _2445_/CLK _2411_/D VGND VGND VPWR VPWR _2411_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1224_ _1224_/A VGND VGND VPWR VPWR _1225_/A sky130_fd_sc_hd__inv_2
X_2342_ M1_CLK_IN VGND VGND VPWR VPWR _2342_/Y sky130_fd_sc_hd__inv_2
X_2273_ _1503_/Y _1649_/B _2270_/X _1945_/B _2263_/X VGND VGND VPWR VPWR _2421_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_25_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1988_ _2477_/Q VGND VGND VPWR VPWR _1992_/A sky130_fd_sc_hd__inv_2
Xclkbuf_2_3_0_m1_clk_local clkbuf_2_3_0_m1_clk_local/A VGND VGND VPWR VPWR clkbuf_3_7_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
X_2609_ _2388_/CLK _1493_/Y VGND VGND VPWR VPWR _2609_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_28_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_2_0_addressalyzerBlock.SPI_CLK clkbuf_2_1_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR clkbuf_4_5_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
X_1842_ _1179_/X _1735_/D _1841_/Y VGND VGND VPWR VPWR _2569_/D sky130_fd_sc_hd__o21a_4
X_1773_ _1773_/A VGND VGND VPWR VPWR _2158_/B sky130_fd_sc_hd__inv_2
XFILLER_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1911_ _1901_/X _1911_/B VGND VGND VPWR VPWR _1911_/Y sky130_fd_sc_hd__nor2_4
XFILLER_6_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1207_ _2647_/Q _1179_/A _1206_/X VGND VGND VPWR VPWR _1207_/Y sky130_fd_sc_hd__o21ai_4
X_2187_ _1611_/A _1373_/B _1656_/A VGND VGND VPWR VPWR _2187_/X sky130_fd_sc_hd__a21o_4
X_2325_ _2324_/X _1688_/Y _1870_/X VGND VGND VPWR VPWR _2325_/X sky130_fd_sc_hd__o21a_4
X_2256_ _2244_/X _2255_/Y _2247_/X _1908_/Y _2249_/X VGND VGND VPWR VPWR _2429_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_40_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2041_ _2040_/X VGND VGND VPWR VPWR _2041_/Y sky130_fd_sc_hd__inv_2
X_2110_ _2108_/A MOSI_fromHost VGND VGND VPWR VPWR _2454_/D sky130_fd_sc_hd__and2_4
XFILLER_47_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1756_ _1753_/X _1754_/X _1755_/Y VGND VGND VPWR VPWR _1756_/Y sky130_fd_sc_hd__a21oi_4
X_1825_ _2573_/Q _2461_/Q _2257_/A VGND VGND VPWR VPWR _1825_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_4_6_0_m1_clk_local clkbuf_4_7_0_m1_clk_local/A VGND VGND VPWR VPWR _2626_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_1687_ _1728_/C VGND VGND VPWR VPWR _2340_/B sky130_fd_sc_hd__inv_2
X_2308_ _2290_/Y _1602_/C _2089_/A VGND VGND VPWR VPWR _2308_/Y sky130_fd_sc_hd__nand3_4
XFILLER_45_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2239_ _2239_/A VGND VGND VPWR VPWR _2239_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2590_ _2590_/CLK _2590_/D VGND VGND VPWR VPWR _1762_/B sky130_fd_sc_hd__dfxtp_4
X_1610_ _1609_/X VGND VGND VPWR VPWR _1611_/A sky130_fd_sc_hd__buf_2
XFILLER_8_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1541_ _1530_/Y VGND VGND VPWR VPWR _1549_/A sky130_fd_sc_hd__buf_2
XFILLER_5_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1472_ _1471_/X VGND VGND VPWR VPWR _1473_/C sky130_fd_sc_hd__buf_2
X_2024_ _2002_/X _2013_/D _1346_/X VGND VGND VPWR VPWR _2024_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_54_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1739_ _1739_/A _1739_/B VGND VGND VPWR VPWR _1739_/Y sky130_fd_sc_hd__nor2_4
X_1808_ _2461_/Q VGND VGND VPWR VPWR _1808_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2642_ _2641_/CLK _1279_/Y VGND VGND VPWR VPWR _1277_/A sky130_fd_sc_hd__dfxtp_4
X_2573_ _2581_/CLK _2573_/D VGND VGND VPWR VPWR _2573_/Q sky130_fd_sc_hd__dfxtp_4
X_1524_ _1473_/C _1429_/Y _1466_/A _2602_/Q _2340_/C VGND VGND VPWR VPWR _1524_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1386_ _1384_/X _1385_/Y VGND VGND VPWR VPWR _1387_/A sky130_fd_sc_hd__nand2_4
X_1455_ _1449_/Y _1453_/Y _1454_/X VGND VGND VPWR VPWR _1455_/Y sky130_fd_sc_hd__a21oi_4
X_2007_ _2006_/Y VGND VGND VPWR VPWR _2493_/D sky130_fd_sc_hd__inv_2
XFILLER_35_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1240_ _2628_/Q _1349_/A VGND VGND VPWR VPWR _1240_/Y sky130_fd_sc_hd__nand2_4
XFILLER_2_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2625_ _2470_/CLK _2625_/D VGND VGND VPWR VPWR _1360_/A sky130_fd_sc_hd__dfxtp_4
X_2487_ _2470_/CLK _2034_/X VGND VGND VPWR VPWR _2017_/C sky130_fd_sc_hd__dfxtp_4
X_2556_ _2562_/CLK _2556_/D VGND VGND VPWR VPWR _2556_/Q sky130_fd_sc_hd__dfxtp_4
X_1507_ _1506_/Y _1449_/B VGND VGND VPWR VPWR _1507_/Y sky130_fd_sc_hd__nand2_4
XFILLER_55_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1369_ _1368_/Y VGND VGND VPWR VPWR _2626_/D sky130_fd_sc_hd__inv_2
X_1438_ _1438_/A _1438_/B _1438_/C _1438_/D VGND VGND VPWR VPWR _1439_/A sky130_fd_sc_hd__and4_4
XFILLER_55_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2341_ EXT_RESET_N_fromHost VGND VGND VPWR VPWR _2341_/Y sky130_fd_sc_hd__inv_2
X_2410_ _2410_/CLK _2410_/D VGND VGND VPWR VPWR _2410_/Q sky130_fd_sc_hd__dfxtp_4
X_1223_ _1216_/Y _1218_/Y _1222_/X VGND VGND VPWR VPWR _2645_/D sky130_fd_sc_hd__a21oi_4
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2272_ _2136_/Y _2262_/X _2270_/X _1942_/B _2264_/X VGND VGND VPWR VPWR _2422_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_52_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1987_ _1987_/A VGND VGND VPWR VPWR _1994_/C sky130_fd_sc_hd__inv_2
XFILLER_20_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2539_ _2519_/CLK _2539_/D VGND VGND VPWR VPWR _2539_/Q sky130_fd_sc_hd__dfxtp_4
X_2608_ _2606_/CLK _1502_/Y VGND VGND VPWR VPWR _1436_/B sky130_fd_sc_hd__dfxtp_4
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1910_ _2428_/Q VGND VGND VPWR VPWR _1911_/B sky130_fd_sc_hd__inv_2
X_1841_ _1841_/A VGND VGND VPWR VPWR _1841_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1772_ _2609_/Q _1751_/B _1436_/C _1771_/Y VGND VGND VPWR VPWR _1777_/A sky130_fd_sc_hd__o22a_4
X_2324_ _1731_/B _1566_/X _1689_/A VGND VGND VPWR VPWR _2324_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_4_14_0_m1_clk_local clkbuf_3_7_0_m1_clk_local/X VGND VGND VPWR VPWR _2498_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_1206_ _1206_/A _1180_/Y VGND VGND VPWR VPWR _1206_/X sky130_fd_sc_hd__or2_4
X_2186_ _1335_/C _1646_/A _1741_/Y VGND VGND VPWR VPWR _2186_/X sky130_fd_sc_hd__o21a_4
X_2255_ _2257_/A _1698_/A _1503_/A VGND VGND VPWR VPWR _2255_/Y sky130_fd_sc_hd__nand3_4
XFILLER_43_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2040_ _1994_/D VGND VGND VPWR VPWR _2040_/X sky130_fd_sc_hd__buf_2
X_1755_ _1280_/Y _1614_/X _1646_/X VGND VGND VPWR VPWR _1755_/Y sky130_fd_sc_hd__o21ai_4
X_1686_ _1678_/Y _1682_/Y _1685_/X VGND VGND VPWR VPWR _1686_/Y sky130_fd_sc_hd__a21oi_4
X_1824_ _1838_/A VGND VGND VPWR VPWR _2257_/A sky130_fd_sc_hd__buf_2
XFILLER_57_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2307_ _2142_/Y _2292_/X _2306_/Y VGND VGND VPWR VPWR _2307_/Y sky130_fd_sc_hd__o21ai_4
X_2238_ _1609_/B _1189_/Y _1583_/X _1696_/A VGND VGND VPWR VPWR _2239_/A sky130_fd_sc_hd__and4_4
XFILLER_54_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2169_ _2546_/Q _1739_/B _2167_/Y _2168_/Y VGND VGND VPWR VPWR _2169_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_5_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1540_ _2266_/A _1527_/Y _1556_/A VGND VGND VPWR VPWR _1540_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_5_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1471_ _2604_/Q VGND VGND VPWR VPWR _1471_/X sky130_fd_sc_hd__buf_2
X_2023_ _2022_/Y VGND VGND VPWR VPWR _2490_/D sky130_fd_sc_hd__inv_2
XFILLER_35_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1807_ _1786_/Y _2572_/Q _1806_/X VGND VGND VPWR VPWR _1807_/X sky130_fd_sc_hd__o21a_4
X_1738_ _1831_/A _1738_/B VGND VGND VPWR VPWR _2591_/D sky130_fd_sc_hd__nor2_4
X_1669_ _1579_/X _1669_/B _1590_/B VGND VGND VPWR VPWR _1669_/Y sky130_fd_sc_hd__nor3_4
XFILLER_45_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1454_ _1222_/A VGND VGND VPWR VPWR _1454_/X sky130_fd_sc_hd__buf_2
X_2641_ _2641_/CLK _1282_/X VGND VGND VPWR VPWR _2641_/Q sky130_fd_sc_hd__dfxtp_4
X_2572_ _2581_/CLK _2572_/D VGND VGND VPWR VPWR _2572_/Q sky130_fd_sc_hd__dfxtp_4
X_1523_ _1519_/Y _1521_/Y _1522_/Y VGND VGND VPWR VPWR _2605_/D sky130_fd_sc_hd__a21oi_4
X_1385_ _1385_/A _1379_/A _2621_/Q _1385_/D VGND VGND VPWR VPWR _1385_/Y sky130_fd_sc_hd__nand4_4
X_2006_ _2001_/Y _2006_/B _2005_/Y VGND VGND VPWR VPWR _2006_/Y sky130_fd_sc_hd__nand3_4
XFILLER_23_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2624_ _2370_/CLK _2624_/D VGND VGND VPWR VPWR _1236_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_9_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2486_ _2483_/CLK _2486_/D VGND VGND VPWR VPWR _2037_/D sky130_fd_sc_hd__dfxtp_4
X_2555_ _2562_/CLK _1885_/X VGND VGND VPWR VPWR _2555_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_4_2_0_addressalyzerBlock.SPI_CLK clkbuf_4_3_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2445_/CLK sky130_fd_sc_hd__clkbuf_1
X_1437_ _1483_/B VGND VGND VPWR VPWR _1438_/D sky130_fd_sc_hd__buf_2
X_1506_ _1503_/Y _1445_/D _1505_/Y VGND VGND VPWR VPWR _1506_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_55_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1368_ _1362_/X _1367_/Y VGND VGND VPWR VPWR _1368_/Y sky130_fd_sc_hd__nand2_4
X_1299_ _1299_/A VGND VGND VPWR VPWR _1300_/B sky130_fd_sc_hd__inv_2
XFILLER_23_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_7_0_addressalyzerBlock.SPI_CLK clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2340_ _2102_/A _2340_/B _2340_/C VGND VGND VPWR VPWR _2393_/D sky130_fd_sc_hd__nor3_4
X_2271_ _1490_/Y _2262_/X _2270_/X _1746_/Y _2264_/X VGND VGND VPWR VPWR _2271_/Y
+ sky130_fd_sc_hd__o32ai_4
X_1222_ _1222_/A VGND VGND VPWR VPWR _1222_/X sky130_fd_sc_hd__buf_2
XFILLER_37_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1986_ _2030_/A VGND VGND VPWR VPWR _1986_/Y sky130_fd_sc_hd__inv_2
X_2607_ _2606_/CLK _2607_/D VGND VGND VPWR VPWR _1436_/C sky130_fd_sc_hd__dfxtp_4
X_2469_ _2641_/CLK _2090_/Y VGND VGND VPWR VPWR _2088_/B sky130_fd_sc_hd__dfxtp_4
X_2538_ _2519_/CLK _1911_/Y VGND VGND VPWR VPWR _2538_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1840_ _1834_/A _1840_/B _1840_/C VGND VGND VPWR VPWR _1841_/A sky130_fd_sc_hd__nand3_4
XFILLER_42_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1771_ _2397_/Q VGND VGND VPWR VPWR _1771_/Y sky130_fd_sc_hd__inv_2
X_2323_ _2322_/Y _1697_/Y _1781_/X VGND VGND VPWR VPWR _2392_/D sky130_fd_sc_hd__a21oi_4
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2254_ _2244_/X _2253_/Y _2247_/X _1906_/Y _2249_/X VGND VGND VPWR VPWR _2254_/Y
+ sky130_fd_sc_hd__o32ai_4
X_1205_ _1203_/Y _1187_/X _1204_/Y VGND VGND VPWR VPWR _1205_/Y sky130_fd_sc_hd__a21oi_4
X_2185_ _2173_/Y _2183_/Y _2184_/Y VGND VGND VPWR VPWR _2185_/Y sky130_fd_sc_hd__o21ai_4
X_1969_ _1969_/A _2505_/Q VGND VGND VPWR VPWR _1969_/X sky130_fd_sc_hd__and2_4
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1823_ _2573_/Q _1808_/Y _1822_/X VGND VGND VPWR VPWR _2574_/D sky130_fd_sc_hd__o21a_4
X_1754_ _1534_/X _2555_/Q _1614_/X VGND VGND VPWR VPWR _1754_/X sky130_fd_sc_hd__o21a_4
X_1685_ _1681_/X _1684_/Y _1500_/X VGND VGND VPWR VPWR _1685_/X sky130_fd_sc_hd__a21o_4
X_2237_ _2235_/Y _1662_/A _2236_/Y VGND VGND VPWR VPWR _2237_/Y sky130_fd_sc_hd__a21oi_4
X_2306_ _2304_/A _1602_/C _2404_/Q VGND VGND VPWR VPWR _2306_/Y sky130_fd_sc_hd__nand3_4
XFILLER_53_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2168_ _1673_/C _1672_/A VGND VGND VPWR VPWR _2168_/Y sky130_fd_sc_hd__nor2_4
XFILLER_38_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2099_ _2104_/A _2098_/Y _2099_/C VGND VGND VPWR VPWR _2099_/X sky130_fd_sc_hd__and3_4
XFILLER_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1470_ _1438_/D VGND VGND VPWR VPWR _1473_/B sky130_fd_sc_hd__buf_2
XFILLER_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2022_ _2022_/A _2006_/B _2021_/Y VGND VGND VPWR VPWR _2022_/Y sky130_fd_sc_hd__nand3_4
X_1806_ _2591_/Q _1520_/X _1799_/X VGND VGND VPWR VPWR _1806_/X sky130_fd_sc_hd__o21a_4
X_1737_ _1831_/B VGND VGND VPWR VPWR _1738_/B sky130_fd_sc_hd__inv_2
X_1668_ _1667_/X VGND VGND VPWR VPWR _1673_/C sky130_fd_sc_hd__buf_2
X_1599_ _1600_/B _1488_/X _1598_/X _1530_/Y VGND VGND VPWR VPWR _1602_/A sky130_fd_sc_hd__a211o_4
XFILLER_45_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_2_0_m1_clk_local clkbuf_4_3_0_m1_clk_local/A VGND VGND VPWR VPWR _2528_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2640_ _2638_/CLK _2640_/D VGND VGND VPWR VPWR _1277_/D sky130_fd_sc_hd__dfxtp_4
X_2571_ _2457_/CLK _2571_/D VGND VGND VPWR VPWR _1829_/A sky130_fd_sc_hd__dfxtp_4
X_1522_ _1473_/B _1448_/A _1213_/X VGND VGND VPWR VPWR _1522_/Y sky130_fd_sc_hd__o21ai_4
X_1453_ _1450_/X _1452_/Y _2335_/B VGND VGND VPWR VPWR _1453_/Y sky130_fd_sc_hd__o21ai_4
X_2005_ _2011_/A _2020_/A _2492_/Q CLK_LED VGND VGND VPWR VPWR _2005_/Y sky130_fd_sc_hd__nand4_4
XFILLER_55_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1384_ _1385_/A _1390_/B _1374_/X VGND VGND VPWR VPWR _1384_/X sky130_fd_sc_hd__o21a_4
XFILLER_35_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2554_ _2554_/CLK _1887_/X VGND VGND VPWR VPWR _2554_/Q sky130_fd_sc_hd__dfxtp_4
X_2623_ _2367_/CLK _2623_/D VGND VGND VPWR VPWR _2623_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_13_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2485_ _2483_/CLK _2044_/X VGND VGND VPWR VPWR _2043_/D sky130_fd_sc_hd__dfxtp_4
X_1367_ _1367_/A _1366_/X _1360_/A _1238_/D VGND VGND VPWR VPWR _1367_/Y sky130_fd_sc_hd__nand4_4
X_1436_ _2609_/Q _1436_/B _1436_/C _1486_/A VGND VGND VPWR VPWR _1438_/A sky130_fd_sc_hd__and4_4
X_1505_ _1505_/A _1505_/B _1505_/C _1435_/Y VGND VGND VPWR VPWR _1505_/Y sky130_fd_sc_hd__nand4_4
X_1298_ _1270_/A VGND VGND VPWR VPWR _2006_/B sky130_fd_sc_hd__buf_2
XFILLER_11_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1221_ _1221_/A VGND VGND VPWR VPWR _1222_/A sky130_fd_sc_hd__buf_2
X_2270_ _2246_/Y VGND VGND VPWR VPWR _2270_/X sky130_fd_sc_hd__buf_2
XFILLER_37_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1985_ _1985_/A VGND VGND VPWR VPWR _1985_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2537_ _2506_/CLK _2537_/D VGND VGND VPWR VPWR _2537_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2606_ _2606_/CLK _2606_/D VGND VGND VPWR VPWR _1486_/A sky130_fd_sc_hd__dfxtp_4
X_1419_ _1419_/A _2010_/B _1419_/C VGND VGND VPWR VPWR _1419_/X sky130_fd_sc_hd__and3_4
X_2468_ _2570_/CLK _2092_/Y VGND VGND VPWR VPWR _2468_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_28_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2399_ _2606_/CLK _2399_/D VGND VGND VPWR VPWR _1750_/A sky130_fd_sc_hd__dfxtp_4
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1770_ _1769_/X VGND VGND VPWR VPWR _1783_/B sky130_fd_sc_hd__inv_2
XFILLER_6_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1204_ _2170_/B _1216_/B _1191_/X VGND VGND VPWR VPWR _1204_/Y sky130_fd_sc_hd__o21ai_4
X_2322_ _2322_/A _2392_/Q VGND VGND VPWR VPWR _2322_/Y sky130_fd_sc_hd__nand2_4
X_2184_ _1225_/A _2148_/X _1651_/X _1649_/Y VGND VGND VPWR VPWR _2184_/Y sky130_fd_sc_hd__a2bb2oi_4
X_2253_ _2257_/A _1698_/A _2253_/C VGND VGND VPWR VPWR _2253_/Y sky130_fd_sc_hd__nand3_4
XFILLER_18_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1899_ _1900_/A _1899_/B VGND VGND VPWR VPWR _1899_/X sky130_fd_sc_hd__and2_4
X_1968_ _1969_/A _1968_/B VGND VGND VPWR VPWR _2502_/D sky130_fd_sc_hd__and2_4
XFILLER_16_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1822_ _2574_/Q _2461_/Q _1813_/X VGND VGND VPWR VPWR _1822_/X sky130_fd_sc_hd__o21a_4
X_1753_ _1749_/X _1752_/X _1471_/X VGND VGND VPWR VPWR _1753_/X sky130_fd_sc_hd__a21o_4
X_1684_ _1575_/Y _1683_/Y _1444_/Y VGND VGND VPWR VPWR _1684_/Y sky130_fd_sc_hd__nand3_4
X_2167_ _2147_/Y _2165_/Y _2166_/Y VGND VGND VPWR VPWR _2167_/Y sky130_fd_sc_hd__o21ai_4
X_2236_ _1662_/A _1218_/A VGND VGND VPWR VPWR _2236_/Y sky130_fd_sc_hd__nor2_4
XFILLER_38_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2305_ _1503_/Y _2292_/X _2304_/Y VGND VGND VPWR VPWR _2305_/Y sky130_fd_sc_hd__o21ai_4
X_2098_ _2452_/Q VGND VGND VPWR VPWR _2098_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_4_10_0_m1_clk_local clkbuf_3_5_0_m1_clk_local/X VGND VGND VPWR VPWR _2513_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2021_ _2002_/X _2013_/D _2003_/Y VGND VGND VPWR VPWR _2021_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_47_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1736_ _1736_/A _2463_/Q VGND VGND VPWR VPWR _1831_/B sky130_fd_sc_hd__nor2_4
X_1805_ _1786_/Y _2573_/Q _1804_/X VGND VGND VPWR VPWR _1805_/X sky130_fd_sc_hd__o21a_4
X_1667_ _1667_/A _1667_/B _1667_/C _1667_/D VGND VGND VPWR VPWR _1667_/X sky130_fd_sc_hd__and4_4
X_1598_ _1443_/A _2390_/Q _1520_/A VGND VGND VPWR VPWR _1598_/X sky130_fd_sc_hd__o21a_4
XFILLER_53_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2219_ _2089_/Y _1624_/X _2218_/Y VGND VGND VPWR VPWR _2219_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_53_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2570_ _2570_/CLK _2570_/D VGND VGND VPWR VPWR _1735_/C sky130_fd_sc_hd__dfxtp_4
X_1383_ _1383_/A _2621_/Q _1383_/C _2619_/Q VGND VGND VPWR VPWR _1390_/B sky130_fd_sc_hd__and4_4
XFILLER_4_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1452_ _1440_/B _1440_/D _1451_/X VGND VGND VPWR VPWR _1452_/Y sky130_fd_sc_hd__a21oi_4
X_1521_ _1520_/X _1460_/X _1462_/X VGND VGND VPWR VPWR _1521_/Y sky130_fd_sc_hd__a21oi_4
X_2004_ _2002_/X _2003_/Y _2008_/A VGND VGND VPWR VPWR _2020_/A sky130_fd_sc_hd__nor3_4
XFILLER_23_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_7_0_addressalyzerBlock.SPI_CLK clkbuf_4_7_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2554_/CLK sky130_fd_sc_hd__clkbuf_1
X_1719_ _1719_/A _1640_/X VGND VGND VPWR VPWR _1719_/X sky130_fd_sc_hd__or2_4
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2553_ _2550_/CLK _2553_/D VGND VGND VPWR VPWR _2553_/Q sky130_fd_sc_hd__dfxtp_4
X_2622_ _2367_/CLK _2622_/D VGND VGND VPWR VPWR _1385_/A sky130_fd_sc_hd__dfxtp_4
X_1504_ _1494_/B VGND VGND VPWR VPWR _1505_/A sky130_fd_sc_hd__inv_2
X_2484_ _2470_/CLK _2046_/Y VGND VGND VPWR VPWR _1987_/A sky130_fd_sc_hd__dfxtp_4
X_1366_ _1365_/X VGND VGND VPWR VPWR _1366_/X sky130_fd_sc_hd__buf_2
X_1435_ _1434_/Y VGND VGND VPWR VPWR _1435_/Y sky130_fd_sc_hd__inv_2
X_1297_ _1296_/Y VGND VGND VPWR VPWR _2638_/D sky130_fd_sc_hd__inv_2
XFILLER_23_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1220_ _1219_/X VGND VGND VPWR VPWR _1221_/A sky130_fd_sc_hd__buf_2
XFILLER_52_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1984_ _1984_/A VGND VGND VPWR VPWR _1998_/A sky130_fd_sc_hd__inv_2
XFILLER_60_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2467_ _2457_/CLK _2467_/D VGND VGND VPWR VPWR _2467_/Q sky130_fd_sc_hd__dfxtp_4
X_2536_ _2519_/CLK _1916_/X VGND VGND VPWR VPWR HASH_ADDR[5] sky130_fd_sc_hd__dfxtp_4
X_2605_ _2388_/CLK _2605_/D VGND VGND VPWR VPWR _1483_/B sky130_fd_sc_hd__dfxtp_4
X_1349_ _1349_/A VGND VGND VPWR VPWR _1349_/Y sky130_fd_sc_hd__inv_2
X_1418_ _1409_/A _1409_/C VGND VGND VPWR VPWR _1419_/A sky130_fd_sc_hd__or2_4
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2398_ _2606_/CLK _2318_/X VGND VGND VPWR VPWR _1773_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_51_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2321_ _2223_/Y _2310_/X _1520_/X _2312_/X VGND VGND VPWR VPWR _2395_/D sky130_fd_sc_hd__a2bb2o_4
X_1203_ _2647_/Q _1194_/B _1202_/X VGND VGND VPWR VPWR _1203_/Y sky130_fd_sc_hd__o21ai_4
X_2252_ _2244_/X _2133_/Y _2247_/X _1905_/B _2249_/X VGND VGND VPWR VPWR _2431_/D
+ sky130_fd_sc_hd__o32ai_4
X_2183_ _2180_/X _2182_/X _1701_/A VGND VGND VPWR VPWR _2183_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_33_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1898_ _2096_/A VGND VGND VPWR VPWR _1900_/A sky130_fd_sc_hd__buf_2
X_1967_ _1284_/X _1966_/Y VGND VGND VPWR VPWR _2503_/D sky130_fd_sc_hd__nor2_4
X_2519_ _2519_/CLK _1940_/Y VGND VGND VPWR VPWR _2519_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1683_ _1683_/A VGND VGND VPWR VPWR _1683_/Y sky130_fd_sc_hd__inv_2
X_1821_ _2574_/Q _1809_/X _1820_/X VGND VGND VPWR VPWR _2575_/D sky130_fd_sc_hd__o21a_4
X_1752_ _2134_/C _1751_/A _1633_/X _1751_/Y VGND VGND VPWR VPWR _1752_/X sky130_fd_sc_hd__a211o_4
X_2304_ _2304_/A _1602_/C _1409_/A VGND VGND VPWR VPWR _2304_/Y sky130_fd_sc_hd__nand3_4
X_2097_ _2108_/A _2097_/B VGND VGND VPWR VPWR _2097_/X sky130_fd_sc_hd__and2_4
XFILLER_57_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2166_ _2166_/A THREAD_COUNT[3] VGND VGND VPWR VPWR _2166_/Y sky130_fd_sc_hd__nand2_4
X_2235_ _2233_/Y _2234_/X VGND VGND VPWR VPWR _2235_/Y sky130_fd_sc_hd__nand2_4
XFILLER_38_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2020_ _2020_/A VGND VGND VPWR VPWR _2022_/A sky130_fd_sc_hd__inv_2
XFILLER_39_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1735_ _1829_/A _1179_/A _1735_/C _1735_/D VGND VGND VPWR VPWR _1831_/A sky130_fd_sc_hd__nand4_4
X_1666_ _2146_/A VGND VGND VPWR VPWR _2166_/A sky130_fd_sc_hd__buf_2
X_1804_ _2591_/Q _1514_/X _1799_/X VGND VGND VPWR VPWR _1804_/X sky130_fd_sc_hd__o21a_4
X_1597_ _1664_/A VGND VGND VPWR VPWR _1600_/B sky130_fd_sc_hd__buf_2
XFILLER_53_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2149_ _1534_/A _2554_/Q _2148_/X VGND VGND VPWR VPWR _2149_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_26_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2218_ _1625_/X _2411_/Q _1617_/Y VGND VGND VPWR VPWR _2218_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_14_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_m1_clk_local clkbuf_0_m1_clk_local/X VGND VGND VPWR VPWR clkbuf_2_3_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
X_1520_ _1520_/A VGND VGND VPWR VPWR _1520_/X sky130_fd_sc_hd__buf_2
X_1382_ _1373_/B _1366_/X _1381_/Y VGND VGND VPWR VPWR _2623_/D sky130_fd_sc_hd__o21a_4
Xclkbuf_4_12_0_addressalyzerBlock.SPI_CLK clkbuf_3_6_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR _2590_/CLK sky130_fd_sc_hd__clkbuf_1
X_1451_ _1434_/Y VGND VGND VPWR VPWR _1451_/X sky130_fd_sc_hd__buf_2
X_2003_ _1999_/A VGND VGND VPWR VPWR _2003_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1649_ _1659_/A _1649_/B VGND VGND VPWR VPWR _1649_/Y sky130_fd_sc_hd__nor2_4
X_1718_ _1702_/Y _1717_/Y _1614_/X VGND VGND VPWR VPWR _1718_/Y sky130_fd_sc_hd__o21ai_4
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2483_ _2483_/CLK _2050_/Y VGND VGND VPWR VPWR _2030_/A sky130_fd_sc_hd__dfxtp_4
X_2621_ _2367_/CLK _1390_/Y VGND VGND VPWR VPWR _2621_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2552_ _2554_/CLK _1889_/X VGND VGND VPWR VPWR _2552_/Q sky130_fd_sc_hd__dfxtp_4
X_1503_ _1503_/A VGND VGND VPWR VPWR _1503_/Y sky130_fd_sc_hd__inv_2
X_1365_ _1383_/A _1383_/C _2619_/Q _1365_/D VGND VGND VPWR VPWR _1365_/X sky130_fd_sc_hd__and4_4
X_1434_ _2386_/Q _1566_/A VGND VGND VPWR VPWR _1434_/Y sky130_fd_sc_hd__nor2_4
X_1296_ _1296_/A _1296_/B VGND VGND VPWR VPWR _1296_/Y sky130_fd_sc_hd__nand2_4
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_4_0_m1_clk_local clkbuf_3_4_0_m1_clk_local/A VGND VGND VPWR VPWR clkbuf_4_9_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1983_ _1222_/X _1983_/B VGND VGND VPWR VPWR _1983_/Y sky130_fd_sc_hd__nor2_4
XFILLER_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2604_ _2598_/CLK _2604_/D VGND VGND VPWR VPWR _2604_/Q sky130_fd_sc_hd__dfxtp_4
X_2466_ _2550_/CLK _2094_/X VGND VGND VPWR VPWR _2351_/C sky130_fd_sc_hd__dfxtp_4
X_1417_ _1417_/A VGND VGND VPWR VPWR _2614_/D sky130_fd_sc_hd__inv_2
X_2535_ _2519_/CLK _1917_/X VGND VGND VPWR VPWR HASH_ADDR[4] sky130_fd_sc_hd__dfxtp_4
X_1348_ _1347_/Y VGND VGND VPWR VPWR _2629_/D sky130_fd_sc_hd__inv_2
XFILLER_36_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1279_ _1279_/A VGND VGND VPWR VPWR _1279_/Y sky130_fd_sc_hd__inv_2
X_2397_ _2410_/CLK _2319_/X VGND VGND VPWR VPWR _2397_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2251_ _2244_/X _2130_/Y _2247_/X _1902_/Y _2249_/X VGND VGND VPWR VPWR _2432_/D
+ sky130_fd_sc_hd__o32ai_4
X_2320_ _1764_/Y _2310_/X _1514_/X _2312_/X VGND VGND VPWR VPWR _2320_/X sky130_fd_sc_hd__a2bb2o_4
X_1202_ _2648_/Q _1179_/A VGND VGND VPWR VPWR _1202_/X sky130_fd_sc_hd__or2_4
X_2182_ _2441_/Q _1635_/X _1632_/Y _2181_/Y VGND VGND VPWR VPWR _2182_/X sky130_fd_sc_hd__a211o_4
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1966_ _1966_/A VGND VGND VPWR VPWR _1966_/Y sky130_fd_sc_hd__inv_2
X_1897_ _1896_/A _1897_/B VGND VGND VPWR VPWR _2545_/D sky130_fd_sc_hd__and2_4
X_2449_ _2598_/CLK _2449_/D VGND VGND VPWR VPWR _2449_/Q sky130_fd_sc_hd__dfxtp_4
X_2518_ _2528_/CLK _2518_/D VGND VGND VPWR VPWR _2518_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1820_ _2575_/Q _1810_/X _1813_/X VGND VGND VPWR VPWR _1820_/X sky130_fd_sc_hd__o21a_4
XFILLER_15_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1682_ _1566_/X _1577_/X _1683_/A _2385_/Q _1681_/X VGND VGND VPWR VPWR _1682_/Y
+ sky130_fd_sc_hd__o41ai_4
X_1751_ _1751_/A _1751_/B VGND VGND VPWR VPWR _1751_/Y sky130_fd_sc_hd__nor2_4
X_2234_ _1860_/B _2543_/Q _1661_/D _2234_/D VGND VGND VPWR VPWR _2234_/X sky130_fd_sc_hd__or4_4
X_2303_ _2136_/Y _2291_/X _2302_/Y VGND VGND VPWR VPWR _2303_/Y sky130_fd_sc_hd__o21ai_4
X_2096_ _2096_/A VGND VGND VPWR VPWR _2108_/A sky130_fd_sc_hd__buf_2
X_2165_ _2162_/Y _2163_/X _2164_/X VGND VGND VPWR VPWR _2165_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_38_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1949_ _1947_/A _1948_/Y VGND VGND VPWR VPWR _1949_/Y sky130_fd_sc_hd__nor2_4
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1803_ _1786_/Y _2574_/Q _1802_/X VGND VGND VPWR VPWR _2582_/D sky130_fd_sc_hd__o21a_4
X_1734_ _1733_/Y VGND VGND VPWR VPWR _2592_/D sky130_fd_sc_hd__inv_2
X_1665_ _1570_/A _1664_/Y _1660_/A VGND VGND VPWR VPWR _2146_/A sky130_fd_sc_hd__nor3_4
X_1596_ _1545_/X _1576_/X _1588_/Y _1593_/Y _1595_/X VGND VGND VPWR VPWR _2598_/D
+ sky130_fd_sc_hd__a41oi_4
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2217_ _1534_/X _2551_/Q _1640_/X VGND VGND VPWR VPWR _2217_/Y sky130_fd_sc_hd__o21ai_4
X_2079_ _2078_/X _1991_/B _1991_/C VGND VGND VPWR VPWR _2084_/C sky130_fd_sc_hd__nand3_4
XFILLER_38_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2148_ _1613_/Y VGND VGND VPWR VPWR _2148_/X sky130_fd_sc_hd__buf_2
XFILLER_55_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1450_ _1446_/Y VGND VGND VPWR VPWR _1450_/X sky130_fd_sc_hd__buf_2
X_1381_ _1373_/B _1379_/X _1385_/D _1365_/D _1275_/X VGND VGND VPWR VPWR _1381_/Y
+ sky130_fd_sc_hd__a41oi_4
X_2002_ _1998_/A VGND VGND VPWR VPWR _2002_/X sky130_fd_sc_hd__buf_2
XFILLER_50_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1648_ _1667_/B VGND VGND VPWR VPWR _1649_/B sky130_fd_sc_hd__inv_2
X_1579_ _1428_/B VGND VGND VPWR VPWR _1579_/X sky130_fd_sc_hd__buf_2
XFILLER_6_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1717_ _1712_/Y _1633_/X _1716_/Y VGND VGND VPWR VPWR _1717_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_58_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2620_ _2367_/CLK _2620_/D VGND VGND VPWR VPWR _2620_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_9_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2482_ _2483_/CLK _2052_/Y VGND VGND VPWR VPWR _1985_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2551_ _2554_/CLK _2551_/D VGND VGND VPWR VPWR _2551_/Q sky130_fd_sc_hd__dfxtp_4
X_1502_ _1496_/Y _1498_/Y _1501_/X VGND VGND VPWR VPWR _1502_/Y sky130_fd_sc_hd__a21oi_4
X_1433_ _1433_/A VGND VGND VPWR VPWR _1440_/B sky130_fd_sc_hd__buf_2
X_1364_ _2620_/Q VGND VGND VPWR VPWR _1383_/C sky130_fd_sc_hd__buf_2
X_1295_ _1295_/A _1308_/A _1299_/A _1292_/C VGND VGND VPWR VPWR _1296_/B sky130_fd_sc_hd__nand4_4
XFILLER_23_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_3_0_addressalyzerBlock.SPI_CLK clkbuf_2_3_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_10_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1982_ _1981_/X VGND VGND VPWR VPWR _2495_/D sky130_fd_sc_hd__inv_2
XFILLER_33_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2534_ _2496_/CLK _1918_/X VGND VGND VPWR VPWR HASH_ADDR[3] sky130_fd_sc_hd__dfxtp_4
XFILLER_9_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2603_ _2598_/CLK _2603_/D VGND VGND VPWR VPWR _2603_/Q sky130_fd_sc_hd__dfxtp_4
X_2465_ _2457_/CLK _2095_/X VGND VGND VPWR VPWR _2094_/B sky130_fd_sc_hd__dfxtp_4
X_1416_ _1413_/Y _1419_/C _1415_/Y VGND VGND VPWR VPWR _1417_/A sky130_fd_sc_hd__o21ai_4
X_1347_ _1344_/X _1345_/Y _1346_/X VGND VGND VPWR VPWR _1347_/Y sky130_fd_sc_hd__nand3_4
XFILLER_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2396_ _2410_/CLK _2320_/X VGND VGND VPWR VPWR _1764_/A sky130_fd_sc_hd__dfxtp_4
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1278_ _1276_/Y _1278_/B VGND VGND VPWR VPWR _1279_/A sky130_fd_sc_hd__nand2_4
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1201_ _1199_/Y _1187_/X _1200_/Y VGND VGND VPWR VPWR _1201_/Y sky130_fd_sc_hd__a21oi_4
X_2250_ _2244_/X _2127_/Y _2247_/X _1710_/B _2249_/X VGND VGND VPWR VPWR _2433_/D
+ sky130_fd_sc_hd__o32ai_4
X_2181_ _2181_/A _1771_/Y VGND VGND VPWR VPWR _2181_/Y sky130_fd_sc_hd__nor2_4
XFILLER_33_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1965_ _1284_/X _1965_/B VGND VGND VPWR VPWR _1965_/Y sky130_fd_sc_hd__nor2_4
X_1896_ _1896_/A _2550_/Q VGND VGND VPWR VPWR _2546_/D sky130_fd_sc_hd__and2_4
X_2517_ _2638_/CLK _1945_/Y VGND VGND VPWR VPWR _1957_/B sky130_fd_sc_hd__dfxtp_4
X_2379_ _2498_/CLK _2379_/D VGND VGND VPWR VPWR _2379_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2448_ _2557_/CLK _2448_/D VGND VGND VPWR VPWR _2448_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_17_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1750_ _1750_/A VGND VGND VPWR VPWR _1751_/B sky130_fd_sc_hd__inv_2
X_1681_ _1679_/Y _1680_/X _1529_/Y VGND VGND VPWR VPWR _1681_/X sky130_fd_sc_hd__o21a_4
X_2233_ _2216_/Y _2231_/Y _2232_/Y VGND VGND VPWR VPWR _2233_/Y sky130_fd_sc_hd__o21ai_4
X_2164_ _1611_/A _1236_/A _1656_/A VGND VGND VPWR VPWR _2164_/X sky130_fd_sc_hd__a21o_4
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2302_ _2304_/A _1602_/C HASH_LED VGND VGND VPWR VPWR _2302_/Y sky130_fd_sc_hd__nand3_4
X_2095_ _1900_/A IRQ_OUT_fromClient VGND VGND VPWR VPWR _2095_/X sky130_fd_sc_hd__and2_4
XFILLER_53_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1879_ _1878_/A DATA_FROM_HASH[1] VGND VGND VPWR VPWR _2560_/D sky130_fd_sc_hd__and2_4
X_1948_ _1948_/A VGND VGND VPWR VPWR _1948_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1733_ _1730_/X _1731_/Y _1732_/Y VGND VGND VPWR VPWR _1733_/Y sky130_fd_sc_hd__o21ai_4
X_1802_ _2591_/Q _1503_/A _1799_/X VGND VGND VPWR VPWR _1802_/X sky130_fd_sc_hd__o21a_4
X_1664_ _1664_/A _1579_/X _1428_/C VGND VGND VPWR VPWR _1664_/Y sky130_fd_sc_hd__nand3_4
X_1595_ _1549_/A _1594_/X _1781_/A VGND VGND VPWR VPWR _1595_/X sky130_fd_sc_hd__a21o_4
X_2147_ _2616_/Q _1571_/A _1661_/C _1661_/D _2146_/Y VGND VGND VPWR VPWR _2147_/Y
+ sky130_fd_sc_hd__o41ai_4
X_2216_ _1409_/C _1860_/B _1661_/C _1661_/D _2146_/Y VGND VGND VPWR VPWR _2216_/Y
+ sky130_fd_sc_hd__o41ai_4
XFILLER_26_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2078_ _1991_/A VGND VGND VPWR VPWR _2078_/X sky130_fd_sc_hd__buf_2
XFILLER_26_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1380_ _1383_/C VGND VGND VPWR VPWR _1385_/D sky130_fd_sc_hd__buf_2
X_2001_ _2010_/C _2001_/B VGND VGND VPWR VPWR _2001_/Y sky130_fd_sc_hd__nand2_4
XFILLER_50_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1716_ _1715_/X _1534_/A VGND VGND VPWR VPWR _1716_/Y sky130_fd_sc_hd__nand2_4
XFILLER_58_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1647_ _1667_/C _1667_/D VGND VGND VPWR VPWR _1659_/A sky130_fd_sc_hd__nand2_4
X_1578_ _1577_/X _1460_/X _1503_/A VGND VGND VPWR VPWR _1578_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_26_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2550_ _2550_/CLK _2550_/D VGND VGND VPWR VPWR _2550_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_13_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2481_ _2483_/CLK _2057_/X VGND VGND VPWR VPWR _1993_/D sky130_fd_sc_hd__dfxtp_4
X_1363_ _1397_/B _1233_/C _1397_/C VGND VGND VPWR VPWR _1383_/A sky130_fd_sc_hd__nor3_4
X_1501_ _1450_/X _1499_/Y _1500_/X VGND VGND VPWR VPWR _1501_/X sky130_fd_sc_hd__a21o_4
X_1432_ _1429_/Y _1701_/A _1466_/A _2602_/Q VGND VGND VPWR VPWR _1433_/A sky130_fd_sc_hd__and4_4
X_1294_ _1301_/A _1293_/Y _1275_/X VGND VGND VPWR VPWR _1296_/A sky130_fd_sc_hd__a21oi_4
XFILLER_54_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1981_ _1979_/A _1976_/A _1976_/B VGND VGND VPWR VPWR _1981_/X sky130_fd_sc_hd__or3_4
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2602_ _2388_/CLK _1551_/Y VGND VGND VPWR VPWR _2602_/Q sky130_fd_sc_hd__dfxtp_4
X_2533_ _2519_/CLK _2533_/D VGND VGND VPWR VPWR HASH_ADDR[2] sky130_fd_sc_hd__dfxtp_4
X_2464_ _2457_/CLK _2097_/X VGND VGND VPWR VPWR _2464_/Q sky130_fd_sc_hd__dfxtp_4
X_1415_ _1419_/C _1413_/Y _1283_/X VGND VGND VPWR VPWR _1415_/Y sky130_fd_sc_hd__a21oi_4
X_1346_ _1270_/A VGND VGND VPWR VPWR _1346_/X sky130_fd_sc_hd__buf_2
XFILLER_3_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2395_ _2410_/CLK _2395_/D VGND VGND VPWR VPWR _1767_/B sky130_fd_sc_hd__dfxtp_4
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1277_ _1277_/A _1277_/B _2641_/Q _1277_/D VGND VGND VPWR VPWR _1278_/B sky130_fd_sc_hd__nand4_4
XFILLER_24_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1200_ _1762_/B _1216_/B _1191_/X VGND VGND VPWR VPWR _1200_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_2_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2180_ _2176_/Y _2179_/Y _2449_/Q VGND VGND VPWR VPWR _2180_/X sky130_fd_sc_hd__a21o_4
XFILLER_18_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1895_ _1896_/A DATA_AVAILABLE[0] VGND VGND VPWR VPWR _2547_/D sky130_fd_sc_hd__and2_4
Xclkbuf_3_0_0_m1_clk_local clkbuf_3_1_0_m1_clk_local/A VGND VGND VPWR VPWR clkbuf_4_1_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
X_1964_ _1964_/A VGND VGND VPWR VPWR _1965_/B sky130_fd_sc_hd__inv_2
X_2447_ _2557_/CLK _2117_/Y VGND VGND VPWR VPWR _2447_/Q sky130_fd_sc_hd__dfxtp_4
X_2516_ _2638_/CLK _1947_/Y VGND VGND VPWR VPWR _1958_/B sky130_fd_sc_hd__dfxtp_4
X_2378_ _2498_/CLK _2377_/Q VGND VGND VPWR VPWR _2379_/D sky130_fd_sc_hd__dfxtp_4
X_1329_ _2629_/Q VGND VGND VPWR VPWR _1329_/X sky130_fd_sc_hd__buf_2
XFILLER_17_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1680_ _1185_/A _1680_/B VGND VGND VPWR VPWR _1680_/X sky130_fd_sc_hd__or2_4
X_2301_ _1490_/Y _2291_/X _2300_/Y VGND VGND VPWR VPWR _2407_/D sky130_fd_sc_hd__o21ai_4
X_2232_ THREAD_COUNT[0] _2166_/A _2168_/Y VGND VGND VPWR VPWR _2232_/Y sky130_fd_sc_hd__a21boi_4
X_2163_ _1335_/A _1646_/X _1741_/Y VGND VGND VPWR VPWR _2163_/X sky130_fd_sc_hd__o21a_4
XFILLER_38_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2094_ _1900_/A _2094_/B VGND VGND VPWR VPWR _2094_/X sky130_fd_sc_hd__and2_4
XFILLER_0_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1878_ _1878_/A DATA_FROM_HASH[2] VGND VGND VPWR VPWR _2561_/D sky130_fd_sc_hd__and2_4
X_1947_ _1947_/A _1947_/B VGND VGND VPWR VPWR _1947_/Y sky130_fd_sc_hd__nor2_4
XFILLER_52_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1732_ _1730_/X _1739_/A _1781_/A VGND VGND VPWR VPWR _1732_/Y sky130_fd_sc_hd__a21oi_4
X_1663_ _1662_/Y VGND VGND VPWR VPWR _1739_/A sky130_fd_sc_hd__buf_2
X_1801_ _1786_/Y _2575_/Q _1800_/X VGND VGND VPWR VPWR _2583_/D sky130_fd_sc_hd__o21a_4
X_1594_ _1590_/B VGND VGND VPWR VPWR _1594_/X sky130_fd_sc_hd__buf_2
X_2146_ _2146_/A VGND VGND VPWR VPWR _2146_/Y sky130_fd_sc_hd__inv_2
X_2077_ _2071_/Y _2060_/B _2076_/Y VGND VGND VPWR VPWR _2475_/D sky130_fd_sc_hd__a21oi_4
X_2215_ _1726_/A _2213_/Y _2214_/Y VGND VGND VPWR VPWR _2215_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_38_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2000_ CLK_LED VGND VGND VPWR VPWR _2001_/B sky130_fd_sc_hd__inv_2
XFILLER_50_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_3_0_addressalyzerBlock.SPI_CLK clkbuf_2_1_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR clkbuf_4_7_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
X_1646_ _1646_/A VGND VGND VPWR VPWR _1646_/X sky130_fd_sc_hd__buf_2
Xclkbuf_4_9_0_m1_clk_local clkbuf_4_9_0_m1_clk_local/A VGND VGND VPWR VPWR _2370_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_1715_ _2445_/Q _1703_/X _1632_/Y _1714_/Y VGND VGND VPWR VPWR _1715_/X sky130_fd_sc_hd__a211o_4
X_1577_ _1443_/A VGND VGND VPWR VPWR _1577_/X sky130_fd_sc_hd__buf_2
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2129_ _2120_/X _2127_/Y _2128_/Y VGND VGND VPWR VPWR _2445_/D sky130_fd_sc_hd__o21ai_4
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2480_ _2483_/CLK _2480_/D VGND VGND VPWR VPWR _1993_/C sky130_fd_sc_hd__dfxtp_4
X_1500_ _1221_/A VGND VGND VPWR VPWR _1500_/X sky130_fd_sc_hd__buf_2
XFILLER_9_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1362_ _1367_/A _1361_/Y _1306_/X VGND VGND VPWR VPWR _1362_/X sky130_fd_sc_hd__o21a_4
X_1293_ _1295_/A VGND VGND VPWR VPWR _1293_/Y sky130_fd_sc_hd__inv_2
X_1431_ _2603_/Q VGND VGND VPWR VPWR _1466_/A sky130_fd_sc_hd__buf_2
XFILLER_51_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1629_ _1621_/X _1627_/Y _1628_/X VGND VGND VPWR VPWR _1629_/X sky130_fd_sc_hd__a21o_4
XFILLER_46_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1980_ _1980_/A _1980_/B _1979_/X VGND VGND VPWR VPWR _2496_/D sky130_fd_sc_hd__and3_4
XFILLER_9_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2532_ _2496_/CLK _1920_/X VGND VGND VPWR VPWR HASH_ADDR[1] sky130_fd_sc_hd__dfxtp_4
X_2463_ _2570_/CLK _2099_/X VGND VGND VPWR VPWR _2463_/Q sky130_fd_sc_hd__dfxtp_4
X_2601_ _2388_/CLK _1557_/X VGND VGND VPWR VPWR _1608_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_9_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1345_ _1333_/Y VGND VGND VPWR VPWR _1345_/Y sky130_fd_sc_hd__inv_2
X_1414_ _1409_/A _1409_/C VGND VGND VPWR VPWR _1419_/C sky130_fd_sc_hd__nand2_4
X_2394_ _2590_/CLK _2325_/X VGND VGND VPWR VPWR _1728_/C sky130_fd_sc_hd__dfxtp_4
X_1276_ _1282_/C _1854_/A _1275_/X VGND VGND VPWR VPWR _1276_/Y sky130_fd_sc_hd__a21oi_4
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1894_ _1896_/A DATA_AVAILABLE[1] VGND VGND VPWR VPWR _1894_/X sky130_fd_sc_hd__and2_4
X_1963_ _1947_/A _1963_/B VGND VGND VPWR VPWR _1963_/Y sky130_fd_sc_hd__nor2_4
X_2446_ _2410_/CLK _2446_/D VGND VGND VPWR VPWR _2125_/C sky130_fd_sc_hd__dfxtp_4
X_2515_ _2638_/CLK _1949_/Y VGND VGND VPWR VPWR _2515_/Q sky130_fd_sc_hd__dfxtp_4
X_2377_ _2498_/CLK _2377_/D VGND VGND VPWR VPWR _2377_/Q sky130_fd_sc_hd__dfxtp_4
X_1328_ _1242_/B VGND VGND VPWR VPWR _1335_/C sky130_fd_sc_hd__buf_2
X_1259_ _1226_/Y VGND VGND VPWR VPWR _1292_/C sky130_fd_sc_hd__inv_2
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2231_ _2228_/Y _2229_/Y _2230_/X VGND VGND VPWR VPWR _2231_/Y sky130_fd_sc_hd__a21oi_4
X_2300_ _2304_/A _2298_/B _2300_/C VGND VGND VPWR VPWR _2300_/Y sky130_fd_sc_hd__nand3_4
X_2093_ _1900_/A _2093_/B VGND VGND VPWR VPWR _2467_/D sky130_fd_sc_hd__and2_4
XFILLER_53_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2162_ _2149_/Y _2160_/Y _2161_/Y VGND VGND VPWR VPWR _2162_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_38_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1877_ _1878_/A DATA_FROM_HASH[3] VGND VGND VPWR VPWR _2562_/D sky130_fd_sc_hd__and2_4
X_1946_ _2420_/Q VGND VGND VPWR VPWR _1947_/B sky130_fd_sc_hd__inv_2
X_2429_ _2428_/CLK _2429_/D VGND VGND VPWR VPWR _2177_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_44_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1800_ _1788_/X _2253_/C _1799_/X VGND VGND VPWR VPWR _1800_/X sky130_fd_sc_hd__o21a_4
XFILLER_18_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1662_ _1662_/A VGND VGND VPWR VPWR _1662_/Y sky130_fd_sc_hd__inv_2
X_1731_ _1697_/A _1731_/B _1689_/A VGND VGND VPWR VPWR _1731_/Y sky130_fd_sc_hd__nor3_4
XFILLER_11_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2214_ _1762_/A _2436_/Q VGND VGND VPWR VPWR _2214_/Y sky130_fd_sc_hd__nand2_4
X_1593_ _1613_/A _1667_/B _1488_/X VGND VGND VPWR VPWR _1593_/Y sky130_fd_sc_hd__o21ai_4
X_2076_ _2071_/Y _2060_/B _1346_/X VGND VGND VPWR VPWR _2076_/Y sky130_fd_sc_hd__o21ai_4
X_2145_ _2144_/Y _2138_/Y _2125_/A _1966_/Y _2139_/X VGND VGND VPWR VPWR _2439_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_34_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1929_ _2411_/Q VGND VGND VPWR VPWR _1929_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1645_ _1645_/A VGND VGND VPWR VPWR _1646_/A sky130_fd_sc_hd__inv_2
X_1576_ _2337_/A _1575_/Y _1445_/A _1445_/D _1185_/A VGND VGND VPWR VPWR _1576_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_6_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1714_ _1630_/X _1713_/Y VGND VGND VPWR VPWR _1714_/Y sky130_fd_sc_hd__nor2_4
XFILLER_54_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2059_ _1992_/D VGND VGND VPWR VPWR _2060_/B sky130_fd_sc_hd__buf_2
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2128_ _2125_/A _2335_/A _2445_/Q VGND VGND VPWR VPWR _2128_/Y sky130_fd_sc_hd__nand3_4
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1430_ _2604_/Q VGND VGND VPWR VPWR _1701_/A sky130_fd_sc_hd__buf_2
X_1361_ _1360_/Y _1350_/X VGND VGND VPWR VPWR _1361_/Y sky130_fd_sc_hd__nor2_4
X_1292_ _1308_/A _1299_/A _1292_/C VGND VGND VPWR VPWR _1301_/A sky130_fd_sc_hd__nand3_4
XFILLER_36_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1559_ _1570_/A _1559_/B VGND VGND VPWR VPWR _1667_/A sky130_fd_sc_hd__nor2_4
X_1628_ _2449_/Q VGND VGND VPWR VPWR _1628_/X sky130_fd_sc_hd__buf_2
XFILLER_54_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2600_ _2590_/CLK _2600_/D VGND VGND VPWR VPWR _2600_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1413_ _1409_/B VGND VGND VPWR VPWR _1413_/Y sky130_fd_sc_hd__inv_2
X_2393_ _2570_/CLK _2393_/D VGND VGND VPWR VPWR _1697_/A sky130_fd_sc_hd__dfxtp_4
X_2462_ _2390_/CLK _2462_/D VGND VGND VPWR VPWR _1680_/B sky130_fd_sc_hd__dfxtp_4
X_2531_ _2513_/CLK _2531_/D VGND VGND VPWR VPWR HASH_ADDR[0] sky130_fd_sc_hd__dfxtp_4
X_1275_ _1274_/X VGND VGND VPWR VPWR _1275_/X sky130_fd_sc_hd__buf_2
X_1344_ _1324_/X _1321_/X _1329_/X VGND VGND VPWR VPWR _1344_/X sky130_fd_sc_hd__a21o_4
XFILLER_59_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1962_ _2441_/Q VGND VGND VPWR VPWR _1963_/B sky130_fd_sc_hd__inv_2
X_1893_ _1896_/A DATA_AVAILABLE[2] VGND VGND VPWR VPWR _2549_/D sky130_fd_sc_hd__and2_4
X_2376_ _2498_/CLK _2376_/D VGND VGND VPWR VPWR _2377_/D sky130_fd_sc_hd__dfxtp_4
X_2514_ _2513_/CLK _1951_/X VGND VGND VPWR VPWR DATA_TO_HASH[7] sky130_fd_sc_hd__dfxtp_4
X_2445_ _2445_/CLK _2445_/D VGND VGND VPWR VPWR _2445_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1258_ _1228_/Y _1240_/Y _1238_/Y VGND VGND VPWR VPWR _1258_/Y sky130_fd_sc_hd__nor3_4
X_1189_ _2384_/Q VGND VGND VPWR VPWR _1189_/Y sky130_fd_sc_hd__inv_2
X_1327_ _1326_/Y VGND VGND VPWR VPWR _2633_/D sky130_fd_sc_hd__inv_2
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2230_ _1612_/A _2621_/Q _1656_/A VGND VGND VPWR VPWR _2230_/X sky130_fd_sc_hd__a21o_4
XFILLER_46_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2092_ _1222_/X _2091_/Y VGND VGND VPWR VPWR _2092_/Y sky130_fd_sc_hd__nor2_4
XFILLER_38_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2161_ _1256_/Y _2148_/X _1651_/X _1856_/A VGND VGND VPWR VPWR _2161_/Y sky130_fd_sc_hd__a2bb2oi_4
XFILLER_0_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1945_ _1947_/A _1945_/B VGND VGND VPWR VPWR _1945_/Y sky130_fd_sc_hd__nor2_4
XFILLER_21_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1876_ _1878_/A DATA_FROM_HASH[4] VGND VGND VPWR VPWR _1876_/X sky130_fd_sc_hd__and2_4
X_2359_ EXT_RESET_N_fromHost VGND VGND VPWR VPWR EXT_RESET_N_toClient sky130_fd_sc_hd__buf_2
XFILLER_56_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2428_ _2428_/CLK _2428_/D VGND VGND VPWR VPWR _2428_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_44_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_3_0_addressalyzerBlock.SPI_CLK clkbuf_4_3_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2410_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_60_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1661_ _1383_/C _1860_/B _1661_/C _1661_/D VGND VGND VPWR VPWR _1661_/X sky130_fd_sc_hd__or4_4
X_1730_ _1728_/C _1434_/Y _1728_/Y _1729_/Y VGND VGND VPWR VPWR _1730_/X sky130_fd_sc_hd__a211o_4
X_1592_ _1426_/A _1664_/A VGND VGND VPWR VPWR _1667_/B sky130_fd_sc_hd__nor2_4
X_2213_ _2544_/Q _1739_/B _2212_/Y _2168_/Y VGND VGND VPWR VPWR _2213_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_38_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2144_ _1520_/X VGND VGND VPWR VPWR _2144_/Y sky130_fd_sc_hd__inv_2
X_2075_ _2075_/A VGND VGND VPWR VPWR _2075_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1859_ _1612_/X _1857_/Y _1858_/Y VGND VGND VPWR VPWR _1859_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1928_ _1930_/A _1927_/Y VGND VGND VPWR VPWR _2528_/D sky130_fd_sc_hd__nor2_4
Xclkbuf_2_2_0_m1_clk_local clkbuf_2_3_0_m1_clk_local/A VGND VGND VPWR VPWR clkbuf_3_4_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1713_ _1768_/B VGND VGND VPWR VPWR _1713_/Y sky130_fd_sc_hd__inv_2
X_1644_ _1643_/X VGND VGND VPWR VPWR _1645_/A sky130_fd_sc_hd__buf_2
X_1575_ _1566_/A VGND VGND VPWR VPWR _1575_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2127_ _1840_/B _2121_/X _1459_/A VGND VGND VPWR VPWR _2127_/Y sky130_fd_sc_hd__nand3_4
X_2058_ _2477_/Q VGND VGND VPWR VPWR _2058_/X sky130_fd_sc_hd__buf_2
XFILLER_41_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1360_ _1360_/A VGND VGND VPWR VPWR _1360_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1291_ _1246_/Y VGND VGND VPWR VPWR _1308_/A sky130_fd_sc_hd__inv_2
XFILLER_63_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1558_ _1428_/B VGND VGND VPWR VPWR _1559_/B sky130_fd_sc_hd__inv_2
X_1627_ _1622_/Y _1624_/X _1626_/Y VGND VGND VPWR VPWR _1627_/Y sky130_fd_sc_hd__o21ai_4
X_1489_ _1487_/Y _1488_/X _1450_/X VGND VGND VPWR VPWR _1489_/X sky130_fd_sc_hd__a21o_4
XFILLER_54_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_5_0_m1_clk_local clkbuf_4_5_0_m1_clk_local/A VGND VGND VPWR VPWR _2483_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2530_ _2528_/CLK _1924_/Y VGND VGND VPWR VPWR _1931_/B sky130_fd_sc_hd__dfxtp_4
X_1412_ _1411_/X _2010_/B _1397_/C VGND VGND VPWR VPWR _1412_/X sky130_fd_sc_hd__and3_4
X_1343_ _1335_/D _1333_/Y _1342_/Y VGND VGND VPWR VPWR _1343_/X sky130_fd_sc_hd__o21a_4
X_2392_ _2570_/CLK _2392_/D VGND VGND VPWR VPWR _2392_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_3_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2461_ _2390_/CLK _2461_/D VGND VGND VPWR VPWR _2461_/Q sky130_fd_sc_hd__dfxtp_4
X_1274_ _2363_/Q VGND VGND VPWR VPWR _1274_/X sky130_fd_sc_hd__buf_2
XFILLER_36_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1892_ _2096_/A VGND VGND VPWR VPWR _1896_/A sky130_fd_sc_hd__buf_2
X_1961_ _1947_/A _1960_/Y VGND VGND VPWR VPWR _2506_/D sky130_fd_sc_hd__nor2_4
X_2513_ _2513_/CLK _1952_/X VGND VGND VPWR VPWR DATA_TO_HASH[6] sky130_fd_sc_hd__dfxtp_4
X_2375_ _2496_/CLK _2375_/D VGND VGND VPWR VPWR _2376_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_56_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1326_ _1316_/B _1323_/Y _1325_/Y VGND VGND VPWR VPWR _1326_/Y sky130_fd_sc_hd__o21ai_4
X_2444_ _2445_/CLK _2444_/D VGND VGND VPWR VPWR _2444_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_64_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1188_ _1188_/A VGND VGND VPWR VPWR _1216_/B sky130_fd_sc_hd__buf_2
X_1257_ _1257_/A VGND VGND VPWR VPWR _1257_/X sky130_fd_sc_hd__buf_2
XFILLER_24_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_0 DATA_AVAILABLE[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2160_ _2157_/X _2159_/X _1701_/A VGND VGND VPWR VPWR _2160_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_61_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2091_ _2467_/Q VGND VGND VPWR VPWR _2091_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1875_ _1878_/A DATA_FROM_HASH[5] VGND VGND VPWR VPWR _2564_/D sky130_fd_sc_hd__and2_4
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1944_ _1944_/A VGND VGND VPWR VPWR _1945_/B sky130_fd_sc_hd__inv_2
X_2427_ _2445_/CLK _2427_/D VGND VGND VPWR VPWR _1913_/A sky130_fd_sc_hd__dfxtp_4
X_1309_ _1307_/X _1308_/Y VGND VGND VPWR VPWR _1309_/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2289_ _1219_/X _1579_/X _1691_/Y _1562_/A VGND VGND VPWR VPWR _2290_/A sky130_fd_sc_hd__nor4_4
X_2358_ VGND VGND VPWR VPWR _2358_/HI zero sky130_fd_sc_hd__conb_1
XFILLER_20_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1660_ _1660_/A VGND VGND VPWR VPWR _1661_/D sky130_fd_sc_hd__buf_2
X_1591_ _1427_/A VGND VGND VPWR VPWR _1664_/A sky130_fd_sc_hd__inv_2
XFILLER_7_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2212_ _2194_/Y _2210_/Y _2211_/Y VGND VGND VPWR VPWR _2212_/Y sky130_fd_sc_hd__o21ai_4
X_2143_ _2142_/Y _2138_/Y _2125_/A _1965_/B _2139_/X VGND VGND VPWR VPWR _2143_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_61_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2074_ _1990_/B _2072_/Y _2073_/Y VGND VGND VPWR VPWR _2075_/A sky130_fd_sc_hd__a21o_4
X_1858_ _1612_/X _1367_/A _1656_/X VGND VGND VPWR VPWR _1858_/Y sky130_fd_sc_hd__a21oi_4
X_1927_ _1927_/A VGND VGND VPWR VPWR _1927_/Y sky130_fd_sc_hd__inv_2
X_1789_ _1189_/Y VGND VGND VPWR VPWR _1838_/A sky130_fd_sc_hd__buf_2
XFILLER_44_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1643_ _1651_/A _1667_/B _1667_/C _1667_/D VGND VGND VPWR VPWR _1643_/X sky130_fd_sc_hd__and4_4
XFILLER_6_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1712_ _1712_/A _1711_/X VGND VGND VPWR VPWR _1712_/Y sky130_fd_sc_hd__nand2_4
X_1574_ _2386_/Q VGND VGND VPWR VPWR _2337_/A sky130_fd_sc_hd__inv_2
XFILLER_6_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_13_0_m1_clk_local clkbuf_3_6_0_m1_clk_local/X VGND VGND VPWR VPWR _2372_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_2057_ _2056_/X _2044_/B _2040_/X VGND VGND VPWR VPWR _2057_/X sky130_fd_sc_hd__and3_4
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2126_ _2120_/X _2122_/Y _2125_/Y VGND VGND VPWR VPWR _2446_/D sky130_fd_sc_hd__o21ai_4
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1290_ _1290_/A VGND VGND VPWR VPWR _1290_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1626_ _1625_/X _2434_/Q _2448_/Q VGND VGND VPWR VPWR _1626_/Y sky130_fd_sc_hd__a21oi_4
X_1557_ _1557_/A _2104_/A _1557_/C VGND VGND VPWR VPWR _1557_/X sky130_fd_sc_hd__and3_4
X_1488_ _1435_/Y VGND VGND VPWR VPWR _1488_/X sky130_fd_sc_hd__buf_2
XFILLER_54_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2109_ _2108_/A _2109_/B VGND VGND VPWR VPWR _2109_/X sky130_fd_sc_hd__and2_4
XFILLER_42_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2460_ _2570_/CLK _2104_/X VGND VGND VPWR VPWR _1178_/A sky130_fd_sc_hd__dfxtp_4
X_1411_ _2615_/Q _1411_/B VGND VGND VPWR VPWR _1411_/X sky130_fd_sc_hd__or2_4
X_1342_ _1335_/D _1324_/X _1329_/X _1321_/X _1339_/X VGND VGND VPWR VPWR _1342_/Y
+ sky130_fd_sc_hd__a41oi_4
X_2391_ _2570_/CLK _2391_/D VGND VGND VPWR VPWR _1689_/A sky130_fd_sc_hd__dfxtp_4
X_1273_ _1277_/A VGND VGND VPWR VPWR _1854_/A sky130_fd_sc_hd__inv_2
XFILLER_51_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1609_ _1651_/A _1609_/B _1667_/C _1667_/D VGND VGND VPWR VPWR _1609_/X sky130_fd_sc_hd__and4_4
X_2589_ _2390_/CLK _1782_/Y VGND VGND VPWR VPWR _1780_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_59_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1891_ _1891_/A DATA_AVAILABLE[3] VGND VGND VPWR VPWR _2550_/D sky130_fd_sc_hd__and2_4
X_1960_ _1960_/A VGND VGND VPWR VPWR _1960_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2443_ _2445_/CLK _2135_/Y VGND VGND VPWR VPWR _2134_/C sky130_fd_sc_hd__dfxtp_4
X_2512_ _2513_/CLK _1953_/X VGND VGND VPWR VPWR DATA_TO_HASH[5] sky130_fd_sc_hd__dfxtp_4
X_2374_ _2496_/CLK _2373_/Q VGND VGND VPWR VPWR _2375_/D sky130_fd_sc_hd__dfxtp_4
X_1325_ _1316_/B _1324_/X _1321_/X _1316_/D _1274_/X VGND VGND VPWR VPWR _1325_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1256_ _1277_/D VGND VGND VPWR VPWR _1256_/Y sky130_fd_sc_hd__inv_2
X_1187_ _1187_/A VGND VGND VPWR VPWR _1187_/X sky130_fd_sc_hd__buf_2
XFILLER_24_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE2_1 DATA_FROM_HASH[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_8_0_addressalyzerBlock.SPI_CLK clkbuf_4_9_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2606_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_23_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2090_ _1284_/X _2089_/Y VGND VGND VPWR VPWR _2090_/Y sky130_fd_sc_hd__nor2_4
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1874_ _1874_/A VGND VGND VPWR VPWR _1878_/A sky130_fd_sc_hd__buf_2
XFILLER_9_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1943_ _1339_/X VGND VGND VPWR VPWR _1947_/A sky130_fd_sc_hd__buf_2
X_2426_ _2428_/CLK _2426_/D VGND VGND VPWR VPWR _2426_/Q sky130_fd_sc_hd__dfxtp_4
X_1239_ _1228_/Y _1238_/Y VGND VGND VPWR VPWR _1239_/Y sky130_fd_sc_hd__nor2_4
X_1308_ _1308_/A _2636_/Q _1308_/C VGND VGND VPWR VPWR _1308_/Y sky130_fd_sc_hd__nand3_4
XFILLER_37_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2288_ _1581_/X _2260_/Y _2278_/A _1929_/Y _2279_/X VGND VGND VPWR VPWR _2411_/D
+ sky130_fd_sc_hd__o32ai_4
X_2357_ VGND VGND VPWR VPWR one _2357_/LO sky130_fd_sc_hd__conb_1
XFILLER_12_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1590_ _1428_/D _1590_/B VGND VGND VPWR VPWR _1613_/A sky130_fd_sc_hd__nor2_4
X_2073_ _1990_/B _2072_/Y _1374_/X VGND VGND VPWR VPWR _2073_/Y sky130_fd_sc_hd__o21ai_4
X_2211_ _2146_/A THREAD_COUNT[1] VGND VGND VPWR VPWR _2211_/Y sky130_fd_sc_hd__nand2_4
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2142_ _1514_/A VGND VGND VPWR VPWR _2142_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1857_ _1855_/Y _1646_/X _1856_/X VGND VGND VPWR VPWR _1857_/Y sky130_fd_sc_hd__a21oi_4
X_1788_ _2591_/Q VGND VGND VPWR VPWR _1788_/X sky130_fd_sc_hd__buf_2
X_1926_ _1930_/A _1925_/Y VGND VGND VPWR VPWR _2529_/D sky130_fd_sc_hd__nor2_4
XFILLER_39_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2409_ _2408_/CLK _2296_/Y VGND VGND VPWR VPWR _2295_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1642_ _1615_/Y _1639_/Y _1641_/X VGND VGND VPWR VPWR _1642_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_6_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1711_ _1937_/A _2181_/A _1708_/X _1710_/Y VGND VGND VPWR VPWR _1711_/X sky130_fd_sc_hd__a211o_4
X_1573_ _1564_/X _1572_/Y _1454_/X VGND VGND VPWR VPWR _2600_/D sky130_fd_sc_hd__a21oi_4
X_2056_ _2053_/Y _2062_/B _2055_/X _1993_/C _1993_/D VGND VGND VPWR VPWR _2056_/X
+ sky130_fd_sc_hd__a41o_4
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2125_ _2125_/A _2335_/A _2125_/C VGND VGND VPWR VPWR _2125_/Y sky130_fd_sc_hd__nand3_4
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1909_ _1901_/X _1908_/Y VGND VGND VPWR VPWR _2539_/D sky130_fd_sc_hd__nor2_4
XFILLER_22_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1556_ _1556_/A _1537_/X VGND VGND VPWR VPWR _1557_/C sky130_fd_sc_hd__nand2_4
X_1625_ _1623_/Y VGND VGND VPWR VPWR _1625_/X sky130_fd_sc_hd__buf_2
X_1487_ _1487_/A _1505_/B _1494_/B _1505_/C VGND VGND VPWR VPWR _1487_/Y sky130_fd_sc_hd__nand4_4
X_2108_ _2108_/A SCLK_fromHost VGND VGND VPWR VPWR _2456_/D sky130_fd_sc_hd__and2_4
XFILLER_54_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2039_ _2039_/A VGND VGND VPWR VPWR _2486_/D sky130_fd_sc_hd__inv_2
XFILLER_45_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1410_ _1409_/Y VGND VGND VPWR VPWR _1411_/B sky130_fd_sc_hd__inv_2
XFILLER_5_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1341_ _1335_/C _1338_/X _1340_/Y VGND VGND VPWR VPWR _1341_/X sky130_fd_sc_hd__o21a_4
X_2390_ _2390_/CLK _2390_/D VGND VGND VPWR VPWR _2390_/Q sky130_fd_sc_hd__dfxtp_4
X_1272_ _2641_/Q _1265_/Y _1277_/D _1224_/A VGND VGND VPWR VPWR _1282_/C sky130_fd_sc_hd__nand4_4
X_1608_ _2602_/Q _1608_/B VGND VGND VPWR VPWR _1667_/D sky130_fd_sc_hd__nor2_4
X_2588_ _2390_/CLK _2588_/D VGND VGND VPWR VPWR _2349_/A sky130_fd_sc_hd__dfxtp_4
X_1539_ _1466_/A _1482_/Y _1538_/X VGND VGND VPWR VPWR _1539_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_59_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_1_0_m1_clk_local clkbuf_4_1_0_m1_clk_local/A VGND VGND VPWR VPWR _2638_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1890_ _1891_/A _2559_/Q VGND VGND VPWR VPWR _2551_/D sky130_fd_sc_hd__and2_4
X_2373_ _2496_/CLK _2373_/D VGND VGND VPWR VPWR _2373_/Q sky130_fd_sc_hd__dfxtp_4
X_2511_ _2483_/CLK _1954_/X VGND VGND VPWR VPWR DATA_TO_HASH[4] sky130_fd_sc_hd__dfxtp_4
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2442_ _2598_/CLK _2442_/D VGND VGND VPWR VPWR _1960_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_4_13_0_addressalyzerBlock.SPI_CLK clkbuf_3_6_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR _2550_/CLK sky130_fd_sc_hd__clkbuf_1
X_1324_ _1239_/Y VGND VGND VPWR VPWR _1324_/X sky130_fd_sc_hd__buf_2
X_1186_ _1188_/A VGND VGND VPWR VPWR _1187_/A sky130_fd_sc_hd__buf_2
X_1255_ _1254_/X VGND VGND VPWR VPWR _1971_/A sky130_fd_sc_hd__buf_2
XFILLER_33_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE2_2 SCLK_fromHost VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_7_0_m1_clk_local clkbuf_3_7_0_m1_clk_local/A VGND VGND VPWR VPWR clkbuf_3_7_0_m1_clk_local/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1942_ _1938_/A _1942_/B VGND VGND VPWR VPWR _2518_/D sky130_fd_sc_hd__nor2_4
X_1873_ _1838_/A VGND VGND VPWR VPWR _1874_/A sky130_fd_sc_hd__buf_2
X_2356_ _2354_/Y _2322_/A _2355_/Y VGND VGND VPWR VPWR _2652_/D sky130_fd_sc_hd__a21oi_4
X_2425_ _2408_/CLK _2425_/D VGND VGND VPWR VPWR _1937_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_56_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1238_ _2620_/Q _1379_/A _1365_/D _1238_/D VGND VGND VPWR VPWR _1238_/Y sky130_fd_sc_hd__nand4_4
X_1307_ _2636_/Q _1305_/X _1306_/X VGND VGND VPWR VPWR _1307_/X sky130_fd_sc_hd__o21a_4
XFILLER_37_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2287_ _1581_/X _2257_/Y _2278_/A _1927_/Y _2279_/X VGND VGND VPWR VPWR _2412_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2210_ _2207_/Y _2208_/X _2209_/X VGND VGND VPWR VPWR _2210_/Y sky130_fd_sc_hd__a21oi_4
X_2072_ _2071_/Y _2060_/B VGND VGND VPWR VPWR _2072_/Y sky130_fd_sc_hd__nor2_4
XFILLER_46_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2141_ _1503_/Y _2138_/Y _2125_/A _1963_/B _2139_/X VGND VGND VPWR VPWR _2441_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_61_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1925_ _2174_/B VGND VGND VPWR VPWR _1925_/Y sky130_fd_sc_hd__inv_2
X_1856_ _1856_/A _1318_/A _1651_/X VGND VGND VPWR VPWR _1856_/X sky130_fd_sc_hd__and3_4
X_1787_ _1786_/Y VGND VGND VPWR VPWR _1983_/B sky130_fd_sc_hd__buf_2
XFILLER_55_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2339_ _1840_/C _2385_/Q _2102_/A _2338_/X VGND VGND VPWR VPWR _2385_/D sky130_fd_sc_hd__a211o_4
X_2408_ _2408_/CLK _2299_/Y VGND VGND VPWR VPWR ID_toHost sky130_fd_sc_hd__dfxtp_4
XFILLER_25_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1572_ _1569_/X _1556_/A _1860_/B VGND VGND VPWR VPWR _1572_/Y sky130_fd_sc_hd__o21ai_4
X_1641_ _1251_/Y _1640_/X VGND VGND VPWR VPWR _1641_/X sky130_fd_sc_hd__or2_4
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1710_ _1630_/X _1710_/B VGND VGND VPWR VPWR _1710_/Y sky130_fd_sc_hd__nor2_4
X_2124_ _1555_/A VGND VGND VPWR VPWR _2335_/A sky130_fd_sc_hd__buf_2
X_2055_ _1993_/A VGND VGND VPWR VPWR _2055_/X sky130_fd_sc_hd__buf_2
XFILLER_34_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1839_ _2463_/Q VGND VGND VPWR VPWR _1840_/C sky130_fd_sc_hd__inv_2
X_1908_ _2177_/B VGND VGND VPWR VPWR _1908_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1624_ _1623_/Y VGND VGND VPWR VPWR _1624_/X sky130_fd_sc_hd__buf_2
X_1555_ _1555_/A VGND VGND VPWR VPWR _2104_/A sky130_fd_sc_hd__buf_2
X_2107_ _2108_/A _2456_/Q VGND VGND VPWR VPWR _2107_/X sky130_fd_sc_hd__and2_4
XFILLER_39_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1486_ _1486_/A VGND VGND VPWR VPWR _1505_/C sky130_fd_sc_hd__buf_2
X_2038_ _2038_/A _2038_/B VGND VGND VPWR VPWR _2039_/A sky130_fd_sc_hd__nand2_4
XFILLER_22_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1340_ _1335_/C _1318_/B _1335_/D _1329_/X _1339_/X VGND VGND VPWR VPWR _1340_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1271_ _1268_/Y _2010_/B _1271_/C VGND VGND VPWR VPWR _2643_/D sky130_fd_sc_hd__and3_4
XFILLER_51_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1538_ _1466_/Y _1467_/Y _1537_/X _1548_/D _1488_/X VGND VGND VPWR VPWR _1538_/X
+ sky130_fd_sc_hd__o41a_4
X_1469_ _1466_/Y _1467_/Y _1424_/Y _1548_/D VGND VGND VPWR VPWR _1469_/Y sky130_fd_sc_hd__nor4_4
X_2587_ _2606_/CLK _1792_/X VGND VGND VPWR VPWR _1420_/A sky130_fd_sc_hd__dfxtp_4
X_1607_ _2604_/Q _2603_/Q VGND VGND VPWR VPWR _1667_/C sky130_fd_sc_hd__nor2_4
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2510_ _2513_/CLK _1955_/X VGND VGND VPWR VPWR DATA_TO_HASH[3] sky130_fd_sc_hd__dfxtp_4
X_2372_ _2372_/CLK _2371_/Q VGND VGND VPWR VPWR _2373_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1323_ _1323_/A VGND VGND VPWR VPWR _1323_/Y sky130_fd_sc_hd__inv_2
X_2441_ _2598_/CLK _2441_/D VGND VGND VPWR VPWR _2441_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_64_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1185_ _1185_/A VGND VGND VPWR VPWR _1188_/A sky130_fd_sc_hd__inv_2
X_1254_ _1374_/A VGND VGND VPWR VPWR _1254_/X sky130_fd_sc_hd__buf_2
XFILLER_32_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2639_ _2638_/CLK _1290_/Y VGND VGND VPWR VPWR _1224_/A sky130_fd_sc_hd__dfxtp_4
XINSDIODE2_3 _1969_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1872_ _1870_/X DATA_FROM_HASH[6] VGND VGND VPWR VPWR _2565_/D sky130_fd_sc_hd__and2_4
XFILLER_14_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1941_ _1941_/A VGND VGND VPWR VPWR _1942_/B sky130_fd_sc_hd__inv_2
X_2355_ _1676_/B _1187_/A _1213_/X VGND VGND VPWR VPWR _2355_/Y sky130_fd_sc_hd__o21ai_4
X_1306_ _1270_/A VGND VGND VPWR VPWR _1306_/X sky130_fd_sc_hd__buf_2
XFILLER_29_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2286_ _1581_/X _2255_/Y _2278_/A _1925_/Y _2279_/X VGND VGND VPWR VPWR _2413_/D
+ sky130_fd_sc_hd__o32ai_4
X_2424_ _2428_/CLK _2424_/D VGND VGND VPWR VPWR _1847_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_56_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1237_ _1237_/A VGND VGND VPWR VPWR _1238_/D sky130_fd_sc_hd__inv_2
XFILLER_18_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2140_ _2136_/Y _2138_/Y _2120_/X _1960_/Y _2139_/X VGND VGND VPWR VPWR _2442_/D
+ sky130_fd_sc_hd__o32ai_4
X_2071_ _2071_/A VGND VGND VPWR VPWR _2071_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1855_ _1843_/Y _1853_/Y _1854_/X VGND VGND VPWR VPWR _1855_/Y sky130_fd_sc_hd__o21ai_4
X_1924_ _1930_/A _1923_/Y VGND VGND VPWR VPWR _1924_/Y sky130_fd_sc_hd__nor2_4
X_1786_ _2591_/Q VGND VGND VPWR VPWR _1786_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2338_ _2338_/A _1188_/A _1680_/B VGND VGND VPWR VPWR _2338_/X sky130_fd_sc_hd__and3_4
X_2269_ _2268_/Y _2262_/X _2258_/X _1847_/Y _2264_/X VGND VGND VPWR VPWR _2424_/D
+ sky130_fd_sc_hd__o32ai_4
X_2407_ _2408_/CLK _2407_/D VGND VGND VPWR VPWR _2300_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1571_ _1571_/A VGND VGND VPWR VPWR _1860_/B sky130_fd_sc_hd__buf_2
X_1640_ _1613_/Y VGND VGND VPWR VPWR _1640_/X sky130_fd_sc_hd__buf_2
XFILLER_6_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2123_ _2123_/A VGND VGND VPWR VPWR _2125_/A sky130_fd_sc_hd__buf_2
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2054_ _2478_/Q VGND VGND VPWR VPWR _2062_/B sky130_fd_sc_hd__buf_2
XFILLER_34_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1838_ _1838_/A VGND VGND VPWR VPWR _1840_/B sky130_fd_sc_hd__buf_2
X_1907_ _1901_/X _1906_/Y VGND VGND VPWR VPWR _2540_/D sky130_fd_sc_hd__nor2_4
X_1769_ _1486_/A _1764_/Y _1766_/Y _1767_/X _1768_/X VGND VGND VPWR VPWR _1769_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_25_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1485_ _1436_/C VGND VGND VPWR VPWR _1494_/B sky130_fd_sc_hd__buf_2
X_1623_ _2447_/Q VGND VGND VPWR VPWR _1623_/Y sky130_fd_sc_hd__inv_2
X_1554_ _1189_/Y VGND VGND VPWR VPWR _1555_/A sky130_fd_sc_hd__buf_2
.ends

