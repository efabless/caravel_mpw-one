magic
tech sky130A
magscale 12 1
timestamp 1598785497
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
