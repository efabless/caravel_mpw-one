magic
tech sky130A
magscale 1 2
timestamp 1624984707
<< obsli1 >>
rect 1104 17 218868 23375
<< obsm1 >>
rect 14 8 219774 23384
<< metal2 >>
rect 202 22600 258 23800
rect 662 22600 718 23800
rect 1122 22600 1178 23800
rect 1582 22600 1638 23800
rect 2042 22600 2098 23800
rect 2502 22600 2558 23800
rect 3054 22600 3110 23800
rect 3514 22600 3570 23800
rect 3974 22600 4030 23800
rect 4434 22600 4490 23800
rect 4894 22600 4950 23800
rect 5446 22600 5502 23800
rect 5906 22600 5962 23800
rect 6366 22600 6422 23800
rect 6826 22600 6882 23800
rect 7286 22600 7342 23800
rect 7746 22600 7802 23800
rect 8298 22600 8354 23800
rect 8758 22600 8814 23800
rect 9218 22600 9274 23800
rect 9678 22600 9734 23800
rect 10138 22600 10194 23800
rect 10690 22600 10746 23800
rect 11150 22600 11206 23800
rect 11610 22600 11666 23800
rect 12070 22600 12126 23800
rect 12530 22600 12586 23800
rect 13082 22600 13138 23800
rect 13542 22600 13598 23800
rect 14002 22600 14058 23800
rect 14462 22600 14518 23800
rect 14922 22600 14978 23800
rect 15382 22600 15438 23800
rect 15934 22600 15990 23800
rect 16394 22600 16450 23800
rect 16854 22600 16910 23800
rect 17314 22600 17370 23800
rect 17774 22600 17830 23800
rect 18326 22600 18382 23800
rect 18786 22600 18842 23800
rect 19246 22600 19302 23800
rect 19706 22600 19762 23800
rect 20166 22600 20222 23800
rect 20718 22600 20774 23800
rect 21178 22600 21234 23800
rect 21638 22600 21694 23800
rect 22098 22600 22154 23800
rect 22558 22600 22614 23800
rect 23018 22600 23074 23800
rect 23570 22600 23626 23800
rect 24030 22600 24086 23800
rect 24490 22600 24546 23800
rect 24950 22600 25006 23800
rect 25410 22600 25466 23800
rect 25962 22600 26018 23800
rect 26422 22600 26478 23800
rect 26882 22600 26938 23800
rect 27342 22600 27398 23800
rect 27802 22600 27858 23800
rect 28354 22600 28410 23800
rect 28814 22600 28870 23800
rect 29274 22600 29330 23800
rect 29734 22600 29790 23800
rect 30194 22600 30250 23800
rect 30654 22600 30710 23800
rect 31206 22600 31262 23800
rect 31666 22600 31722 23800
rect 32126 22600 32182 23800
rect 32586 22600 32642 23800
rect 33046 22600 33102 23800
rect 33598 22600 33654 23800
rect 34058 22600 34114 23800
rect 34518 22600 34574 23800
rect 34978 22600 35034 23800
rect 35438 22600 35494 23800
rect 35898 22600 35954 23800
rect 36450 22600 36506 23800
rect 36910 22600 36966 23800
rect 37370 22600 37426 23800
rect 37830 22600 37886 23800
rect 38290 22600 38346 23800
rect 38842 22600 38898 23800
rect 39302 22600 39358 23800
rect 39762 22600 39818 23800
rect 40222 22600 40278 23800
rect 40682 22600 40738 23800
rect 41234 22600 41290 23800
rect 41694 22600 41750 23800
rect 42154 22600 42210 23800
rect 42614 22600 42670 23800
rect 43074 22600 43130 23800
rect 43534 22600 43590 23800
rect 44086 22600 44142 23800
rect 44546 22600 44602 23800
rect 45006 22600 45062 23800
rect 45466 22600 45522 23800
rect 45926 22600 45982 23800
rect 46478 22600 46534 23800
rect 46938 22600 46994 23800
rect 47398 22600 47454 23800
rect 47858 22600 47914 23800
rect 48318 22600 48374 23800
rect 48870 22600 48926 23800
rect 49330 22600 49386 23800
rect 49790 22600 49846 23800
rect 50250 22600 50306 23800
rect 50710 22600 50766 23800
rect 51170 22600 51226 23800
rect 51722 22600 51778 23800
rect 52182 22600 52238 23800
rect 52642 22600 52698 23800
rect 53102 22600 53158 23800
rect 53562 22600 53618 23800
rect 54114 22600 54170 23800
rect 54574 22600 54630 23800
rect 55034 22600 55090 23800
rect 55494 22600 55550 23800
rect 55954 22600 56010 23800
rect 56506 22600 56562 23800
rect 56966 22600 57022 23800
rect 57426 22600 57482 23800
rect 57886 22600 57942 23800
rect 58346 22600 58402 23800
rect 58806 22600 58862 23800
rect 59358 22600 59414 23800
rect 59818 22600 59874 23800
rect 60278 22600 60334 23800
rect 60738 22600 60794 23800
rect 61198 22600 61254 23800
rect 61750 22600 61806 23800
rect 62210 22600 62266 23800
rect 62670 22600 62726 23800
rect 63130 22600 63186 23800
rect 63590 22600 63646 23800
rect 64050 22600 64106 23800
rect 64602 22600 64658 23800
rect 65062 22600 65118 23800
rect 65522 22600 65578 23800
rect 65982 22600 66038 23800
rect 66442 22600 66498 23800
rect 66994 22600 67050 23800
rect 67454 22600 67510 23800
rect 67914 22600 67970 23800
rect 68374 22600 68430 23800
rect 68834 22600 68890 23800
rect 69386 22600 69442 23800
rect 69846 22600 69902 23800
rect 70306 22600 70362 23800
rect 70766 22600 70822 23800
rect 71226 22600 71282 23800
rect 71686 22600 71742 23800
rect 72238 22600 72294 23800
rect 72698 22600 72754 23800
rect 73158 22600 73214 23800
rect 73618 22600 73674 23800
rect 74078 22600 74134 23800
rect 74630 22600 74686 23800
rect 75090 22600 75146 23800
rect 75550 22600 75606 23800
rect 76010 22600 76066 23800
rect 76470 22600 76526 23800
rect 77022 22600 77078 23800
rect 77482 22600 77538 23800
rect 77942 22600 77998 23800
rect 78402 22600 78458 23800
rect 78862 22600 78918 23800
rect 79322 22600 79378 23800
rect 79874 22600 79930 23800
rect 80334 22600 80390 23800
rect 80794 22600 80850 23800
rect 81254 22600 81310 23800
rect 81714 22600 81770 23800
rect 82266 22600 82322 23800
rect 82726 22600 82782 23800
rect 83186 22600 83242 23800
rect 83646 22600 83702 23800
rect 84106 22600 84162 23800
rect 84658 22600 84714 23800
rect 85118 22600 85174 23800
rect 85578 22600 85634 23800
rect 86038 22600 86094 23800
rect 86498 22600 86554 23800
rect 86958 22600 87014 23800
rect 87510 22600 87566 23800
rect 87970 22600 88026 23800
rect 88430 22600 88486 23800
rect 88890 22600 88946 23800
rect 89350 22600 89406 23800
rect 89902 22600 89958 23800
rect 90362 22600 90418 23800
rect 90822 22600 90878 23800
rect 91282 22600 91338 23800
rect 91742 22600 91798 23800
rect 92294 22600 92350 23800
rect 92754 22600 92810 23800
rect 93214 22600 93270 23800
rect 93674 22600 93730 23800
rect 94134 22600 94190 23800
rect 94594 22600 94650 23800
rect 95146 22600 95202 23800
rect 95606 22600 95662 23800
rect 96066 22600 96122 23800
rect 96526 22600 96582 23800
rect 96986 22600 97042 23800
rect 97538 22600 97594 23800
rect 97998 22600 98054 23800
rect 98458 22600 98514 23800
rect 98918 22600 98974 23800
rect 99378 22600 99434 23800
rect 99838 22600 99894 23800
rect 100390 22600 100446 23800
rect 100850 22600 100906 23800
rect 101310 22600 101366 23800
rect 101770 22600 101826 23800
rect 102230 22600 102286 23800
rect 102782 22600 102838 23800
rect 103242 22600 103298 23800
rect 103702 22600 103758 23800
rect 104162 22600 104218 23800
rect 104622 22600 104678 23800
rect 105174 22600 105230 23800
rect 105634 22600 105690 23800
rect 106094 22600 106150 23800
rect 106554 22600 106610 23800
rect 107014 22600 107070 23800
rect 107474 22600 107530 23800
rect 108026 22600 108082 23800
rect 108486 22600 108542 23800
rect 108946 22600 109002 23800
rect 109406 22600 109462 23800
rect 109866 22600 109922 23800
rect 110418 22600 110474 23800
rect 110878 22600 110934 23800
rect 111338 22600 111394 23800
rect 111798 22600 111854 23800
rect 112258 22600 112314 23800
rect 112810 22600 112866 23800
rect 113270 22600 113326 23800
rect 113730 22600 113786 23800
rect 114190 22600 114246 23800
rect 114650 22600 114706 23800
rect 115110 22600 115166 23800
rect 115662 22600 115718 23800
rect 116122 22600 116178 23800
rect 116582 22600 116638 23800
rect 117042 22600 117098 23800
rect 117502 22600 117558 23800
rect 118054 22600 118110 23800
rect 118514 22600 118570 23800
rect 118974 22600 119030 23800
rect 119434 22600 119490 23800
rect 119894 22600 119950 23800
rect 120446 22600 120502 23800
rect 120906 22600 120962 23800
rect 121366 22600 121422 23800
rect 121826 22600 121882 23800
rect 122286 22600 122342 23800
rect 122746 22600 122802 23800
rect 123298 22600 123354 23800
rect 123758 22600 123814 23800
rect 124218 22600 124274 23800
rect 124678 22600 124734 23800
rect 125138 22600 125194 23800
rect 125690 22600 125746 23800
rect 126150 22600 126206 23800
rect 126610 22600 126666 23800
rect 127070 22600 127126 23800
rect 127530 22600 127586 23800
rect 127990 22600 128046 23800
rect 128542 22600 128598 23800
rect 129002 22600 129058 23800
rect 129462 22600 129518 23800
rect 129922 22600 129978 23800
rect 130382 22600 130438 23800
rect 130934 22600 130990 23800
rect 131394 22600 131450 23800
rect 131854 22600 131910 23800
rect 132314 22600 132370 23800
rect 132774 22600 132830 23800
rect 133326 22600 133382 23800
rect 133786 22600 133842 23800
rect 134246 22600 134302 23800
rect 134706 22600 134762 23800
rect 135166 22600 135222 23800
rect 135626 22600 135682 23800
rect 136178 22600 136234 23800
rect 136638 22600 136694 23800
rect 137098 22600 137154 23800
rect 137558 22600 137614 23800
rect 138018 22600 138074 23800
rect 138570 22600 138626 23800
rect 139030 22600 139086 23800
rect 139490 22600 139546 23800
rect 139950 22600 140006 23800
rect 140410 22600 140466 23800
rect 140962 22600 141018 23800
rect 141422 22600 141478 23800
rect 141882 22600 141938 23800
rect 142342 22600 142398 23800
rect 142802 22600 142858 23800
rect 143262 22600 143318 23800
rect 143814 22600 143870 23800
rect 144274 22600 144330 23800
rect 144734 22600 144790 23800
rect 145194 22600 145250 23800
rect 145654 22600 145710 23800
rect 146206 22600 146262 23800
rect 146666 22600 146722 23800
rect 147126 22600 147182 23800
rect 147586 22600 147642 23800
rect 148046 22600 148102 23800
rect 148598 22600 148654 23800
rect 149058 22600 149114 23800
rect 149518 22600 149574 23800
rect 149978 22600 150034 23800
rect 150438 22600 150494 23800
rect 150898 22600 150954 23800
rect 151450 22600 151506 23800
rect 151910 22600 151966 23800
rect 152370 22600 152426 23800
rect 152830 22600 152886 23800
rect 153290 22600 153346 23800
rect 153842 22600 153898 23800
rect 154302 22600 154358 23800
rect 154762 22600 154818 23800
rect 155222 22600 155278 23800
rect 155682 22600 155738 23800
rect 156234 22600 156290 23800
rect 156694 22600 156750 23800
rect 157154 22600 157210 23800
rect 157614 22600 157670 23800
rect 158074 22600 158130 23800
rect 158534 22600 158590 23800
rect 159086 22600 159142 23800
rect 159546 22600 159602 23800
rect 160006 22600 160062 23800
rect 160466 22600 160522 23800
rect 160926 22600 160982 23800
rect 161478 22600 161534 23800
rect 161938 22600 161994 23800
rect 162398 22600 162454 23800
rect 162858 22600 162914 23800
rect 163318 22600 163374 23800
rect 163778 22600 163834 23800
rect 164330 22600 164386 23800
rect 164790 22600 164846 23800
rect 165250 22600 165306 23800
rect 165710 22600 165766 23800
rect 166170 22600 166226 23800
rect 166722 22600 166778 23800
rect 167182 22600 167238 23800
rect 167642 22600 167698 23800
rect 168102 22600 168158 23800
rect 168562 22600 168618 23800
rect 169114 22600 169170 23800
rect 169574 22600 169630 23800
rect 170034 22600 170090 23800
rect 170494 22600 170550 23800
rect 170954 22600 171010 23800
rect 171414 22600 171470 23800
rect 171966 22600 172022 23800
rect 172426 22600 172482 23800
rect 172886 22600 172942 23800
rect 173346 22600 173402 23800
rect 173806 22600 173862 23800
rect 174358 22600 174414 23800
rect 174818 22600 174874 23800
rect 175278 22600 175334 23800
rect 175738 22600 175794 23800
rect 176198 22600 176254 23800
rect 176750 22600 176806 23800
rect 177210 22600 177266 23800
rect 177670 22600 177726 23800
rect 178130 22600 178186 23800
rect 178590 22600 178646 23800
rect 179050 22600 179106 23800
rect 179602 22600 179658 23800
rect 180062 22600 180118 23800
rect 180522 22600 180578 23800
rect 180982 22600 181038 23800
rect 181442 22600 181498 23800
rect 181994 22600 182050 23800
rect 182454 22600 182510 23800
rect 182914 22600 182970 23800
rect 183374 22600 183430 23800
rect 183834 22600 183890 23800
rect 184386 22600 184442 23800
rect 184846 22600 184902 23800
rect 185306 22600 185362 23800
rect 185766 22600 185822 23800
rect 186226 22600 186282 23800
rect 186686 22600 186742 23800
rect 187238 22600 187294 23800
rect 187698 22600 187754 23800
rect 188158 22600 188214 23800
rect 188618 22600 188674 23800
rect 189078 22600 189134 23800
rect 189630 22600 189686 23800
rect 190090 22600 190146 23800
rect 190550 22600 190606 23800
rect 191010 22600 191066 23800
rect 191470 22600 191526 23800
rect 191930 22600 191986 23800
rect 192482 22600 192538 23800
rect 192942 22600 192998 23800
rect 193402 22600 193458 23800
rect 193862 22600 193918 23800
rect 194322 22600 194378 23800
rect 194874 22600 194930 23800
rect 195334 22600 195390 23800
rect 195794 22600 195850 23800
rect 196254 22600 196310 23800
rect 196714 22600 196770 23800
rect 197266 22600 197322 23800
rect 197726 22600 197782 23800
rect 198186 22600 198242 23800
rect 198646 22600 198702 23800
rect 199106 22600 199162 23800
rect 199566 22600 199622 23800
rect 200118 22600 200174 23800
rect 200578 22600 200634 23800
rect 201038 22600 201094 23800
rect 201498 22600 201554 23800
rect 201958 22600 202014 23800
rect 202510 22600 202566 23800
rect 202970 22600 203026 23800
rect 203430 22600 203486 23800
rect 203890 22600 203946 23800
rect 204350 22600 204406 23800
rect 204902 22600 204958 23800
rect 205362 22600 205418 23800
rect 205822 22600 205878 23800
rect 206282 22600 206338 23800
rect 206742 22600 206798 23800
rect 207202 22600 207258 23800
rect 207754 22600 207810 23800
rect 208214 22600 208270 23800
rect 208674 22600 208730 23800
rect 209134 22600 209190 23800
rect 209594 22600 209650 23800
rect 210146 22600 210202 23800
rect 210606 22600 210662 23800
rect 211066 22600 211122 23800
rect 211526 22600 211582 23800
rect 211986 22600 212042 23800
rect 212538 22600 212594 23800
rect 212998 22600 213054 23800
rect 213458 22600 213514 23800
rect 213918 22600 213974 23800
rect 214378 22600 214434 23800
rect 214838 22600 214894 23800
rect 215390 22600 215446 23800
rect 215850 22600 215906 23800
rect 216310 22600 216366 23800
rect 216770 22600 216826 23800
rect 217230 22600 217286 23800
rect 217782 22600 217838 23800
rect 218242 22600 218298 23800
rect 218702 22600 218758 23800
rect 219162 22600 219218 23800
rect 219622 22600 219678 23800
rect 202 -400 258 800
rect 570 -400 626 800
rect 938 -400 994 800
rect 1306 -400 1362 800
rect 1674 -400 1730 800
rect 2042 -400 2098 800
rect 2410 -400 2466 800
rect 2778 -400 2834 800
rect 3146 -400 3202 800
rect 3514 -400 3570 800
rect 3974 -400 4030 800
rect 4342 -400 4398 800
rect 4710 -400 4766 800
rect 5078 -400 5134 800
rect 5446 -400 5502 800
rect 5814 -400 5870 800
rect 6182 -400 6238 800
rect 6550 -400 6606 800
rect 6918 -400 6974 800
rect 7286 -400 7342 800
rect 7746 -400 7802 800
rect 8114 -400 8170 800
rect 8482 -400 8538 800
rect 8850 -400 8906 800
rect 9218 -400 9274 800
rect 9586 -400 9642 800
rect 9954 -400 10010 800
rect 10322 -400 10378 800
rect 10690 -400 10746 800
rect 11058 -400 11114 800
rect 11518 -400 11574 800
rect 11886 -400 11942 800
rect 12254 -400 12310 800
rect 12622 -400 12678 800
rect 12990 -400 13046 800
rect 13358 -400 13414 800
rect 13726 -400 13782 800
rect 14094 -400 14150 800
rect 14462 -400 14518 800
rect 14830 -400 14886 800
rect 15290 -400 15346 800
rect 15658 -400 15714 800
rect 16026 -400 16082 800
rect 16394 -400 16450 800
rect 16762 -400 16818 800
rect 17130 -400 17186 800
rect 17498 -400 17554 800
rect 17866 -400 17922 800
rect 18234 -400 18290 800
rect 18602 -400 18658 800
rect 19062 -400 19118 800
rect 19430 -400 19486 800
rect 19798 -400 19854 800
rect 20166 -400 20222 800
rect 20534 -400 20590 800
rect 20902 -400 20958 800
rect 21270 -400 21326 800
rect 21638 -400 21694 800
rect 22006 -400 22062 800
rect 22374 -400 22430 800
rect 22834 -400 22890 800
rect 23202 -400 23258 800
rect 23570 -400 23626 800
rect 23938 -400 23994 800
rect 24306 -400 24362 800
rect 24674 -400 24730 800
rect 25042 -400 25098 800
rect 25410 -400 25466 800
rect 25778 -400 25834 800
rect 26146 -400 26202 800
rect 26606 -400 26662 800
rect 26974 -400 27030 800
rect 27342 -400 27398 800
rect 27710 -400 27766 800
rect 28078 -400 28134 800
rect 28446 -400 28502 800
rect 28814 -400 28870 800
rect 29182 -400 29238 800
rect 29550 -400 29606 800
rect 29918 -400 29974 800
rect 30378 -400 30434 800
rect 30746 -400 30802 800
rect 31114 -400 31170 800
rect 31482 -400 31538 800
rect 31850 -400 31906 800
rect 32218 -400 32274 800
rect 32586 -400 32642 800
rect 32954 -400 33010 800
rect 33322 -400 33378 800
rect 33782 -400 33838 800
rect 34150 -400 34206 800
rect 34518 -400 34574 800
rect 34886 -400 34942 800
rect 35254 -400 35310 800
rect 35622 -400 35678 800
rect 35990 -400 36046 800
rect 36358 -400 36414 800
rect 36726 -400 36782 800
rect 37094 -400 37150 800
rect 37554 -400 37610 800
rect 37922 -400 37978 800
rect 38290 -400 38346 800
rect 38658 -400 38714 800
rect 39026 -400 39082 800
rect 39394 -400 39450 800
rect 39762 -400 39818 800
rect 40130 -400 40186 800
rect 40498 -400 40554 800
rect 40866 -400 40922 800
rect 41326 -400 41382 800
rect 41694 -400 41750 800
rect 42062 -400 42118 800
rect 42430 -400 42486 800
rect 42798 -400 42854 800
rect 43166 -400 43222 800
rect 43534 -400 43590 800
rect 43902 -400 43958 800
rect 44270 -400 44326 800
rect 44638 -400 44694 800
rect 45098 -400 45154 800
rect 45466 -400 45522 800
rect 45834 -400 45890 800
rect 46202 -400 46258 800
rect 46570 -400 46626 800
rect 46938 -400 46994 800
rect 47306 -400 47362 800
rect 47674 -400 47730 800
rect 48042 -400 48098 800
rect 48410 -400 48466 800
rect 48870 -400 48926 800
rect 49238 -400 49294 800
rect 49606 -400 49662 800
rect 49974 -400 50030 800
rect 50342 -400 50398 800
rect 50710 -400 50766 800
rect 51078 -400 51134 800
rect 51446 -400 51502 800
rect 51814 -400 51870 800
rect 52182 -400 52238 800
rect 52642 -400 52698 800
rect 53010 -400 53066 800
rect 53378 -400 53434 800
rect 53746 -400 53802 800
rect 54114 -400 54170 800
rect 54482 -400 54538 800
rect 54850 -400 54906 800
rect 55218 -400 55274 800
rect 55586 -400 55642 800
rect 55954 -400 56010 800
rect 56414 -400 56470 800
rect 56782 -400 56838 800
rect 57150 -400 57206 800
rect 57518 -400 57574 800
rect 57886 -400 57942 800
rect 58254 -400 58310 800
rect 58622 -400 58678 800
rect 58990 -400 59046 800
rect 59358 -400 59414 800
rect 59726 -400 59782 800
rect 60186 -400 60242 800
rect 60554 -400 60610 800
rect 60922 -400 60978 800
rect 61290 -400 61346 800
rect 61658 -400 61714 800
rect 62026 -400 62082 800
rect 62394 -400 62450 800
rect 62762 -400 62818 800
rect 63130 -400 63186 800
rect 63590 -400 63646 800
rect 63958 -400 64014 800
rect 64326 -400 64382 800
rect 64694 -400 64750 800
rect 65062 -400 65118 800
rect 65430 -400 65486 800
rect 65798 -400 65854 800
rect 66166 -400 66222 800
rect 66534 -400 66590 800
rect 66902 -400 66958 800
rect 67362 -400 67418 800
rect 67730 -400 67786 800
rect 68098 -400 68154 800
rect 68466 -400 68522 800
rect 68834 -400 68890 800
rect 69202 -400 69258 800
rect 69570 -400 69626 800
rect 69938 -400 69994 800
rect 70306 -400 70362 800
rect 70674 -400 70730 800
rect 71134 -400 71190 800
rect 71502 -400 71558 800
rect 71870 -400 71926 800
rect 72238 -400 72294 800
rect 72606 -400 72662 800
rect 72974 -400 73030 800
rect 73342 -400 73398 800
rect 73710 -400 73766 800
rect 74078 -400 74134 800
rect 74446 -400 74502 800
rect 74906 -400 74962 800
rect 75274 -400 75330 800
rect 75642 -400 75698 800
rect 76010 -400 76066 800
rect 76378 -400 76434 800
rect 76746 -400 76802 800
rect 77114 -400 77170 800
rect 77482 -400 77538 800
rect 77850 -400 77906 800
rect 78218 -400 78274 800
rect 78678 -400 78734 800
rect 79046 -400 79102 800
rect 79414 -400 79470 800
rect 79782 -400 79838 800
rect 80150 -400 80206 800
rect 80518 -400 80574 800
rect 80886 -400 80942 800
rect 81254 -400 81310 800
rect 81622 -400 81678 800
rect 81990 -400 82046 800
rect 82450 -400 82506 800
rect 82818 -400 82874 800
rect 83186 -400 83242 800
rect 83554 -400 83610 800
rect 83922 -400 83978 800
rect 84290 -400 84346 800
rect 84658 -400 84714 800
rect 85026 -400 85082 800
rect 85394 -400 85450 800
rect 85762 -400 85818 800
rect 86222 -400 86278 800
rect 86590 -400 86646 800
rect 86958 -400 87014 800
rect 87326 -400 87382 800
rect 87694 -400 87750 800
rect 88062 -400 88118 800
rect 88430 -400 88486 800
rect 88798 -400 88854 800
rect 89166 -400 89222 800
rect 89534 -400 89590 800
rect 89994 -400 90050 800
rect 90362 -400 90418 800
rect 90730 -400 90786 800
rect 91098 -400 91154 800
rect 91466 -400 91522 800
rect 91834 -400 91890 800
rect 92202 -400 92258 800
rect 92570 -400 92626 800
rect 92938 -400 92994 800
rect 93306 -400 93362 800
rect 93766 -400 93822 800
rect 94134 -400 94190 800
rect 94502 -400 94558 800
rect 94870 -400 94926 800
rect 95238 -400 95294 800
rect 95606 -400 95662 800
rect 95974 -400 96030 800
rect 96342 -400 96398 800
rect 96710 -400 96766 800
rect 97170 -400 97226 800
rect 97538 -400 97594 800
rect 97906 -400 97962 800
rect 98274 -400 98330 800
rect 98642 -400 98698 800
rect 99010 -400 99066 800
rect 99378 -400 99434 800
rect 99746 -400 99802 800
rect 100114 -400 100170 800
rect 100482 -400 100538 800
rect 100942 -400 100998 800
rect 101310 -400 101366 800
rect 101678 -400 101734 800
rect 102046 -400 102102 800
rect 102414 -400 102470 800
rect 102782 -400 102838 800
rect 103150 -400 103206 800
rect 103518 -400 103574 800
rect 103886 -400 103942 800
rect 104254 -400 104310 800
rect 104714 -400 104770 800
rect 105082 -400 105138 800
rect 105450 -400 105506 800
rect 105818 -400 105874 800
rect 106186 -400 106242 800
rect 106554 -400 106610 800
rect 106922 -400 106978 800
rect 107290 -400 107346 800
rect 107658 -400 107714 800
rect 108026 -400 108082 800
rect 108486 -400 108542 800
rect 108854 -400 108910 800
rect 109222 -400 109278 800
rect 109590 -400 109646 800
rect 109958 -400 110014 800
rect 110326 -400 110382 800
rect 110694 -400 110750 800
rect 111062 -400 111118 800
rect 111430 -400 111486 800
rect 111798 -400 111854 800
rect 112258 -400 112314 800
rect 112626 -400 112682 800
rect 112994 -400 113050 800
rect 113362 -400 113418 800
rect 113730 -400 113786 800
rect 114098 -400 114154 800
rect 114466 -400 114522 800
rect 114834 -400 114890 800
rect 115202 -400 115258 800
rect 115570 -400 115626 800
rect 116030 -400 116086 800
rect 116398 -400 116454 800
rect 116766 -400 116822 800
rect 117134 -400 117190 800
rect 117502 -400 117558 800
rect 117870 -400 117926 800
rect 118238 -400 118294 800
rect 118606 -400 118662 800
rect 118974 -400 119030 800
rect 119342 -400 119398 800
rect 119802 -400 119858 800
rect 120170 -400 120226 800
rect 120538 -400 120594 800
rect 120906 -400 120962 800
rect 121274 -400 121330 800
rect 121642 -400 121698 800
rect 122010 -400 122066 800
rect 122378 -400 122434 800
rect 122746 -400 122802 800
rect 123114 -400 123170 800
rect 123574 -400 123630 800
rect 123942 -400 123998 800
rect 124310 -400 124366 800
rect 124678 -400 124734 800
rect 125046 -400 125102 800
rect 125414 -400 125470 800
rect 125782 -400 125838 800
rect 126150 -400 126206 800
rect 126518 -400 126574 800
rect 126978 -400 127034 800
rect 127346 -400 127402 800
rect 127714 -400 127770 800
rect 128082 -400 128138 800
rect 128450 -400 128506 800
rect 128818 -400 128874 800
rect 129186 -400 129242 800
rect 129554 -400 129610 800
rect 129922 -400 129978 800
rect 130290 -400 130346 800
rect 130750 -400 130806 800
rect 131118 -400 131174 800
rect 131486 -400 131542 800
rect 131854 -400 131910 800
rect 132222 -400 132278 800
rect 132590 -400 132646 800
rect 132958 -400 133014 800
rect 133326 -400 133382 800
rect 133694 -400 133750 800
rect 134062 -400 134118 800
rect 134522 -400 134578 800
rect 134890 -400 134946 800
rect 135258 -400 135314 800
rect 135626 -400 135682 800
rect 135994 -400 136050 800
rect 136362 -400 136418 800
rect 136730 -400 136786 800
rect 137098 -400 137154 800
rect 137466 -400 137522 800
rect 137834 -400 137890 800
rect 138294 -400 138350 800
rect 138662 -400 138718 800
rect 139030 -400 139086 800
rect 139398 -400 139454 800
rect 139766 -400 139822 800
rect 140134 -400 140190 800
rect 140502 -400 140558 800
rect 140870 -400 140926 800
rect 141238 -400 141294 800
rect 141606 -400 141662 800
rect 142066 -400 142122 800
rect 142434 -400 142490 800
rect 142802 -400 142858 800
rect 143170 -400 143226 800
rect 143538 -400 143594 800
rect 143906 -400 143962 800
rect 144274 -400 144330 800
rect 144642 -400 144698 800
rect 145010 -400 145066 800
rect 145378 -400 145434 800
rect 145838 -400 145894 800
rect 146206 -400 146262 800
rect 146574 -400 146630 800
rect 146942 -400 146998 800
rect 147310 -400 147366 800
rect 147678 -400 147734 800
rect 148046 -400 148102 800
rect 148414 -400 148470 800
rect 148782 -400 148838 800
rect 149150 -400 149206 800
rect 149610 -400 149666 800
rect 149978 -400 150034 800
rect 150346 -400 150402 800
rect 150714 -400 150770 800
rect 151082 -400 151138 800
rect 151450 -400 151506 800
rect 151818 -400 151874 800
rect 152186 -400 152242 800
rect 152554 -400 152610 800
rect 152922 -400 152978 800
rect 153382 -400 153438 800
rect 153750 -400 153806 800
rect 154118 -400 154174 800
rect 154486 -400 154542 800
rect 154854 -400 154910 800
rect 155222 -400 155278 800
rect 155590 -400 155646 800
rect 155958 -400 156014 800
rect 156326 -400 156382 800
rect 156694 -400 156750 800
rect 157154 -400 157210 800
rect 157522 -400 157578 800
rect 157890 -400 157946 800
rect 158258 -400 158314 800
rect 158626 -400 158682 800
rect 158994 -400 159050 800
rect 159362 -400 159418 800
rect 159730 -400 159786 800
rect 160098 -400 160154 800
rect 160558 -400 160614 800
rect 160926 -400 160982 800
rect 161294 -400 161350 800
rect 161662 -400 161718 800
rect 162030 -400 162086 800
rect 162398 -400 162454 800
rect 162766 -400 162822 800
rect 163134 -400 163190 800
rect 163502 -400 163558 800
rect 163870 -400 163926 800
rect 164330 -400 164386 800
rect 164698 -400 164754 800
rect 165066 -400 165122 800
rect 165434 -400 165490 800
rect 165802 -400 165858 800
rect 166170 -400 166226 800
rect 166538 -400 166594 800
rect 166906 -400 166962 800
rect 167274 -400 167330 800
rect 167642 -400 167698 800
rect 168102 -400 168158 800
rect 168470 -400 168526 800
rect 168838 -400 168894 800
rect 169206 -400 169262 800
rect 169574 -400 169630 800
rect 169942 -400 169998 800
rect 170310 -400 170366 800
rect 170678 -400 170734 800
rect 171046 -400 171102 800
rect 171414 -400 171470 800
rect 171874 -400 171930 800
rect 172242 -400 172298 800
rect 172610 -400 172666 800
rect 172978 -400 173034 800
rect 173346 -400 173402 800
rect 173714 -400 173770 800
rect 174082 -400 174138 800
rect 174450 -400 174506 800
rect 174818 -400 174874 800
rect 175186 -400 175242 800
rect 175646 -400 175702 800
rect 176014 -400 176070 800
rect 176382 -400 176438 800
rect 176750 -400 176806 800
rect 177118 -400 177174 800
rect 177486 -400 177542 800
rect 177854 -400 177910 800
rect 178222 -400 178278 800
rect 178590 -400 178646 800
rect 178958 -400 179014 800
rect 179418 -400 179474 800
rect 179786 -400 179842 800
rect 180154 -400 180210 800
rect 180522 -400 180578 800
rect 180890 -400 180946 800
rect 181258 -400 181314 800
rect 181626 -400 181682 800
rect 181994 -400 182050 800
rect 182362 -400 182418 800
rect 182730 -400 182786 800
rect 183190 -400 183246 800
rect 183558 -400 183614 800
rect 183926 -400 183982 800
rect 184294 -400 184350 800
rect 184662 -400 184718 800
rect 185030 -400 185086 800
rect 185398 -400 185454 800
rect 185766 -400 185822 800
rect 186134 -400 186190 800
rect 186502 -400 186558 800
rect 186962 -400 187018 800
rect 187330 -400 187386 800
rect 187698 -400 187754 800
rect 188066 -400 188122 800
rect 188434 -400 188490 800
rect 188802 -400 188858 800
rect 189170 -400 189226 800
rect 189538 -400 189594 800
rect 189906 -400 189962 800
rect 190366 -400 190422 800
rect 190734 -400 190790 800
rect 191102 -400 191158 800
rect 191470 -400 191526 800
rect 191838 -400 191894 800
rect 192206 -400 192262 800
rect 192574 -400 192630 800
rect 192942 -400 192998 800
rect 193310 -400 193366 800
rect 193678 -400 193734 800
rect 194138 -400 194194 800
rect 194506 -400 194562 800
rect 194874 -400 194930 800
rect 195242 -400 195298 800
rect 195610 -400 195666 800
rect 195978 -400 196034 800
rect 196346 -400 196402 800
rect 196714 -400 196770 800
rect 197082 -400 197138 800
rect 197450 -400 197506 800
rect 197910 -400 197966 800
rect 198278 -400 198334 800
rect 198646 -400 198702 800
rect 199014 -400 199070 800
rect 199382 -400 199438 800
rect 199750 -400 199806 800
rect 200118 -400 200174 800
rect 200486 -400 200542 800
rect 200854 -400 200910 800
rect 201222 -400 201278 800
rect 201682 -400 201738 800
rect 202050 -400 202106 800
rect 202418 -400 202474 800
rect 202786 -400 202842 800
rect 203154 -400 203210 800
rect 203522 -400 203578 800
rect 203890 -400 203946 800
rect 204258 -400 204314 800
rect 204626 -400 204682 800
rect 204994 -400 205050 800
rect 205454 -400 205510 800
rect 205822 -400 205878 800
rect 206190 -400 206246 800
rect 206558 -400 206614 800
rect 206926 -400 206982 800
rect 207294 -400 207350 800
rect 207662 -400 207718 800
rect 208030 -400 208086 800
rect 208398 -400 208454 800
rect 208766 -400 208822 800
rect 209226 -400 209282 800
rect 209594 -400 209650 800
rect 209962 -400 210018 800
rect 210330 -400 210386 800
rect 210698 -400 210754 800
rect 211066 -400 211122 800
rect 211434 -400 211490 800
rect 211802 -400 211858 800
rect 212170 -400 212226 800
rect 212538 -400 212594 800
rect 212998 -400 213054 800
rect 213366 -400 213422 800
rect 213734 -400 213790 800
rect 214102 -400 214158 800
rect 214470 -400 214526 800
rect 214838 -400 214894 800
rect 215206 -400 215262 800
rect 215574 -400 215630 800
rect 215942 -400 215998 800
rect 216310 -400 216366 800
rect 216770 -400 216826 800
rect 217138 -400 217194 800
rect 217506 -400 217562 800
rect 217874 -400 217930 800
rect 218242 -400 218298 800
rect 218610 -400 218666 800
rect 218978 -400 219034 800
rect 219346 -400 219402 800
rect 219714 -400 219770 800
<< obsm2 >>
rect 20 22544 146 23390
rect 314 22544 606 23390
rect 774 22544 1066 23390
rect 1234 22544 1526 23390
rect 1694 22544 1986 23390
rect 2154 22544 2446 23390
rect 2614 22544 2998 23390
rect 3166 22544 3458 23390
rect 3626 22544 3918 23390
rect 4086 22544 4378 23390
rect 4546 22544 4838 23390
rect 5006 22544 5390 23390
rect 5558 22544 5850 23390
rect 6018 22544 6310 23390
rect 6478 22544 6770 23390
rect 6938 22544 7230 23390
rect 7398 22544 7690 23390
rect 7858 22544 8242 23390
rect 8410 22544 8702 23390
rect 8870 22544 9162 23390
rect 9330 22544 9622 23390
rect 9790 22544 10082 23390
rect 10250 22544 10634 23390
rect 10802 22544 11094 23390
rect 11262 22544 11554 23390
rect 11722 22544 12014 23390
rect 12182 22544 12474 23390
rect 12642 22544 13026 23390
rect 13194 22544 13486 23390
rect 13654 22544 13946 23390
rect 14114 22544 14406 23390
rect 14574 22544 14866 23390
rect 15034 22544 15326 23390
rect 15494 22544 15878 23390
rect 16046 22544 16338 23390
rect 16506 22544 16798 23390
rect 16966 22544 17258 23390
rect 17426 22544 17718 23390
rect 17886 22544 18270 23390
rect 18438 22544 18730 23390
rect 18898 22544 19190 23390
rect 19358 22544 19650 23390
rect 19818 22544 20110 23390
rect 20278 22544 20662 23390
rect 20830 22544 21122 23390
rect 21290 22544 21582 23390
rect 21750 22544 22042 23390
rect 22210 22544 22502 23390
rect 22670 22544 22962 23390
rect 23130 22544 23514 23390
rect 23682 22544 23974 23390
rect 24142 22544 24434 23390
rect 24602 22544 24894 23390
rect 25062 22544 25354 23390
rect 25522 22544 25906 23390
rect 26074 22544 26366 23390
rect 26534 22544 26826 23390
rect 26994 22544 27286 23390
rect 27454 22544 27746 23390
rect 27914 22544 28298 23390
rect 28466 22544 28758 23390
rect 28926 22544 29218 23390
rect 29386 22544 29678 23390
rect 29846 22544 30138 23390
rect 30306 22544 30598 23390
rect 30766 22544 31150 23390
rect 31318 22544 31610 23390
rect 31778 22544 32070 23390
rect 32238 22544 32530 23390
rect 32698 22544 32990 23390
rect 33158 22544 33542 23390
rect 33710 22544 34002 23390
rect 34170 22544 34462 23390
rect 34630 22544 34922 23390
rect 35090 22544 35382 23390
rect 35550 22544 35842 23390
rect 36010 22544 36394 23390
rect 36562 22544 36854 23390
rect 37022 22544 37314 23390
rect 37482 22544 37774 23390
rect 37942 22544 38234 23390
rect 38402 22544 38786 23390
rect 38954 22544 39246 23390
rect 39414 22544 39706 23390
rect 39874 22544 40166 23390
rect 40334 22544 40626 23390
rect 40794 22544 41178 23390
rect 41346 22544 41638 23390
rect 41806 22544 42098 23390
rect 42266 22544 42558 23390
rect 42726 22544 43018 23390
rect 43186 22544 43478 23390
rect 43646 22544 44030 23390
rect 44198 22544 44490 23390
rect 44658 22544 44950 23390
rect 45118 22544 45410 23390
rect 45578 22544 45870 23390
rect 46038 22544 46422 23390
rect 46590 22544 46882 23390
rect 47050 22544 47342 23390
rect 47510 22544 47802 23390
rect 47970 22544 48262 23390
rect 48430 22544 48814 23390
rect 48982 22544 49274 23390
rect 49442 22544 49734 23390
rect 49902 22544 50194 23390
rect 50362 22544 50654 23390
rect 50822 22544 51114 23390
rect 51282 22544 51666 23390
rect 51834 22544 52126 23390
rect 52294 22544 52586 23390
rect 52754 22544 53046 23390
rect 53214 22544 53506 23390
rect 53674 22544 54058 23390
rect 54226 22544 54518 23390
rect 54686 22544 54978 23390
rect 55146 22544 55438 23390
rect 55606 22544 55898 23390
rect 56066 22544 56450 23390
rect 56618 22544 56910 23390
rect 57078 22544 57370 23390
rect 57538 22544 57830 23390
rect 57998 22544 58290 23390
rect 58458 22544 58750 23390
rect 58918 22544 59302 23390
rect 59470 22544 59762 23390
rect 59930 22544 60222 23390
rect 60390 22544 60682 23390
rect 60850 22544 61142 23390
rect 61310 22544 61694 23390
rect 61862 22544 62154 23390
rect 62322 22544 62614 23390
rect 62782 22544 63074 23390
rect 63242 22544 63534 23390
rect 63702 22544 63994 23390
rect 64162 22544 64546 23390
rect 64714 22544 65006 23390
rect 65174 22544 65466 23390
rect 65634 22544 65926 23390
rect 66094 22544 66386 23390
rect 66554 22544 66938 23390
rect 67106 22544 67398 23390
rect 67566 22544 67858 23390
rect 68026 22544 68318 23390
rect 68486 22544 68778 23390
rect 68946 22544 69330 23390
rect 69498 22544 69790 23390
rect 69958 22544 70250 23390
rect 70418 22544 70710 23390
rect 70878 22544 71170 23390
rect 71338 22544 71630 23390
rect 71798 22544 72182 23390
rect 72350 22544 72642 23390
rect 72810 22544 73102 23390
rect 73270 22544 73562 23390
rect 73730 22544 74022 23390
rect 74190 22544 74574 23390
rect 74742 22544 75034 23390
rect 75202 22544 75494 23390
rect 75662 22544 75954 23390
rect 76122 22544 76414 23390
rect 76582 22544 76966 23390
rect 77134 22544 77426 23390
rect 77594 22544 77886 23390
rect 78054 22544 78346 23390
rect 78514 22544 78806 23390
rect 78974 22544 79266 23390
rect 79434 22544 79818 23390
rect 79986 22544 80278 23390
rect 80446 22544 80738 23390
rect 80906 22544 81198 23390
rect 81366 22544 81658 23390
rect 81826 22544 82210 23390
rect 82378 22544 82670 23390
rect 82838 22544 83130 23390
rect 83298 22544 83590 23390
rect 83758 22544 84050 23390
rect 84218 22544 84602 23390
rect 84770 22544 85062 23390
rect 85230 22544 85522 23390
rect 85690 22544 85982 23390
rect 86150 22544 86442 23390
rect 86610 22544 86902 23390
rect 87070 22544 87454 23390
rect 87622 22544 87914 23390
rect 88082 22544 88374 23390
rect 88542 22544 88834 23390
rect 89002 22544 89294 23390
rect 89462 22544 89846 23390
rect 90014 22544 90306 23390
rect 90474 22544 90766 23390
rect 90934 22544 91226 23390
rect 91394 22544 91686 23390
rect 91854 22544 92238 23390
rect 92406 22544 92698 23390
rect 92866 22544 93158 23390
rect 93326 22544 93618 23390
rect 93786 22544 94078 23390
rect 94246 22544 94538 23390
rect 94706 22544 95090 23390
rect 95258 22544 95550 23390
rect 95718 22544 96010 23390
rect 96178 22544 96470 23390
rect 96638 22544 96930 23390
rect 97098 22544 97482 23390
rect 97650 22544 97942 23390
rect 98110 22544 98402 23390
rect 98570 22544 98862 23390
rect 99030 22544 99322 23390
rect 99490 22544 99782 23390
rect 99950 22544 100334 23390
rect 100502 22544 100794 23390
rect 100962 22544 101254 23390
rect 101422 22544 101714 23390
rect 101882 22544 102174 23390
rect 102342 22544 102726 23390
rect 102894 22544 103186 23390
rect 103354 22544 103646 23390
rect 103814 22544 104106 23390
rect 104274 22544 104566 23390
rect 104734 22544 105118 23390
rect 105286 22544 105578 23390
rect 105746 22544 106038 23390
rect 106206 22544 106498 23390
rect 106666 22544 106958 23390
rect 107126 22544 107418 23390
rect 107586 22544 107970 23390
rect 108138 22544 108430 23390
rect 108598 22544 108890 23390
rect 109058 22544 109350 23390
rect 109518 22544 109810 23390
rect 109978 22544 110362 23390
rect 110530 22544 110822 23390
rect 110990 22544 111282 23390
rect 111450 22544 111742 23390
rect 111910 22544 112202 23390
rect 112370 22544 112754 23390
rect 112922 22544 113214 23390
rect 113382 22544 113674 23390
rect 113842 22544 114134 23390
rect 114302 22544 114594 23390
rect 114762 22544 115054 23390
rect 115222 22544 115606 23390
rect 115774 22544 116066 23390
rect 116234 22544 116526 23390
rect 116694 22544 116986 23390
rect 117154 22544 117446 23390
rect 117614 22544 117998 23390
rect 118166 22544 118458 23390
rect 118626 22544 118918 23390
rect 119086 22544 119378 23390
rect 119546 22544 119838 23390
rect 120006 22544 120390 23390
rect 120558 22544 120850 23390
rect 121018 22544 121310 23390
rect 121478 22544 121770 23390
rect 121938 22544 122230 23390
rect 122398 22544 122690 23390
rect 122858 22544 123242 23390
rect 123410 22544 123702 23390
rect 123870 22544 124162 23390
rect 124330 22544 124622 23390
rect 124790 22544 125082 23390
rect 125250 22544 125634 23390
rect 125802 22544 126094 23390
rect 126262 22544 126554 23390
rect 126722 22544 127014 23390
rect 127182 22544 127474 23390
rect 127642 22544 127934 23390
rect 128102 22544 128486 23390
rect 128654 22544 128946 23390
rect 129114 22544 129406 23390
rect 129574 22544 129866 23390
rect 130034 22544 130326 23390
rect 130494 22544 130878 23390
rect 131046 22544 131338 23390
rect 131506 22544 131798 23390
rect 131966 22544 132258 23390
rect 132426 22544 132718 23390
rect 132886 22544 133270 23390
rect 133438 22544 133730 23390
rect 133898 22544 134190 23390
rect 134358 22544 134650 23390
rect 134818 22544 135110 23390
rect 135278 22544 135570 23390
rect 135738 22544 136122 23390
rect 136290 22544 136582 23390
rect 136750 22544 137042 23390
rect 137210 22544 137502 23390
rect 137670 22544 137962 23390
rect 138130 22544 138514 23390
rect 138682 22544 138974 23390
rect 139142 22544 139434 23390
rect 139602 22544 139894 23390
rect 140062 22544 140354 23390
rect 140522 22544 140906 23390
rect 141074 22544 141366 23390
rect 141534 22544 141826 23390
rect 141994 22544 142286 23390
rect 142454 22544 142746 23390
rect 142914 22544 143206 23390
rect 143374 22544 143758 23390
rect 143926 22544 144218 23390
rect 144386 22544 144678 23390
rect 144846 22544 145138 23390
rect 145306 22544 145598 23390
rect 145766 22544 146150 23390
rect 146318 22544 146610 23390
rect 146778 22544 147070 23390
rect 147238 22544 147530 23390
rect 147698 22544 147990 23390
rect 148158 22544 148542 23390
rect 148710 22544 149002 23390
rect 149170 22544 149462 23390
rect 149630 22544 149922 23390
rect 150090 22544 150382 23390
rect 150550 22544 150842 23390
rect 151010 22544 151394 23390
rect 151562 22544 151854 23390
rect 152022 22544 152314 23390
rect 152482 22544 152774 23390
rect 152942 22544 153234 23390
rect 153402 22544 153786 23390
rect 153954 22544 154246 23390
rect 154414 22544 154706 23390
rect 154874 22544 155166 23390
rect 155334 22544 155626 23390
rect 155794 22544 156178 23390
rect 156346 22544 156638 23390
rect 156806 22544 157098 23390
rect 157266 22544 157558 23390
rect 157726 22544 158018 23390
rect 158186 22544 158478 23390
rect 158646 22544 159030 23390
rect 159198 22544 159490 23390
rect 159658 22544 159950 23390
rect 160118 22544 160410 23390
rect 160578 22544 160870 23390
rect 161038 22544 161422 23390
rect 161590 22544 161882 23390
rect 162050 22544 162342 23390
rect 162510 22544 162802 23390
rect 162970 22544 163262 23390
rect 163430 22544 163722 23390
rect 163890 22544 164274 23390
rect 164442 22544 164734 23390
rect 164902 22544 165194 23390
rect 165362 22544 165654 23390
rect 165822 22544 166114 23390
rect 166282 22544 166666 23390
rect 166834 22544 167126 23390
rect 167294 22544 167586 23390
rect 167754 22544 168046 23390
rect 168214 22544 168506 23390
rect 168674 22544 169058 23390
rect 169226 22544 169518 23390
rect 169686 22544 169978 23390
rect 170146 22544 170438 23390
rect 170606 22544 170898 23390
rect 171066 22544 171358 23390
rect 171526 22544 171910 23390
rect 172078 22544 172370 23390
rect 172538 22544 172830 23390
rect 172998 22544 173290 23390
rect 173458 22544 173750 23390
rect 173918 22544 174302 23390
rect 174470 22544 174762 23390
rect 174930 22544 175222 23390
rect 175390 22544 175682 23390
rect 175850 22544 176142 23390
rect 176310 22544 176694 23390
rect 176862 22544 177154 23390
rect 177322 22544 177614 23390
rect 177782 22544 178074 23390
rect 178242 22544 178534 23390
rect 178702 22544 178994 23390
rect 179162 22544 179546 23390
rect 179714 22544 180006 23390
rect 180174 22544 180466 23390
rect 180634 22544 180926 23390
rect 181094 22544 181386 23390
rect 181554 22544 181938 23390
rect 182106 22544 182398 23390
rect 182566 22544 182858 23390
rect 183026 22544 183318 23390
rect 183486 22544 183778 23390
rect 183946 22544 184330 23390
rect 184498 22544 184790 23390
rect 184958 22544 185250 23390
rect 185418 22544 185710 23390
rect 185878 22544 186170 23390
rect 186338 22544 186630 23390
rect 186798 22544 187182 23390
rect 187350 22544 187642 23390
rect 187810 22544 188102 23390
rect 188270 22544 188562 23390
rect 188730 22544 189022 23390
rect 189190 22544 189574 23390
rect 189742 22544 190034 23390
rect 190202 22544 190494 23390
rect 190662 22544 190954 23390
rect 191122 22544 191414 23390
rect 191582 22544 191874 23390
rect 192042 22544 192426 23390
rect 192594 22544 192886 23390
rect 193054 22544 193346 23390
rect 193514 22544 193806 23390
rect 193974 22544 194266 23390
rect 194434 22544 194818 23390
rect 194986 22544 195278 23390
rect 195446 22544 195738 23390
rect 195906 22544 196198 23390
rect 196366 22544 196658 23390
rect 196826 22544 197210 23390
rect 197378 22544 197670 23390
rect 197838 22544 198130 23390
rect 198298 22544 198590 23390
rect 198758 22544 199050 23390
rect 199218 22544 199510 23390
rect 199678 22544 200062 23390
rect 200230 22544 200522 23390
rect 200690 22544 200982 23390
rect 201150 22544 201442 23390
rect 201610 22544 201902 23390
rect 202070 22544 202454 23390
rect 202622 22544 202914 23390
rect 203082 22544 203374 23390
rect 203542 22544 203834 23390
rect 204002 22544 204294 23390
rect 204462 22544 204846 23390
rect 205014 22544 205306 23390
rect 205474 22544 205766 23390
rect 205934 22544 206226 23390
rect 206394 22544 206686 23390
rect 206854 22544 207146 23390
rect 207314 22544 207698 23390
rect 207866 22544 208158 23390
rect 208326 22544 208618 23390
rect 208786 22544 209078 23390
rect 209246 22544 209538 23390
rect 209706 22544 210090 23390
rect 210258 22544 210550 23390
rect 210718 22544 211010 23390
rect 211178 22544 211470 23390
rect 211638 22544 211930 23390
rect 212098 22544 212482 23390
rect 212650 22544 212942 23390
rect 213110 22544 213402 23390
rect 213570 22544 213862 23390
rect 214030 22544 214322 23390
rect 214490 22544 214782 23390
rect 214950 22544 215334 23390
rect 215502 22544 215794 23390
rect 215962 22544 216254 23390
rect 216422 22544 216714 23390
rect 216882 22544 217174 23390
rect 217342 22544 217726 23390
rect 217894 22544 218186 23390
rect 218354 22544 218646 23390
rect 218814 22544 219106 23390
rect 219274 22544 219566 23390
rect 219734 22544 219768 23390
rect 20 856 219768 22544
rect 20 2 146 856
rect 314 2 514 856
rect 682 2 882 856
rect 1050 2 1250 856
rect 1418 2 1618 856
rect 1786 2 1986 856
rect 2154 2 2354 856
rect 2522 2 2722 856
rect 2890 2 3090 856
rect 3258 2 3458 856
rect 3626 2 3918 856
rect 4086 2 4286 856
rect 4454 2 4654 856
rect 4822 2 5022 856
rect 5190 2 5390 856
rect 5558 2 5758 856
rect 5926 2 6126 856
rect 6294 2 6494 856
rect 6662 2 6862 856
rect 7030 2 7230 856
rect 7398 2 7690 856
rect 7858 2 8058 856
rect 8226 2 8426 856
rect 8594 2 8794 856
rect 8962 2 9162 856
rect 9330 2 9530 856
rect 9698 2 9898 856
rect 10066 2 10266 856
rect 10434 2 10634 856
rect 10802 2 11002 856
rect 11170 2 11462 856
rect 11630 2 11830 856
rect 11998 2 12198 856
rect 12366 2 12566 856
rect 12734 2 12934 856
rect 13102 2 13302 856
rect 13470 2 13670 856
rect 13838 2 14038 856
rect 14206 2 14406 856
rect 14574 2 14774 856
rect 14942 2 15234 856
rect 15402 2 15602 856
rect 15770 2 15970 856
rect 16138 2 16338 856
rect 16506 2 16706 856
rect 16874 2 17074 856
rect 17242 2 17442 856
rect 17610 2 17810 856
rect 17978 2 18178 856
rect 18346 2 18546 856
rect 18714 2 19006 856
rect 19174 2 19374 856
rect 19542 2 19742 856
rect 19910 2 20110 856
rect 20278 2 20478 856
rect 20646 2 20846 856
rect 21014 2 21214 856
rect 21382 2 21582 856
rect 21750 2 21950 856
rect 22118 2 22318 856
rect 22486 2 22778 856
rect 22946 2 23146 856
rect 23314 2 23514 856
rect 23682 2 23882 856
rect 24050 2 24250 856
rect 24418 2 24618 856
rect 24786 2 24986 856
rect 25154 2 25354 856
rect 25522 2 25722 856
rect 25890 2 26090 856
rect 26258 2 26550 856
rect 26718 2 26918 856
rect 27086 2 27286 856
rect 27454 2 27654 856
rect 27822 2 28022 856
rect 28190 2 28390 856
rect 28558 2 28758 856
rect 28926 2 29126 856
rect 29294 2 29494 856
rect 29662 2 29862 856
rect 30030 2 30322 856
rect 30490 2 30690 856
rect 30858 2 31058 856
rect 31226 2 31426 856
rect 31594 2 31794 856
rect 31962 2 32162 856
rect 32330 2 32530 856
rect 32698 2 32898 856
rect 33066 2 33266 856
rect 33434 2 33726 856
rect 33894 2 34094 856
rect 34262 2 34462 856
rect 34630 2 34830 856
rect 34998 2 35198 856
rect 35366 2 35566 856
rect 35734 2 35934 856
rect 36102 2 36302 856
rect 36470 2 36670 856
rect 36838 2 37038 856
rect 37206 2 37498 856
rect 37666 2 37866 856
rect 38034 2 38234 856
rect 38402 2 38602 856
rect 38770 2 38970 856
rect 39138 2 39338 856
rect 39506 2 39706 856
rect 39874 2 40074 856
rect 40242 2 40442 856
rect 40610 2 40810 856
rect 40978 2 41270 856
rect 41438 2 41638 856
rect 41806 2 42006 856
rect 42174 2 42374 856
rect 42542 2 42742 856
rect 42910 2 43110 856
rect 43278 2 43478 856
rect 43646 2 43846 856
rect 44014 2 44214 856
rect 44382 2 44582 856
rect 44750 2 45042 856
rect 45210 2 45410 856
rect 45578 2 45778 856
rect 45946 2 46146 856
rect 46314 2 46514 856
rect 46682 2 46882 856
rect 47050 2 47250 856
rect 47418 2 47618 856
rect 47786 2 47986 856
rect 48154 2 48354 856
rect 48522 2 48814 856
rect 48982 2 49182 856
rect 49350 2 49550 856
rect 49718 2 49918 856
rect 50086 2 50286 856
rect 50454 2 50654 856
rect 50822 2 51022 856
rect 51190 2 51390 856
rect 51558 2 51758 856
rect 51926 2 52126 856
rect 52294 2 52586 856
rect 52754 2 52954 856
rect 53122 2 53322 856
rect 53490 2 53690 856
rect 53858 2 54058 856
rect 54226 2 54426 856
rect 54594 2 54794 856
rect 54962 2 55162 856
rect 55330 2 55530 856
rect 55698 2 55898 856
rect 56066 2 56358 856
rect 56526 2 56726 856
rect 56894 2 57094 856
rect 57262 2 57462 856
rect 57630 2 57830 856
rect 57998 2 58198 856
rect 58366 2 58566 856
rect 58734 2 58934 856
rect 59102 2 59302 856
rect 59470 2 59670 856
rect 59838 2 60130 856
rect 60298 2 60498 856
rect 60666 2 60866 856
rect 61034 2 61234 856
rect 61402 2 61602 856
rect 61770 2 61970 856
rect 62138 2 62338 856
rect 62506 2 62706 856
rect 62874 2 63074 856
rect 63242 2 63534 856
rect 63702 2 63902 856
rect 64070 2 64270 856
rect 64438 2 64638 856
rect 64806 2 65006 856
rect 65174 2 65374 856
rect 65542 2 65742 856
rect 65910 2 66110 856
rect 66278 2 66478 856
rect 66646 2 66846 856
rect 67014 2 67306 856
rect 67474 2 67674 856
rect 67842 2 68042 856
rect 68210 2 68410 856
rect 68578 2 68778 856
rect 68946 2 69146 856
rect 69314 2 69514 856
rect 69682 2 69882 856
rect 70050 2 70250 856
rect 70418 2 70618 856
rect 70786 2 71078 856
rect 71246 2 71446 856
rect 71614 2 71814 856
rect 71982 2 72182 856
rect 72350 2 72550 856
rect 72718 2 72918 856
rect 73086 2 73286 856
rect 73454 2 73654 856
rect 73822 2 74022 856
rect 74190 2 74390 856
rect 74558 2 74850 856
rect 75018 2 75218 856
rect 75386 2 75586 856
rect 75754 2 75954 856
rect 76122 2 76322 856
rect 76490 2 76690 856
rect 76858 2 77058 856
rect 77226 2 77426 856
rect 77594 2 77794 856
rect 77962 2 78162 856
rect 78330 2 78622 856
rect 78790 2 78990 856
rect 79158 2 79358 856
rect 79526 2 79726 856
rect 79894 2 80094 856
rect 80262 2 80462 856
rect 80630 2 80830 856
rect 80998 2 81198 856
rect 81366 2 81566 856
rect 81734 2 81934 856
rect 82102 2 82394 856
rect 82562 2 82762 856
rect 82930 2 83130 856
rect 83298 2 83498 856
rect 83666 2 83866 856
rect 84034 2 84234 856
rect 84402 2 84602 856
rect 84770 2 84970 856
rect 85138 2 85338 856
rect 85506 2 85706 856
rect 85874 2 86166 856
rect 86334 2 86534 856
rect 86702 2 86902 856
rect 87070 2 87270 856
rect 87438 2 87638 856
rect 87806 2 88006 856
rect 88174 2 88374 856
rect 88542 2 88742 856
rect 88910 2 89110 856
rect 89278 2 89478 856
rect 89646 2 89938 856
rect 90106 2 90306 856
rect 90474 2 90674 856
rect 90842 2 91042 856
rect 91210 2 91410 856
rect 91578 2 91778 856
rect 91946 2 92146 856
rect 92314 2 92514 856
rect 92682 2 92882 856
rect 93050 2 93250 856
rect 93418 2 93710 856
rect 93878 2 94078 856
rect 94246 2 94446 856
rect 94614 2 94814 856
rect 94982 2 95182 856
rect 95350 2 95550 856
rect 95718 2 95918 856
rect 96086 2 96286 856
rect 96454 2 96654 856
rect 96822 2 97114 856
rect 97282 2 97482 856
rect 97650 2 97850 856
rect 98018 2 98218 856
rect 98386 2 98586 856
rect 98754 2 98954 856
rect 99122 2 99322 856
rect 99490 2 99690 856
rect 99858 2 100058 856
rect 100226 2 100426 856
rect 100594 2 100886 856
rect 101054 2 101254 856
rect 101422 2 101622 856
rect 101790 2 101990 856
rect 102158 2 102358 856
rect 102526 2 102726 856
rect 102894 2 103094 856
rect 103262 2 103462 856
rect 103630 2 103830 856
rect 103998 2 104198 856
rect 104366 2 104658 856
rect 104826 2 105026 856
rect 105194 2 105394 856
rect 105562 2 105762 856
rect 105930 2 106130 856
rect 106298 2 106498 856
rect 106666 2 106866 856
rect 107034 2 107234 856
rect 107402 2 107602 856
rect 107770 2 107970 856
rect 108138 2 108430 856
rect 108598 2 108798 856
rect 108966 2 109166 856
rect 109334 2 109534 856
rect 109702 2 109902 856
rect 110070 2 110270 856
rect 110438 2 110638 856
rect 110806 2 111006 856
rect 111174 2 111374 856
rect 111542 2 111742 856
rect 111910 2 112202 856
rect 112370 2 112570 856
rect 112738 2 112938 856
rect 113106 2 113306 856
rect 113474 2 113674 856
rect 113842 2 114042 856
rect 114210 2 114410 856
rect 114578 2 114778 856
rect 114946 2 115146 856
rect 115314 2 115514 856
rect 115682 2 115974 856
rect 116142 2 116342 856
rect 116510 2 116710 856
rect 116878 2 117078 856
rect 117246 2 117446 856
rect 117614 2 117814 856
rect 117982 2 118182 856
rect 118350 2 118550 856
rect 118718 2 118918 856
rect 119086 2 119286 856
rect 119454 2 119746 856
rect 119914 2 120114 856
rect 120282 2 120482 856
rect 120650 2 120850 856
rect 121018 2 121218 856
rect 121386 2 121586 856
rect 121754 2 121954 856
rect 122122 2 122322 856
rect 122490 2 122690 856
rect 122858 2 123058 856
rect 123226 2 123518 856
rect 123686 2 123886 856
rect 124054 2 124254 856
rect 124422 2 124622 856
rect 124790 2 124990 856
rect 125158 2 125358 856
rect 125526 2 125726 856
rect 125894 2 126094 856
rect 126262 2 126462 856
rect 126630 2 126922 856
rect 127090 2 127290 856
rect 127458 2 127658 856
rect 127826 2 128026 856
rect 128194 2 128394 856
rect 128562 2 128762 856
rect 128930 2 129130 856
rect 129298 2 129498 856
rect 129666 2 129866 856
rect 130034 2 130234 856
rect 130402 2 130694 856
rect 130862 2 131062 856
rect 131230 2 131430 856
rect 131598 2 131798 856
rect 131966 2 132166 856
rect 132334 2 132534 856
rect 132702 2 132902 856
rect 133070 2 133270 856
rect 133438 2 133638 856
rect 133806 2 134006 856
rect 134174 2 134466 856
rect 134634 2 134834 856
rect 135002 2 135202 856
rect 135370 2 135570 856
rect 135738 2 135938 856
rect 136106 2 136306 856
rect 136474 2 136674 856
rect 136842 2 137042 856
rect 137210 2 137410 856
rect 137578 2 137778 856
rect 137946 2 138238 856
rect 138406 2 138606 856
rect 138774 2 138974 856
rect 139142 2 139342 856
rect 139510 2 139710 856
rect 139878 2 140078 856
rect 140246 2 140446 856
rect 140614 2 140814 856
rect 140982 2 141182 856
rect 141350 2 141550 856
rect 141718 2 142010 856
rect 142178 2 142378 856
rect 142546 2 142746 856
rect 142914 2 143114 856
rect 143282 2 143482 856
rect 143650 2 143850 856
rect 144018 2 144218 856
rect 144386 2 144586 856
rect 144754 2 144954 856
rect 145122 2 145322 856
rect 145490 2 145782 856
rect 145950 2 146150 856
rect 146318 2 146518 856
rect 146686 2 146886 856
rect 147054 2 147254 856
rect 147422 2 147622 856
rect 147790 2 147990 856
rect 148158 2 148358 856
rect 148526 2 148726 856
rect 148894 2 149094 856
rect 149262 2 149554 856
rect 149722 2 149922 856
rect 150090 2 150290 856
rect 150458 2 150658 856
rect 150826 2 151026 856
rect 151194 2 151394 856
rect 151562 2 151762 856
rect 151930 2 152130 856
rect 152298 2 152498 856
rect 152666 2 152866 856
rect 153034 2 153326 856
rect 153494 2 153694 856
rect 153862 2 154062 856
rect 154230 2 154430 856
rect 154598 2 154798 856
rect 154966 2 155166 856
rect 155334 2 155534 856
rect 155702 2 155902 856
rect 156070 2 156270 856
rect 156438 2 156638 856
rect 156806 2 157098 856
rect 157266 2 157466 856
rect 157634 2 157834 856
rect 158002 2 158202 856
rect 158370 2 158570 856
rect 158738 2 158938 856
rect 159106 2 159306 856
rect 159474 2 159674 856
rect 159842 2 160042 856
rect 160210 2 160502 856
rect 160670 2 160870 856
rect 161038 2 161238 856
rect 161406 2 161606 856
rect 161774 2 161974 856
rect 162142 2 162342 856
rect 162510 2 162710 856
rect 162878 2 163078 856
rect 163246 2 163446 856
rect 163614 2 163814 856
rect 163982 2 164274 856
rect 164442 2 164642 856
rect 164810 2 165010 856
rect 165178 2 165378 856
rect 165546 2 165746 856
rect 165914 2 166114 856
rect 166282 2 166482 856
rect 166650 2 166850 856
rect 167018 2 167218 856
rect 167386 2 167586 856
rect 167754 2 168046 856
rect 168214 2 168414 856
rect 168582 2 168782 856
rect 168950 2 169150 856
rect 169318 2 169518 856
rect 169686 2 169886 856
rect 170054 2 170254 856
rect 170422 2 170622 856
rect 170790 2 170990 856
rect 171158 2 171358 856
rect 171526 2 171818 856
rect 171986 2 172186 856
rect 172354 2 172554 856
rect 172722 2 172922 856
rect 173090 2 173290 856
rect 173458 2 173658 856
rect 173826 2 174026 856
rect 174194 2 174394 856
rect 174562 2 174762 856
rect 174930 2 175130 856
rect 175298 2 175590 856
rect 175758 2 175958 856
rect 176126 2 176326 856
rect 176494 2 176694 856
rect 176862 2 177062 856
rect 177230 2 177430 856
rect 177598 2 177798 856
rect 177966 2 178166 856
rect 178334 2 178534 856
rect 178702 2 178902 856
rect 179070 2 179362 856
rect 179530 2 179730 856
rect 179898 2 180098 856
rect 180266 2 180466 856
rect 180634 2 180834 856
rect 181002 2 181202 856
rect 181370 2 181570 856
rect 181738 2 181938 856
rect 182106 2 182306 856
rect 182474 2 182674 856
rect 182842 2 183134 856
rect 183302 2 183502 856
rect 183670 2 183870 856
rect 184038 2 184238 856
rect 184406 2 184606 856
rect 184774 2 184974 856
rect 185142 2 185342 856
rect 185510 2 185710 856
rect 185878 2 186078 856
rect 186246 2 186446 856
rect 186614 2 186906 856
rect 187074 2 187274 856
rect 187442 2 187642 856
rect 187810 2 188010 856
rect 188178 2 188378 856
rect 188546 2 188746 856
rect 188914 2 189114 856
rect 189282 2 189482 856
rect 189650 2 189850 856
rect 190018 2 190310 856
rect 190478 2 190678 856
rect 190846 2 191046 856
rect 191214 2 191414 856
rect 191582 2 191782 856
rect 191950 2 192150 856
rect 192318 2 192518 856
rect 192686 2 192886 856
rect 193054 2 193254 856
rect 193422 2 193622 856
rect 193790 2 194082 856
rect 194250 2 194450 856
rect 194618 2 194818 856
rect 194986 2 195186 856
rect 195354 2 195554 856
rect 195722 2 195922 856
rect 196090 2 196290 856
rect 196458 2 196658 856
rect 196826 2 197026 856
rect 197194 2 197394 856
rect 197562 2 197854 856
rect 198022 2 198222 856
rect 198390 2 198590 856
rect 198758 2 198958 856
rect 199126 2 199326 856
rect 199494 2 199694 856
rect 199862 2 200062 856
rect 200230 2 200430 856
rect 200598 2 200798 856
rect 200966 2 201166 856
rect 201334 2 201626 856
rect 201794 2 201994 856
rect 202162 2 202362 856
rect 202530 2 202730 856
rect 202898 2 203098 856
rect 203266 2 203466 856
rect 203634 2 203834 856
rect 204002 2 204202 856
rect 204370 2 204570 856
rect 204738 2 204938 856
rect 205106 2 205398 856
rect 205566 2 205766 856
rect 205934 2 206134 856
rect 206302 2 206502 856
rect 206670 2 206870 856
rect 207038 2 207238 856
rect 207406 2 207606 856
rect 207774 2 207974 856
rect 208142 2 208342 856
rect 208510 2 208710 856
rect 208878 2 209170 856
rect 209338 2 209538 856
rect 209706 2 209906 856
rect 210074 2 210274 856
rect 210442 2 210642 856
rect 210810 2 211010 856
rect 211178 2 211378 856
rect 211546 2 211746 856
rect 211914 2 212114 856
rect 212282 2 212482 856
rect 212650 2 212942 856
rect 213110 2 213310 856
rect 213478 2 213678 856
rect 213846 2 214046 856
rect 214214 2 214414 856
rect 214582 2 214782 856
rect 214950 2 215150 856
rect 215318 2 215518 856
rect 215686 2 215886 856
rect 216054 2 216254 856
rect 216422 2 216714 856
rect 216882 2 217082 856
rect 217250 2 217450 856
rect 217618 2 217818 856
rect 217986 2 218186 856
rect 218354 2 218554 856
rect 218722 2 218922 856
rect 219090 2 219290 856
rect 219458 2 219658 856
<< metal3 >>
rect -2762 25990 222734 26170
rect -2498 25726 222470 25906
rect -2234 25462 222206 25642
rect -1970 25198 221942 25378
rect -1706 24934 221678 25114
rect -1442 24670 221414 24850
rect -1178 24406 221150 24586
rect -914 24142 220886 24322
rect -650 23878 220622 24058
rect -386 23614 220358 23794
rect 219200 22040 220400 22160
rect 219200 19728 220400 19848
rect -400 19320 800 19440
rect 219200 17416 220400 17536
rect 219200 15104 220400 15224
rect 219200 12792 220400 12912
rect -400 11568 800 11688
rect 219200 10344 220400 10464
rect 219200 8032 220400 8152
rect 219200 5720 220400 5840
rect -400 3816 800 3936
rect 219200 3408 220400 3528
rect 219200 1096 220400 1216
rect -386 -402 220358 -222
rect -650 -666 220622 -486
rect -914 -930 220886 -750
rect -1178 -1194 221150 -1014
rect -1442 -1458 221414 -1278
rect -1706 -1722 221678 -1542
rect -1970 -1986 221942 -1806
rect -2234 -2250 222206 -2070
rect -2498 -2514 222470 -2334
rect -2762 -2778 222734 -2598
<< obsm3 >>
rect 800 22240 219407 22813
rect 800 21960 219120 22240
rect 800 19928 219407 21960
rect 800 19648 219120 19928
rect 800 19520 219407 19648
rect 880 19240 219407 19520
rect 800 17616 219407 19240
rect 800 17336 219120 17616
rect 800 15304 219407 17336
rect 800 15024 219120 15304
rect 800 12992 219407 15024
rect 800 12712 219120 12992
rect 800 11768 219407 12712
rect 880 11488 219407 11768
rect 800 10544 219407 11488
rect 800 10264 219120 10544
rect 800 8232 219407 10264
rect 800 7952 219120 8232
rect 800 5920 219407 7952
rect 800 5640 219120 5920
rect 800 4016 219407 5640
rect 880 3736 219407 4016
rect 800 3608 219407 3736
rect 800 3328 219120 3608
rect 800 1296 219407 3328
rect 800 1016 219120 1296
rect 800 35 219407 1016
<< metal4 >>
rect -2762 -2778 -2582 26170
rect -2498 -2514 -2318 25906
rect -2234 -2250 -2054 25642
rect -1970 -1986 -1790 25378
rect -1706 -1722 -1526 25114
rect -1442 -1458 -1262 24850
rect -1178 -1194 -998 24586
rect -914 -930 -734 24322
rect -650 -666 -470 24058
rect -386 -402 -206 23794
rect 4014 -666 4194 24058
rect 4834 -1194 5014 24586
rect 5654 -1722 5834 25114
rect 6474 -2250 6654 25642
rect 7294 -2778 7474 26170
rect 19064 -666 19244 24058
rect 19884 -1194 20064 24586
rect 20704 -1722 20884 25114
rect 21524 -2250 21704 25642
rect 22344 -2778 22524 26170
rect 34114 -666 34294 24058
rect 34934 -1194 35114 24586
rect 35754 -1722 35934 25114
rect 36574 -2250 36754 25642
rect 37394 -2778 37574 26170
rect 49164 -666 49344 24058
rect 49984 -1194 50164 24586
rect 50804 -1722 50984 25114
rect 51624 -2250 51804 25642
rect 52444 -2778 52624 26170
rect 64214 -666 64394 24058
rect 65034 -1194 65214 24586
rect 65854 -1722 66034 25114
rect 66674 -2250 66854 25642
rect 67494 -2778 67674 26170
rect 79264 -666 79444 24058
rect 80084 -1194 80264 24586
rect 80904 -1722 81084 25114
rect 81724 -2250 81904 25642
rect 82544 -2778 82724 26170
rect 94314 -666 94494 24058
rect 95134 -1194 95314 24586
rect 95954 -1722 96134 25114
rect 96774 -2250 96954 25642
rect 97594 -2778 97774 26170
rect 109364 -666 109544 24058
rect 110184 -1194 110364 24586
rect 111004 -1722 111184 25114
rect 111824 -2250 112004 25642
rect 112644 -2778 112824 26170
rect 124414 -666 124594 24058
rect 125234 -1194 125414 24586
rect 126054 -1722 126234 25114
rect 126874 -2250 127054 25642
rect 127694 -2778 127874 26170
rect 139464 -666 139644 24058
rect 140284 -1194 140464 24586
rect 141104 -1722 141284 25114
rect 141924 -2250 142104 25642
rect 142744 -2778 142924 26170
rect 154514 -666 154694 24058
rect 155334 -1194 155514 24586
rect 156154 -1722 156334 25114
rect 156974 -2250 157154 25642
rect 157794 -2778 157974 26170
rect 169564 -666 169744 24058
rect 170384 -1194 170564 24586
rect 171204 -1722 171384 25114
rect 172024 -2250 172204 25642
rect 172844 -2778 173024 26170
rect 184614 -666 184794 24058
rect 185434 -1194 185614 24586
rect 186254 -1722 186434 25114
rect 187074 -2250 187254 25642
rect 187894 -2778 188074 26170
rect 199664 -666 199844 24058
rect 200484 -1194 200664 24586
rect 201304 -1722 201484 25114
rect 202124 -2250 202304 25642
rect 202944 -2778 203124 26170
rect 214714 -666 214894 24058
rect 215534 -1194 215714 24586
rect 216354 -1722 216534 25114
rect 217174 -2250 217354 25642
rect 217994 -2778 218174 26170
rect 220178 -402 220358 23794
rect 220442 -666 220622 24058
rect 220706 -930 220886 24322
rect 220970 -1194 221150 24586
rect 221234 -1458 221414 24850
rect 221498 -1722 221678 25114
rect 221762 -1986 221942 25378
rect 222026 -2250 222206 25642
rect 222290 -2514 222470 25906
rect 222554 -2778 222734 26170
<< obsm4 >>
rect 5395 35 5574 22405
rect 5914 9303 6394 22405
rect 5914 7662 6369 9303
rect 5914 35 6394 7662
rect 6734 19308 7214 22405
rect 6734 17657 7088 19308
rect 6734 35 7214 17657
rect 7554 19308 18984 22405
rect 7683 17657 18984 19308
rect 7554 35 18984 17657
rect 19324 11821 19804 22405
rect 19324 10153 19712 11821
rect 19324 35 19804 10153
rect 20144 11821 20624 22405
rect 20226 10153 20624 11821
rect 20144 35 20624 10153
rect 20964 6829 21444 22405
rect 20964 5157 21361 6829
rect 20964 35 21444 5157
rect 21784 16822 22264 22405
rect 21784 15160 22180 16822
rect 21784 6829 22264 15160
rect 21865 5157 22264 6829
rect 21784 35 22264 5157
rect 22604 16822 34034 22405
rect 22679 15160 34034 16822
rect 22604 35 34034 15160
rect 34374 35 34854 22405
rect 35194 35 35674 22405
rect 36014 9325 36494 22405
rect 36014 7648 36456 9325
rect 36014 35 36494 7648
rect 36834 19308 37314 22405
rect 36834 17657 37188 19308
rect 36834 9325 37314 17657
rect 36948 7648 37314 9325
rect 36834 35 37314 7648
rect 37654 19308 49084 22405
rect 37783 17657 49084 19308
rect 37654 35 49084 17657
rect 49424 11821 49904 22405
rect 49424 10153 49812 11821
rect 49424 35 49904 10153
rect 50244 11821 50724 22405
rect 50326 10153 50724 11821
rect 50244 35 50724 10153
rect 51064 6829 51544 22405
rect 51064 5157 51461 6829
rect 51064 35 51544 5157
rect 51884 16822 52364 22405
rect 51884 15160 52280 16822
rect 51884 6829 52364 15160
rect 51965 5157 52364 6829
rect 51884 35 52364 5157
rect 52704 16822 64134 22405
rect 52779 15160 64134 16822
rect 52704 35 64134 15160
rect 64474 35 64954 22405
rect 65294 35 65774 22405
rect 66114 9325 66594 22405
rect 66114 7648 66556 9325
rect 66114 35 66594 7648
rect 66934 19308 67414 22405
rect 66934 17657 67288 19308
rect 66934 9325 67414 17657
rect 67048 7648 67414 9325
rect 66934 35 67414 7648
rect 67754 19308 79184 22405
rect 67883 17657 79184 19308
rect 67754 35 79184 17657
rect 79524 11803 80004 22405
rect 79524 10166 79981 11803
rect 79524 35 80004 10166
rect 80344 35 80824 22405
rect 81164 35 81644 22405
rect 81984 16822 82464 22405
rect 81984 15160 82380 16822
rect 81984 35 82464 15160
rect 82804 16822 94234 22405
rect 82879 15160 94234 16822
rect 82804 4325 94234 15160
rect 82804 2645 94077 4325
rect 82804 35 94234 2645
rect 94574 4325 95054 22405
rect 94628 2645 95054 4325
rect 94574 35 95054 2645
rect 95394 35 95874 22405
rect 96214 35 96694 22405
rect 97034 19308 97514 22405
rect 97034 17657 97448 19308
rect 97034 35 97514 17657
rect 97854 19308 109284 22405
rect 97963 17657 109284 19308
rect 97854 35 109284 17657
rect 109624 35 110104 22405
rect 110444 35 110924 22405
rect 111264 35 111744 22405
rect 112084 16822 112564 22405
rect 112084 15160 112480 16822
rect 112084 6806 112564 15160
rect 112102 5174 112564 6806
rect 112084 35 112564 5174
rect 112904 16822 124334 22405
rect 112979 15160 124334 16822
rect 112904 4309 124334 15160
rect 112904 2690 124308 4309
rect 112904 35 124334 2690
rect 124674 14318 125154 22405
rect 124674 12648 125068 14318
rect 124674 35 125154 12648
rect 125494 14318 125974 22405
rect 125546 12648 125974 14318
rect 125494 35 125974 12648
rect 126314 9307 126794 22405
rect 126314 7662 126774 9307
rect 126314 35 126794 7662
rect 127134 19308 127614 22405
rect 127134 18057 127368 19308
rect 127134 35 127614 18057
rect 127954 19308 139384 22405
rect 127963 18057 139384 19308
rect 127954 35 139384 18057
rect 139724 11821 140204 22405
rect 139724 10153 140112 11821
rect 139724 35 140204 10153
rect 140544 11821 141024 22405
rect 140626 10153 141024 11821
rect 140544 35 141024 10153
rect 141364 6829 141844 22405
rect 141364 5157 141761 6829
rect 141364 35 141844 5157
rect 142184 16822 142664 22405
rect 142184 15160 142580 16822
rect 142184 6829 142664 15160
rect 142265 5157 142664 6829
rect 142184 35 142664 5157
rect 143004 16822 154434 22405
rect 143079 15160 154434 16822
rect 143004 35 154434 15160
rect 154774 35 155254 22405
rect 155594 35 156074 22405
rect 156414 9357 156894 22405
rect 156414 7612 156823 9357
rect 156414 35 156894 7612
rect 157234 19308 157714 22405
rect 157234 17657 157588 19308
rect 157234 9357 157714 17657
rect 157274 7612 157714 9357
rect 157234 35 157714 7612
rect 158054 19308 169484 22405
rect 158183 17657 169484 19308
rect 158054 35 169484 17657
rect 169824 11821 170304 22405
rect 169824 10153 170212 11821
rect 169824 35 170304 10153
rect 170644 11821 171124 22405
rect 170726 10153 171124 11821
rect 170644 35 171124 10153
rect 171464 6829 171944 22405
rect 171464 5157 171861 6829
rect 171464 35 171944 5157
rect 172284 16822 172764 22405
rect 172284 15160 172680 16822
rect 172284 6829 172764 15160
rect 172365 5157 172764 6829
rect 172284 35 172764 5157
rect 173104 16822 184534 22405
rect 173179 15160 184534 16822
rect 173104 35 184534 15160
rect 184874 35 185354 22405
rect 185694 35 186174 22405
rect 186514 9325 186994 22405
rect 186514 7648 186956 9325
rect 186514 35 186994 7648
rect 187334 19308 187814 22405
rect 187334 17657 187688 19308
rect 187334 9325 187814 17657
rect 187448 7648 187814 9325
rect 187334 35 187814 7648
rect 188154 19308 199584 22405
rect 188283 17657 199584 19308
rect 188154 35 199584 17657
rect 199924 11821 200404 22405
rect 199924 10153 200312 11821
rect 199924 35 200404 10153
rect 200744 11821 201224 22405
rect 200826 10153 201224 11821
rect 200744 35 201224 10153
rect 201564 6829 202044 22405
rect 201564 5157 201961 6829
rect 201564 35 202044 5157
rect 202384 16822 202864 22405
rect 202384 15160 202780 16822
rect 202384 6829 202864 15160
rect 202465 5157 202864 6829
rect 202384 35 202864 5157
rect 203204 16822 214634 22405
rect 203279 15160 214634 16822
rect 203204 35 214634 15160
rect 214974 35 215454 22405
rect 215794 35 216141 22405
<< labels >>
rlabel metal3 s -400 3816 800 3936 6 caravel_clk
port 1 nsew signal input
rlabel metal3 s -400 11568 800 11688 6 caravel_clk2
port 2 nsew signal input
rlabel metal3 s -400 19320 800 19440 6 caravel_rstn
port 3 nsew signal input
rlabel metal2 s 34978 22600 35034 23800 6 la_data_in_core[0]
port 4 nsew signal output
rlabel metal2 s 178130 22600 178186 23800 6 la_data_in_core[100]
port 5 nsew signal output
rlabel metal2 s 179602 22600 179658 23800 6 la_data_in_core[101]
port 6 nsew signal output
rlabel metal2 s 180982 22600 181038 23800 6 la_data_in_core[102]
port 7 nsew signal output
rlabel metal2 s 182454 22600 182510 23800 6 la_data_in_core[103]
port 8 nsew signal output
rlabel metal2 s 183834 22600 183890 23800 6 la_data_in_core[104]
port 9 nsew signal output
rlabel metal2 s 185306 22600 185362 23800 6 la_data_in_core[105]
port 10 nsew signal output
rlabel metal2 s 186686 22600 186742 23800 6 la_data_in_core[106]
port 11 nsew signal output
rlabel metal2 s 188158 22600 188214 23800 6 la_data_in_core[107]
port 12 nsew signal output
rlabel metal2 s 189630 22600 189686 23800 6 la_data_in_core[108]
port 13 nsew signal output
rlabel metal2 s 191010 22600 191066 23800 6 la_data_in_core[109]
port 14 nsew signal output
rlabel metal2 s 49330 22600 49386 23800 6 la_data_in_core[10]
port 15 nsew signal output
rlabel metal2 s 192482 22600 192538 23800 6 la_data_in_core[110]
port 16 nsew signal output
rlabel metal2 s 193862 22600 193918 23800 6 la_data_in_core[111]
port 17 nsew signal output
rlabel metal2 s 195334 22600 195390 23800 6 la_data_in_core[112]
port 18 nsew signal output
rlabel metal2 s 196714 22600 196770 23800 6 la_data_in_core[113]
port 19 nsew signal output
rlabel metal2 s 198186 22600 198242 23800 6 la_data_in_core[114]
port 20 nsew signal output
rlabel metal2 s 199566 22600 199622 23800 6 la_data_in_core[115]
port 21 nsew signal output
rlabel metal2 s 201038 22600 201094 23800 6 la_data_in_core[116]
port 22 nsew signal output
rlabel metal2 s 202510 22600 202566 23800 6 la_data_in_core[117]
port 23 nsew signal output
rlabel metal2 s 203890 22600 203946 23800 6 la_data_in_core[118]
port 24 nsew signal output
rlabel metal2 s 205362 22600 205418 23800 6 la_data_in_core[119]
port 25 nsew signal output
rlabel metal2 s 50710 22600 50766 23800 6 la_data_in_core[11]
port 26 nsew signal output
rlabel metal2 s 206742 22600 206798 23800 6 la_data_in_core[120]
port 27 nsew signal output
rlabel metal2 s 208214 22600 208270 23800 6 la_data_in_core[121]
port 28 nsew signal output
rlabel metal2 s 209594 22600 209650 23800 6 la_data_in_core[122]
port 29 nsew signal output
rlabel metal2 s 211066 22600 211122 23800 6 la_data_in_core[123]
port 30 nsew signal output
rlabel metal2 s 212538 22600 212594 23800 6 la_data_in_core[124]
port 31 nsew signal output
rlabel metal2 s 213918 22600 213974 23800 6 la_data_in_core[125]
port 32 nsew signal output
rlabel metal2 s 215390 22600 215446 23800 6 la_data_in_core[126]
port 33 nsew signal output
rlabel metal2 s 216770 22600 216826 23800 6 la_data_in_core[127]
port 34 nsew signal output
rlabel metal2 s 52182 22600 52238 23800 6 la_data_in_core[12]
port 35 nsew signal output
rlabel metal2 s 53562 22600 53618 23800 6 la_data_in_core[13]
port 36 nsew signal output
rlabel metal2 s 55034 22600 55090 23800 6 la_data_in_core[14]
port 37 nsew signal output
rlabel metal2 s 56506 22600 56562 23800 6 la_data_in_core[15]
port 38 nsew signal output
rlabel metal2 s 57886 22600 57942 23800 6 la_data_in_core[16]
port 39 nsew signal output
rlabel metal2 s 59358 22600 59414 23800 6 la_data_in_core[17]
port 40 nsew signal output
rlabel metal2 s 60738 22600 60794 23800 6 la_data_in_core[18]
port 41 nsew signal output
rlabel metal2 s 62210 22600 62266 23800 6 la_data_in_core[19]
port 42 nsew signal output
rlabel metal2 s 36450 22600 36506 23800 6 la_data_in_core[1]
port 43 nsew signal output
rlabel metal2 s 63590 22600 63646 23800 6 la_data_in_core[20]
port 44 nsew signal output
rlabel metal2 s 65062 22600 65118 23800 6 la_data_in_core[21]
port 45 nsew signal output
rlabel metal2 s 66442 22600 66498 23800 6 la_data_in_core[22]
port 46 nsew signal output
rlabel metal2 s 67914 22600 67970 23800 6 la_data_in_core[23]
port 47 nsew signal output
rlabel metal2 s 69386 22600 69442 23800 6 la_data_in_core[24]
port 48 nsew signal output
rlabel metal2 s 70766 22600 70822 23800 6 la_data_in_core[25]
port 49 nsew signal output
rlabel metal2 s 72238 22600 72294 23800 6 la_data_in_core[26]
port 50 nsew signal output
rlabel metal2 s 73618 22600 73674 23800 6 la_data_in_core[27]
port 51 nsew signal output
rlabel metal2 s 75090 22600 75146 23800 6 la_data_in_core[28]
port 52 nsew signal output
rlabel metal2 s 76470 22600 76526 23800 6 la_data_in_core[29]
port 53 nsew signal output
rlabel metal2 s 37830 22600 37886 23800 6 la_data_in_core[2]
port 54 nsew signal output
rlabel metal2 s 77942 22600 77998 23800 6 la_data_in_core[30]
port 55 nsew signal output
rlabel metal2 s 79322 22600 79378 23800 6 la_data_in_core[31]
port 56 nsew signal output
rlabel metal2 s 80794 22600 80850 23800 6 la_data_in_core[32]
port 57 nsew signal output
rlabel metal2 s 82266 22600 82322 23800 6 la_data_in_core[33]
port 58 nsew signal output
rlabel metal2 s 83646 22600 83702 23800 6 la_data_in_core[34]
port 59 nsew signal output
rlabel metal2 s 85118 22600 85174 23800 6 la_data_in_core[35]
port 60 nsew signal output
rlabel metal2 s 86498 22600 86554 23800 6 la_data_in_core[36]
port 61 nsew signal output
rlabel metal2 s 87970 22600 88026 23800 6 la_data_in_core[37]
port 62 nsew signal output
rlabel metal2 s 89350 22600 89406 23800 6 la_data_in_core[38]
port 63 nsew signal output
rlabel metal2 s 90822 22600 90878 23800 6 la_data_in_core[39]
port 64 nsew signal output
rlabel metal2 s 39302 22600 39358 23800 6 la_data_in_core[3]
port 65 nsew signal output
rlabel metal2 s 92294 22600 92350 23800 6 la_data_in_core[40]
port 66 nsew signal output
rlabel metal2 s 93674 22600 93730 23800 6 la_data_in_core[41]
port 67 nsew signal output
rlabel metal2 s 95146 22600 95202 23800 6 la_data_in_core[42]
port 68 nsew signal output
rlabel metal2 s 96526 22600 96582 23800 6 la_data_in_core[43]
port 69 nsew signal output
rlabel metal2 s 97998 22600 98054 23800 6 la_data_in_core[44]
port 70 nsew signal output
rlabel metal2 s 99378 22600 99434 23800 6 la_data_in_core[45]
port 71 nsew signal output
rlabel metal2 s 100850 22600 100906 23800 6 la_data_in_core[46]
port 72 nsew signal output
rlabel metal2 s 102230 22600 102286 23800 6 la_data_in_core[47]
port 73 nsew signal output
rlabel metal2 s 103702 22600 103758 23800 6 la_data_in_core[48]
port 74 nsew signal output
rlabel metal2 s 105174 22600 105230 23800 6 la_data_in_core[49]
port 75 nsew signal output
rlabel metal2 s 40682 22600 40738 23800 6 la_data_in_core[4]
port 76 nsew signal output
rlabel metal2 s 106554 22600 106610 23800 6 la_data_in_core[50]
port 77 nsew signal output
rlabel metal2 s 108026 22600 108082 23800 6 la_data_in_core[51]
port 78 nsew signal output
rlabel metal2 s 109406 22600 109462 23800 6 la_data_in_core[52]
port 79 nsew signal output
rlabel metal2 s 110878 22600 110934 23800 6 la_data_in_core[53]
port 80 nsew signal output
rlabel metal2 s 112258 22600 112314 23800 6 la_data_in_core[54]
port 81 nsew signal output
rlabel metal2 s 113730 22600 113786 23800 6 la_data_in_core[55]
port 82 nsew signal output
rlabel metal2 s 115110 22600 115166 23800 6 la_data_in_core[56]
port 83 nsew signal output
rlabel metal2 s 116582 22600 116638 23800 6 la_data_in_core[57]
port 84 nsew signal output
rlabel metal2 s 118054 22600 118110 23800 6 la_data_in_core[58]
port 85 nsew signal output
rlabel metal2 s 119434 22600 119490 23800 6 la_data_in_core[59]
port 86 nsew signal output
rlabel metal2 s 42154 22600 42210 23800 6 la_data_in_core[5]
port 87 nsew signal output
rlabel metal2 s 120906 22600 120962 23800 6 la_data_in_core[60]
port 88 nsew signal output
rlabel metal2 s 122286 22600 122342 23800 6 la_data_in_core[61]
port 89 nsew signal output
rlabel metal2 s 123758 22600 123814 23800 6 la_data_in_core[62]
port 90 nsew signal output
rlabel metal2 s 125138 22600 125194 23800 6 la_data_in_core[63]
port 91 nsew signal output
rlabel metal2 s 126610 22600 126666 23800 6 la_data_in_core[64]
port 92 nsew signal output
rlabel metal2 s 127990 22600 128046 23800 6 la_data_in_core[65]
port 93 nsew signal output
rlabel metal2 s 129462 22600 129518 23800 6 la_data_in_core[66]
port 94 nsew signal output
rlabel metal2 s 130934 22600 130990 23800 6 la_data_in_core[67]
port 95 nsew signal output
rlabel metal2 s 132314 22600 132370 23800 6 la_data_in_core[68]
port 96 nsew signal output
rlabel metal2 s 133786 22600 133842 23800 6 la_data_in_core[69]
port 97 nsew signal output
rlabel metal2 s 43534 22600 43590 23800 6 la_data_in_core[6]
port 98 nsew signal output
rlabel metal2 s 135166 22600 135222 23800 6 la_data_in_core[70]
port 99 nsew signal output
rlabel metal2 s 136638 22600 136694 23800 6 la_data_in_core[71]
port 100 nsew signal output
rlabel metal2 s 138018 22600 138074 23800 6 la_data_in_core[72]
port 101 nsew signal output
rlabel metal2 s 139490 22600 139546 23800 6 la_data_in_core[73]
port 102 nsew signal output
rlabel metal2 s 140962 22600 141018 23800 6 la_data_in_core[74]
port 103 nsew signal output
rlabel metal2 s 142342 22600 142398 23800 6 la_data_in_core[75]
port 104 nsew signal output
rlabel metal2 s 143814 22600 143870 23800 6 la_data_in_core[76]
port 105 nsew signal output
rlabel metal2 s 145194 22600 145250 23800 6 la_data_in_core[77]
port 106 nsew signal output
rlabel metal2 s 146666 22600 146722 23800 6 la_data_in_core[78]
port 107 nsew signal output
rlabel metal2 s 148046 22600 148102 23800 6 la_data_in_core[79]
port 108 nsew signal output
rlabel metal2 s 45006 22600 45062 23800 6 la_data_in_core[7]
port 109 nsew signal output
rlabel metal2 s 149518 22600 149574 23800 6 la_data_in_core[80]
port 110 nsew signal output
rlabel metal2 s 150898 22600 150954 23800 6 la_data_in_core[81]
port 111 nsew signal output
rlabel metal2 s 152370 22600 152426 23800 6 la_data_in_core[82]
port 112 nsew signal output
rlabel metal2 s 153842 22600 153898 23800 6 la_data_in_core[83]
port 113 nsew signal output
rlabel metal2 s 155222 22600 155278 23800 6 la_data_in_core[84]
port 114 nsew signal output
rlabel metal2 s 156694 22600 156750 23800 6 la_data_in_core[85]
port 115 nsew signal output
rlabel metal2 s 158074 22600 158130 23800 6 la_data_in_core[86]
port 116 nsew signal output
rlabel metal2 s 159546 22600 159602 23800 6 la_data_in_core[87]
port 117 nsew signal output
rlabel metal2 s 160926 22600 160982 23800 6 la_data_in_core[88]
port 118 nsew signal output
rlabel metal2 s 162398 22600 162454 23800 6 la_data_in_core[89]
port 119 nsew signal output
rlabel metal2 s 46478 22600 46534 23800 6 la_data_in_core[8]
port 120 nsew signal output
rlabel metal2 s 163778 22600 163834 23800 6 la_data_in_core[90]
port 121 nsew signal output
rlabel metal2 s 165250 22600 165306 23800 6 la_data_in_core[91]
port 122 nsew signal output
rlabel metal2 s 166722 22600 166778 23800 6 la_data_in_core[92]
port 123 nsew signal output
rlabel metal2 s 168102 22600 168158 23800 6 la_data_in_core[93]
port 124 nsew signal output
rlabel metal2 s 169574 22600 169630 23800 6 la_data_in_core[94]
port 125 nsew signal output
rlabel metal2 s 170954 22600 171010 23800 6 la_data_in_core[95]
port 126 nsew signal output
rlabel metal2 s 172426 22600 172482 23800 6 la_data_in_core[96]
port 127 nsew signal output
rlabel metal2 s 173806 22600 173862 23800 6 la_data_in_core[97]
port 128 nsew signal output
rlabel metal2 s 175278 22600 175334 23800 6 la_data_in_core[98]
port 129 nsew signal output
rlabel metal2 s 176750 22600 176806 23800 6 la_data_in_core[99]
port 130 nsew signal output
rlabel metal2 s 47858 22600 47914 23800 6 la_data_in_core[9]
port 131 nsew signal output
rlabel metal2 s 202 -400 258 800 6 la_data_in_mprj[0]
port 132 nsew signal output
rlabel metal2 s 151082 -400 151138 800 6 la_data_in_mprj[100]
port 133 nsew signal output
rlabel metal2 s 152554 -400 152610 800 6 la_data_in_mprj[101]
port 134 nsew signal output
rlabel metal2 s 154118 -400 154174 800 6 la_data_in_mprj[102]
port 135 nsew signal output
rlabel metal2 s 155590 -400 155646 800 6 la_data_in_mprj[103]
port 136 nsew signal output
rlabel metal2 s 157154 -400 157210 800 6 la_data_in_mprj[104]
port 137 nsew signal output
rlabel metal2 s 158626 -400 158682 800 6 la_data_in_mprj[105]
port 138 nsew signal output
rlabel metal2 s 160098 -400 160154 800 6 la_data_in_mprj[106]
port 139 nsew signal output
rlabel metal2 s 161662 -400 161718 800 6 la_data_in_mprj[107]
port 140 nsew signal output
rlabel metal2 s 163134 -400 163190 800 6 la_data_in_mprj[108]
port 141 nsew signal output
rlabel metal2 s 164698 -400 164754 800 6 la_data_in_mprj[109]
port 142 nsew signal output
rlabel metal2 s 15290 -400 15346 800 6 la_data_in_mprj[10]
port 143 nsew signal output
rlabel metal2 s 166170 -400 166226 800 6 la_data_in_mprj[110]
port 144 nsew signal output
rlabel metal2 s 167642 -400 167698 800 6 la_data_in_mprj[111]
port 145 nsew signal output
rlabel metal2 s 169206 -400 169262 800 6 la_data_in_mprj[112]
port 146 nsew signal output
rlabel metal2 s 170678 -400 170734 800 6 la_data_in_mprj[113]
port 147 nsew signal output
rlabel metal2 s 172242 -400 172298 800 6 la_data_in_mprj[114]
port 148 nsew signal output
rlabel metal2 s 173714 -400 173770 800 6 la_data_in_mprj[115]
port 149 nsew signal output
rlabel metal2 s 175186 -400 175242 800 6 la_data_in_mprj[116]
port 150 nsew signal output
rlabel metal2 s 176750 -400 176806 800 6 la_data_in_mprj[117]
port 151 nsew signal output
rlabel metal2 s 178222 -400 178278 800 6 la_data_in_mprj[118]
port 152 nsew signal output
rlabel metal2 s 179786 -400 179842 800 6 la_data_in_mprj[119]
port 153 nsew signal output
rlabel metal2 s 16762 -400 16818 800 6 la_data_in_mprj[11]
port 154 nsew signal output
rlabel metal2 s 181258 -400 181314 800 6 la_data_in_mprj[120]
port 155 nsew signal output
rlabel metal2 s 182730 -400 182786 800 6 la_data_in_mprj[121]
port 156 nsew signal output
rlabel metal2 s 184294 -400 184350 800 6 la_data_in_mprj[122]
port 157 nsew signal output
rlabel metal2 s 185766 -400 185822 800 6 la_data_in_mprj[123]
port 158 nsew signal output
rlabel metal2 s 187330 -400 187386 800 6 la_data_in_mprj[124]
port 159 nsew signal output
rlabel metal2 s 188802 -400 188858 800 6 la_data_in_mprj[125]
port 160 nsew signal output
rlabel metal2 s 190366 -400 190422 800 6 la_data_in_mprj[126]
port 161 nsew signal output
rlabel metal2 s 191838 -400 191894 800 6 la_data_in_mprj[127]
port 162 nsew signal output
rlabel metal2 s 18234 -400 18290 800 6 la_data_in_mprj[12]
port 163 nsew signal output
rlabel metal2 s 19798 -400 19854 800 6 la_data_in_mprj[13]
port 164 nsew signal output
rlabel metal2 s 21270 -400 21326 800 6 la_data_in_mprj[14]
port 165 nsew signal output
rlabel metal2 s 22834 -400 22890 800 6 la_data_in_mprj[15]
port 166 nsew signal output
rlabel metal2 s 24306 -400 24362 800 6 la_data_in_mprj[16]
port 167 nsew signal output
rlabel metal2 s 25778 -400 25834 800 6 la_data_in_mprj[17]
port 168 nsew signal output
rlabel metal2 s 27342 -400 27398 800 6 la_data_in_mprj[18]
port 169 nsew signal output
rlabel metal2 s 28814 -400 28870 800 6 la_data_in_mprj[19]
port 170 nsew signal output
rlabel metal2 s 1674 -400 1730 800 6 la_data_in_mprj[1]
port 171 nsew signal output
rlabel metal2 s 30378 -400 30434 800 6 la_data_in_mprj[20]
port 172 nsew signal output
rlabel metal2 s 31850 -400 31906 800 6 la_data_in_mprj[21]
port 173 nsew signal output
rlabel metal2 s 33322 -400 33378 800 6 la_data_in_mprj[22]
port 174 nsew signal output
rlabel metal2 s 34886 -400 34942 800 6 la_data_in_mprj[23]
port 175 nsew signal output
rlabel metal2 s 36358 -400 36414 800 6 la_data_in_mprj[24]
port 176 nsew signal output
rlabel metal2 s 37922 -400 37978 800 6 la_data_in_mprj[25]
port 177 nsew signal output
rlabel metal2 s 39394 -400 39450 800 6 la_data_in_mprj[26]
port 178 nsew signal output
rlabel metal2 s 40866 -400 40922 800 6 la_data_in_mprj[27]
port 179 nsew signal output
rlabel metal2 s 42430 -400 42486 800 6 la_data_in_mprj[28]
port 180 nsew signal output
rlabel metal2 s 43902 -400 43958 800 6 la_data_in_mprj[29]
port 181 nsew signal output
rlabel metal2 s 3146 -400 3202 800 6 la_data_in_mprj[2]
port 182 nsew signal output
rlabel metal2 s 45466 -400 45522 800 6 la_data_in_mprj[30]
port 183 nsew signal output
rlabel metal2 s 46938 -400 46994 800 6 la_data_in_mprj[31]
port 184 nsew signal output
rlabel metal2 s 48410 -400 48466 800 6 la_data_in_mprj[32]
port 185 nsew signal output
rlabel metal2 s 49974 -400 50030 800 6 la_data_in_mprj[33]
port 186 nsew signal output
rlabel metal2 s 51446 -400 51502 800 6 la_data_in_mprj[34]
port 187 nsew signal output
rlabel metal2 s 53010 -400 53066 800 6 la_data_in_mprj[35]
port 188 nsew signal output
rlabel metal2 s 54482 -400 54538 800 6 la_data_in_mprj[36]
port 189 nsew signal output
rlabel metal2 s 55954 -400 56010 800 6 la_data_in_mprj[37]
port 190 nsew signal output
rlabel metal2 s 57518 -400 57574 800 6 la_data_in_mprj[38]
port 191 nsew signal output
rlabel metal2 s 58990 -400 59046 800 6 la_data_in_mprj[39]
port 192 nsew signal output
rlabel metal2 s 4710 -400 4766 800 6 la_data_in_mprj[3]
port 193 nsew signal output
rlabel metal2 s 60554 -400 60610 800 6 la_data_in_mprj[40]
port 194 nsew signal output
rlabel metal2 s 62026 -400 62082 800 6 la_data_in_mprj[41]
port 195 nsew signal output
rlabel metal2 s 63590 -400 63646 800 6 la_data_in_mprj[42]
port 196 nsew signal output
rlabel metal2 s 65062 -400 65118 800 6 la_data_in_mprj[43]
port 197 nsew signal output
rlabel metal2 s 66534 -400 66590 800 6 la_data_in_mprj[44]
port 198 nsew signal output
rlabel metal2 s 68098 -400 68154 800 6 la_data_in_mprj[45]
port 199 nsew signal output
rlabel metal2 s 69570 -400 69626 800 6 la_data_in_mprj[46]
port 200 nsew signal output
rlabel metal2 s 71134 -400 71190 800 6 la_data_in_mprj[47]
port 201 nsew signal output
rlabel metal2 s 72606 -400 72662 800 6 la_data_in_mprj[48]
port 202 nsew signal output
rlabel metal2 s 74078 -400 74134 800 6 la_data_in_mprj[49]
port 203 nsew signal output
rlabel metal2 s 6182 -400 6238 800 6 la_data_in_mprj[4]
port 204 nsew signal output
rlabel metal2 s 75642 -400 75698 800 6 la_data_in_mprj[50]
port 205 nsew signal output
rlabel metal2 s 77114 -400 77170 800 6 la_data_in_mprj[51]
port 206 nsew signal output
rlabel metal2 s 78678 -400 78734 800 6 la_data_in_mprj[52]
port 207 nsew signal output
rlabel metal2 s 80150 -400 80206 800 6 la_data_in_mprj[53]
port 208 nsew signal output
rlabel metal2 s 81622 -400 81678 800 6 la_data_in_mprj[54]
port 209 nsew signal output
rlabel metal2 s 83186 -400 83242 800 6 la_data_in_mprj[55]
port 210 nsew signal output
rlabel metal2 s 84658 -400 84714 800 6 la_data_in_mprj[56]
port 211 nsew signal output
rlabel metal2 s 86222 -400 86278 800 6 la_data_in_mprj[57]
port 212 nsew signal output
rlabel metal2 s 87694 -400 87750 800 6 la_data_in_mprj[58]
port 213 nsew signal output
rlabel metal2 s 89166 -400 89222 800 6 la_data_in_mprj[59]
port 214 nsew signal output
rlabel metal2 s 7746 -400 7802 800 6 la_data_in_mprj[5]
port 215 nsew signal output
rlabel metal2 s 90730 -400 90786 800 6 la_data_in_mprj[60]
port 216 nsew signal output
rlabel metal2 s 92202 -400 92258 800 6 la_data_in_mprj[61]
port 217 nsew signal output
rlabel metal2 s 93766 -400 93822 800 6 la_data_in_mprj[62]
port 218 nsew signal output
rlabel metal2 s 95238 -400 95294 800 6 la_data_in_mprj[63]
port 219 nsew signal output
rlabel metal2 s 96710 -400 96766 800 6 la_data_in_mprj[64]
port 220 nsew signal output
rlabel metal2 s 98274 -400 98330 800 6 la_data_in_mprj[65]
port 221 nsew signal output
rlabel metal2 s 99746 -400 99802 800 6 la_data_in_mprj[66]
port 222 nsew signal output
rlabel metal2 s 101310 -400 101366 800 6 la_data_in_mprj[67]
port 223 nsew signal output
rlabel metal2 s 102782 -400 102838 800 6 la_data_in_mprj[68]
port 224 nsew signal output
rlabel metal2 s 104254 -400 104310 800 6 la_data_in_mprj[69]
port 225 nsew signal output
rlabel metal2 s 9218 -400 9274 800 6 la_data_in_mprj[6]
port 226 nsew signal output
rlabel metal2 s 105818 -400 105874 800 6 la_data_in_mprj[70]
port 227 nsew signal output
rlabel metal2 s 107290 -400 107346 800 6 la_data_in_mprj[71]
port 228 nsew signal output
rlabel metal2 s 108854 -400 108910 800 6 la_data_in_mprj[72]
port 229 nsew signal output
rlabel metal2 s 110326 -400 110382 800 6 la_data_in_mprj[73]
port 230 nsew signal output
rlabel metal2 s 111798 -400 111854 800 6 la_data_in_mprj[74]
port 231 nsew signal output
rlabel metal2 s 113362 -400 113418 800 6 la_data_in_mprj[75]
port 232 nsew signal output
rlabel metal2 s 114834 -400 114890 800 6 la_data_in_mprj[76]
port 233 nsew signal output
rlabel metal2 s 116398 -400 116454 800 6 la_data_in_mprj[77]
port 234 nsew signal output
rlabel metal2 s 117870 -400 117926 800 6 la_data_in_mprj[78]
port 235 nsew signal output
rlabel metal2 s 119342 -400 119398 800 6 la_data_in_mprj[79]
port 236 nsew signal output
rlabel metal2 s 10690 -400 10746 800 6 la_data_in_mprj[7]
port 237 nsew signal output
rlabel metal2 s 120906 -400 120962 800 6 la_data_in_mprj[80]
port 238 nsew signal output
rlabel metal2 s 122378 -400 122434 800 6 la_data_in_mprj[81]
port 239 nsew signal output
rlabel metal2 s 123942 -400 123998 800 6 la_data_in_mprj[82]
port 240 nsew signal output
rlabel metal2 s 125414 -400 125470 800 6 la_data_in_mprj[83]
port 241 nsew signal output
rlabel metal2 s 126978 -400 127034 800 6 la_data_in_mprj[84]
port 242 nsew signal output
rlabel metal2 s 128450 -400 128506 800 6 la_data_in_mprj[85]
port 243 nsew signal output
rlabel metal2 s 129922 -400 129978 800 6 la_data_in_mprj[86]
port 244 nsew signal output
rlabel metal2 s 131486 -400 131542 800 6 la_data_in_mprj[87]
port 245 nsew signal output
rlabel metal2 s 132958 -400 133014 800 6 la_data_in_mprj[88]
port 246 nsew signal output
rlabel metal2 s 134522 -400 134578 800 6 la_data_in_mprj[89]
port 247 nsew signal output
rlabel metal2 s 12254 -400 12310 800 6 la_data_in_mprj[8]
port 248 nsew signal output
rlabel metal2 s 135994 -400 136050 800 6 la_data_in_mprj[90]
port 249 nsew signal output
rlabel metal2 s 137466 -400 137522 800 6 la_data_in_mprj[91]
port 250 nsew signal output
rlabel metal2 s 139030 -400 139086 800 6 la_data_in_mprj[92]
port 251 nsew signal output
rlabel metal2 s 140502 -400 140558 800 6 la_data_in_mprj[93]
port 252 nsew signal output
rlabel metal2 s 142066 -400 142122 800 6 la_data_in_mprj[94]
port 253 nsew signal output
rlabel metal2 s 143538 -400 143594 800 6 la_data_in_mprj[95]
port 254 nsew signal output
rlabel metal2 s 145010 -400 145066 800 6 la_data_in_mprj[96]
port 255 nsew signal output
rlabel metal2 s 146574 -400 146630 800 6 la_data_in_mprj[97]
port 256 nsew signal output
rlabel metal2 s 148046 -400 148102 800 6 la_data_in_mprj[98]
port 257 nsew signal output
rlabel metal2 s 149610 -400 149666 800 6 la_data_in_mprj[99]
port 258 nsew signal output
rlabel metal2 s 13726 -400 13782 800 6 la_data_in_mprj[9]
port 259 nsew signal output
rlabel metal2 s 35438 22600 35494 23800 6 la_data_out_core[0]
port 260 nsew signal input
rlabel metal2 s 178590 22600 178646 23800 6 la_data_out_core[100]
port 261 nsew signal input
rlabel metal2 s 180062 22600 180118 23800 6 la_data_out_core[101]
port 262 nsew signal input
rlabel metal2 s 181442 22600 181498 23800 6 la_data_out_core[102]
port 263 nsew signal input
rlabel metal2 s 182914 22600 182970 23800 6 la_data_out_core[103]
port 264 nsew signal input
rlabel metal2 s 184386 22600 184442 23800 6 la_data_out_core[104]
port 265 nsew signal input
rlabel metal2 s 185766 22600 185822 23800 6 la_data_out_core[105]
port 266 nsew signal input
rlabel metal2 s 187238 22600 187294 23800 6 la_data_out_core[106]
port 267 nsew signal input
rlabel metal2 s 188618 22600 188674 23800 6 la_data_out_core[107]
port 268 nsew signal input
rlabel metal2 s 190090 22600 190146 23800 6 la_data_out_core[108]
port 269 nsew signal input
rlabel metal2 s 191470 22600 191526 23800 6 la_data_out_core[109]
port 270 nsew signal input
rlabel metal2 s 49790 22600 49846 23800 6 la_data_out_core[10]
port 271 nsew signal input
rlabel metal2 s 192942 22600 192998 23800 6 la_data_out_core[110]
port 272 nsew signal input
rlabel metal2 s 194322 22600 194378 23800 6 la_data_out_core[111]
port 273 nsew signal input
rlabel metal2 s 195794 22600 195850 23800 6 la_data_out_core[112]
port 274 nsew signal input
rlabel metal2 s 197266 22600 197322 23800 6 la_data_out_core[113]
port 275 nsew signal input
rlabel metal2 s 198646 22600 198702 23800 6 la_data_out_core[114]
port 276 nsew signal input
rlabel metal2 s 200118 22600 200174 23800 6 la_data_out_core[115]
port 277 nsew signal input
rlabel metal2 s 201498 22600 201554 23800 6 la_data_out_core[116]
port 278 nsew signal input
rlabel metal2 s 202970 22600 203026 23800 6 la_data_out_core[117]
port 279 nsew signal input
rlabel metal2 s 204350 22600 204406 23800 6 la_data_out_core[118]
port 280 nsew signal input
rlabel metal2 s 205822 22600 205878 23800 6 la_data_out_core[119]
port 281 nsew signal input
rlabel metal2 s 51170 22600 51226 23800 6 la_data_out_core[11]
port 282 nsew signal input
rlabel metal2 s 207202 22600 207258 23800 6 la_data_out_core[120]
port 283 nsew signal input
rlabel metal2 s 208674 22600 208730 23800 6 la_data_out_core[121]
port 284 nsew signal input
rlabel metal2 s 210146 22600 210202 23800 6 la_data_out_core[122]
port 285 nsew signal input
rlabel metal2 s 211526 22600 211582 23800 6 la_data_out_core[123]
port 286 nsew signal input
rlabel metal2 s 212998 22600 213054 23800 6 la_data_out_core[124]
port 287 nsew signal input
rlabel metal2 s 214378 22600 214434 23800 6 la_data_out_core[125]
port 288 nsew signal input
rlabel metal2 s 215850 22600 215906 23800 6 la_data_out_core[126]
port 289 nsew signal input
rlabel metal2 s 217230 22600 217286 23800 6 la_data_out_core[127]
port 290 nsew signal input
rlabel metal2 s 52642 22600 52698 23800 6 la_data_out_core[12]
port 291 nsew signal input
rlabel metal2 s 54114 22600 54170 23800 6 la_data_out_core[13]
port 292 nsew signal input
rlabel metal2 s 55494 22600 55550 23800 6 la_data_out_core[14]
port 293 nsew signal input
rlabel metal2 s 56966 22600 57022 23800 6 la_data_out_core[15]
port 294 nsew signal input
rlabel metal2 s 58346 22600 58402 23800 6 la_data_out_core[16]
port 295 nsew signal input
rlabel metal2 s 59818 22600 59874 23800 6 la_data_out_core[17]
port 296 nsew signal input
rlabel metal2 s 61198 22600 61254 23800 6 la_data_out_core[18]
port 297 nsew signal input
rlabel metal2 s 62670 22600 62726 23800 6 la_data_out_core[19]
port 298 nsew signal input
rlabel metal2 s 36910 22600 36966 23800 6 la_data_out_core[1]
port 299 nsew signal input
rlabel metal2 s 64050 22600 64106 23800 6 la_data_out_core[20]
port 300 nsew signal input
rlabel metal2 s 65522 22600 65578 23800 6 la_data_out_core[21]
port 301 nsew signal input
rlabel metal2 s 66994 22600 67050 23800 6 la_data_out_core[22]
port 302 nsew signal input
rlabel metal2 s 68374 22600 68430 23800 6 la_data_out_core[23]
port 303 nsew signal input
rlabel metal2 s 69846 22600 69902 23800 6 la_data_out_core[24]
port 304 nsew signal input
rlabel metal2 s 71226 22600 71282 23800 6 la_data_out_core[25]
port 305 nsew signal input
rlabel metal2 s 72698 22600 72754 23800 6 la_data_out_core[26]
port 306 nsew signal input
rlabel metal2 s 74078 22600 74134 23800 6 la_data_out_core[27]
port 307 nsew signal input
rlabel metal2 s 75550 22600 75606 23800 6 la_data_out_core[28]
port 308 nsew signal input
rlabel metal2 s 77022 22600 77078 23800 6 la_data_out_core[29]
port 309 nsew signal input
rlabel metal2 s 38290 22600 38346 23800 6 la_data_out_core[2]
port 310 nsew signal input
rlabel metal2 s 78402 22600 78458 23800 6 la_data_out_core[30]
port 311 nsew signal input
rlabel metal2 s 79874 22600 79930 23800 6 la_data_out_core[31]
port 312 nsew signal input
rlabel metal2 s 81254 22600 81310 23800 6 la_data_out_core[32]
port 313 nsew signal input
rlabel metal2 s 82726 22600 82782 23800 6 la_data_out_core[33]
port 314 nsew signal input
rlabel metal2 s 84106 22600 84162 23800 6 la_data_out_core[34]
port 315 nsew signal input
rlabel metal2 s 85578 22600 85634 23800 6 la_data_out_core[35]
port 316 nsew signal input
rlabel metal2 s 86958 22600 87014 23800 6 la_data_out_core[36]
port 317 nsew signal input
rlabel metal2 s 88430 22600 88486 23800 6 la_data_out_core[37]
port 318 nsew signal input
rlabel metal2 s 89902 22600 89958 23800 6 la_data_out_core[38]
port 319 nsew signal input
rlabel metal2 s 91282 22600 91338 23800 6 la_data_out_core[39]
port 320 nsew signal input
rlabel metal2 s 39762 22600 39818 23800 6 la_data_out_core[3]
port 321 nsew signal input
rlabel metal2 s 92754 22600 92810 23800 6 la_data_out_core[40]
port 322 nsew signal input
rlabel metal2 s 94134 22600 94190 23800 6 la_data_out_core[41]
port 323 nsew signal input
rlabel metal2 s 95606 22600 95662 23800 6 la_data_out_core[42]
port 324 nsew signal input
rlabel metal2 s 96986 22600 97042 23800 6 la_data_out_core[43]
port 325 nsew signal input
rlabel metal2 s 98458 22600 98514 23800 6 la_data_out_core[44]
port 326 nsew signal input
rlabel metal2 s 99838 22600 99894 23800 6 la_data_out_core[45]
port 327 nsew signal input
rlabel metal2 s 101310 22600 101366 23800 6 la_data_out_core[46]
port 328 nsew signal input
rlabel metal2 s 102782 22600 102838 23800 6 la_data_out_core[47]
port 329 nsew signal input
rlabel metal2 s 104162 22600 104218 23800 6 la_data_out_core[48]
port 330 nsew signal input
rlabel metal2 s 105634 22600 105690 23800 6 la_data_out_core[49]
port 331 nsew signal input
rlabel metal2 s 41234 22600 41290 23800 6 la_data_out_core[4]
port 332 nsew signal input
rlabel metal2 s 107014 22600 107070 23800 6 la_data_out_core[50]
port 333 nsew signal input
rlabel metal2 s 108486 22600 108542 23800 6 la_data_out_core[51]
port 334 nsew signal input
rlabel metal2 s 109866 22600 109922 23800 6 la_data_out_core[52]
port 335 nsew signal input
rlabel metal2 s 111338 22600 111394 23800 6 la_data_out_core[53]
port 336 nsew signal input
rlabel metal2 s 112810 22600 112866 23800 6 la_data_out_core[54]
port 337 nsew signal input
rlabel metal2 s 114190 22600 114246 23800 6 la_data_out_core[55]
port 338 nsew signal input
rlabel metal2 s 115662 22600 115718 23800 6 la_data_out_core[56]
port 339 nsew signal input
rlabel metal2 s 117042 22600 117098 23800 6 la_data_out_core[57]
port 340 nsew signal input
rlabel metal2 s 118514 22600 118570 23800 6 la_data_out_core[58]
port 341 nsew signal input
rlabel metal2 s 119894 22600 119950 23800 6 la_data_out_core[59]
port 342 nsew signal input
rlabel metal2 s 42614 22600 42670 23800 6 la_data_out_core[5]
port 343 nsew signal input
rlabel metal2 s 121366 22600 121422 23800 6 la_data_out_core[60]
port 344 nsew signal input
rlabel metal2 s 122746 22600 122802 23800 6 la_data_out_core[61]
port 345 nsew signal input
rlabel metal2 s 124218 22600 124274 23800 6 la_data_out_core[62]
port 346 nsew signal input
rlabel metal2 s 125690 22600 125746 23800 6 la_data_out_core[63]
port 347 nsew signal input
rlabel metal2 s 127070 22600 127126 23800 6 la_data_out_core[64]
port 348 nsew signal input
rlabel metal2 s 128542 22600 128598 23800 6 la_data_out_core[65]
port 349 nsew signal input
rlabel metal2 s 129922 22600 129978 23800 6 la_data_out_core[66]
port 350 nsew signal input
rlabel metal2 s 131394 22600 131450 23800 6 la_data_out_core[67]
port 351 nsew signal input
rlabel metal2 s 132774 22600 132830 23800 6 la_data_out_core[68]
port 352 nsew signal input
rlabel metal2 s 134246 22600 134302 23800 6 la_data_out_core[69]
port 353 nsew signal input
rlabel metal2 s 44086 22600 44142 23800 6 la_data_out_core[6]
port 354 nsew signal input
rlabel metal2 s 135626 22600 135682 23800 6 la_data_out_core[70]
port 355 nsew signal input
rlabel metal2 s 137098 22600 137154 23800 6 la_data_out_core[71]
port 356 nsew signal input
rlabel metal2 s 138570 22600 138626 23800 6 la_data_out_core[72]
port 357 nsew signal input
rlabel metal2 s 139950 22600 140006 23800 6 la_data_out_core[73]
port 358 nsew signal input
rlabel metal2 s 141422 22600 141478 23800 6 la_data_out_core[74]
port 359 nsew signal input
rlabel metal2 s 142802 22600 142858 23800 6 la_data_out_core[75]
port 360 nsew signal input
rlabel metal2 s 144274 22600 144330 23800 6 la_data_out_core[76]
port 361 nsew signal input
rlabel metal2 s 145654 22600 145710 23800 6 la_data_out_core[77]
port 362 nsew signal input
rlabel metal2 s 147126 22600 147182 23800 6 la_data_out_core[78]
port 363 nsew signal input
rlabel metal2 s 148598 22600 148654 23800 6 la_data_out_core[79]
port 364 nsew signal input
rlabel metal2 s 45466 22600 45522 23800 6 la_data_out_core[7]
port 365 nsew signal input
rlabel metal2 s 149978 22600 150034 23800 6 la_data_out_core[80]
port 366 nsew signal input
rlabel metal2 s 151450 22600 151506 23800 6 la_data_out_core[81]
port 367 nsew signal input
rlabel metal2 s 152830 22600 152886 23800 6 la_data_out_core[82]
port 368 nsew signal input
rlabel metal2 s 154302 22600 154358 23800 6 la_data_out_core[83]
port 369 nsew signal input
rlabel metal2 s 155682 22600 155738 23800 6 la_data_out_core[84]
port 370 nsew signal input
rlabel metal2 s 157154 22600 157210 23800 6 la_data_out_core[85]
port 371 nsew signal input
rlabel metal2 s 158534 22600 158590 23800 6 la_data_out_core[86]
port 372 nsew signal input
rlabel metal2 s 160006 22600 160062 23800 6 la_data_out_core[87]
port 373 nsew signal input
rlabel metal2 s 161478 22600 161534 23800 6 la_data_out_core[88]
port 374 nsew signal input
rlabel metal2 s 162858 22600 162914 23800 6 la_data_out_core[89]
port 375 nsew signal input
rlabel metal2 s 46938 22600 46994 23800 6 la_data_out_core[8]
port 376 nsew signal input
rlabel metal2 s 164330 22600 164386 23800 6 la_data_out_core[90]
port 377 nsew signal input
rlabel metal2 s 165710 22600 165766 23800 6 la_data_out_core[91]
port 378 nsew signal input
rlabel metal2 s 167182 22600 167238 23800 6 la_data_out_core[92]
port 379 nsew signal input
rlabel metal2 s 168562 22600 168618 23800 6 la_data_out_core[93]
port 380 nsew signal input
rlabel metal2 s 170034 22600 170090 23800 6 la_data_out_core[94]
port 381 nsew signal input
rlabel metal2 s 171414 22600 171470 23800 6 la_data_out_core[95]
port 382 nsew signal input
rlabel metal2 s 172886 22600 172942 23800 6 la_data_out_core[96]
port 383 nsew signal input
rlabel metal2 s 174358 22600 174414 23800 6 la_data_out_core[97]
port 384 nsew signal input
rlabel metal2 s 175738 22600 175794 23800 6 la_data_out_core[98]
port 385 nsew signal input
rlabel metal2 s 177210 22600 177266 23800 6 la_data_out_core[99]
port 386 nsew signal input
rlabel metal2 s 48318 22600 48374 23800 6 la_data_out_core[9]
port 387 nsew signal input
rlabel metal2 s 570 -400 626 800 6 la_data_out_mprj[0]
port 388 nsew signal input
rlabel metal2 s 151450 -400 151506 800 6 la_data_out_mprj[100]
port 389 nsew signal input
rlabel metal2 s 152922 -400 152978 800 6 la_data_out_mprj[101]
port 390 nsew signal input
rlabel metal2 s 154486 -400 154542 800 6 la_data_out_mprj[102]
port 391 nsew signal input
rlabel metal2 s 155958 -400 156014 800 6 la_data_out_mprj[103]
port 392 nsew signal input
rlabel metal2 s 157522 -400 157578 800 6 la_data_out_mprj[104]
port 393 nsew signal input
rlabel metal2 s 158994 -400 159050 800 6 la_data_out_mprj[105]
port 394 nsew signal input
rlabel metal2 s 160558 -400 160614 800 6 la_data_out_mprj[106]
port 395 nsew signal input
rlabel metal2 s 162030 -400 162086 800 6 la_data_out_mprj[107]
port 396 nsew signal input
rlabel metal2 s 163502 -400 163558 800 6 la_data_out_mprj[108]
port 397 nsew signal input
rlabel metal2 s 165066 -400 165122 800 6 la_data_out_mprj[109]
port 398 nsew signal input
rlabel metal2 s 15658 -400 15714 800 6 la_data_out_mprj[10]
port 399 nsew signal input
rlabel metal2 s 166538 -400 166594 800 6 la_data_out_mprj[110]
port 400 nsew signal input
rlabel metal2 s 168102 -400 168158 800 6 la_data_out_mprj[111]
port 401 nsew signal input
rlabel metal2 s 169574 -400 169630 800 6 la_data_out_mprj[112]
port 402 nsew signal input
rlabel metal2 s 171046 -400 171102 800 6 la_data_out_mprj[113]
port 403 nsew signal input
rlabel metal2 s 172610 -400 172666 800 6 la_data_out_mprj[114]
port 404 nsew signal input
rlabel metal2 s 174082 -400 174138 800 6 la_data_out_mprj[115]
port 405 nsew signal input
rlabel metal2 s 175646 -400 175702 800 6 la_data_out_mprj[116]
port 406 nsew signal input
rlabel metal2 s 177118 -400 177174 800 6 la_data_out_mprj[117]
port 407 nsew signal input
rlabel metal2 s 178590 -400 178646 800 6 la_data_out_mprj[118]
port 408 nsew signal input
rlabel metal2 s 180154 -400 180210 800 6 la_data_out_mprj[119]
port 409 nsew signal input
rlabel metal2 s 17130 -400 17186 800 6 la_data_out_mprj[11]
port 410 nsew signal input
rlabel metal2 s 181626 -400 181682 800 6 la_data_out_mprj[120]
port 411 nsew signal input
rlabel metal2 s 183190 -400 183246 800 6 la_data_out_mprj[121]
port 412 nsew signal input
rlabel metal2 s 184662 -400 184718 800 6 la_data_out_mprj[122]
port 413 nsew signal input
rlabel metal2 s 186134 -400 186190 800 6 la_data_out_mprj[123]
port 414 nsew signal input
rlabel metal2 s 187698 -400 187754 800 6 la_data_out_mprj[124]
port 415 nsew signal input
rlabel metal2 s 189170 -400 189226 800 6 la_data_out_mprj[125]
port 416 nsew signal input
rlabel metal2 s 190734 -400 190790 800 6 la_data_out_mprj[126]
port 417 nsew signal input
rlabel metal2 s 192206 -400 192262 800 6 la_data_out_mprj[127]
port 418 nsew signal input
rlabel metal2 s 18602 -400 18658 800 6 la_data_out_mprj[12]
port 419 nsew signal input
rlabel metal2 s 20166 -400 20222 800 6 la_data_out_mprj[13]
port 420 nsew signal input
rlabel metal2 s 21638 -400 21694 800 6 la_data_out_mprj[14]
port 421 nsew signal input
rlabel metal2 s 23202 -400 23258 800 6 la_data_out_mprj[15]
port 422 nsew signal input
rlabel metal2 s 24674 -400 24730 800 6 la_data_out_mprj[16]
port 423 nsew signal input
rlabel metal2 s 26146 -400 26202 800 6 la_data_out_mprj[17]
port 424 nsew signal input
rlabel metal2 s 27710 -400 27766 800 6 la_data_out_mprj[18]
port 425 nsew signal input
rlabel metal2 s 29182 -400 29238 800 6 la_data_out_mprj[19]
port 426 nsew signal input
rlabel metal2 s 2042 -400 2098 800 6 la_data_out_mprj[1]
port 427 nsew signal input
rlabel metal2 s 30746 -400 30802 800 6 la_data_out_mprj[20]
port 428 nsew signal input
rlabel metal2 s 32218 -400 32274 800 6 la_data_out_mprj[21]
port 429 nsew signal input
rlabel metal2 s 33782 -400 33838 800 6 la_data_out_mprj[22]
port 430 nsew signal input
rlabel metal2 s 35254 -400 35310 800 6 la_data_out_mprj[23]
port 431 nsew signal input
rlabel metal2 s 36726 -400 36782 800 6 la_data_out_mprj[24]
port 432 nsew signal input
rlabel metal2 s 38290 -400 38346 800 6 la_data_out_mprj[25]
port 433 nsew signal input
rlabel metal2 s 39762 -400 39818 800 6 la_data_out_mprj[26]
port 434 nsew signal input
rlabel metal2 s 41326 -400 41382 800 6 la_data_out_mprj[27]
port 435 nsew signal input
rlabel metal2 s 42798 -400 42854 800 6 la_data_out_mprj[28]
port 436 nsew signal input
rlabel metal2 s 44270 -400 44326 800 6 la_data_out_mprj[29]
port 437 nsew signal input
rlabel metal2 s 3514 -400 3570 800 6 la_data_out_mprj[2]
port 438 nsew signal input
rlabel metal2 s 45834 -400 45890 800 6 la_data_out_mprj[30]
port 439 nsew signal input
rlabel metal2 s 47306 -400 47362 800 6 la_data_out_mprj[31]
port 440 nsew signal input
rlabel metal2 s 48870 -400 48926 800 6 la_data_out_mprj[32]
port 441 nsew signal input
rlabel metal2 s 50342 -400 50398 800 6 la_data_out_mprj[33]
port 442 nsew signal input
rlabel metal2 s 51814 -400 51870 800 6 la_data_out_mprj[34]
port 443 nsew signal input
rlabel metal2 s 53378 -400 53434 800 6 la_data_out_mprj[35]
port 444 nsew signal input
rlabel metal2 s 54850 -400 54906 800 6 la_data_out_mprj[36]
port 445 nsew signal input
rlabel metal2 s 56414 -400 56470 800 6 la_data_out_mprj[37]
port 446 nsew signal input
rlabel metal2 s 57886 -400 57942 800 6 la_data_out_mprj[38]
port 447 nsew signal input
rlabel metal2 s 59358 -400 59414 800 6 la_data_out_mprj[39]
port 448 nsew signal input
rlabel metal2 s 5078 -400 5134 800 6 la_data_out_mprj[3]
port 449 nsew signal input
rlabel metal2 s 60922 -400 60978 800 6 la_data_out_mprj[40]
port 450 nsew signal input
rlabel metal2 s 62394 -400 62450 800 6 la_data_out_mprj[41]
port 451 nsew signal input
rlabel metal2 s 63958 -400 64014 800 6 la_data_out_mprj[42]
port 452 nsew signal input
rlabel metal2 s 65430 -400 65486 800 6 la_data_out_mprj[43]
port 453 nsew signal input
rlabel metal2 s 66902 -400 66958 800 6 la_data_out_mprj[44]
port 454 nsew signal input
rlabel metal2 s 68466 -400 68522 800 6 la_data_out_mprj[45]
port 455 nsew signal input
rlabel metal2 s 69938 -400 69994 800 6 la_data_out_mprj[46]
port 456 nsew signal input
rlabel metal2 s 71502 -400 71558 800 6 la_data_out_mprj[47]
port 457 nsew signal input
rlabel metal2 s 72974 -400 73030 800 6 la_data_out_mprj[48]
port 458 nsew signal input
rlabel metal2 s 74446 -400 74502 800 6 la_data_out_mprj[49]
port 459 nsew signal input
rlabel metal2 s 6550 -400 6606 800 6 la_data_out_mprj[4]
port 460 nsew signal input
rlabel metal2 s 76010 -400 76066 800 6 la_data_out_mprj[50]
port 461 nsew signal input
rlabel metal2 s 77482 -400 77538 800 6 la_data_out_mprj[51]
port 462 nsew signal input
rlabel metal2 s 79046 -400 79102 800 6 la_data_out_mprj[52]
port 463 nsew signal input
rlabel metal2 s 80518 -400 80574 800 6 la_data_out_mprj[53]
port 464 nsew signal input
rlabel metal2 s 81990 -400 82046 800 6 la_data_out_mprj[54]
port 465 nsew signal input
rlabel metal2 s 83554 -400 83610 800 6 la_data_out_mprj[55]
port 466 nsew signal input
rlabel metal2 s 85026 -400 85082 800 6 la_data_out_mprj[56]
port 467 nsew signal input
rlabel metal2 s 86590 -400 86646 800 6 la_data_out_mprj[57]
port 468 nsew signal input
rlabel metal2 s 88062 -400 88118 800 6 la_data_out_mprj[58]
port 469 nsew signal input
rlabel metal2 s 89534 -400 89590 800 6 la_data_out_mprj[59]
port 470 nsew signal input
rlabel metal2 s 8114 -400 8170 800 6 la_data_out_mprj[5]
port 471 nsew signal input
rlabel metal2 s 91098 -400 91154 800 6 la_data_out_mprj[60]
port 472 nsew signal input
rlabel metal2 s 92570 -400 92626 800 6 la_data_out_mprj[61]
port 473 nsew signal input
rlabel metal2 s 94134 -400 94190 800 6 la_data_out_mprj[62]
port 474 nsew signal input
rlabel metal2 s 95606 -400 95662 800 6 la_data_out_mprj[63]
port 475 nsew signal input
rlabel metal2 s 97170 -400 97226 800 6 la_data_out_mprj[64]
port 476 nsew signal input
rlabel metal2 s 98642 -400 98698 800 6 la_data_out_mprj[65]
port 477 nsew signal input
rlabel metal2 s 100114 -400 100170 800 6 la_data_out_mprj[66]
port 478 nsew signal input
rlabel metal2 s 101678 -400 101734 800 6 la_data_out_mprj[67]
port 479 nsew signal input
rlabel metal2 s 103150 -400 103206 800 6 la_data_out_mprj[68]
port 480 nsew signal input
rlabel metal2 s 104714 -400 104770 800 6 la_data_out_mprj[69]
port 481 nsew signal input
rlabel metal2 s 9586 -400 9642 800 6 la_data_out_mprj[6]
port 482 nsew signal input
rlabel metal2 s 106186 -400 106242 800 6 la_data_out_mprj[70]
port 483 nsew signal input
rlabel metal2 s 107658 -400 107714 800 6 la_data_out_mprj[71]
port 484 nsew signal input
rlabel metal2 s 109222 -400 109278 800 6 la_data_out_mprj[72]
port 485 nsew signal input
rlabel metal2 s 110694 -400 110750 800 6 la_data_out_mprj[73]
port 486 nsew signal input
rlabel metal2 s 112258 -400 112314 800 6 la_data_out_mprj[74]
port 487 nsew signal input
rlabel metal2 s 113730 -400 113786 800 6 la_data_out_mprj[75]
port 488 nsew signal input
rlabel metal2 s 115202 -400 115258 800 6 la_data_out_mprj[76]
port 489 nsew signal input
rlabel metal2 s 116766 -400 116822 800 6 la_data_out_mprj[77]
port 490 nsew signal input
rlabel metal2 s 118238 -400 118294 800 6 la_data_out_mprj[78]
port 491 nsew signal input
rlabel metal2 s 119802 -400 119858 800 6 la_data_out_mprj[79]
port 492 nsew signal input
rlabel metal2 s 11058 -400 11114 800 6 la_data_out_mprj[7]
port 493 nsew signal input
rlabel metal2 s 121274 -400 121330 800 6 la_data_out_mprj[80]
port 494 nsew signal input
rlabel metal2 s 122746 -400 122802 800 6 la_data_out_mprj[81]
port 495 nsew signal input
rlabel metal2 s 124310 -400 124366 800 6 la_data_out_mprj[82]
port 496 nsew signal input
rlabel metal2 s 125782 -400 125838 800 6 la_data_out_mprj[83]
port 497 nsew signal input
rlabel metal2 s 127346 -400 127402 800 6 la_data_out_mprj[84]
port 498 nsew signal input
rlabel metal2 s 128818 -400 128874 800 6 la_data_out_mprj[85]
port 499 nsew signal input
rlabel metal2 s 130290 -400 130346 800 6 la_data_out_mprj[86]
port 500 nsew signal input
rlabel metal2 s 131854 -400 131910 800 6 la_data_out_mprj[87]
port 501 nsew signal input
rlabel metal2 s 133326 -400 133382 800 6 la_data_out_mprj[88]
port 502 nsew signal input
rlabel metal2 s 134890 -400 134946 800 6 la_data_out_mprj[89]
port 503 nsew signal input
rlabel metal2 s 12622 -400 12678 800 6 la_data_out_mprj[8]
port 504 nsew signal input
rlabel metal2 s 136362 -400 136418 800 6 la_data_out_mprj[90]
port 505 nsew signal input
rlabel metal2 s 137834 -400 137890 800 6 la_data_out_mprj[91]
port 506 nsew signal input
rlabel metal2 s 139398 -400 139454 800 6 la_data_out_mprj[92]
port 507 nsew signal input
rlabel metal2 s 140870 -400 140926 800 6 la_data_out_mprj[93]
port 508 nsew signal input
rlabel metal2 s 142434 -400 142490 800 6 la_data_out_mprj[94]
port 509 nsew signal input
rlabel metal2 s 143906 -400 143962 800 6 la_data_out_mprj[95]
port 510 nsew signal input
rlabel metal2 s 145378 -400 145434 800 6 la_data_out_mprj[96]
port 511 nsew signal input
rlabel metal2 s 146942 -400 146998 800 6 la_data_out_mprj[97]
port 512 nsew signal input
rlabel metal2 s 148414 -400 148470 800 6 la_data_out_mprj[98]
port 513 nsew signal input
rlabel metal2 s 149978 -400 150034 800 6 la_data_out_mprj[99]
port 514 nsew signal input
rlabel metal2 s 14094 -400 14150 800 6 la_data_out_mprj[9]
port 515 nsew signal input
rlabel metal2 s 938 -400 994 800 6 la_iena_mprj[0]
port 516 nsew signal input
rlabel metal2 s 151818 -400 151874 800 6 la_iena_mprj[100]
port 517 nsew signal input
rlabel metal2 s 153382 -400 153438 800 6 la_iena_mprj[101]
port 518 nsew signal input
rlabel metal2 s 154854 -400 154910 800 6 la_iena_mprj[102]
port 519 nsew signal input
rlabel metal2 s 156326 -400 156382 800 6 la_iena_mprj[103]
port 520 nsew signal input
rlabel metal2 s 157890 -400 157946 800 6 la_iena_mprj[104]
port 521 nsew signal input
rlabel metal2 s 159362 -400 159418 800 6 la_iena_mprj[105]
port 522 nsew signal input
rlabel metal2 s 160926 -400 160982 800 6 la_iena_mprj[106]
port 523 nsew signal input
rlabel metal2 s 162398 -400 162454 800 6 la_iena_mprj[107]
port 524 nsew signal input
rlabel metal2 s 163870 -400 163926 800 6 la_iena_mprj[108]
port 525 nsew signal input
rlabel metal2 s 165434 -400 165490 800 6 la_iena_mprj[109]
port 526 nsew signal input
rlabel metal2 s 16026 -400 16082 800 6 la_iena_mprj[10]
port 527 nsew signal input
rlabel metal2 s 166906 -400 166962 800 6 la_iena_mprj[110]
port 528 nsew signal input
rlabel metal2 s 168470 -400 168526 800 6 la_iena_mprj[111]
port 529 nsew signal input
rlabel metal2 s 169942 -400 169998 800 6 la_iena_mprj[112]
port 530 nsew signal input
rlabel metal2 s 171414 -400 171470 800 6 la_iena_mprj[113]
port 531 nsew signal input
rlabel metal2 s 172978 -400 173034 800 6 la_iena_mprj[114]
port 532 nsew signal input
rlabel metal2 s 174450 -400 174506 800 6 la_iena_mprj[115]
port 533 nsew signal input
rlabel metal2 s 176014 -400 176070 800 6 la_iena_mprj[116]
port 534 nsew signal input
rlabel metal2 s 177486 -400 177542 800 6 la_iena_mprj[117]
port 535 nsew signal input
rlabel metal2 s 178958 -400 179014 800 6 la_iena_mprj[118]
port 536 nsew signal input
rlabel metal2 s 180522 -400 180578 800 6 la_iena_mprj[119]
port 537 nsew signal input
rlabel metal2 s 17498 -400 17554 800 6 la_iena_mprj[11]
port 538 nsew signal input
rlabel metal2 s 181994 -400 182050 800 6 la_iena_mprj[120]
port 539 nsew signal input
rlabel metal2 s 183558 -400 183614 800 6 la_iena_mprj[121]
port 540 nsew signal input
rlabel metal2 s 185030 -400 185086 800 6 la_iena_mprj[122]
port 541 nsew signal input
rlabel metal2 s 186502 -400 186558 800 6 la_iena_mprj[123]
port 542 nsew signal input
rlabel metal2 s 188066 -400 188122 800 6 la_iena_mprj[124]
port 543 nsew signal input
rlabel metal2 s 189538 -400 189594 800 6 la_iena_mprj[125]
port 544 nsew signal input
rlabel metal2 s 191102 -400 191158 800 6 la_iena_mprj[126]
port 545 nsew signal input
rlabel metal2 s 192574 -400 192630 800 6 la_iena_mprj[127]
port 546 nsew signal input
rlabel metal2 s 19062 -400 19118 800 6 la_iena_mprj[12]
port 547 nsew signal input
rlabel metal2 s 20534 -400 20590 800 6 la_iena_mprj[13]
port 548 nsew signal input
rlabel metal2 s 22006 -400 22062 800 6 la_iena_mprj[14]
port 549 nsew signal input
rlabel metal2 s 23570 -400 23626 800 6 la_iena_mprj[15]
port 550 nsew signal input
rlabel metal2 s 25042 -400 25098 800 6 la_iena_mprj[16]
port 551 nsew signal input
rlabel metal2 s 26606 -400 26662 800 6 la_iena_mprj[17]
port 552 nsew signal input
rlabel metal2 s 28078 -400 28134 800 6 la_iena_mprj[18]
port 553 nsew signal input
rlabel metal2 s 29550 -400 29606 800 6 la_iena_mprj[19]
port 554 nsew signal input
rlabel metal2 s 2410 -400 2466 800 6 la_iena_mprj[1]
port 555 nsew signal input
rlabel metal2 s 31114 -400 31170 800 6 la_iena_mprj[20]
port 556 nsew signal input
rlabel metal2 s 32586 -400 32642 800 6 la_iena_mprj[21]
port 557 nsew signal input
rlabel metal2 s 34150 -400 34206 800 6 la_iena_mprj[22]
port 558 nsew signal input
rlabel metal2 s 35622 -400 35678 800 6 la_iena_mprj[23]
port 559 nsew signal input
rlabel metal2 s 37094 -400 37150 800 6 la_iena_mprj[24]
port 560 nsew signal input
rlabel metal2 s 38658 -400 38714 800 6 la_iena_mprj[25]
port 561 nsew signal input
rlabel metal2 s 40130 -400 40186 800 6 la_iena_mprj[26]
port 562 nsew signal input
rlabel metal2 s 41694 -400 41750 800 6 la_iena_mprj[27]
port 563 nsew signal input
rlabel metal2 s 43166 -400 43222 800 6 la_iena_mprj[28]
port 564 nsew signal input
rlabel metal2 s 44638 -400 44694 800 6 la_iena_mprj[29]
port 565 nsew signal input
rlabel metal2 s 3974 -400 4030 800 6 la_iena_mprj[2]
port 566 nsew signal input
rlabel metal2 s 46202 -400 46258 800 6 la_iena_mprj[30]
port 567 nsew signal input
rlabel metal2 s 47674 -400 47730 800 6 la_iena_mprj[31]
port 568 nsew signal input
rlabel metal2 s 49238 -400 49294 800 6 la_iena_mprj[32]
port 569 nsew signal input
rlabel metal2 s 50710 -400 50766 800 6 la_iena_mprj[33]
port 570 nsew signal input
rlabel metal2 s 52182 -400 52238 800 6 la_iena_mprj[34]
port 571 nsew signal input
rlabel metal2 s 53746 -400 53802 800 6 la_iena_mprj[35]
port 572 nsew signal input
rlabel metal2 s 55218 -400 55274 800 6 la_iena_mprj[36]
port 573 nsew signal input
rlabel metal2 s 56782 -400 56838 800 6 la_iena_mprj[37]
port 574 nsew signal input
rlabel metal2 s 58254 -400 58310 800 6 la_iena_mprj[38]
port 575 nsew signal input
rlabel metal2 s 59726 -400 59782 800 6 la_iena_mprj[39]
port 576 nsew signal input
rlabel metal2 s 5446 -400 5502 800 6 la_iena_mprj[3]
port 577 nsew signal input
rlabel metal2 s 61290 -400 61346 800 6 la_iena_mprj[40]
port 578 nsew signal input
rlabel metal2 s 62762 -400 62818 800 6 la_iena_mprj[41]
port 579 nsew signal input
rlabel metal2 s 64326 -400 64382 800 6 la_iena_mprj[42]
port 580 nsew signal input
rlabel metal2 s 65798 -400 65854 800 6 la_iena_mprj[43]
port 581 nsew signal input
rlabel metal2 s 67362 -400 67418 800 6 la_iena_mprj[44]
port 582 nsew signal input
rlabel metal2 s 68834 -400 68890 800 6 la_iena_mprj[45]
port 583 nsew signal input
rlabel metal2 s 70306 -400 70362 800 6 la_iena_mprj[46]
port 584 nsew signal input
rlabel metal2 s 71870 -400 71926 800 6 la_iena_mprj[47]
port 585 nsew signal input
rlabel metal2 s 73342 -400 73398 800 6 la_iena_mprj[48]
port 586 nsew signal input
rlabel metal2 s 74906 -400 74962 800 6 la_iena_mprj[49]
port 587 nsew signal input
rlabel metal2 s 6918 -400 6974 800 6 la_iena_mprj[4]
port 588 nsew signal input
rlabel metal2 s 76378 -400 76434 800 6 la_iena_mprj[50]
port 589 nsew signal input
rlabel metal2 s 77850 -400 77906 800 6 la_iena_mprj[51]
port 590 nsew signal input
rlabel metal2 s 79414 -400 79470 800 6 la_iena_mprj[52]
port 591 nsew signal input
rlabel metal2 s 80886 -400 80942 800 6 la_iena_mprj[53]
port 592 nsew signal input
rlabel metal2 s 82450 -400 82506 800 6 la_iena_mprj[54]
port 593 nsew signal input
rlabel metal2 s 83922 -400 83978 800 6 la_iena_mprj[55]
port 594 nsew signal input
rlabel metal2 s 85394 -400 85450 800 6 la_iena_mprj[56]
port 595 nsew signal input
rlabel metal2 s 86958 -400 87014 800 6 la_iena_mprj[57]
port 596 nsew signal input
rlabel metal2 s 88430 -400 88486 800 6 la_iena_mprj[58]
port 597 nsew signal input
rlabel metal2 s 89994 -400 90050 800 6 la_iena_mprj[59]
port 598 nsew signal input
rlabel metal2 s 8482 -400 8538 800 6 la_iena_mprj[5]
port 599 nsew signal input
rlabel metal2 s 91466 -400 91522 800 6 la_iena_mprj[60]
port 600 nsew signal input
rlabel metal2 s 92938 -400 92994 800 6 la_iena_mprj[61]
port 601 nsew signal input
rlabel metal2 s 94502 -400 94558 800 6 la_iena_mprj[62]
port 602 nsew signal input
rlabel metal2 s 95974 -400 96030 800 6 la_iena_mprj[63]
port 603 nsew signal input
rlabel metal2 s 97538 -400 97594 800 6 la_iena_mprj[64]
port 604 nsew signal input
rlabel metal2 s 99010 -400 99066 800 6 la_iena_mprj[65]
port 605 nsew signal input
rlabel metal2 s 100482 -400 100538 800 6 la_iena_mprj[66]
port 606 nsew signal input
rlabel metal2 s 102046 -400 102102 800 6 la_iena_mprj[67]
port 607 nsew signal input
rlabel metal2 s 103518 -400 103574 800 6 la_iena_mprj[68]
port 608 nsew signal input
rlabel metal2 s 105082 -400 105138 800 6 la_iena_mprj[69]
port 609 nsew signal input
rlabel metal2 s 9954 -400 10010 800 6 la_iena_mprj[6]
port 610 nsew signal input
rlabel metal2 s 106554 -400 106610 800 6 la_iena_mprj[70]
port 611 nsew signal input
rlabel metal2 s 108026 -400 108082 800 6 la_iena_mprj[71]
port 612 nsew signal input
rlabel metal2 s 109590 -400 109646 800 6 la_iena_mprj[72]
port 613 nsew signal input
rlabel metal2 s 111062 -400 111118 800 6 la_iena_mprj[73]
port 614 nsew signal input
rlabel metal2 s 112626 -400 112682 800 6 la_iena_mprj[74]
port 615 nsew signal input
rlabel metal2 s 114098 -400 114154 800 6 la_iena_mprj[75]
port 616 nsew signal input
rlabel metal2 s 115570 -400 115626 800 6 la_iena_mprj[76]
port 617 nsew signal input
rlabel metal2 s 117134 -400 117190 800 6 la_iena_mprj[77]
port 618 nsew signal input
rlabel metal2 s 118606 -400 118662 800 6 la_iena_mprj[78]
port 619 nsew signal input
rlabel metal2 s 120170 -400 120226 800 6 la_iena_mprj[79]
port 620 nsew signal input
rlabel metal2 s 11518 -400 11574 800 6 la_iena_mprj[7]
port 621 nsew signal input
rlabel metal2 s 121642 -400 121698 800 6 la_iena_mprj[80]
port 622 nsew signal input
rlabel metal2 s 123114 -400 123170 800 6 la_iena_mprj[81]
port 623 nsew signal input
rlabel metal2 s 124678 -400 124734 800 6 la_iena_mprj[82]
port 624 nsew signal input
rlabel metal2 s 126150 -400 126206 800 6 la_iena_mprj[83]
port 625 nsew signal input
rlabel metal2 s 127714 -400 127770 800 6 la_iena_mprj[84]
port 626 nsew signal input
rlabel metal2 s 129186 -400 129242 800 6 la_iena_mprj[85]
port 627 nsew signal input
rlabel metal2 s 130750 -400 130806 800 6 la_iena_mprj[86]
port 628 nsew signal input
rlabel metal2 s 132222 -400 132278 800 6 la_iena_mprj[87]
port 629 nsew signal input
rlabel metal2 s 133694 -400 133750 800 6 la_iena_mprj[88]
port 630 nsew signal input
rlabel metal2 s 135258 -400 135314 800 6 la_iena_mprj[89]
port 631 nsew signal input
rlabel metal2 s 12990 -400 13046 800 6 la_iena_mprj[8]
port 632 nsew signal input
rlabel metal2 s 136730 -400 136786 800 6 la_iena_mprj[90]
port 633 nsew signal input
rlabel metal2 s 138294 -400 138350 800 6 la_iena_mprj[91]
port 634 nsew signal input
rlabel metal2 s 139766 -400 139822 800 6 la_iena_mprj[92]
port 635 nsew signal input
rlabel metal2 s 141238 -400 141294 800 6 la_iena_mprj[93]
port 636 nsew signal input
rlabel metal2 s 142802 -400 142858 800 6 la_iena_mprj[94]
port 637 nsew signal input
rlabel metal2 s 144274 -400 144330 800 6 la_iena_mprj[95]
port 638 nsew signal input
rlabel metal2 s 145838 -400 145894 800 6 la_iena_mprj[96]
port 639 nsew signal input
rlabel metal2 s 147310 -400 147366 800 6 la_iena_mprj[97]
port 640 nsew signal input
rlabel metal2 s 148782 -400 148838 800 6 la_iena_mprj[98]
port 641 nsew signal input
rlabel metal2 s 150346 -400 150402 800 6 la_iena_mprj[99]
port 642 nsew signal input
rlabel metal2 s 14462 -400 14518 800 6 la_iena_mprj[9]
port 643 nsew signal input
rlabel metal2 s 35898 22600 35954 23800 6 la_oenb_core[0]
port 644 nsew signal output
rlabel metal2 s 179050 22600 179106 23800 6 la_oenb_core[100]
port 645 nsew signal output
rlabel metal2 s 180522 22600 180578 23800 6 la_oenb_core[101]
port 646 nsew signal output
rlabel metal2 s 181994 22600 182050 23800 6 la_oenb_core[102]
port 647 nsew signal output
rlabel metal2 s 183374 22600 183430 23800 6 la_oenb_core[103]
port 648 nsew signal output
rlabel metal2 s 184846 22600 184902 23800 6 la_oenb_core[104]
port 649 nsew signal output
rlabel metal2 s 186226 22600 186282 23800 6 la_oenb_core[105]
port 650 nsew signal output
rlabel metal2 s 187698 22600 187754 23800 6 la_oenb_core[106]
port 651 nsew signal output
rlabel metal2 s 189078 22600 189134 23800 6 la_oenb_core[107]
port 652 nsew signal output
rlabel metal2 s 190550 22600 190606 23800 6 la_oenb_core[108]
port 653 nsew signal output
rlabel metal2 s 191930 22600 191986 23800 6 la_oenb_core[109]
port 654 nsew signal output
rlabel metal2 s 50250 22600 50306 23800 6 la_oenb_core[10]
port 655 nsew signal output
rlabel metal2 s 193402 22600 193458 23800 6 la_oenb_core[110]
port 656 nsew signal output
rlabel metal2 s 194874 22600 194930 23800 6 la_oenb_core[111]
port 657 nsew signal output
rlabel metal2 s 196254 22600 196310 23800 6 la_oenb_core[112]
port 658 nsew signal output
rlabel metal2 s 197726 22600 197782 23800 6 la_oenb_core[113]
port 659 nsew signal output
rlabel metal2 s 199106 22600 199162 23800 6 la_oenb_core[114]
port 660 nsew signal output
rlabel metal2 s 200578 22600 200634 23800 6 la_oenb_core[115]
port 661 nsew signal output
rlabel metal2 s 201958 22600 202014 23800 6 la_oenb_core[116]
port 662 nsew signal output
rlabel metal2 s 203430 22600 203486 23800 6 la_oenb_core[117]
port 663 nsew signal output
rlabel metal2 s 204902 22600 204958 23800 6 la_oenb_core[118]
port 664 nsew signal output
rlabel metal2 s 206282 22600 206338 23800 6 la_oenb_core[119]
port 665 nsew signal output
rlabel metal2 s 51722 22600 51778 23800 6 la_oenb_core[11]
port 666 nsew signal output
rlabel metal2 s 207754 22600 207810 23800 6 la_oenb_core[120]
port 667 nsew signal output
rlabel metal2 s 209134 22600 209190 23800 6 la_oenb_core[121]
port 668 nsew signal output
rlabel metal2 s 210606 22600 210662 23800 6 la_oenb_core[122]
port 669 nsew signal output
rlabel metal2 s 211986 22600 212042 23800 6 la_oenb_core[123]
port 670 nsew signal output
rlabel metal2 s 213458 22600 213514 23800 6 la_oenb_core[124]
port 671 nsew signal output
rlabel metal2 s 214838 22600 214894 23800 6 la_oenb_core[125]
port 672 nsew signal output
rlabel metal2 s 216310 22600 216366 23800 6 la_oenb_core[126]
port 673 nsew signal output
rlabel metal2 s 217782 22600 217838 23800 6 la_oenb_core[127]
port 674 nsew signal output
rlabel metal2 s 53102 22600 53158 23800 6 la_oenb_core[12]
port 675 nsew signal output
rlabel metal2 s 54574 22600 54630 23800 6 la_oenb_core[13]
port 676 nsew signal output
rlabel metal2 s 55954 22600 56010 23800 6 la_oenb_core[14]
port 677 nsew signal output
rlabel metal2 s 57426 22600 57482 23800 6 la_oenb_core[15]
port 678 nsew signal output
rlabel metal2 s 58806 22600 58862 23800 6 la_oenb_core[16]
port 679 nsew signal output
rlabel metal2 s 60278 22600 60334 23800 6 la_oenb_core[17]
port 680 nsew signal output
rlabel metal2 s 61750 22600 61806 23800 6 la_oenb_core[18]
port 681 nsew signal output
rlabel metal2 s 63130 22600 63186 23800 6 la_oenb_core[19]
port 682 nsew signal output
rlabel metal2 s 37370 22600 37426 23800 6 la_oenb_core[1]
port 683 nsew signal output
rlabel metal2 s 64602 22600 64658 23800 6 la_oenb_core[20]
port 684 nsew signal output
rlabel metal2 s 65982 22600 66038 23800 6 la_oenb_core[21]
port 685 nsew signal output
rlabel metal2 s 67454 22600 67510 23800 6 la_oenb_core[22]
port 686 nsew signal output
rlabel metal2 s 68834 22600 68890 23800 6 la_oenb_core[23]
port 687 nsew signal output
rlabel metal2 s 70306 22600 70362 23800 6 la_oenb_core[24]
port 688 nsew signal output
rlabel metal2 s 71686 22600 71742 23800 6 la_oenb_core[25]
port 689 nsew signal output
rlabel metal2 s 73158 22600 73214 23800 6 la_oenb_core[26]
port 690 nsew signal output
rlabel metal2 s 74630 22600 74686 23800 6 la_oenb_core[27]
port 691 nsew signal output
rlabel metal2 s 76010 22600 76066 23800 6 la_oenb_core[28]
port 692 nsew signal output
rlabel metal2 s 77482 22600 77538 23800 6 la_oenb_core[29]
port 693 nsew signal output
rlabel metal2 s 38842 22600 38898 23800 6 la_oenb_core[2]
port 694 nsew signal output
rlabel metal2 s 78862 22600 78918 23800 6 la_oenb_core[30]
port 695 nsew signal output
rlabel metal2 s 80334 22600 80390 23800 6 la_oenb_core[31]
port 696 nsew signal output
rlabel metal2 s 81714 22600 81770 23800 6 la_oenb_core[32]
port 697 nsew signal output
rlabel metal2 s 83186 22600 83242 23800 6 la_oenb_core[33]
port 698 nsew signal output
rlabel metal2 s 84658 22600 84714 23800 6 la_oenb_core[34]
port 699 nsew signal output
rlabel metal2 s 86038 22600 86094 23800 6 la_oenb_core[35]
port 700 nsew signal output
rlabel metal2 s 87510 22600 87566 23800 6 la_oenb_core[36]
port 701 nsew signal output
rlabel metal2 s 88890 22600 88946 23800 6 la_oenb_core[37]
port 702 nsew signal output
rlabel metal2 s 90362 22600 90418 23800 6 la_oenb_core[38]
port 703 nsew signal output
rlabel metal2 s 91742 22600 91798 23800 6 la_oenb_core[39]
port 704 nsew signal output
rlabel metal2 s 40222 22600 40278 23800 6 la_oenb_core[3]
port 705 nsew signal output
rlabel metal2 s 93214 22600 93270 23800 6 la_oenb_core[40]
port 706 nsew signal output
rlabel metal2 s 94594 22600 94650 23800 6 la_oenb_core[41]
port 707 nsew signal output
rlabel metal2 s 96066 22600 96122 23800 6 la_oenb_core[42]
port 708 nsew signal output
rlabel metal2 s 97538 22600 97594 23800 6 la_oenb_core[43]
port 709 nsew signal output
rlabel metal2 s 98918 22600 98974 23800 6 la_oenb_core[44]
port 710 nsew signal output
rlabel metal2 s 100390 22600 100446 23800 6 la_oenb_core[45]
port 711 nsew signal output
rlabel metal2 s 101770 22600 101826 23800 6 la_oenb_core[46]
port 712 nsew signal output
rlabel metal2 s 103242 22600 103298 23800 6 la_oenb_core[47]
port 713 nsew signal output
rlabel metal2 s 104622 22600 104678 23800 6 la_oenb_core[48]
port 714 nsew signal output
rlabel metal2 s 106094 22600 106150 23800 6 la_oenb_core[49]
port 715 nsew signal output
rlabel metal2 s 41694 22600 41750 23800 6 la_oenb_core[4]
port 716 nsew signal output
rlabel metal2 s 107474 22600 107530 23800 6 la_oenb_core[50]
port 717 nsew signal output
rlabel metal2 s 108946 22600 109002 23800 6 la_oenb_core[51]
port 718 nsew signal output
rlabel metal2 s 110418 22600 110474 23800 6 la_oenb_core[52]
port 719 nsew signal output
rlabel metal2 s 111798 22600 111854 23800 6 la_oenb_core[53]
port 720 nsew signal output
rlabel metal2 s 113270 22600 113326 23800 6 la_oenb_core[54]
port 721 nsew signal output
rlabel metal2 s 114650 22600 114706 23800 6 la_oenb_core[55]
port 722 nsew signal output
rlabel metal2 s 116122 22600 116178 23800 6 la_oenb_core[56]
port 723 nsew signal output
rlabel metal2 s 117502 22600 117558 23800 6 la_oenb_core[57]
port 724 nsew signal output
rlabel metal2 s 118974 22600 119030 23800 6 la_oenb_core[58]
port 725 nsew signal output
rlabel metal2 s 120446 22600 120502 23800 6 la_oenb_core[59]
port 726 nsew signal output
rlabel metal2 s 43074 22600 43130 23800 6 la_oenb_core[5]
port 727 nsew signal output
rlabel metal2 s 121826 22600 121882 23800 6 la_oenb_core[60]
port 728 nsew signal output
rlabel metal2 s 123298 22600 123354 23800 6 la_oenb_core[61]
port 729 nsew signal output
rlabel metal2 s 124678 22600 124734 23800 6 la_oenb_core[62]
port 730 nsew signal output
rlabel metal2 s 126150 22600 126206 23800 6 la_oenb_core[63]
port 731 nsew signal output
rlabel metal2 s 127530 22600 127586 23800 6 la_oenb_core[64]
port 732 nsew signal output
rlabel metal2 s 129002 22600 129058 23800 6 la_oenb_core[65]
port 733 nsew signal output
rlabel metal2 s 130382 22600 130438 23800 6 la_oenb_core[66]
port 734 nsew signal output
rlabel metal2 s 131854 22600 131910 23800 6 la_oenb_core[67]
port 735 nsew signal output
rlabel metal2 s 133326 22600 133382 23800 6 la_oenb_core[68]
port 736 nsew signal output
rlabel metal2 s 134706 22600 134762 23800 6 la_oenb_core[69]
port 737 nsew signal output
rlabel metal2 s 44546 22600 44602 23800 6 la_oenb_core[6]
port 738 nsew signal output
rlabel metal2 s 136178 22600 136234 23800 6 la_oenb_core[70]
port 739 nsew signal output
rlabel metal2 s 137558 22600 137614 23800 6 la_oenb_core[71]
port 740 nsew signal output
rlabel metal2 s 139030 22600 139086 23800 6 la_oenb_core[72]
port 741 nsew signal output
rlabel metal2 s 140410 22600 140466 23800 6 la_oenb_core[73]
port 742 nsew signal output
rlabel metal2 s 141882 22600 141938 23800 6 la_oenb_core[74]
port 743 nsew signal output
rlabel metal2 s 143262 22600 143318 23800 6 la_oenb_core[75]
port 744 nsew signal output
rlabel metal2 s 144734 22600 144790 23800 6 la_oenb_core[76]
port 745 nsew signal output
rlabel metal2 s 146206 22600 146262 23800 6 la_oenb_core[77]
port 746 nsew signal output
rlabel metal2 s 147586 22600 147642 23800 6 la_oenb_core[78]
port 747 nsew signal output
rlabel metal2 s 149058 22600 149114 23800 6 la_oenb_core[79]
port 748 nsew signal output
rlabel metal2 s 45926 22600 45982 23800 6 la_oenb_core[7]
port 749 nsew signal output
rlabel metal2 s 150438 22600 150494 23800 6 la_oenb_core[80]
port 750 nsew signal output
rlabel metal2 s 151910 22600 151966 23800 6 la_oenb_core[81]
port 751 nsew signal output
rlabel metal2 s 153290 22600 153346 23800 6 la_oenb_core[82]
port 752 nsew signal output
rlabel metal2 s 154762 22600 154818 23800 6 la_oenb_core[83]
port 753 nsew signal output
rlabel metal2 s 156234 22600 156290 23800 6 la_oenb_core[84]
port 754 nsew signal output
rlabel metal2 s 157614 22600 157670 23800 6 la_oenb_core[85]
port 755 nsew signal output
rlabel metal2 s 159086 22600 159142 23800 6 la_oenb_core[86]
port 756 nsew signal output
rlabel metal2 s 160466 22600 160522 23800 6 la_oenb_core[87]
port 757 nsew signal output
rlabel metal2 s 161938 22600 161994 23800 6 la_oenb_core[88]
port 758 nsew signal output
rlabel metal2 s 163318 22600 163374 23800 6 la_oenb_core[89]
port 759 nsew signal output
rlabel metal2 s 47398 22600 47454 23800 6 la_oenb_core[8]
port 760 nsew signal output
rlabel metal2 s 164790 22600 164846 23800 6 la_oenb_core[90]
port 761 nsew signal output
rlabel metal2 s 166170 22600 166226 23800 6 la_oenb_core[91]
port 762 nsew signal output
rlabel metal2 s 167642 22600 167698 23800 6 la_oenb_core[92]
port 763 nsew signal output
rlabel metal2 s 169114 22600 169170 23800 6 la_oenb_core[93]
port 764 nsew signal output
rlabel metal2 s 170494 22600 170550 23800 6 la_oenb_core[94]
port 765 nsew signal output
rlabel metal2 s 171966 22600 172022 23800 6 la_oenb_core[95]
port 766 nsew signal output
rlabel metal2 s 173346 22600 173402 23800 6 la_oenb_core[96]
port 767 nsew signal output
rlabel metal2 s 174818 22600 174874 23800 6 la_oenb_core[97]
port 768 nsew signal output
rlabel metal2 s 176198 22600 176254 23800 6 la_oenb_core[98]
port 769 nsew signal output
rlabel metal2 s 177670 22600 177726 23800 6 la_oenb_core[99]
port 770 nsew signal output
rlabel metal2 s 48870 22600 48926 23800 6 la_oenb_core[9]
port 771 nsew signal output
rlabel metal2 s 1306 -400 1362 800 6 la_oenb_mprj[0]
port 772 nsew signal input
rlabel metal2 s 152186 -400 152242 800 6 la_oenb_mprj[100]
port 773 nsew signal input
rlabel metal2 s 153750 -400 153806 800 6 la_oenb_mprj[101]
port 774 nsew signal input
rlabel metal2 s 155222 -400 155278 800 6 la_oenb_mprj[102]
port 775 nsew signal input
rlabel metal2 s 156694 -400 156750 800 6 la_oenb_mprj[103]
port 776 nsew signal input
rlabel metal2 s 158258 -400 158314 800 6 la_oenb_mprj[104]
port 777 nsew signal input
rlabel metal2 s 159730 -400 159786 800 6 la_oenb_mprj[105]
port 778 nsew signal input
rlabel metal2 s 161294 -400 161350 800 6 la_oenb_mprj[106]
port 779 nsew signal input
rlabel metal2 s 162766 -400 162822 800 6 la_oenb_mprj[107]
port 780 nsew signal input
rlabel metal2 s 164330 -400 164386 800 6 la_oenb_mprj[108]
port 781 nsew signal input
rlabel metal2 s 165802 -400 165858 800 6 la_oenb_mprj[109]
port 782 nsew signal input
rlabel metal2 s 16394 -400 16450 800 6 la_oenb_mprj[10]
port 783 nsew signal input
rlabel metal2 s 167274 -400 167330 800 6 la_oenb_mprj[110]
port 784 nsew signal input
rlabel metal2 s 168838 -400 168894 800 6 la_oenb_mprj[111]
port 785 nsew signal input
rlabel metal2 s 170310 -400 170366 800 6 la_oenb_mprj[112]
port 786 nsew signal input
rlabel metal2 s 171874 -400 171930 800 6 la_oenb_mprj[113]
port 787 nsew signal input
rlabel metal2 s 173346 -400 173402 800 6 la_oenb_mprj[114]
port 788 nsew signal input
rlabel metal2 s 174818 -400 174874 800 6 la_oenb_mprj[115]
port 789 nsew signal input
rlabel metal2 s 176382 -400 176438 800 6 la_oenb_mprj[116]
port 790 nsew signal input
rlabel metal2 s 177854 -400 177910 800 6 la_oenb_mprj[117]
port 791 nsew signal input
rlabel metal2 s 179418 -400 179474 800 6 la_oenb_mprj[118]
port 792 nsew signal input
rlabel metal2 s 180890 -400 180946 800 6 la_oenb_mprj[119]
port 793 nsew signal input
rlabel metal2 s 17866 -400 17922 800 6 la_oenb_mprj[11]
port 794 nsew signal input
rlabel metal2 s 182362 -400 182418 800 6 la_oenb_mprj[120]
port 795 nsew signal input
rlabel metal2 s 183926 -400 183982 800 6 la_oenb_mprj[121]
port 796 nsew signal input
rlabel metal2 s 185398 -400 185454 800 6 la_oenb_mprj[122]
port 797 nsew signal input
rlabel metal2 s 186962 -400 187018 800 6 la_oenb_mprj[123]
port 798 nsew signal input
rlabel metal2 s 188434 -400 188490 800 6 la_oenb_mprj[124]
port 799 nsew signal input
rlabel metal2 s 189906 -400 189962 800 6 la_oenb_mprj[125]
port 800 nsew signal input
rlabel metal2 s 191470 -400 191526 800 6 la_oenb_mprj[126]
port 801 nsew signal input
rlabel metal2 s 192942 -400 192998 800 6 la_oenb_mprj[127]
port 802 nsew signal input
rlabel metal2 s 19430 -400 19486 800 6 la_oenb_mprj[12]
port 803 nsew signal input
rlabel metal2 s 20902 -400 20958 800 6 la_oenb_mprj[13]
port 804 nsew signal input
rlabel metal2 s 22374 -400 22430 800 6 la_oenb_mprj[14]
port 805 nsew signal input
rlabel metal2 s 23938 -400 23994 800 6 la_oenb_mprj[15]
port 806 nsew signal input
rlabel metal2 s 25410 -400 25466 800 6 la_oenb_mprj[16]
port 807 nsew signal input
rlabel metal2 s 26974 -400 27030 800 6 la_oenb_mprj[17]
port 808 nsew signal input
rlabel metal2 s 28446 -400 28502 800 6 la_oenb_mprj[18]
port 809 nsew signal input
rlabel metal2 s 29918 -400 29974 800 6 la_oenb_mprj[19]
port 810 nsew signal input
rlabel metal2 s 2778 -400 2834 800 6 la_oenb_mprj[1]
port 811 nsew signal input
rlabel metal2 s 31482 -400 31538 800 6 la_oenb_mprj[20]
port 812 nsew signal input
rlabel metal2 s 32954 -400 33010 800 6 la_oenb_mprj[21]
port 813 nsew signal input
rlabel metal2 s 34518 -400 34574 800 6 la_oenb_mprj[22]
port 814 nsew signal input
rlabel metal2 s 35990 -400 36046 800 6 la_oenb_mprj[23]
port 815 nsew signal input
rlabel metal2 s 37554 -400 37610 800 6 la_oenb_mprj[24]
port 816 nsew signal input
rlabel metal2 s 39026 -400 39082 800 6 la_oenb_mprj[25]
port 817 nsew signal input
rlabel metal2 s 40498 -400 40554 800 6 la_oenb_mprj[26]
port 818 nsew signal input
rlabel metal2 s 42062 -400 42118 800 6 la_oenb_mprj[27]
port 819 nsew signal input
rlabel metal2 s 43534 -400 43590 800 6 la_oenb_mprj[28]
port 820 nsew signal input
rlabel metal2 s 45098 -400 45154 800 6 la_oenb_mprj[29]
port 821 nsew signal input
rlabel metal2 s 4342 -400 4398 800 6 la_oenb_mprj[2]
port 822 nsew signal input
rlabel metal2 s 46570 -400 46626 800 6 la_oenb_mprj[30]
port 823 nsew signal input
rlabel metal2 s 48042 -400 48098 800 6 la_oenb_mprj[31]
port 824 nsew signal input
rlabel metal2 s 49606 -400 49662 800 6 la_oenb_mprj[32]
port 825 nsew signal input
rlabel metal2 s 51078 -400 51134 800 6 la_oenb_mprj[33]
port 826 nsew signal input
rlabel metal2 s 52642 -400 52698 800 6 la_oenb_mprj[34]
port 827 nsew signal input
rlabel metal2 s 54114 -400 54170 800 6 la_oenb_mprj[35]
port 828 nsew signal input
rlabel metal2 s 55586 -400 55642 800 6 la_oenb_mprj[36]
port 829 nsew signal input
rlabel metal2 s 57150 -400 57206 800 6 la_oenb_mprj[37]
port 830 nsew signal input
rlabel metal2 s 58622 -400 58678 800 6 la_oenb_mprj[38]
port 831 nsew signal input
rlabel metal2 s 60186 -400 60242 800 6 la_oenb_mprj[39]
port 832 nsew signal input
rlabel metal2 s 5814 -400 5870 800 6 la_oenb_mprj[3]
port 833 nsew signal input
rlabel metal2 s 61658 -400 61714 800 6 la_oenb_mprj[40]
port 834 nsew signal input
rlabel metal2 s 63130 -400 63186 800 6 la_oenb_mprj[41]
port 835 nsew signal input
rlabel metal2 s 64694 -400 64750 800 6 la_oenb_mprj[42]
port 836 nsew signal input
rlabel metal2 s 66166 -400 66222 800 6 la_oenb_mprj[43]
port 837 nsew signal input
rlabel metal2 s 67730 -400 67786 800 6 la_oenb_mprj[44]
port 838 nsew signal input
rlabel metal2 s 69202 -400 69258 800 6 la_oenb_mprj[45]
port 839 nsew signal input
rlabel metal2 s 70674 -400 70730 800 6 la_oenb_mprj[46]
port 840 nsew signal input
rlabel metal2 s 72238 -400 72294 800 6 la_oenb_mprj[47]
port 841 nsew signal input
rlabel metal2 s 73710 -400 73766 800 6 la_oenb_mprj[48]
port 842 nsew signal input
rlabel metal2 s 75274 -400 75330 800 6 la_oenb_mprj[49]
port 843 nsew signal input
rlabel metal2 s 7286 -400 7342 800 6 la_oenb_mprj[4]
port 844 nsew signal input
rlabel metal2 s 76746 -400 76802 800 6 la_oenb_mprj[50]
port 845 nsew signal input
rlabel metal2 s 78218 -400 78274 800 6 la_oenb_mprj[51]
port 846 nsew signal input
rlabel metal2 s 79782 -400 79838 800 6 la_oenb_mprj[52]
port 847 nsew signal input
rlabel metal2 s 81254 -400 81310 800 6 la_oenb_mprj[53]
port 848 nsew signal input
rlabel metal2 s 82818 -400 82874 800 6 la_oenb_mprj[54]
port 849 nsew signal input
rlabel metal2 s 84290 -400 84346 800 6 la_oenb_mprj[55]
port 850 nsew signal input
rlabel metal2 s 85762 -400 85818 800 6 la_oenb_mprj[56]
port 851 nsew signal input
rlabel metal2 s 87326 -400 87382 800 6 la_oenb_mprj[57]
port 852 nsew signal input
rlabel metal2 s 88798 -400 88854 800 6 la_oenb_mprj[58]
port 853 nsew signal input
rlabel metal2 s 90362 -400 90418 800 6 la_oenb_mprj[59]
port 854 nsew signal input
rlabel metal2 s 8850 -400 8906 800 6 la_oenb_mprj[5]
port 855 nsew signal input
rlabel metal2 s 91834 -400 91890 800 6 la_oenb_mprj[60]
port 856 nsew signal input
rlabel metal2 s 93306 -400 93362 800 6 la_oenb_mprj[61]
port 857 nsew signal input
rlabel metal2 s 94870 -400 94926 800 6 la_oenb_mprj[62]
port 858 nsew signal input
rlabel metal2 s 96342 -400 96398 800 6 la_oenb_mprj[63]
port 859 nsew signal input
rlabel metal2 s 97906 -400 97962 800 6 la_oenb_mprj[64]
port 860 nsew signal input
rlabel metal2 s 99378 -400 99434 800 6 la_oenb_mprj[65]
port 861 nsew signal input
rlabel metal2 s 100942 -400 100998 800 6 la_oenb_mprj[66]
port 862 nsew signal input
rlabel metal2 s 102414 -400 102470 800 6 la_oenb_mprj[67]
port 863 nsew signal input
rlabel metal2 s 103886 -400 103942 800 6 la_oenb_mprj[68]
port 864 nsew signal input
rlabel metal2 s 105450 -400 105506 800 6 la_oenb_mprj[69]
port 865 nsew signal input
rlabel metal2 s 10322 -400 10378 800 6 la_oenb_mprj[6]
port 866 nsew signal input
rlabel metal2 s 106922 -400 106978 800 6 la_oenb_mprj[70]
port 867 nsew signal input
rlabel metal2 s 108486 -400 108542 800 6 la_oenb_mprj[71]
port 868 nsew signal input
rlabel metal2 s 109958 -400 110014 800 6 la_oenb_mprj[72]
port 869 nsew signal input
rlabel metal2 s 111430 -400 111486 800 6 la_oenb_mprj[73]
port 870 nsew signal input
rlabel metal2 s 112994 -400 113050 800 6 la_oenb_mprj[74]
port 871 nsew signal input
rlabel metal2 s 114466 -400 114522 800 6 la_oenb_mprj[75]
port 872 nsew signal input
rlabel metal2 s 116030 -400 116086 800 6 la_oenb_mprj[76]
port 873 nsew signal input
rlabel metal2 s 117502 -400 117558 800 6 la_oenb_mprj[77]
port 874 nsew signal input
rlabel metal2 s 118974 -400 119030 800 6 la_oenb_mprj[78]
port 875 nsew signal input
rlabel metal2 s 120538 -400 120594 800 6 la_oenb_mprj[79]
port 876 nsew signal input
rlabel metal2 s 11886 -400 11942 800 6 la_oenb_mprj[7]
port 877 nsew signal input
rlabel metal2 s 122010 -400 122066 800 6 la_oenb_mprj[80]
port 878 nsew signal input
rlabel metal2 s 123574 -400 123630 800 6 la_oenb_mprj[81]
port 879 nsew signal input
rlabel metal2 s 125046 -400 125102 800 6 la_oenb_mprj[82]
port 880 nsew signal input
rlabel metal2 s 126518 -400 126574 800 6 la_oenb_mprj[83]
port 881 nsew signal input
rlabel metal2 s 128082 -400 128138 800 6 la_oenb_mprj[84]
port 882 nsew signal input
rlabel metal2 s 129554 -400 129610 800 6 la_oenb_mprj[85]
port 883 nsew signal input
rlabel metal2 s 131118 -400 131174 800 6 la_oenb_mprj[86]
port 884 nsew signal input
rlabel metal2 s 132590 -400 132646 800 6 la_oenb_mprj[87]
port 885 nsew signal input
rlabel metal2 s 134062 -400 134118 800 6 la_oenb_mprj[88]
port 886 nsew signal input
rlabel metal2 s 135626 -400 135682 800 6 la_oenb_mprj[89]
port 887 nsew signal input
rlabel metal2 s 13358 -400 13414 800 6 la_oenb_mprj[8]
port 888 nsew signal input
rlabel metal2 s 137098 -400 137154 800 6 la_oenb_mprj[90]
port 889 nsew signal input
rlabel metal2 s 138662 -400 138718 800 6 la_oenb_mprj[91]
port 890 nsew signal input
rlabel metal2 s 140134 -400 140190 800 6 la_oenb_mprj[92]
port 891 nsew signal input
rlabel metal2 s 141606 -400 141662 800 6 la_oenb_mprj[93]
port 892 nsew signal input
rlabel metal2 s 143170 -400 143226 800 6 la_oenb_mprj[94]
port 893 nsew signal input
rlabel metal2 s 144642 -400 144698 800 6 la_oenb_mprj[95]
port 894 nsew signal input
rlabel metal2 s 146206 -400 146262 800 6 la_oenb_mprj[96]
port 895 nsew signal input
rlabel metal2 s 147678 -400 147734 800 6 la_oenb_mprj[97]
port 896 nsew signal input
rlabel metal2 s 149150 -400 149206 800 6 la_oenb_mprj[98]
port 897 nsew signal input
rlabel metal2 s 150714 -400 150770 800 6 la_oenb_mprj[99]
port 898 nsew signal input
rlabel metal2 s 14830 -400 14886 800 6 la_oenb_mprj[9]
port 899 nsew signal input
rlabel metal2 s 194506 -400 194562 800 6 mprj_adr_o_core[0]
port 900 nsew signal input
rlabel metal2 s 203522 -400 203578 800 6 mprj_adr_o_core[10]
port 901 nsew signal input
rlabel metal2 s 204258 -400 204314 800 6 mprj_adr_o_core[11]
port 902 nsew signal input
rlabel metal2 s 204994 -400 205050 800 6 mprj_adr_o_core[12]
port 903 nsew signal input
rlabel metal2 s 205822 -400 205878 800 6 mprj_adr_o_core[13]
port 904 nsew signal input
rlabel metal2 s 206558 -400 206614 800 6 mprj_adr_o_core[14]
port 905 nsew signal input
rlabel metal2 s 207294 -400 207350 800 6 mprj_adr_o_core[15]
port 906 nsew signal input
rlabel metal2 s 208030 -400 208086 800 6 mprj_adr_o_core[16]
port 907 nsew signal input
rlabel metal2 s 208766 -400 208822 800 6 mprj_adr_o_core[17]
port 908 nsew signal input
rlabel metal2 s 209594 -400 209650 800 6 mprj_adr_o_core[18]
port 909 nsew signal input
rlabel metal2 s 210330 -400 210386 800 6 mprj_adr_o_core[19]
port 910 nsew signal input
rlabel metal2 s 195610 -400 195666 800 6 mprj_adr_o_core[1]
port 911 nsew signal input
rlabel metal2 s 211066 -400 211122 800 6 mprj_adr_o_core[20]
port 912 nsew signal input
rlabel metal2 s 211802 -400 211858 800 6 mprj_adr_o_core[21]
port 913 nsew signal input
rlabel metal2 s 212538 -400 212594 800 6 mprj_adr_o_core[22]
port 914 nsew signal input
rlabel metal2 s 213366 -400 213422 800 6 mprj_adr_o_core[23]
port 915 nsew signal input
rlabel metal2 s 214102 -400 214158 800 6 mprj_adr_o_core[24]
port 916 nsew signal input
rlabel metal2 s 214838 -400 214894 800 6 mprj_adr_o_core[25]
port 917 nsew signal input
rlabel metal2 s 215574 -400 215630 800 6 mprj_adr_o_core[26]
port 918 nsew signal input
rlabel metal2 s 216310 -400 216366 800 6 mprj_adr_o_core[27]
port 919 nsew signal input
rlabel metal2 s 217138 -400 217194 800 6 mprj_adr_o_core[28]
port 920 nsew signal input
rlabel metal2 s 217874 -400 217930 800 6 mprj_adr_o_core[29]
port 921 nsew signal input
rlabel metal2 s 196714 -400 196770 800 6 mprj_adr_o_core[2]
port 922 nsew signal input
rlabel metal2 s 218610 -400 218666 800 6 mprj_adr_o_core[30]
port 923 nsew signal input
rlabel metal2 s 219346 -400 219402 800 6 mprj_adr_o_core[31]
port 924 nsew signal input
rlabel metal2 s 197910 -400 197966 800 6 mprj_adr_o_core[3]
port 925 nsew signal input
rlabel metal2 s 199014 -400 199070 800 6 mprj_adr_o_core[4]
port 926 nsew signal input
rlabel metal2 s 199750 -400 199806 800 6 mprj_adr_o_core[5]
port 927 nsew signal input
rlabel metal2 s 200486 -400 200542 800 6 mprj_adr_o_core[6]
port 928 nsew signal input
rlabel metal2 s 201222 -400 201278 800 6 mprj_adr_o_core[7]
port 929 nsew signal input
rlabel metal2 s 202050 -400 202106 800 6 mprj_adr_o_core[8]
port 930 nsew signal input
rlabel metal2 s 202786 -400 202842 800 6 mprj_adr_o_core[9]
port 931 nsew signal input
rlabel metal2 s 2502 22600 2558 23800 6 mprj_adr_o_user[0]
port 932 nsew signal output
rlabel metal2 s 14002 22600 14058 23800 6 mprj_adr_o_user[10]
port 933 nsew signal output
rlabel metal2 s 14922 22600 14978 23800 6 mprj_adr_o_user[11]
port 934 nsew signal output
rlabel metal2 s 15934 22600 15990 23800 6 mprj_adr_o_user[12]
port 935 nsew signal output
rlabel metal2 s 16854 22600 16910 23800 6 mprj_adr_o_user[13]
port 936 nsew signal output
rlabel metal2 s 17774 22600 17830 23800 6 mprj_adr_o_user[14]
port 937 nsew signal output
rlabel metal2 s 18786 22600 18842 23800 6 mprj_adr_o_user[15]
port 938 nsew signal output
rlabel metal2 s 19706 22600 19762 23800 6 mprj_adr_o_user[16]
port 939 nsew signal output
rlabel metal2 s 20718 22600 20774 23800 6 mprj_adr_o_user[17]
port 940 nsew signal output
rlabel metal2 s 21638 22600 21694 23800 6 mprj_adr_o_user[18]
port 941 nsew signal output
rlabel metal2 s 22558 22600 22614 23800 6 mprj_adr_o_user[19]
port 942 nsew signal output
rlabel metal2 s 3974 22600 4030 23800 6 mprj_adr_o_user[1]
port 943 nsew signal output
rlabel metal2 s 23570 22600 23626 23800 6 mprj_adr_o_user[20]
port 944 nsew signal output
rlabel metal2 s 24490 22600 24546 23800 6 mprj_adr_o_user[21]
port 945 nsew signal output
rlabel metal2 s 25410 22600 25466 23800 6 mprj_adr_o_user[22]
port 946 nsew signal output
rlabel metal2 s 26422 22600 26478 23800 6 mprj_adr_o_user[23]
port 947 nsew signal output
rlabel metal2 s 27342 22600 27398 23800 6 mprj_adr_o_user[24]
port 948 nsew signal output
rlabel metal2 s 28354 22600 28410 23800 6 mprj_adr_o_user[25]
port 949 nsew signal output
rlabel metal2 s 29274 22600 29330 23800 6 mprj_adr_o_user[26]
port 950 nsew signal output
rlabel metal2 s 30194 22600 30250 23800 6 mprj_adr_o_user[27]
port 951 nsew signal output
rlabel metal2 s 31206 22600 31262 23800 6 mprj_adr_o_user[28]
port 952 nsew signal output
rlabel metal2 s 32126 22600 32182 23800 6 mprj_adr_o_user[29]
port 953 nsew signal output
rlabel metal2 s 5446 22600 5502 23800 6 mprj_adr_o_user[2]
port 954 nsew signal output
rlabel metal2 s 33046 22600 33102 23800 6 mprj_adr_o_user[30]
port 955 nsew signal output
rlabel metal2 s 34058 22600 34114 23800 6 mprj_adr_o_user[31]
port 956 nsew signal output
rlabel metal2 s 6826 22600 6882 23800 6 mprj_adr_o_user[3]
port 957 nsew signal output
rlabel metal2 s 8298 22600 8354 23800 6 mprj_adr_o_user[4]
port 958 nsew signal output
rlabel metal2 s 9218 22600 9274 23800 6 mprj_adr_o_user[5]
port 959 nsew signal output
rlabel metal2 s 10138 22600 10194 23800 6 mprj_adr_o_user[6]
port 960 nsew signal output
rlabel metal2 s 11150 22600 11206 23800 6 mprj_adr_o_user[7]
port 961 nsew signal output
rlabel metal2 s 12070 22600 12126 23800 6 mprj_adr_o_user[8]
port 962 nsew signal output
rlabel metal2 s 13082 22600 13138 23800 6 mprj_adr_o_user[9]
port 963 nsew signal output
rlabel metal2 s 193310 -400 193366 800 6 mprj_cyc_o_core
port 964 nsew signal input
rlabel metal2 s 1122 22600 1178 23800 6 mprj_cyc_o_user
port 965 nsew signal output
rlabel metal2 s 194874 -400 194930 800 6 mprj_dat_o_core[0]
port 966 nsew signal input
rlabel metal2 s 203890 -400 203946 800 6 mprj_dat_o_core[10]
port 967 nsew signal input
rlabel metal2 s 204626 -400 204682 800 6 mprj_dat_o_core[11]
port 968 nsew signal input
rlabel metal2 s 205454 -400 205510 800 6 mprj_dat_o_core[12]
port 969 nsew signal input
rlabel metal2 s 206190 -400 206246 800 6 mprj_dat_o_core[13]
port 970 nsew signal input
rlabel metal2 s 206926 -400 206982 800 6 mprj_dat_o_core[14]
port 971 nsew signal input
rlabel metal2 s 207662 -400 207718 800 6 mprj_dat_o_core[15]
port 972 nsew signal input
rlabel metal2 s 208398 -400 208454 800 6 mprj_dat_o_core[16]
port 973 nsew signal input
rlabel metal2 s 209226 -400 209282 800 6 mprj_dat_o_core[17]
port 974 nsew signal input
rlabel metal2 s 209962 -400 210018 800 6 mprj_dat_o_core[18]
port 975 nsew signal input
rlabel metal2 s 210698 -400 210754 800 6 mprj_dat_o_core[19]
port 976 nsew signal input
rlabel metal2 s 195978 -400 196034 800 6 mprj_dat_o_core[1]
port 977 nsew signal input
rlabel metal2 s 211434 -400 211490 800 6 mprj_dat_o_core[20]
port 978 nsew signal input
rlabel metal2 s 212170 -400 212226 800 6 mprj_dat_o_core[21]
port 979 nsew signal input
rlabel metal2 s 212998 -400 213054 800 6 mprj_dat_o_core[22]
port 980 nsew signal input
rlabel metal2 s 213734 -400 213790 800 6 mprj_dat_o_core[23]
port 981 nsew signal input
rlabel metal2 s 214470 -400 214526 800 6 mprj_dat_o_core[24]
port 982 nsew signal input
rlabel metal2 s 215206 -400 215262 800 6 mprj_dat_o_core[25]
port 983 nsew signal input
rlabel metal2 s 215942 -400 215998 800 6 mprj_dat_o_core[26]
port 984 nsew signal input
rlabel metal2 s 216770 -400 216826 800 6 mprj_dat_o_core[27]
port 985 nsew signal input
rlabel metal2 s 217506 -400 217562 800 6 mprj_dat_o_core[28]
port 986 nsew signal input
rlabel metal2 s 218242 -400 218298 800 6 mprj_dat_o_core[29]
port 987 nsew signal input
rlabel metal2 s 197082 -400 197138 800 6 mprj_dat_o_core[2]
port 988 nsew signal input
rlabel metal2 s 218978 -400 219034 800 6 mprj_dat_o_core[30]
port 989 nsew signal input
rlabel metal2 s 219714 -400 219770 800 6 mprj_dat_o_core[31]
port 990 nsew signal input
rlabel metal2 s 198278 -400 198334 800 6 mprj_dat_o_core[3]
port 991 nsew signal input
rlabel metal2 s 199382 -400 199438 800 6 mprj_dat_o_core[4]
port 992 nsew signal input
rlabel metal2 s 200118 -400 200174 800 6 mprj_dat_o_core[5]
port 993 nsew signal input
rlabel metal2 s 200854 -400 200910 800 6 mprj_dat_o_core[6]
port 994 nsew signal input
rlabel metal2 s 201682 -400 201738 800 6 mprj_dat_o_core[7]
port 995 nsew signal input
rlabel metal2 s 202418 -400 202474 800 6 mprj_dat_o_core[8]
port 996 nsew signal input
rlabel metal2 s 203154 -400 203210 800 6 mprj_dat_o_core[9]
port 997 nsew signal input
rlabel metal2 s 3054 22600 3110 23800 6 mprj_dat_o_user[0]
port 998 nsew signal output
rlabel metal2 s 14462 22600 14518 23800 6 mprj_dat_o_user[10]
port 999 nsew signal output
rlabel metal2 s 15382 22600 15438 23800 6 mprj_dat_o_user[11]
port 1000 nsew signal output
rlabel metal2 s 16394 22600 16450 23800 6 mprj_dat_o_user[12]
port 1001 nsew signal output
rlabel metal2 s 17314 22600 17370 23800 6 mprj_dat_o_user[13]
port 1002 nsew signal output
rlabel metal2 s 18326 22600 18382 23800 6 mprj_dat_o_user[14]
port 1003 nsew signal output
rlabel metal2 s 19246 22600 19302 23800 6 mprj_dat_o_user[15]
port 1004 nsew signal output
rlabel metal2 s 20166 22600 20222 23800 6 mprj_dat_o_user[16]
port 1005 nsew signal output
rlabel metal2 s 21178 22600 21234 23800 6 mprj_dat_o_user[17]
port 1006 nsew signal output
rlabel metal2 s 22098 22600 22154 23800 6 mprj_dat_o_user[18]
port 1007 nsew signal output
rlabel metal2 s 23018 22600 23074 23800 6 mprj_dat_o_user[19]
port 1008 nsew signal output
rlabel metal2 s 4434 22600 4490 23800 6 mprj_dat_o_user[1]
port 1009 nsew signal output
rlabel metal2 s 24030 22600 24086 23800 6 mprj_dat_o_user[20]
port 1010 nsew signal output
rlabel metal2 s 24950 22600 25006 23800 6 mprj_dat_o_user[21]
port 1011 nsew signal output
rlabel metal2 s 25962 22600 26018 23800 6 mprj_dat_o_user[22]
port 1012 nsew signal output
rlabel metal2 s 26882 22600 26938 23800 6 mprj_dat_o_user[23]
port 1013 nsew signal output
rlabel metal2 s 27802 22600 27858 23800 6 mprj_dat_o_user[24]
port 1014 nsew signal output
rlabel metal2 s 28814 22600 28870 23800 6 mprj_dat_o_user[25]
port 1015 nsew signal output
rlabel metal2 s 29734 22600 29790 23800 6 mprj_dat_o_user[26]
port 1016 nsew signal output
rlabel metal2 s 30654 22600 30710 23800 6 mprj_dat_o_user[27]
port 1017 nsew signal output
rlabel metal2 s 31666 22600 31722 23800 6 mprj_dat_o_user[28]
port 1018 nsew signal output
rlabel metal2 s 32586 22600 32642 23800 6 mprj_dat_o_user[29]
port 1019 nsew signal output
rlabel metal2 s 5906 22600 5962 23800 6 mprj_dat_o_user[2]
port 1020 nsew signal output
rlabel metal2 s 33598 22600 33654 23800 6 mprj_dat_o_user[30]
port 1021 nsew signal output
rlabel metal2 s 34518 22600 34574 23800 6 mprj_dat_o_user[31]
port 1022 nsew signal output
rlabel metal2 s 7286 22600 7342 23800 6 mprj_dat_o_user[3]
port 1023 nsew signal output
rlabel metal2 s 8758 22600 8814 23800 6 mprj_dat_o_user[4]
port 1024 nsew signal output
rlabel metal2 s 9678 22600 9734 23800 6 mprj_dat_o_user[5]
port 1025 nsew signal output
rlabel metal2 s 10690 22600 10746 23800 6 mprj_dat_o_user[6]
port 1026 nsew signal output
rlabel metal2 s 11610 22600 11666 23800 6 mprj_dat_o_user[7]
port 1027 nsew signal output
rlabel metal2 s 12530 22600 12586 23800 6 mprj_dat_o_user[8]
port 1028 nsew signal output
rlabel metal2 s 13542 22600 13598 23800 6 mprj_dat_o_user[9]
port 1029 nsew signal output
rlabel metal2 s 195242 -400 195298 800 6 mprj_sel_o_core[0]
port 1030 nsew signal input
rlabel metal2 s 196346 -400 196402 800 6 mprj_sel_o_core[1]
port 1031 nsew signal input
rlabel metal2 s 197450 -400 197506 800 6 mprj_sel_o_core[2]
port 1032 nsew signal input
rlabel metal2 s 198646 -400 198702 800 6 mprj_sel_o_core[3]
port 1033 nsew signal input
rlabel metal2 s 3514 22600 3570 23800 6 mprj_sel_o_user[0]
port 1034 nsew signal output
rlabel metal2 s 4894 22600 4950 23800 6 mprj_sel_o_user[1]
port 1035 nsew signal output
rlabel metal2 s 6366 22600 6422 23800 6 mprj_sel_o_user[2]
port 1036 nsew signal output
rlabel metal2 s 7746 22600 7802 23800 6 mprj_sel_o_user[3]
port 1037 nsew signal output
rlabel metal2 s 193678 -400 193734 800 6 mprj_stb_o_core
port 1038 nsew signal input
rlabel metal2 s 1582 22600 1638 23800 6 mprj_stb_o_user
port 1039 nsew signal output
rlabel metal2 s 194138 -400 194194 800 6 mprj_we_o_core
port 1040 nsew signal input
rlabel metal2 s 2042 22600 2098 23800 6 mprj_we_o_user
port 1041 nsew signal output
rlabel metal3 s 219200 1096 220400 1216 6 user1_vcc_powergood
port 1042 nsew signal output
rlabel metal3 s 219200 3408 220400 3528 6 user1_vdd_powergood
port 1043 nsew signal output
rlabel metal3 s 219200 5720 220400 5840 6 user2_vcc_powergood
port 1044 nsew signal output
rlabel metal3 s 219200 8032 220400 8152 6 user2_vdd_powergood
port 1045 nsew signal output
rlabel metal2 s 202 22600 258 23800 6 user_clock
port 1046 nsew signal output
rlabel metal2 s 218242 22600 218298 23800 6 user_clock2
port 1047 nsew signal output
rlabel metal3 s 219200 10344 220400 10464 6 user_irq[0]
port 1048 nsew signal output
rlabel metal3 s 219200 12792 220400 12912 6 user_irq[1]
port 1049 nsew signal output
rlabel metal3 s 219200 15104 220400 15224 6 user_irq[2]
port 1050 nsew signal output
rlabel metal2 s 218702 22600 218758 23800 6 user_irq_core[0]
port 1051 nsew signal input
rlabel metal2 s 219162 22600 219218 23800 6 user_irq_core[1]
port 1052 nsew signal input
rlabel metal2 s 219622 22600 219678 23800 6 user_irq_core[2]
port 1053 nsew signal input
rlabel metal3 s 219200 17416 220400 17536 6 user_irq_ena[0]
port 1054 nsew signal input
rlabel metal3 s 219200 19728 220400 19848 6 user_irq_ena[1]
port 1055 nsew signal input
rlabel metal3 s 219200 22040 220400 22160 6 user_irq_ena[2]
port 1056 nsew signal input
rlabel metal2 s 662 22600 718 23800 6 user_reset
port 1057 nsew signal output
rlabel metal3 s -386 23614 220358 23794 6 vccd
port 1058 nsew power bidirectional
rlabel metal3 s -386 -402 220358 -222 8 vccd
port 1059 nsew power bidirectional
rlabel metal4 s 214714 -666 214894 24058 6 vccd
port 1060 nsew power bidirectional
rlabel metal4 s 184614 -666 184794 24058 6 vccd
port 1061 nsew power bidirectional
rlabel metal4 s 154514 -666 154694 24058 6 vccd
port 1062 nsew power bidirectional
rlabel metal4 s 124414 -666 124594 24058 6 vccd
port 1063 nsew power bidirectional
rlabel metal4 s 94314 -666 94494 24058 6 vccd
port 1064 nsew power bidirectional
rlabel metal4 s 64214 -666 64394 24058 6 vccd
port 1065 nsew power bidirectional
rlabel metal4 s 34114 -666 34294 24058 6 vccd
port 1066 nsew power bidirectional
rlabel metal4 s 4014 -666 4194 24058 6 vccd
port 1067 nsew power bidirectional
rlabel metal4 s 220178 -402 220358 23794 6 vccd
port 1068 nsew power bidirectional
rlabel metal4 s -386 -402 -206 23794 4 vccd
port 1069 nsew power bidirectional
rlabel metal3 s -650 23878 220622 24058 6 vssd
port 1070 nsew ground bidirectional
rlabel metal3 s -650 -666 220622 -486 8 vssd
port 1071 nsew ground bidirectional
rlabel metal4 s 220442 -666 220622 24058 6 vssd
port 1072 nsew ground bidirectional
rlabel metal4 s 199664 -666 199844 24058 6 vssd
port 1073 nsew ground bidirectional
rlabel metal4 s 169564 -666 169744 24058 6 vssd
port 1074 nsew ground bidirectional
rlabel metal4 s 139464 -666 139644 24058 6 vssd
port 1075 nsew ground bidirectional
rlabel metal4 s 109364 -666 109544 24058 6 vssd
port 1076 nsew ground bidirectional
rlabel metal4 s 79264 -666 79444 24058 6 vssd
port 1077 nsew ground bidirectional
rlabel metal4 s 49164 -666 49344 24058 6 vssd
port 1078 nsew ground bidirectional
rlabel metal4 s 19064 -666 19244 24058 6 vssd
port 1079 nsew ground bidirectional
rlabel metal4 s -650 -666 -470 24058 4 vssd
port 1080 nsew ground bidirectional
rlabel metal3 s -914 24142 220886 24322 6 vccd1
port 1081 nsew power bidirectional
rlabel metal3 s -914 -930 220886 -750 8 vccd1
port 1082 nsew power bidirectional
rlabel metal4 s 215534 -1194 215714 24586 6 vccd1
port 1083 nsew power bidirectional
rlabel metal4 s 185434 -1194 185614 24586 6 vccd1
port 1084 nsew power bidirectional
rlabel metal4 s 155334 -1194 155514 24586 6 vccd1
port 1085 nsew power bidirectional
rlabel metal4 s 125234 -1194 125414 24586 6 vccd1
port 1086 nsew power bidirectional
rlabel metal4 s 95134 -1194 95314 24586 6 vccd1
port 1087 nsew power bidirectional
rlabel metal4 s 65034 -1194 65214 24586 6 vccd1
port 1088 nsew power bidirectional
rlabel metal4 s 34934 -1194 35114 24586 6 vccd1
port 1089 nsew power bidirectional
rlabel metal4 s 4834 -1194 5014 24586 6 vccd1
port 1090 nsew power bidirectional
rlabel metal4 s 220706 -930 220886 24322 6 vccd1
port 1091 nsew power bidirectional
rlabel metal4 s -914 -930 -734 24322 4 vccd1
port 1092 nsew power bidirectional
rlabel metal3 s -1178 24406 221150 24586 6 vssd1
port 1093 nsew ground bidirectional
rlabel metal3 s -1178 -1194 221150 -1014 8 vssd1
port 1094 nsew ground bidirectional
rlabel metal4 s 220970 -1194 221150 24586 6 vssd1
port 1095 nsew ground bidirectional
rlabel metal4 s 200484 -1194 200664 24586 6 vssd1
port 1096 nsew ground bidirectional
rlabel metal4 s 170384 -1194 170564 24586 6 vssd1
port 1097 nsew ground bidirectional
rlabel metal4 s 140284 -1194 140464 24586 6 vssd1
port 1098 nsew ground bidirectional
rlabel metal4 s 110184 -1194 110364 24586 6 vssd1
port 1099 nsew ground bidirectional
rlabel metal4 s 80084 -1194 80264 24586 6 vssd1
port 1100 nsew ground bidirectional
rlabel metal4 s 49984 -1194 50164 24586 6 vssd1
port 1101 nsew ground bidirectional
rlabel metal4 s 19884 -1194 20064 24586 6 vssd1
port 1102 nsew ground bidirectional
rlabel metal4 s -1178 -1194 -998 24586 4 vssd1
port 1103 nsew ground bidirectional
rlabel metal3 s -1442 24670 221414 24850 6 vccd2
port 1104 nsew power bidirectional
rlabel metal3 s -1442 -1458 221414 -1278 8 vccd2
port 1105 nsew power bidirectional
rlabel metal4 s 216354 -1722 216534 25114 6 vccd2
port 1106 nsew power bidirectional
rlabel metal4 s 186254 -1722 186434 25114 6 vccd2
port 1107 nsew power bidirectional
rlabel metal4 s 156154 -1722 156334 25114 6 vccd2
port 1108 nsew power bidirectional
rlabel metal4 s 126054 -1722 126234 25114 6 vccd2
port 1109 nsew power bidirectional
rlabel metal4 s 95954 -1722 96134 25114 6 vccd2
port 1110 nsew power bidirectional
rlabel metal4 s 65854 -1722 66034 25114 6 vccd2
port 1111 nsew power bidirectional
rlabel metal4 s 35754 -1722 35934 25114 6 vccd2
port 1112 nsew power bidirectional
rlabel metal4 s 5654 -1722 5834 25114 6 vccd2
port 1113 nsew power bidirectional
rlabel metal4 s 221234 -1458 221414 24850 6 vccd2
port 1114 nsew power bidirectional
rlabel metal4 s -1442 -1458 -1262 24850 4 vccd2
port 1115 nsew power bidirectional
rlabel metal3 s -1706 24934 221678 25114 6 vssd2
port 1116 nsew ground bidirectional
rlabel metal3 s -1706 -1722 221678 -1542 8 vssd2
port 1117 nsew ground bidirectional
rlabel metal4 s 221498 -1722 221678 25114 6 vssd2
port 1118 nsew ground bidirectional
rlabel metal4 s 201304 -1722 201484 25114 6 vssd2
port 1119 nsew ground bidirectional
rlabel metal4 s 171204 -1722 171384 25114 6 vssd2
port 1120 nsew ground bidirectional
rlabel metal4 s 141104 -1722 141284 25114 6 vssd2
port 1121 nsew ground bidirectional
rlabel metal4 s 111004 -1722 111184 25114 6 vssd2
port 1122 nsew ground bidirectional
rlabel metal4 s 80904 -1722 81084 25114 6 vssd2
port 1123 nsew ground bidirectional
rlabel metal4 s 50804 -1722 50984 25114 6 vssd2
port 1124 nsew ground bidirectional
rlabel metal4 s 20704 -1722 20884 25114 6 vssd2
port 1125 nsew ground bidirectional
rlabel metal4 s -1706 -1722 -1526 25114 4 vssd2
port 1126 nsew ground bidirectional
rlabel metal3 s -1970 25198 221942 25378 6 vdda1
port 1127 nsew power bidirectional
rlabel metal3 s -1970 -1986 221942 -1806 8 vdda1
port 1128 nsew power bidirectional
rlabel metal4 s 217174 -2250 217354 25642 6 vdda1
port 1129 nsew power bidirectional
rlabel metal4 s 187074 -2250 187254 25642 6 vdda1
port 1130 nsew power bidirectional
rlabel metal4 s 156974 -2250 157154 25642 6 vdda1
port 1131 nsew power bidirectional
rlabel metal4 s 126874 -2250 127054 25642 6 vdda1
port 1132 nsew power bidirectional
rlabel metal4 s 96774 -2250 96954 25642 6 vdda1
port 1133 nsew power bidirectional
rlabel metal4 s 66674 -2250 66854 25642 6 vdda1
port 1134 nsew power bidirectional
rlabel metal4 s 36574 -2250 36754 25642 6 vdda1
port 1135 nsew power bidirectional
rlabel metal4 s 6474 -2250 6654 25642 6 vdda1
port 1136 nsew power bidirectional
rlabel metal4 s 221762 -1986 221942 25378 6 vdda1
port 1137 nsew power bidirectional
rlabel metal4 s -1970 -1986 -1790 25378 4 vdda1
port 1138 nsew power bidirectional
rlabel metal3 s -2234 25462 222206 25642 6 vssa1
port 1139 nsew ground bidirectional
rlabel metal3 s -2234 -2250 222206 -2070 8 vssa1
port 1140 nsew ground bidirectional
rlabel metal4 s 222026 -2250 222206 25642 6 vssa1
port 1141 nsew ground bidirectional
rlabel metal4 s 202124 -2250 202304 25642 6 vssa1
port 1142 nsew ground bidirectional
rlabel metal4 s 172024 -2250 172204 25642 6 vssa1
port 1143 nsew ground bidirectional
rlabel metal4 s 141924 -2250 142104 25642 6 vssa1
port 1144 nsew ground bidirectional
rlabel metal4 s 111824 -2250 112004 25642 6 vssa1
port 1145 nsew ground bidirectional
rlabel metal4 s 81724 -2250 81904 25642 6 vssa1
port 1146 nsew ground bidirectional
rlabel metal4 s 51624 -2250 51804 25642 6 vssa1
port 1147 nsew ground bidirectional
rlabel metal4 s 21524 -2250 21704 25642 6 vssa1
port 1148 nsew ground bidirectional
rlabel metal4 s -2234 -2250 -2054 25642 4 vssa1
port 1149 nsew ground bidirectional
rlabel metal3 s -2498 25726 222470 25906 6 vdda2
port 1150 nsew power bidirectional
rlabel metal3 s -2498 -2514 222470 -2334 8 vdda2
port 1151 nsew power bidirectional
rlabel metal4 s 217994 -2778 218174 26170 6 vdda2
port 1152 nsew power bidirectional
rlabel metal4 s 187894 -2778 188074 26170 6 vdda2
port 1153 nsew power bidirectional
rlabel metal4 s 157794 -2778 157974 26170 6 vdda2
port 1154 nsew power bidirectional
rlabel metal4 s 127694 -2778 127874 26170 6 vdda2
port 1155 nsew power bidirectional
rlabel metal4 s 97594 -2778 97774 26170 6 vdda2
port 1156 nsew power bidirectional
rlabel metal4 s 67494 -2778 67674 26170 6 vdda2
port 1157 nsew power bidirectional
rlabel metal4 s 37394 -2778 37574 26170 6 vdda2
port 1158 nsew power bidirectional
rlabel metal4 s 7294 -2778 7474 26170 6 vdda2
port 1159 nsew power bidirectional
rlabel metal4 s 222290 -2514 222470 25906 6 vdda2
port 1160 nsew power bidirectional
rlabel metal4 s -2498 -2514 -2318 25906 4 vdda2
port 1161 nsew power bidirectional
rlabel metal3 s -2762 25990 222734 26170 6 vssa2
port 1162 nsew ground bidirectional
rlabel metal3 s -2762 -2778 222734 -2598 8 vssa2
port 1163 nsew ground bidirectional
rlabel metal4 s 222554 -2778 222734 26170 6 vssa2
port 1164 nsew ground bidirectional
rlabel metal4 s 202944 -2778 203124 26170 6 vssa2
port 1165 nsew ground bidirectional
rlabel metal4 s 172844 -2778 173024 26170 6 vssa2
port 1166 nsew ground bidirectional
rlabel metal4 s 142744 -2778 142924 26170 6 vssa2
port 1167 nsew ground bidirectional
rlabel metal4 s 112644 -2778 112824 26170 6 vssa2
port 1168 nsew ground bidirectional
rlabel metal4 s 82544 -2778 82724 26170 6 vssa2
port 1169 nsew ground bidirectional
rlabel metal4 s 52444 -2778 52624 26170 6 vssa2
port 1170 nsew ground bidirectional
rlabel metal4 s 22344 -2778 22524 26170 6 vssa2
port 1171 nsew ground bidirectional
rlabel metal4 s -2762 -2778 -2582 26170 4 vssa2
port 1172 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 220000 23400
string GDS_FILE /project/openlane/mgmt_protect/runs/mgmt_protect/results/magic/mgmt_protect.gds
string GDS_END 8297048
string GDS_START 620638
string LEFview TRUE
<< end >>
