magic
tech sky130A
magscale 12 1
timestamp 1598766293
<< metal5 >>
rect 0 80 15 105
rect 30 80 45 105
rect 0 70 45 80
rect 0 60 40 70
rect 0 45 35 60
rect 0 35 40 45
rect 0 25 45 35
rect 0 0 15 25
rect 30 0 45 25
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
