VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mgmt_core
  CLASS BLOCK ;
  FOREIGN mgmt_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 2150.000 BY 850.000 ;
  PIN clock
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 2.400 ;
    END
  END clock
  PIN core_clk
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2147.600 346.840 2150.000 347.440 ;
    END
  END core_clk
  PIN core_rstn
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2147.600 424.360 2150.000 424.960 ;
    END
  END core_rstn
  PIN flash_clk
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 537.370 0.000 537.650 2.400 ;
    END
  END flash_clk
  PIN flash_clk_ieb
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 634.890 0.000 635.170 2.400 ;
    END
  END flash_clk_ieb
  PIN flash_clk_oeb
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 732.870 0.000 733.150 2.400 ;
    END
  END flash_clk_oeb
  PIN flash_csb
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 2.400 ;
    END
  END flash_csb
  PIN flash_csb_ieb
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 341.870 0.000 342.150 2.400 ;
    END
  END flash_csb_ieb
  PIN flash_csb_oeb
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 439.390 0.000 439.670 2.400 ;
    END
  END flash_csb_oeb
  PIN flash_io0_di
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 830.390 0.000 830.670 2.400 ;
    END
  END flash_io0_di
  PIN flash_io0_do
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 928.370 0.000 928.650 2.400 ;
    END
  END flash_io0_do
  PIN flash_io0_ieb
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1025.890 0.000 1026.170 2.400 ;
    END
  END flash_io0_ieb
  PIN flash_io0_oeb
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1123.870 0.000 1124.150 2.400 ;
    END
  END flash_io0_oeb
  PIN flash_io1_di
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1221.390 0.000 1221.670 2.400 ;
    END
  END flash_io1_di
  PIN flash_io1_do
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1318.910 0.000 1319.190 2.400 ;
    END
  END flash_io1_do
  PIN flash_io1_ieb
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1416.890 0.000 1417.170 2.400 ;
    END
  END flash_io1_ieb
  PIN flash_io1_oeb
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1514.410 0.000 1514.690 2.400 ;
    END
  END flash_io1_oeb
  PIN gpio_in_pad
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1612.390 0.000 1612.670 2.400 ;
    END
  END gpio_in_pad
  PIN gpio_inenb_pad
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1709.910 0.000 1710.190 2.400 ;
    END
  END gpio_inenb_pad
  PIN gpio_mode0_pad
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1807.890 0.000 1808.170 2.400 ;
    END
  END gpio_mode0_pad
  PIN gpio_mode1_pad
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1905.410 0.000 1905.690 2.400 ;
    END
  END gpio_mode1_pad
  PIN gpio_out_pad
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2003.390 0.000 2003.670 2.400 ;
    END
  END gpio_out_pad
  PIN gpio_outenb_pad
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2100.910 0.000 2101.190 2.400 ;
    END
  END gpio_outenb_pad
  PIN jtag_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2147.600 501.200 2150.000 501.800 ;
    END
  END jtag_out
  PIN jtag_outenb
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2147.600 578.720 2150.000 579.320 ;
    END
  END jtag_outenb
  PIN la_input[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.470 847.600 1.750 850.000 ;
    END
  END la_input[0]
  PIN la_input[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 940.330 847.600 940.610 850.000 ;
    END
  END la_input[100]
  PIN la_input[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 949.530 847.600 949.810 850.000 ;
    END
  END la_input[101]
  PIN la_input[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 958.730 847.600 959.010 850.000 ;
    END
  END la_input[102]
  PIN la_input[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 968.390 847.600 968.670 850.000 ;
    END
  END la_input[103]
  PIN la_input[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 977.590 847.600 977.870 850.000 ;
    END
  END la_input[104]
  PIN la_input[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 987.250 847.600 987.530 850.000 ;
    END
  END la_input[105]
  PIN la_input[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 996.450 847.600 996.730 850.000 ;
    END
  END la_input[106]
  PIN la_input[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1005.650 847.600 1005.930 850.000 ;
    END
  END la_input[107]
  PIN la_input[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1015.310 847.600 1015.590 850.000 ;
    END
  END la_input[108]
  PIN la_input[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1024.510 847.600 1024.790 850.000 ;
    END
  END la_input[109]
  PIN la_input[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 95.310 847.600 95.590 850.000 ;
    END
  END la_input[10]
  PIN la_input[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1034.170 847.600 1034.450 850.000 ;
    END
  END la_input[110]
  PIN la_input[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1043.370 847.600 1043.650 850.000 ;
    END
  END la_input[111]
  PIN la_input[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1052.570 847.600 1052.850 850.000 ;
    END
  END la_input[112]
  PIN la_input[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1062.230 847.600 1062.510 850.000 ;
    END
  END la_input[113]
  PIN la_input[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1071.430 847.600 1071.710 850.000 ;
    END
  END la_input[114]
  PIN la_input[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1081.090 847.600 1081.370 850.000 ;
    END
  END la_input[115]
  PIN la_input[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1090.290 847.600 1090.570 850.000 ;
    END
  END la_input[116]
  PIN la_input[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1099.950 847.600 1100.230 850.000 ;
    END
  END la_input[117]
  PIN la_input[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1109.150 847.600 1109.430 850.000 ;
    END
  END la_input[118]
  PIN la_input[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1118.350 847.600 1118.630 850.000 ;
    END
  END la_input[119]
  PIN la_input[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.510 847.600 104.790 850.000 ;
    END
  END la_input[11]
  PIN la_input[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1128.010 847.600 1128.290 850.000 ;
    END
  END la_input[120]
  PIN la_input[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1137.210 847.600 1137.490 850.000 ;
    END
  END la_input[121]
  PIN la_input[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1146.870 847.600 1147.150 850.000 ;
    END
  END la_input[122]
  PIN la_input[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1156.070 847.600 1156.350 850.000 ;
    END
  END la_input[123]
  PIN la_input[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1165.270 847.600 1165.550 850.000 ;
    END
  END la_input[124]
  PIN la_input[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1174.930 847.600 1175.210 850.000 ;
    END
  END la_input[125]
  PIN la_input[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1184.130 847.600 1184.410 850.000 ;
    END
  END la_input[126]
  PIN la_input[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1193.790 847.600 1194.070 850.000 ;
    END
  END la_input[127]
  PIN la_input[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 113.710 847.600 113.990 850.000 ;
    END
  END la_input[12]
  PIN la_input[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 123.370 847.600 123.650 850.000 ;
    END
  END la_input[13]
  PIN la_input[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 132.570 847.600 132.850 850.000 ;
    END
  END la_input[14]
  PIN la_input[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 142.230 847.600 142.510 850.000 ;
    END
  END la_input[15]
  PIN la_input[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 151.430 847.600 151.710 850.000 ;
    END
  END la_input[16]
  PIN la_input[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 160.630 847.600 160.910 850.000 ;
    END
  END la_input[17]
  PIN la_input[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 170.290 847.600 170.570 850.000 ;
    END
  END la_input[18]
  PIN la_input[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 179.490 847.600 179.770 850.000 ;
    END
  END la_input[19]
  PIN la_input[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.670 847.600 10.950 850.000 ;
    END
  END la_input[1]
  PIN la_input[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 189.150 847.600 189.430 850.000 ;
    END
  END la_input[20]
  PIN la_input[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 198.350 847.600 198.630 850.000 ;
    END
  END la_input[21]
  PIN la_input[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 208.010 847.600 208.290 850.000 ;
    END
  END la_input[22]
  PIN la_input[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 217.210 847.600 217.490 850.000 ;
    END
  END la_input[23]
  PIN la_input[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 226.410 847.600 226.690 850.000 ;
    END
  END la_input[24]
  PIN la_input[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 236.070 847.600 236.350 850.000 ;
    END
  END la_input[25]
  PIN la_input[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 245.270 847.600 245.550 850.000 ;
    END
  END la_input[26]
  PIN la_input[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 254.930 847.600 255.210 850.000 ;
    END
  END la_input[27]
  PIN la_input[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 264.130 847.600 264.410 850.000 ;
    END
  END la_input[28]
  PIN la_input[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 273.330 847.600 273.610 850.000 ;
    END
  END la_input[29]
  PIN la_input[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.870 847.600 20.150 850.000 ;
    END
  END la_input[2]
  PIN la_input[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 282.990 847.600 283.270 850.000 ;
    END
  END la_input[30]
  PIN la_input[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 292.190 847.600 292.470 850.000 ;
    END
  END la_input[31]
  PIN la_input[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 301.850 847.600 302.130 850.000 ;
    END
  END la_input[32]
  PIN la_input[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 311.050 847.600 311.330 850.000 ;
    END
  END la_input[33]
  PIN la_input[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 320.250 847.600 320.530 850.000 ;
    END
  END la_input[34]
  PIN la_input[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 329.910 847.600 330.190 850.000 ;
    END
  END la_input[35]
  PIN la_input[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 339.110 847.600 339.390 850.000 ;
    END
  END la_input[36]
  PIN la_input[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 348.770 847.600 349.050 850.000 ;
    END
  END la_input[37]
  PIN la_input[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 357.970 847.600 358.250 850.000 ;
    END
  END la_input[38]
  PIN la_input[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 367.630 847.600 367.910 850.000 ;
    END
  END la_input[39]
  PIN la_input[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.530 847.600 29.810 850.000 ;
    END
  END la_input[3]
  PIN la_input[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 376.830 847.600 377.110 850.000 ;
    END
  END la_input[40]
  PIN la_input[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 386.030 847.600 386.310 850.000 ;
    END
  END la_input[41]
  PIN la_input[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 395.690 847.600 395.970 850.000 ;
    END
  END la_input[42]
  PIN la_input[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 404.890 847.600 405.170 850.000 ;
    END
  END la_input[43]
  PIN la_input[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 414.550 847.600 414.830 850.000 ;
    END
  END la_input[44]
  PIN la_input[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 423.750 847.600 424.030 850.000 ;
    END
  END la_input[45]
  PIN la_input[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 432.950 847.600 433.230 850.000 ;
    END
  END la_input[46]
  PIN la_input[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 442.610 847.600 442.890 850.000 ;
    END
  END la_input[47]
  PIN la_input[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 451.810 847.600 452.090 850.000 ;
    END
  END la_input[48]
  PIN la_input[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 461.470 847.600 461.750 850.000 ;
    END
  END la_input[49]
  PIN la_input[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.730 847.600 39.010 850.000 ;
    END
  END la_input[4]
  PIN la_input[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 470.670 847.600 470.950 850.000 ;
    END
  END la_input[50]
  PIN la_input[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 479.870 847.600 480.150 850.000 ;
    END
  END la_input[51]
  PIN la_input[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 489.530 847.600 489.810 850.000 ;
    END
  END la_input[52]
  PIN la_input[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 498.730 847.600 499.010 850.000 ;
    END
  END la_input[53]
  PIN la_input[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 508.390 847.600 508.670 850.000 ;
    END
  END la_input[54]
  PIN la_input[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 517.590 847.600 517.870 850.000 ;
    END
  END la_input[55]
  PIN la_input[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 526.790 847.600 527.070 850.000 ;
    END
  END la_input[56]
  PIN la_input[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 536.450 847.600 536.730 850.000 ;
    END
  END la_input[57]
  PIN la_input[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 545.650 847.600 545.930 850.000 ;
    END
  END la_input[58]
  PIN la_input[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 555.310 847.600 555.590 850.000 ;
    END
  END la_input[59]
  PIN la_input[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.390 847.600 48.670 850.000 ;
    END
  END la_input[5]
  PIN la_input[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 564.510 847.600 564.790 850.000 ;
    END
  END la_input[60]
  PIN la_input[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 574.170 847.600 574.450 850.000 ;
    END
  END la_input[61]
  PIN la_input[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 583.370 847.600 583.650 850.000 ;
    END
  END la_input[62]
  PIN la_input[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 592.570 847.600 592.850 850.000 ;
    END
  END la_input[63]
  PIN la_input[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 602.230 847.600 602.510 850.000 ;
    END
  END la_input[64]
  PIN la_input[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 611.430 847.600 611.710 850.000 ;
    END
  END la_input[65]
  PIN la_input[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 621.090 847.600 621.370 850.000 ;
    END
  END la_input[66]
  PIN la_input[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 630.290 847.600 630.570 850.000 ;
    END
  END la_input[67]
  PIN la_input[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 639.490 847.600 639.770 850.000 ;
    END
  END la_input[68]
  PIN la_input[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 649.150 847.600 649.430 850.000 ;
    END
  END la_input[69]
  PIN la_input[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.590 847.600 57.870 850.000 ;
    END
  END la_input[6]
  PIN la_input[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 658.350 847.600 658.630 850.000 ;
    END
  END la_input[70]
  PIN la_input[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.010 847.600 668.290 850.000 ;
    END
  END la_input[71]
  PIN la_input[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 677.210 847.600 677.490 850.000 ;
    END
  END la_input[72]
  PIN la_input[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 686.410 847.600 686.690 850.000 ;
    END
  END la_input[73]
  PIN la_input[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 696.070 847.600 696.350 850.000 ;
    END
  END la_input[74]
  PIN la_input[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 705.270 847.600 705.550 850.000 ;
    END
  END la_input[75]
  PIN la_input[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 714.930 847.600 715.210 850.000 ;
    END
  END la_input[76]
  PIN la_input[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 724.130 847.600 724.410 850.000 ;
    END
  END la_input[77]
  PIN la_input[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 733.790 847.600 734.070 850.000 ;
    END
  END la_input[78]
  PIN la_input[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 742.990 847.600 743.270 850.000 ;
    END
  END la_input[79]
  PIN la_input[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.790 847.600 67.070 850.000 ;
    END
  END la_input[7]
  PIN la_input[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 752.190 847.600 752.470 850.000 ;
    END
  END la_input[80]
  PIN la_input[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 761.850 847.600 762.130 850.000 ;
    END
  END la_input[81]
  PIN la_input[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 771.050 847.600 771.330 850.000 ;
    END
  END la_input[82]
  PIN la_input[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 780.710 847.600 780.990 850.000 ;
    END
  END la_input[83]
  PIN la_input[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 789.910 847.600 790.190 850.000 ;
    END
  END la_input[84]
  PIN la_input[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 799.110 847.600 799.390 850.000 ;
    END
  END la_input[85]
  PIN la_input[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 808.770 847.600 809.050 850.000 ;
    END
  END la_input[86]
  PIN la_input[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 817.970 847.600 818.250 850.000 ;
    END
  END la_input[87]
  PIN la_input[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 827.630 847.600 827.910 850.000 ;
    END
  END la_input[88]
  PIN la_input[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 836.830 847.600 837.110 850.000 ;
    END
  END la_input[89]
  PIN la_input[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.450 847.600 76.730 850.000 ;
    END
  END la_input[8]
  PIN la_input[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 846.030 847.600 846.310 850.000 ;
    END
  END la_input[90]
  PIN la_input[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 855.690 847.600 855.970 850.000 ;
    END
  END la_input[91]
  PIN la_input[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 864.890 847.600 865.170 850.000 ;
    END
  END la_input[92]
  PIN la_input[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 874.550 847.600 874.830 850.000 ;
    END
  END la_input[93]
  PIN la_input[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 883.750 847.600 884.030 850.000 ;
    END
  END la_input[94]
  PIN la_input[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 892.950 847.600 893.230 850.000 ;
    END
  END la_input[95]
  PIN la_input[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 902.610 847.600 902.890 850.000 ;
    END
  END la_input[96]
  PIN la_input[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 911.810 847.600 912.090 850.000 ;
    END
  END la_input[97]
  PIN la_input[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 921.470 847.600 921.750 850.000 ;
    END
  END la_input[98]
  PIN la_input[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 930.670 847.600 930.950 850.000 ;
    END
  END la_input[99]
  PIN la_input[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.650 847.600 85.930 850.000 ;
    END
  END la_input[9]
  PIN la_oen[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4.230 847.600 4.510 850.000 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 943.090 847.600 943.370 850.000 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 952.750 847.600 953.030 850.000 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 961.950 847.600 962.230 850.000 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 971.610 847.600 971.890 850.000 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 980.810 847.600 981.090 850.000 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 990.010 847.600 990.290 850.000 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 999.670 847.600 999.950 850.000 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1008.870 847.600 1009.150 850.000 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1018.530 847.600 1018.810 850.000 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1027.730 847.600 1028.010 850.000 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.070 847.600 98.350 850.000 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1036.930 847.600 1037.210 850.000 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1046.590 847.600 1046.870 850.000 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1055.790 847.600 1056.070 850.000 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1065.450 847.600 1065.730 850.000 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1074.650 847.600 1074.930 850.000 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1084.310 847.600 1084.590 850.000 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1093.510 847.600 1093.790 850.000 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1102.710 847.600 1102.990 850.000 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1112.370 847.600 1112.650 850.000 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1121.570 847.600 1121.850 850.000 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 107.730 847.600 108.010 850.000 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1131.230 847.600 1131.510 850.000 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1140.430 847.600 1140.710 850.000 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1149.630 847.600 1149.910 850.000 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1159.290 847.600 1159.570 850.000 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1168.490 847.600 1168.770 850.000 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1178.150 847.600 1178.430 850.000 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1187.350 847.600 1187.630 850.000 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1196.550 847.600 1196.830 850.000 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 116.930 847.600 117.210 850.000 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 126.590 847.600 126.870 850.000 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 135.790 847.600 136.070 850.000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 144.990 847.600 145.270 850.000 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 154.650 847.600 154.930 850.000 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 163.850 847.600 164.130 850.000 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 173.510 847.600 173.790 850.000 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 182.710 847.600 182.990 850.000 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 13.890 847.600 14.170 850.000 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 192.370 847.600 192.650 850.000 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 201.570 847.600 201.850 850.000 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 210.770 847.600 211.050 850.000 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 220.430 847.600 220.710 850.000 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 229.630 847.600 229.910 850.000 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 239.290 847.600 239.570 850.000 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 248.490 847.600 248.770 850.000 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 257.690 847.600 257.970 850.000 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 267.350 847.600 267.630 850.000 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 276.550 847.600 276.830 850.000 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 23.090 847.600 23.370 850.000 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 286.210 847.600 286.490 850.000 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 295.410 847.600 295.690 850.000 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 304.610 847.600 304.890 850.000 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 314.270 847.600 314.550 850.000 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 323.470 847.600 323.750 850.000 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 333.130 847.600 333.410 850.000 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 342.330 847.600 342.610 850.000 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 351.530 847.600 351.810 850.000 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 361.190 847.600 361.470 850.000 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 370.390 847.600 370.670 850.000 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 32.750 847.600 33.030 850.000 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 380.050 847.600 380.330 850.000 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 389.250 847.600 389.530 850.000 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 398.910 847.600 399.190 850.000 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 408.110 847.600 408.390 850.000 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 417.310 847.600 417.590 850.000 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 426.970 847.600 427.250 850.000 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 436.170 847.600 436.450 850.000 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 445.830 847.600 446.110 850.000 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 455.030 847.600 455.310 850.000 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 464.230 847.600 464.510 850.000 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.950 847.600 42.230 850.000 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 473.890 847.600 474.170 850.000 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 483.090 847.600 483.370 850.000 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 492.750 847.600 493.030 850.000 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 501.950 847.600 502.230 850.000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 511.150 847.600 511.430 850.000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 520.810 847.600 521.090 850.000 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 530.010 847.600 530.290 850.000 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 539.670 847.600 539.950 850.000 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 548.870 847.600 549.150 850.000 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 558.530 847.600 558.810 850.000 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 51.150 847.600 51.430 850.000 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 567.730 847.600 568.010 850.000 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 576.930 847.600 577.210 850.000 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 586.590 847.600 586.870 850.000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 595.790 847.600 596.070 850.000 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 605.450 847.600 605.730 850.000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 614.650 847.600 614.930 850.000 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 623.850 847.600 624.130 850.000 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 633.510 847.600 633.790 850.000 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 642.710 847.600 642.990 850.000 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 652.370 847.600 652.650 850.000 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 60.810 847.600 61.090 850.000 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 661.570 847.600 661.850 850.000 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 670.770 847.600 671.050 850.000 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 680.430 847.600 680.710 850.000 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 689.630 847.600 689.910 850.000 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 699.290 847.600 699.570 850.000 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 708.490 847.600 708.770 850.000 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 718.150 847.600 718.430 850.000 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 727.350 847.600 727.630 850.000 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 736.550 847.600 736.830 850.000 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 746.210 847.600 746.490 850.000 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 70.010 847.600 70.290 850.000 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 755.410 847.600 755.690 850.000 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 765.070 847.600 765.350 850.000 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 774.270 847.600 774.550 850.000 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 783.470 847.600 783.750 850.000 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 793.130 847.600 793.410 850.000 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 802.330 847.600 802.610 850.000 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 811.990 847.600 812.270 850.000 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 821.190 847.600 821.470 850.000 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 830.390 847.600 830.670 850.000 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 840.050 847.600 840.330 850.000 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.670 847.600 79.950 850.000 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 849.250 847.600 849.530 850.000 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 858.910 847.600 859.190 850.000 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 868.110 847.600 868.390 850.000 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 877.310 847.600 877.590 850.000 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 886.970 847.600 887.250 850.000 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 896.170 847.600 896.450 850.000 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 905.830 847.600 906.110 850.000 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 915.030 847.600 915.310 850.000 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 924.690 847.600 924.970 850.000 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 933.890 847.600 934.170 850.000 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.870 847.600 89.150 850.000 ;
    END
  END la_oen[9]
  PIN la_output[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 7.450 847.600 7.730 850.000 ;
    END
  END la_output[0]
  PIN la_output[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 946.310 847.600 946.590 850.000 ;
    END
  END la_output[100]
  PIN la_output[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 955.970 847.600 956.250 850.000 ;
    END
  END la_output[101]
  PIN la_output[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 965.170 847.600 965.450 850.000 ;
    END
  END la_output[102]
  PIN la_output[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 974.370 847.600 974.650 850.000 ;
    END
  END la_output[103]
  PIN la_output[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 984.030 847.600 984.310 850.000 ;
    END
  END la_output[104]
  PIN la_output[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 993.230 847.600 993.510 850.000 ;
    END
  END la_output[105]
  PIN la_output[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1002.890 847.600 1003.170 850.000 ;
    END
  END la_output[106]
  PIN la_output[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1012.090 847.600 1012.370 850.000 ;
    END
  END la_output[107]
  PIN la_output[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1021.290 847.600 1021.570 850.000 ;
    END
  END la_output[108]
  PIN la_output[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1030.950 847.600 1031.230 850.000 ;
    END
  END la_output[109]
  PIN la_output[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.290 847.600 101.570 850.000 ;
    END
  END la_output[10]
  PIN la_output[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1040.150 847.600 1040.430 850.000 ;
    END
  END la_output[110]
  PIN la_output[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1049.810 847.600 1050.090 850.000 ;
    END
  END la_output[111]
  PIN la_output[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1059.010 847.600 1059.290 850.000 ;
    END
  END la_output[112]
  PIN la_output[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1068.210 847.600 1068.490 850.000 ;
    END
  END la_output[113]
  PIN la_output[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1077.870 847.600 1078.150 850.000 ;
    END
  END la_output[114]
  PIN la_output[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1087.070 847.600 1087.350 850.000 ;
    END
  END la_output[115]
  PIN la_output[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1096.730 847.600 1097.010 850.000 ;
    END
  END la_output[116]
  PIN la_output[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1105.930 847.600 1106.210 850.000 ;
    END
  END la_output[117]
  PIN la_output[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1115.590 847.600 1115.870 850.000 ;
    END
  END la_output[118]
  PIN la_output[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1124.790 847.600 1125.070 850.000 ;
    END
  END la_output[119]
  PIN la_output[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.950 847.600 111.230 850.000 ;
    END
  END la_output[11]
  PIN la_output[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1133.990 847.600 1134.270 850.000 ;
    END
  END la_output[120]
  PIN la_output[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1143.650 847.600 1143.930 850.000 ;
    END
  END la_output[121]
  PIN la_output[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1152.850 847.600 1153.130 850.000 ;
    END
  END la_output[122]
  PIN la_output[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1162.510 847.600 1162.790 850.000 ;
    END
  END la_output[123]
  PIN la_output[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1171.710 847.600 1171.990 850.000 ;
    END
  END la_output[124]
  PIN la_output[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1180.910 847.600 1181.190 850.000 ;
    END
  END la_output[125]
  PIN la_output[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1190.570 847.600 1190.850 850.000 ;
    END
  END la_output[126]
  PIN la_output[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1199.770 847.600 1200.050 850.000 ;
    END
  END la_output[127]
  PIN la_output[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 120.150 847.600 120.430 850.000 ;
    END
  END la_output[12]
  PIN la_output[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.350 847.600 129.630 850.000 ;
    END
  END la_output[13]
  PIN la_output[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 139.010 847.600 139.290 850.000 ;
    END
  END la_output[14]
  PIN la_output[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 148.210 847.600 148.490 850.000 ;
    END
  END la_output[15]
  PIN la_output[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 157.870 847.600 158.150 850.000 ;
    END
  END la_output[16]
  PIN la_output[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 167.070 847.600 167.350 850.000 ;
    END
  END la_output[17]
  PIN la_output[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 176.270 847.600 176.550 850.000 ;
    END
  END la_output[18]
  PIN la_output[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 185.930 847.600 186.210 850.000 ;
    END
  END la_output[19]
  PIN la_output[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 17.110 847.600 17.390 850.000 ;
    END
  END la_output[1]
  PIN la_output[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 195.130 847.600 195.410 850.000 ;
    END
  END la_output[20]
  PIN la_output[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 204.790 847.600 205.070 850.000 ;
    END
  END la_output[21]
  PIN la_output[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 213.990 847.600 214.270 850.000 ;
    END
  END la_output[22]
  PIN la_output[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 223.650 847.600 223.930 850.000 ;
    END
  END la_output[23]
  PIN la_output[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 232.850 847.600 233.130 850.000 ;
    END
  END la_output[24]
  PIN la_output[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 242.050 847.600 242.330 850.000 ;
    END
  END la_output[25]
  PIN la_output[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 251.710 847.600 251.990 850.000 ;
    END
  END la_output[26]
  PIN la_output[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 260.910 847.600 261.190 850.000 ;
    END
  END la_output[27]
  PIN la_output[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 270.570 847.600 270.850 850.000 ;
    END
  END la_output[28]
  PIN la_output[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 279.770 847.600 280.050 850.000 ;
    END
  END la_output[29]
  PIN la_output[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 26.310 847.600 26.590 850.000 ;
    END
  END la_output[2]
  PIN la_output[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 288.970 847.600 289.250 850.000 ;
    END
  END la_output[30]
  PIN la_output[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 298.630 847.600 298.910 850.000 ;
    END
  END la_output[31]
  PIN la_output[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 307.830 847.600 308.110 850.000 ;
    END
  END la_output[32]
  PIN la_output[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 317.490 847.600 317.770 850.000 ;
    END
  END la_output[33]
  PIN la_output[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 326.690 847.600 326.970 850.000 ;
    END
  END la_output[34]
  PIN la_output[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 335.890 847.600 336.170 850.000 ;
    END
  END la_output[35]
  PIN la_output[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 345.550 847.600 345.830 850.000 ;
    END
  END la_output[36]
  PIN la_output[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 354.750 847.600 355.030 850.000 ;
    END
  END la_output[37]
  PIN la_output[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 364.410 847.600 364.690 850.000 ;
    END
  END la_output[38]
  PIN la_output[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 373.610 847.600 373.890 850.000 ;
    END
  END la_output[39]
  PIN la_output[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 35.510 847.600 35.790 850.000 ;
    END
  END la_output[3]
  PIN la_output[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 383.270 847.600 383.550 850.000 ;
    END
  END la_output[40]
  PIN la_output[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 392.470 847.600 392.750 850.000 ;
    END
  END la_output[41]
  PIN la_output[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 401.670 847.600 401.950 850.000 ;
    END
  END la_output[42]
  PIN la_output[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 411.330 847.600 411.610 850.000 ;
    END
  END la_output[43]
  PIN la_output[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 420.530 847.600 420.810 850.000 ;
    END
  END la_output[44]
  PIN la_output[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 430.190 847.600 430.470 850.000 ;
    END
  END la_output[45]
  PIN la_output[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 439.390 847.600 439.670 850.000 ;
    END
  END la_output[46]
  PIN la_output[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 448.590 847.600 448.870 850.000 ;
    END
  END la_output[47]
  PIN la_output[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 458.250 847.600 458.530 850.000 ;
    END
  END la_output[48]
  PIN la_output[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 467.450 847.600 467.730 850.000 ;
    END
  END la_output[49]
  PIN la_output[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 45.170 847.600 45.450 850.000 ;
    END
  END la_output[4]
  PIN la_output[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 477.110 847.600 477.390 850.000 ;
    END
  END la_output[50]
  PIN la_output[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 486.310 847.600 486.590 850.000 ;
    END
  END la_output[51]
  PIN la_output[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 495.510 847.600 495.790 850.000 ;
    END
  END la_output[52]
  PIN la_output[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 505.170 847.600 505.450 850.000 ;
    END
  END la_output[53]
  PIN la_output[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 514.370 847.600 514.650 850.000 ;
    END
  END la_output[54]
  PIN la_output[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 524.030 847.600 524.310 850.000 ;
    END
  END la_output[55]
  PIN la_output[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 533.230 847.600 533.510 850.000 ;
    END
  END la_output[56]
  PIN la_output[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 542.890 847.600 543.170 850.000 ;
    END
  END la_output[57]
  PIN la_output[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 552.090 847.600 552.370 850.000 ;
    END
  END la_output[58]
  PIN la_output[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 561.290 847.600 561.570 850.000 ;
    END
  END la_output[59]
  PIN la_output[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 54.370 847.600 54.650 850.000 ;
    END
  END la_output[5]
  PIN la_output[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 570.950 847.600 571.230 850.000 ;
    END
  END la_output[60]
  PIN la_output[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 580.150 847.600 580.430 850.000 ;
    END
  END la_output[61]
  PIN la_output[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 589.810 847.600 590.090 850.000 ;
    END
  END la_output[62]
  PIN la_output[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 599.010 847.600 599.290 850.000 ;
    END
  END la_output[63]
  PIN la_output[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 608.210 847.600 608.490 850.000 ;
    END
  END la_output[64]
  PIN la_output[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 617.870 847.600 618.150 850.000 ;
    END
  END la_output[65]
  PIN la_output[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 627.070 847.600 627.350 850.000 ;
    END
  END la_output[66]
  PIN la_output[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 636.730 847.600 637.010 850.000 ;
    END
  END la_output[67]
  PIN la_output[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 645.930 847.600 646.210 850.000 ;
    END
  END la_output[68]
  PIN la_output[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 655.130 847.600 655.410 850.000 ;
    END
  END la_output[69]
  PIN la_output[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 64.030 847.600 64.310 850.000 ;
    END
  END la_output[6]
  PIN la_output[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 664.790 847.600 665.070 850.000 ;
    END
  END la_output[70]
  PIN la_output[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 673.990 847.600 674.270 850.000 ;
    END
  END la_output[71]
  PIN la_output[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 683.650 847.600 683.930 850.000 ;
    END
  END la_output[72]
  PIN la_output[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 692.850 847.600 693.130 850.000 ;
    END
  END la_output[73]
  PIN la_output[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 702.050 847.600 702.330 850.000 ;
    END
  END la_output[74]
  PIN la_output[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 711.710 847.600 711.990 850.000 ;
    END
  END la_output[75]
  PIN la_output[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 720.910 847.600 721.190 850.000 ;
    END
  END la_output[76]
  PIN la_output[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 730.570 847.600 730.850 850.000 ;
    END
  END la_output[77]
  PIN la_output[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 739.770 847.600 740.050 850.000 ;
    END
  END la_output[78]
  PIN la_output[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 749.430 847.600 749.710 850.000 ;
    END
  END la_output[79]
  PIN la_output[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.230 847.600 73.510 850.000 ;
    END
  END la_output[7]
  PIN la_output[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 758.630 847.600 758.910 850.000 ;
    END
  END la_output[80]
  PIN la_output[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 767.830 847.600 768.110 850.000 ;
    END
  END la_output[81]
  PIN la_output[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 777.490 847.600 777.770 850.000 ;
    END
  END la_output[82]
  PIN la_output[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 786.690 847.600 786.970 850.000 ;
    END
  END la_output[83]
  PIN la_output[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 796.350 847.600 796.630 850.000 ;
    END
  END la_output[84]
  PIN la_output[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 805.550 847.600 805.830 850.000 ;
    END
  END la_output[85]
  PIN la_output[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 814.750 847.600 815.030 850.000 ;
    END
  END la_output[86]
  PIN la_output[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 824.410 847.600 824.690 850.000 ;
    END
  END la_output[87]
  PIN la_output[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 833.610 847.600 833.890 850.000 ;
    END
  END la_output[88]
  PIN la_output[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 843.270 847.600 843.550 850.000 ;
    END
  END la_output[89]
  PIN la_output[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.430 847.600 82.710 850.000 ;
    END
  END la_output[8]
  PIN la_output[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 852.470 847.600 852.750 850.000 ;
    END
  END la_output[90]
  PIN la_output[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 861.670 847.600 861.950 850.000 ;
    END
  END la_output[91]
  PIN la_output[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 871.330 847.600 871.610 850.000 ;
    END
  END la_output[92]
  PIN la_output[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 880.530 847.600 880.810 850.000 ;
    END
  END la_output[93]
  PIN la_output[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 890.190 847.600 890.470 850.000 ;
    END
  END la_output[94]
  PIN la_output[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 899.390 847.600 899.670 850.000 ;
    END
  END la_output[95]
  PIN la_output[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 909.050 847.600 909.330 850.000 ;
    END
  END la_output[96]
  PIN la_output[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 918.250 847.600 918.530 850.000 ;
    END
  END la_output[97]
  PIN la_output[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 927.450 847.600 927.730 850.000 ;
    END
  END la_output[98]
  PIN la_output[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 937.110 847.600 937.390 850.000 ;
    END
  END la_output[99]
  PIN la_output[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.090 847.600 92.370 850.000 ;
    END
  END la_output[9]
  PIN mask_rev[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.160 2.400 737.760 ;
    END
  END mask_rev[0]
  PIN mask_rev[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 772.520 2.400 773.120 ;
    END
  END mask_rev[10]
  PIN mask_rev[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 776.600 2.400 777.200 ;
    END
  END mask_rev[11]
  PIN mask_rev[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 780.000 2.400 780.600 ;
    END
  END mask_rev[12]
  PIN mask_rev[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 783.400 2.400 784.000 ;
    END
  END mask_rev[13]
  PIN mask_rev[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 786.800 2.400 787.400 ;
    END
  END mask_rev[14]
  PIN mask_rev[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 790.880 2.400 791.480 ;
    END
  END mask_rev[15]
  PIN mask_rev[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 794.280 2.400 794.880 ;
    END
  END mask_rev[16]
  PIN mask_rev[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 797.680 2.400 798.280 ;
    END
  END mask_rev[17]
  PIN mask_rev[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 801.080 2.400 801.680 ;
    END
  END mask_rev[18]
  PIN mask_rev[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.160 2.400 805.760 ;
    END
  END mask_rev[19]
  PIN mask_rev[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 740.560 2.400 741.160 ;
    END
  END mask_rev[1]
  PIN mask_rev[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 808.560 2.400 809.160 ;
    END
  END mask_rev[20]
  PIN mask_rev[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 811.960 2.400 812.560 ;
    END
  END mask_rev[21]
  PIN mask_rev[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 815.360 2.400 815.960 ;
    END
  END mask_rev[22]
  PIN mask_rev[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 818.760 2.400 819.360 ;
    END
  END mask_rev[23]
  PIN mask_rev[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.840 2.400 823.440 ;
    END
  END mask_rev[24]
  PIN mask_rev[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 826.240 2.400 826.840 ;
    END
  END mask_rev[25]
  PIN mask_rev[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.640 2.400 830.240 ;
    END
  END mask_rev[26]
  PIN mask_rev[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 833.040 2.400 833.640 ;
    END
  END mask_rev[27]
  PIN mask_rev[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 837.120 2.400 837.720 ;
    END
  END mask_rev[28]
  PIN mask_rev[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 840.520 2.400 841.120 ;
    END
  END mask_rev[29]
  PIN mask_rev[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 744.640 2.400 745.240 ;
    END
  END mask_rev[2]
  PIN mask_rev[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.920 2.400 844.520 ;
    END
  END mask_rev[30]
  PIN mask_rev[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 847.320 2.400 847.920 ;
    END
  END mask_rev[31]
  PIN mask_rev[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.040 2.400 748.640 ;
    END
  END mask_rev[3]
  PIN mask_rev[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 751.440 2.400 752.040 ;
    END
  END mask_rev[4]
  PIN mask_rev[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 2.400 755.440 ;
    END
  END mask_rev[5]
  PIN mask_rev[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.920 2.400 759.520 ;
    END
  END mask_rev[6]
  PIN mask_rev[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 762.320 2.400 762.920 ;
    END
  END mask_rev[7]
  PIN mask_rev[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.720 2.400 766.320 ;
    END
  END mask_rev[8]
  PIN mask_rev[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 769.120 2.400 769.720 ;
    END
  END mask_rev[9]
  PIN mgmt_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1202.990 847.600 1203.270 850.000 ;
    END
  END mgmt_addr[0]
  PIN mgmt_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1227.830 847.600 1228.110 850.000 ;
    END
  END mgmt_addr[1]
  PIN mgmt_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1253.130 847.600 1253.410 850.000 ;
    END
  END mgmt_addr[2]
  PIN mgmt_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1271.990 847.600 1272.270 850.000 ;
    END
  END mgmt_addr[3]
  PIN mgmt_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1290.850 847.600 1291.130 850.000 ;
    END
  END mgmt_addr[4]
  PIN mgmt_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1309.250 847.600 1309.530 850.000 ;
    END
  END mgmt_addr[5]
  PIN mgmt_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1328.110 847.600 1328.390 850.000 ;
    END
  END mgmt_addr[6]
  PIN mgmt_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1346.970 847.600 1347.250 850.000 ;
    END
  END mgmt_addr[7]
  PIN mgmt_ena[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1206.210 847.600 1206.490 850.000 ;
    END
  END mgmt_ena[0]
  PIN mgmt_ena[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1231.050 847.600 1231.330 850.000 ;
    END
  END mgmt_ena[1]
  PIN mgmt_in_data[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1209.430 847.600 1209.710 850.000 ;
    END
  END mgmt_in_data[0]
  PIN mgmt_in_data[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1390.670 847.600 1390.950 850.000 ;
    END
  END mgmt_in_data[10]
  PIN mgmt_in_data[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1403.090 847.600 1403.370 850.000 ;
    END
  END mgmt_in_data[11]
  PIN mgmt_in_data[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1415.970 847.600 1416.250 850.000 ;
    END
  END mgmt_in_data[12]
  PIN mgmt_in_data[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1428.390 847.600 1428.670 850.000 ;
    END
  END mgmt_in_data[13]
  PIN mgmt_in_data[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1440.810 847.600 1441.090 850.000 ;
    END
  END mgmt_in_data[14]
  PIN mgmt_in_data[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1453.230 847.600 1453.510 850.000 ;
    END
  END mgmt_in_data[15]
  PIN mgmt_in_data[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1466.110 847.600 1466.390 850.000 ;
    END
  END mgmt_in_data[16]
  PIN mgmt_in_data[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1478.530 847.600 1478.810 850.000 ;
    END
  END mgmt_in_data[17]
  PIN mgmt_in_data[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1490.950 847.600 1491.230 850.000 ;
    END
  END mgmt_in_data[18]
  PIN mgmt_in_data[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1503.370 847.600 1503.650 850.000 ;
    END
  END mgmt_in_data[19]
  PIN mgmt_in_data[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1234.270 847.600 1234.550 850.000 ;
    END
  END mgmt_in_data[1]
  PIN mgmt_in_data[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1515.790 847.600 1516.070 850.000 ;
    END
  END mgmt_in_data[20]
  PIN mgmt_in_data[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1528.670 847.600 1528.950 850.000 ;
    END
  END mgmt_in_data[21]
  PIN mgmt_in_data[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1541.090 847.600 1541.370 850.000 ;
    END
  END mgmt_in_data[22]
  PIN mgmt_in_data[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1553.510 847.600 1553.790 850.000 ;
    END
  END mgmt_in_data[23]
  PIN mgmt_in_data[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1565.930 847.600 1566.210 850.000 ;
    END
  END mgmt_in_data[24]
  PIN mgmt_in_data[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1578.350 847.600 1578.630 850.000 ;
    END
  END mgmt_in_data[25]
  PIN mgmt_in_data[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1591.230 847.600 1591.510 850.000 ;
    END
  END mgmt_in_data[26]
  PIN mgmt_in_data[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1603.650 847.600 1603.930 850.000 ;
    END
  END mgmt_in_data[27]
  PIN mgmt_in_data[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1616.070 847.600 1616.350 850.000 ;
    END
  END mgmt_in_data[28]
  PIN mgmt_in_data[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1628.490 847.600 1628.770 850.000 ;
    END
  END mgmt_in_data[29]
  PIN mgmt_in_data[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1256.350 847.600 1256.630 850.000 ;
    END
  END mgmt_in_data[2]
  PIN mgmt_in_data[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1641.370 847.600 1641.650 850.000 ;
    END
  END mgmt_in_data[30]
  PIN mgmt_in_data[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1653.790 847.600 1654.070 850.000 ;
    END
  END mgmt_in_data[31]
  PIN mgmt_in_data[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1666.210 847.600 1666.490 850.000 ;
    END
  END mgmt_in_data[32]
  PIN mgmt_in_data[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1675.410 847.600 1675.690 850.000 ;
    END
  END mgmt_in_data[33]
  PIN mgmt_in_data[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1685.070 847.600 1685.350 850.000 ;
    END
  END mgmt_in_data[34]
  PIN mgmt_in_data[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1694.270 847.600 1694.550 850.000 ;
    END
  END mgmt_in_data[35]
  PIN mgmt_in_data[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1703.930 847.600 1704.210 850.000 ;
    END
  END mgmt_in_data[36]
  PIN mgmt_in_data[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1713.130 847.600 1713.410 850.000 ;
    END
  END mgmt_in_data[37]
  PIN mgmt_in_data[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1275.210 847.600 1275.490 850.000 ;
    END
  END mgmt_in_data[3]
  PIN mgmt_in_data[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1293.610 847.600 1293.890 850.000 ;
    END
  END mgmt_in_data[4]
  PIN mgmt_in_data[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1312.470 847.600 1312.750 850.000 ;
    END
  END mgmt_in_data[5]
  PIN mgmt_in_data[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1331.330 847.600 1331.610 850.000 ;
    END
  END mgmt_in_data[6]
  PIN mgmt_in_data[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1350.190 847.600 1350.470 850.000 ;
    END
  END mgmt_in_data[7]
  PIN mgmt_in_data[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1365.830 847.600 1366.110 850.000 ;
    END
  END mgmt_in_data[8]
  PIN mgmt_in_data[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1378.250 847.600 1378.530 850.000 ;
    END
  END mgmt_in_data[9]
  PIN mgmt_out_data[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1212.190 847.600 1212.470 850.000 ;
    END
  END mgmt_out_data[0]
  PIN mgmt_out_data[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1393.890 847.600 1394.170 850.000 ;
    END
  END mgmt_out_data[10]
  PIN mgmt_out_data[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1406.310 847.600 1406.590 850.000 ;
    END
  END mgmt_out_data[11]
  PIN mgmt_out_data[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1418.730 847.600 1419.010 850.000 ;
    END
  END mgmt_out_data[12]
  PIN mgmt_out_data[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1431.610 847.600 1431.890 850.000 ;
    END
  END mgmt_out_data[13]
  PIN mgmt_out_data[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1444.030 847.600 1444.310 850.000 ;
    END
  END mgmt_out_data[14]
  PIN mgmt_out_data[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1456.450 847.600 1456.730 850.000 ;
    END
  END mgmt_out_data[15]
  PIN mgmt_out_data[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1468.870 847.600 1469.150 850.000 ;
    END
  END mgmt_out_data[16]
  PIN mgmt_out_data[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1481.750 847.600 1482.030 850.000 ;
    END
  END mgmt_out_data[17]
  PIN mgmt_out_data[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1494.170 847.600 1494.450 850.000 ;
    END
  END mgmt_out_data[18]
  PIN mgmt_out_data[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1506.590 847.600 1506.870 850.000 ;
    END
  END mgmt_out_data[19]
  PIN mgmt_out_data[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1237.490 847.600 1237.770 850.000 ;
    END
  END mgmt_out_data[1]
  PIN mgmt_out_data[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1519.010 847.600 1519.290 850.000 ;
    END
  END mgmt_out_data[20]
  PIN mgmt_out_data[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1531.430 847.600 1531.710 850.000 ;
    END
  END mgmt_out_data[21]
  PIN mgmt_out_data[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1544.310 847.600 1544.590 850.000 ;
    END
  END mgmt_out_data[22]
  PIN mgmt_out_data[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1556.730 847.600 1557.010 850.000 ;
    END
  END mgmt_out_data[23]
  PIN mgmt_out_data[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1569.150 847.600 1569.430 850.000 ;
    END
  END mgmt_out_data[24]
  PIN mgmt_out_data[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1581.570 847.600 1581.850 850.000 ;
    END
  END mgmt_out_data[25]
  PIN mgmt_out_data[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1593.990 847.600 1594.270 850.000 ;
    END
  END mgmt_out_data[26]
  PIN mgmt_out_data[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1606.870 847.600 1607.150 850.000 ;
    END
  END mgmt_out_data[27]
  PIN mgmt_out_data[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1619.290 847.600 1619.570 850.000 ;
    END
  END mgmt_out_data[28]
  PIN mgmt_out_data[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1631.710 847.600 1631.990 850.000 ;
    END
  END mgmt_out_data[29]
  PIN mgmt_out_data[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1259.570 847.600 1259.850 850.000 ;
    END
  END mgmt_out_data[2]
  PIN mgmt_out_data[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1644.130 847.600 1644.410 850.000 ;
    END
  END mgmt_out_data[30]
  PIN mgmt_out_data[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1657.010 847.600 1657.290 850.000 ;
    END
  END mgmt_out_data[31]
  PIN mgmt_out_data[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1669.430 847.600 1669.710 850.000 ;
    END
  END mgmt_out_data[32]
  PIN mgmt_out_data[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1678.630 847.600 1678.910 850.000 ;
    END
  END mgmt_out_data[33]
  PIN mgmt_out_data[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1688.290 847.600 1688.570 850.000 ;
    END
  END mgmt_out_data[34]
  PIN mgmt_out_data[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1697.490 847.600 1697.770 850.000 ;
    END
  END mgmt_out_data[35]
  PIN mgmt_out_data[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1706.690 847.600 1706.970 850.000 ;
    END
  END mgmt_out_data[36]
  PIN mgmt_out_data[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1716.350 847.600 1716.630 850.000 ;
    END
  END mgmt_out_data[37]
  PIN mgmt_out_data[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1277.970 847.600 1278.250 850.000 ;
    END
  END mgmt_out_data[3]
  PIN mgmt_out_data[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1296.830 847.600 1297.110 850.000 ;
    END
  END mgmt_out_data[4]
  PIN mgmt_out_data[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1315.690 847.600 1315.970 850.000 ;
    END
  END mgmt_out_data[5]
  PIN mgmt_out_data[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1334.550 847.600 1334.830 850.000 ;
    END
  END mgmt_out_data[6]
  PIN mgmt_out_data[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1353.410 847.600 1353.690 850.000 ;
    END
  END mgmt_out_data[7]
  PIN mgmt_out_data[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1369.050 847.600 1369.330 850.000 ;
    END
  END mgmt_out_data[8]
  PIN mgmt_out_data[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1381.470 847.600 1381.750 850.000 ;
    END
  END mgmt_out_data[9]
  PIN mgmt_rdata[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1215.410 847.600 1215.690 850.000 ;
    END
  END mgmt_rdata[0]
  PIN mgmt_rdata[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1397.110 847.600 1397.390 850.000 ;
    END
  END mgmt_rdata[10]
  PIN mgmt_rdata[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1409.530 847.600 1409.810 850.000 ;
    END
  END mgmt_rdata[11]
  PIN mgmt_rdata[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1421.950 847.600 1422.230 850.000 ;
    END
  END mgmt_rdata[12]
  PIN mgmt_rdata[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1434.830 847.600 1435.110 850.000 ;
    END
  END mgmt_rdata[13]
  PIN mgmt_rdata[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1447.250 847.600 1447.530 850.000 ;
    END
  END mgmt_rdata[14]
  PIN mgmt_rdata[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1459.670 847.600 1459.950 850.000 ;
    END
  END mgmt_rdata[15]
  PIN mgmt_rdata[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1472.090 847.600 1472.370 850.000 ;
    END
  END mgmt_rdata[16]
  PIN mgmt_rdata[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1484.510 847.600 1484.790 850.000 ;
    END
  END mgmt_rdata[17]
  PIN mgmt_rdata[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1497.390 847.600 1497.670 850.000 ;
    END
  END mgmt_rdata[18]
  PIN mgmt_rdata[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1509.810 847.600 1510.090 850.000 ;
    END
  END mgmt_rdata[19]
  PIN mgmt_rdata[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1240.710 847.600 1240.990 850.000 ;
    END
  END mgmt_rdata[1]
  PIN mgmt_rdata[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1522.230 847.600 1522.510 850.000 ;
    END
  END mgmt_rdata[20]
  PIN mgmt_rdata[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1534.650 847.600 1534.930 850.000 ;
    END
  END mgmt_rdata[21]
  PIN mgmt_rdata[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1547.070 847.600 1547.350 850.000 ;
    END
  END mgmt_rdata[22]
  PIN mgmt_rdata[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1559.950 847.600 1560.230 850.000 ;
    END
  END mgmt_rdata[23]
  PIN mgmt_rdata[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1572.370 847.600 1572.650 850.000 ;
    END
  END mgmt_rdata[24]
  PIN mgmt_rdata[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1584.790 847.600 1585.070 850.000 ;
    END
  END mgmt_rdata[25]
  PIN mgmt_rdata[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1597.210 847.600 1597.490 850.000 ;
    END
  END mgmt_rdata[26]
  PIN mgmt_rdata[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1609.630 847.600 1609.910 850.000 ;
    END
  END mgmt_rdata[27]
  PIN mgmt_rdata[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1622.510 847.600 1622.790 850.000 ;
    END
  END mgmt_rdata[28]
  PIN mgmt_rdata[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1634.930 847.600 1635.210 850.000 ;
    END
  END mgmt_rdata[29]
  PIN mgmt_rdata[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1262.330 847.600 1262.610 850.000 ;
    END
  END mgmt_rdata[2]
  PIN mgmt_rdata[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1647.350 847.600 1647.630 850.000 ;
    END
  END mgmt_rdata[30]
  PIN mgmt_rdata[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1659.770 847.600 1660.050 850.000 ;
    END
  END mgmt_rdata[31]
  PIN mgmt_rdata[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1672.650 847.600 1672.930 850.000 ;
    END
  END mgmt_rdata[32]
  PIN mgmt_rdata[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1681.850 847.600 1682.130 850.000 ;
    END
  END mgmt_rdata[33]
  PIN mgmt_rdata[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1691.050 847.600 1691.330 850.000 ;
    END
  END mgmt_rdata[34]
  PIN mgmt_rdata[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1700.710 847.600 1700.990 850.000 ;
    END
  END mgmt_rdata[35]
  PIN mgmt_rdata[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1709.910 847.600 1710.190 850.000 ;
    END
  END mgmt_rdata[36]
  PIN mgmt_rdata[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1719.570 847.600 1719.850 850.000 ;
    END
  END mgmt_rdata[37]
  PIN mgmt_rdata[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1722.330 847.600 1722.610 850.000 ;
    END
  END mgmt_rdata[38]
  PIN mgmt_rdata[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1725.550 847.600 1725.830 850.000 ;
    END
  END mgmt_rdata[39]
  PIN mgmt_rdata[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1281.190 847.600 1281.470 850.000 ;
    END
  END mgmt_rdata[3]
  PIN mgmt_rdata[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1728.770 847.600 1729.050 850.000 ;
    END
  END mgmt_rdata[40]
  PIN mgmt_rdata[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1731.990 847.600 1732.270 850.000 ;
    END
  END mgmt_rdata[41]
  PIN mgmt_rdata[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1735.210 847.600 1735.490 850.000 ;
    END
  END mgmt_rdata[42]
  PIN mgmt_rdata[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1737.970 847.600 1738.250 850.000 ;
    END
  END mgmt_rdata[43]
  PIN mgmt_rdata[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1741.190 847.600 1741.470 850.000 ;
    END
  END mgmt_rdata[44]
  PIN mgmt_rdata[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1744.410 847.600 1744.690 850.000 ;
    END
  END mgmt_rdata[45]
  PIN mgmt_rdata[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1747.630 847.600 1747.910 850.000 ;
    END
  END mgmt_rdata[46]
  PIN mgmt_rdata[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1750.850 847.600 1751.130 850.000 ;
    END
  END mgmt_rdata[47]
  PIN mgmt_rdata[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1753.610 847.600 1753.890 850.000 ;
    END
  END mgmt_rdata[48]
  PIN mgmt_rdata[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1756.830 847.600 1757.110 850.000 ;
    END
  END mgmt_rdata[49]
  PIN mgmt_rdata[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1300.050 847.600 1300.330 850.000 ;
    END
  END mgmt_rdata[4]
  PIN mgmt_rdata[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1760.050 847.600 1760.330 850.000 ;
    END
  END mgmt_rdata[50]
  PIN mgmt_rdata[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1763.270 847.600 1763.550 850.000 ;
    END
  END mgmt_rdata[51]
  PIN mgmt_rdata[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1766.490 847.600 1766.770 850.000 ;
    END
  END mgmt_rdata[52]
  PIN mgmt_rdata[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1769.250 847.600 1769.530 850.000 ;
    END
  END mgmt_rdata[53]
  PIN mgmt_rdata[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1772.470 847.600 1772.750 850.000 ;
    END
  END mgmt_rdata[54]
  PIN mgmt_rdata[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1775.690 847.600 1775.970 850.000 ;
    END
  END mgmt_rdata[55]
  PIN mgmt_rdata[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1778.910 847.600 1779.190 850.000 ;
    END
  END mgmt_rdata[56]
  PIN mgmt_rdata[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1782.130 847.600 1782.410 850.000 ;
    END
  END mgmt_rdata[57]
  PIN mgmt_rdata[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1784.890 847.600 1785.170 850.000 ;
    END
  END mgmt_rdata[58]
  PIN mgmt_rdata[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1788.110 847.600 1788.390 850.000 ;
    END
  END mgmt_rdata[59]
  PIN mgmt_rdata[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1318.910 847.600 1319.190 850.000 ;
    END
  END mgmt_rdata[5]
  PIN mgmt_rdata[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1791.330 847.600 1791.610 850.000 ;
    END
  END mgmt_rdata[60]
  PIN mgmt_rdata[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1794.550 847.600 1794.830 850.000 ;
    END
  END mgmt_rdata[61]
  PIN mgmt_rdata[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1797.770 847.600 1798.050 850.000 ;
    END
  END mgmt_rdata[62]
  PIN mgmt_rdata[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1800.990 847.600 1801.270 850.000 ;
    END
  END mgmt_rdata[63]
  PIN mgmt_rdata[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1337.770 847.600 1338.050 850.000 ;
    END
  END mgmt_rdata[6]
  PIN mgmt_rdata[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1356.170 847.600 1356.450 850.000 ;
    END
  END mgmt_rdata[7]
  PIN mgmt_rdata[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1371.810 847.600 1372.090 850.000 ;
    END
  END mgmt_rdata[8]
  PIN mgmt_rdata[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1384.690 847.600 1384.970 850.000 ;
    END
  END mgmt_rdata[9]
  PIN mgmt_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1218.630 847.600 1218.910 850.000 ;
    END
  END mgmt_wdata[0]
  PIN mgmt_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1400.330 847.600 1400.610 850.000 ;
    END
  END mgmt_wdata[10]
  PIN mgmt_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1412.750 847.600 1413.030 850.000 ;
    END
  END mgmt_wdata[11]
  PIN mgmt_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1425.170 847.600 1425.450 850.000 ;
    END
  END mgmt_wdata[12]
  PIN mgmt_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1437.590 847.600 1437.870 850.000 ;
    END
  END mgmt_wdata[13]
  PIN mgmt_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1450.470 847.600 1450.750 850.000 ;
    END
  END mgmt_wdata[14]
  PIN mgmt_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1462.890 847.600 1463.170 850.000 ;
    END
  END mgmt_wdata[15]
  PIN mgmt_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1475.310 847.600 1475.590 850.000 ;
    END
  END mgmt_wdata[16]
  PIN mgmt_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1487.730 847.600 1488.010 850.000 ;
    END
  END mgmt_wdata[17]
  PIN mgmt_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1500.150 847.600 1500.430 850.000 ;
    END
  END mgmt_wdata[18]
  PIN mgmt_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1513.030 847.600 1513.310 850.000 ;
    END
  END mgmt_wdata[19]
  PIN mgmt_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1243.470 847.600 1243.750 850.000 ;
    END
  END mgmt_wdata[1]
  PIN mgmt_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1525.450 847.600 1525.730 850.000 ;
    END
  END mgmt_wdata[20]
  PIN mgmt_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1537.870 847.600 1538.150 850.000 ;
    END
  END mgmt_wdata[21]
  PIN mgmt_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1550.290 847.600 1550.570 850.000 ;
    END
  END mgmt_wdata[22]
  PIN mgmt_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1562.710 847.600 1562.990 850.000 ;
    END
  END mgmt_wdata[23]
  PIN mgmt_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1575.590 847.600 1575.870 850.000 ;
    END
  END mgmt_wdata[24]
  PIN mgmt_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1588.010 847.600 1588.290 850.000 ;
    END
  END mgmt_wdata[25]
  PIN mgmt_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1600.430 847.600 1600.710 850.000 ;
    END
  END mgmt_wdata[26]
  PIN mgmt_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1612.850 847.600 1613.130 850.000 ;
    END
  END mgmt_wdata[27]
  PIN mgmt_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1625.730 847.600 1626.010 850.000 ;
    END
  END mgmt_wdata[28]
  PIN mgmt_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1638.150 847.600 1638.430 850.000 ;
    END
  END mgmt_wdata[29]
  PIN mgmt_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1265.550 847.600 1265.830 850.000 ;
    END
  END mgmt_wdata[2]
  PIN mgmt_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1650.570 847.600 1650.850 850.000 ;
    END
  END mgmt_wdata[30]
  PIN mgmt_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1662.990 847.600 1663.270 850.000 ;
    END
  END mgmt_wdata[31]
  PIN mgmt_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1284.410 847.600 1284.690 850.000 ;
    END
  END mgmt_wdata[3]
  PIN mgmt_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1303.270 847.600 1303.550 850.000 ;
    END
  END mgmt_wdata[4]
  PIN mgmt_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1322.130 847.600 1322.410 850.000 ;
    END
  END mgmt_wdata[5]
  PIN mgmt_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1340.530 847.600 1340.810 850.000 ;
    END
  END mgmt_wdata[6]
  PIN mgmt_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1359.390 847.600 1359.670 850.000 ;
    END
  END mgmt_wdata[7]
  PIN mgmt_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1375.030 847.600 1375.310 850.000 ;
    END
  END mgmt_wdata[8]
  PIN mgmt_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1387.450 847.600 1387.730 850.000 ;
    END
  END mgmt_wdata[9]
  PIN mgmt_wen[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1221.850 847.600 1222.130 850.000 ;
    END
  END mgmt_wen[0]
  PIN mgmt_wen[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1246.690 847.600 1246.970 850.000 ;
    END
  END mgmt_wen[1]
  PIN mgmt_wen_mask[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1225.070 847.600 1225.350 850.000 ;
    END
  END mgmt_wen_mask[0]
  PIN mgmt_wen_mask[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1249.910 847.600 1250.190 850.000 ;
    END
  END mgmt_wen_mask[1]
  PIN mgmt_wen_mask[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1268.770 847.600 1269.050 850.000 ;
    END
  END mgmt_wen_mask[2]
  PIN mgmt_wen_mask[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1287.630 847.600 1287.910 850.000 ;
    END
  END mgmt_wen_mask[3]
  PIN mgmt_wen_mask[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1306.490 847.600 1306.770 850.000 ;
    END
  END mgmt_wen_mask[4]
  PIN mgmt_wen_mask[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1324.890 847.600 1325.170 850.000 ;
    END
  END mgmt_wen_mask[5]
  PIN mgmt_wen_mask[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1343.750 847.600 1344.030 850.000 ;
    END
  END mgmt_wen_mask[6]
  PIN mgmt_wen_mask[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1362.610 847.600 1362.890 850.000 ;
    END
  END mgmt_wen_mask[7]
  PIN mprj2_vcc_pwrgood
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1803.750 847.600 1804.030 850.000 ;
    END
  END mprj2_vcc_pwrgood
  PIN mprj2_vdd_pwrgood
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1806.970 847.600 1807.250 850.000 ;
    END
  END mprj2_vdd_pwrgood
  PIN mprj_ack_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1810.190 847.600 1810.470 850.000 ;
    END
  END mprj_ack_i
  PIN mprj_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1838.250 847.600 1838.530 850.000 ;
    END
  END mprj_adr_o[0]
  PIN mprj_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1944.510 847.600 1944.790 850.000 ;
    END
  END mprj_adr_o[10]
  PIN mprj_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1954.170 847.600 1954.450 850.000 ;
    END
  END mprj_adr_o[11]
  PIN mprj_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1963.370 847.600 1963.650 850.000 ;
    END
  END mprj_adr_o[12]
  PIN mprj_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1973.030 847.600 1973.310 850.000 ;
    END
  END mprj_adr_o[13]
  PIN mprj_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1982.230 847.600 1982.510 850.000 ;
    END
  END mprj_adr_o[14]
  PIN mprj_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1991.890 847.600 1992.170 850.000 ;
    END
  END mprj_adr_o[15]
  PIN mprj_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2001.090 847.600 2001.370 850.000 ;
    END
  END mprj_adr_o[16]
  PIN mprj_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2010.290 847.600 2010.570 850.000 ;
    END
  END mprj_adr_o[17]
  PIN mprj_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2019.950 847.600 2020.230 850.000 ;
    END
  END mprj_adr_o[18]
  PIN mprj_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2029.150 847.600 2029.430 850.000 ;
    END
  END mprj_adr_o[19]
  PIN mprj_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1850.670 847.600 1850.950 850.000 ;
    END
  END mprj_adr_o[1]
  PIN mprj_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2038.810 847.600 2039.090 850.000 ;
    END
  END mprj_adr_o[20]
  PIN mprj_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2048.010 847.600 2048.290 850.000 ;
    END
  END mprj_adr_o[21]
  PIN mprj_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2057.210 847.600 2057.490 850.000 ;
    END
  END mprj_adr_o[22]
  PIN mprj_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2066.870 847.600 2067.150 850.000 ;
    END
  END mprj_adr_o[23]
  PIN mprj_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2076.070 847.600 2076.350 850.000 ;
    END
  END mprj_adr_o[24]
  PIN mprj_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2085.730 847.600 2086.010 850.000 ;
    END
  END mprj_adr_o[25]
  PIN mprj_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2094.930 847.600 2095.210 850.000 ;
    END
  END mprj_adr_o[26]
  PIN mprj_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2104.130 847.600 2104.410 850.000 ;
    END
  END mprj_adr_o[27]
  PIN mprj_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2113.790 847.600 2114.070 850.000 ;
    END
  END mprj_adr_o[28]
  PIN mprj_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2122.990 847.600 2123.270 850.000 ;
    END
  END mprj_adr_o[29]
  PIN mprj_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1863.550 847.600 1863.830 850.000 ;
    END
  END mprj_adr_o[2]
  PIN mprj_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2132.650 847.600 2132.930 850.000 ;
    END
  END mprj_adr_o[30]
  PIN mprj_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2141.850 847.600 2142.130 850.000 ;
    END
  END mprj_adr_o[31]
  PIN mprj_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1875.970 847.600 1876.250 850.000 ;
    END
  END mprj_adr_o[3]
  PIN mprj_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1888.390 847.600 1888.670 850.000 ;
    END
  END mprj_adr_o[4]
  PIN mprj_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1897.590 847.600 1897.870 850.000 ;
    END
  END mprj_adr_o[5]
  PIN mprj_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1907.250 847.600 1907.530 850.000 ;
    END
  END mprj_adr_o[6]
  PIN mprj_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1916.450 847.600 1916.730 850.000 ;
    END
  END mprj_adr_o[7]
  PIN mprj_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1926.110 847.600 1926.390 850.000 ;
    END
  END mprj_adr_o[8]
  PIN mprj_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1935.310 847.600 1935.590 850.000 ;
    END
  END mprj_adr_o[9]
  PIN mprj_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1813.410 847.600 1813.690 850.000 ;
    END
  END mprj_cyc_o
  PIN mprj_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1841.470 847.600 1841.750 850.000 ;
    END
  END mprj_dat_i[0]
  PIN mprj_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1947.730 847.600 1948.010 850.000 ;
    END
  END mprj_dat_i[10]
  PIN mprj_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1957.390 847.600 1957.670 850.000 ;
    END
  END mprj_dat_i[11]
  PIN mprj_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1966.590 847.600 1966.870 850.000 ;
    END
  END mprj_dat_i[12]
  PIN mprj_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1976.250 847.600 1976.530 850.000 ;
    END
  END mprj_dat_i[13]
  PIN mprj_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1985.450 847.600 1985.730 850.000 ;
    END
  END mprj_dat_i[14]
  PIN mprj_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1994.650 847.600 1994.930 850.000 ;
    END
  END mprj_dat_i[15]
  PIN mprj_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2004.310 847.600 2004.590 850.000 ;
    END
  END mprj_dat_i[16]
  PIN mprj_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2013.510 847.600 2013.790 850.000 ;
    END
  END mprj_dat_i[17]
  PIN mprj_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2023.170 847.600 2023.450 850.000 ;
    END
  END mprj_dat_i[18]
  PIN mprj_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2032.370 847.600 2032.650 850.000 ;
    END
  END mprj_dat_i[19]
  PIN mprj_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1853.890 847.600 1854.170 850.000 ;
    END
  END mprj_dat_i[1]
  PIN mprj_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2041.570 847.600 2041.850 850.000 ;
    END
  END mprj_dat_i[20]
  PIN mprj_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2051.230 847.600 2051.510 850.000 ;
    END
  END mprj_dat_i[21]
  PIN mprj_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2060.430 847.600 2060.710 850.000 ;
    END
  END mprj_dat_i[22]
  PIN mprj_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2070.090 847.600 2070.370 850.000 ;
    END
  END mprj_dat_i[23]
  PIN mprj_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2079.290 847.600 2079.570 850.000 ;
    END
  END mprj_dat_i[24]
  PIN mprj_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2088.490 847.600 2088.770 850.000 ;
    END
  END mprj_dat_i[25]
  PIN mprj_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2098.150 847.600 2098.430 850.000 ;
    END
  END mprj_dat_i[26]
  PIN mprj_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2107.350 847.600 2107.630 850.000 ;
    END
  END mprj_dat_i[27]
  PIN mprj_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2117.010 847.600 2117.290 850.000 ;
    END
  END mprj_dat_i[28]
  PIN mprj_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2126.210 847.600 2126.490 850.000 ;
    END
  END mprj_dat_i[29]
  PIN mprj_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1866.310 847.600 1866.590 850.000 ;
    END
  END mprj_dat_i[2]
  PIN mprj_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2135.410 847.600 2135.690 850.000 ;
    END
  END mprj_dat_i[30]
  PIN mprj_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2145.070 847.600 2145.350 850.000 ;
    END
  END mprj_dat_i[31]
  PIN mprj_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1879.190 847.600 1879.470 850.000 ;
    END
  END mprj_dat_i[3]
  PIN mprj_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1891.610 847.600 1891.890 850.000 ;
    END
  END mprj_dat_i[4]
  PIN mprj_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1900.810 847.600 1901.090 850.000 ;
    END
  END mprj_dat_i[5]
  PIN mprj_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1910.470 847.600 1910.750 850.000 ;
    END
  END mprj_dat_i[6]
  PIN mprj_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1919.670 847.600 1919.950 850.000 ;
    END
  END mprj_dat_i[7]
  PIN mprj_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1928.870 847.600 1929.150 850.000 ;
    END
  END mprj_dat_i[8]
  PIN mprj_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1938.530 847.600 1938.810 850.000 ;
    END
  END mprj_dat_i[9]
  PIN mprj_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1844.690 847.600 1844.970 850.000 ;
    END
  END mprj_dat_o[0]
  PIN mprj_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1950.950 847.600 1951.230 850.000 ;
    END
  END mprj_dat_o[10]
  PIN mprj_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1960.150 847.600 1960.430 850.000 ;
    END
  END mprj_dat_o[11]
  PIN mprj_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1969.810 847.600 1970.090 850.000 ;
    END
  END mprj_dat_o[12]
  PIN mprj_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1979.010 847.600 1979.290 850.000 ;
    END
  END mprj_dat_o[13]
  PIN mprj_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1988.670 847.600 1988.950 850.000 ;
    END
  END mprj_dat_o[14]
  PIN mprj_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1997.870 847.600 1998.150 850.000 ;
    END
  END mprj_dat_o[15]
  PIN mprj_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2007.530 847.600 2007.810 850.000 ;
    END
  END mprj_dat_o[16]
  PIN mprj_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2016.730 847.600 2017.010 850.000 ;
    END
  END mprj_dat_o[17]
  PIN mprj_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2025.930 847.600 2026.210 850.000 ;
    END
  END mprj_dat_o[18]
  PIN mprj_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2035.590 847.600 2035.870 850.000 ;
    END
  END mprj_dat_o[19]
  PIN mprj_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1857.110 847.600 1857.390 850.000 ;
    END
  END mprj_dat_o[1]
  PIN mprj_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2044.790 847.600 2045.070 850.000 ;
    END
  END mprj_dat_o[20]
  PIN mprj_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2054.450 847.600 2054.730 850.000 ;
    END
  END mprj_dat_o[21]
  PIN mprj_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2063.650 847.600 2063.930 850.000 ;
    END
  END mprj_dat_o[22]
  PIN mprj_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2072.850 847.600 2073.130 850.000 ;
    END
  END mprj_dat_o[23]
  PIN mprj_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2082.510 847.600 2082.790 850.000 ;
    END
  END mprj_dat_o[24]
  PIN mprj_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2091.710 847.600 2091.990 850.000 ;
    END
  END mprj_dat_o[25]
  PIN mprj_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2101.370 847.600 2101.650 850.000 ;
    END
  END mprj_dat_o[26]
  PIN mprj_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2110.570 847.600 2110.850 850.000 ;
    END
  END mprj_dat_o[27]
  PIN mprj_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2119.770 847.600 2120.050 850.000 ;
    END
  END mprj_dat_o[28]
  PIN mprj_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2129.430 847.600 2129.710 850.000 ;
    END
  END mprj_dat_o[29]
  PIN mprj_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1869.530 847.600 1869.810 850.000 ;
    END
  END mprj_dat_o[2]
  PIN mprj_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2138.630 847.600 2138.910 850.000 ;
    END
  END mprj_dat_o[30]
  PIN mprj_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2148.290 847.600 2148.570 850.000 ;
    END
  END mprj_dat_o[31]
  PIN mprj_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1881.950 847.600 1882.230 850.000 ;
    END
  END mprj_dat_o[3]
  PIN mprj_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1894.830 847.600 1895.110 850.000 ;
    END
  END mprj_dat_o[4]
  PIN mprj_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1904.030 847.600 1904.310 850.000 ;
    END
  END mprj_dat_o[5]
  PIN mprj_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1913.230 847.600 1913.510 850.000 ;
    END
  END mprj_dat_o[6]
  PIN mprj_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1922.890 847.600 1923.170 850.000 ;
    END
  END mprj_dat_o[7]
  PIN mprj_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1932.090 847.600 1932.370 850.000 ;
    END
  END mprj_dat_o[8]
  PIN mprj_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1941.750 847.600 1942.030 850.000 ;
    END
  END mprj_dat_o[9]
  PIN mprj_io_loader_clock
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1816.630 847.600 1816.910 850.000 ;
    END
  END mprj_io_loader_clock
  PIN mprj_io_loader_data
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1819.390 847.600 1819.670 850.000 ;
    END
  END mprj_io_loader_data
  PIN mprj_io_loader_resetn
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1822.610 847.600 1822.890 850.000 ;
    END
  END mprj_io_loader_resetn
  PIN mprj_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1847.910 847.600 1848.190 850.000 ;
    END
  END mprj_sel_o[0]
  PIN mprj_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1860.330 847.600 1860.610 850.000 ;
    END
  END mprj_sel_o[1]
  PIN mprj_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1872.750 847.600 1873.030 850.000 ;
    END
  END mprj_sel_o[2]
  PIN mprj_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1885.170 847.600 1885.450 850.000 ;
    END
  END mprj_sel_o[3]
  PIN mprj_stb_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1825.830 847.600 1826.110 850.000 ;
    END
  END mprj_stb_o
  PIN mprj_vcc_pwrgood
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1829.050 847.600 1829.330 850.000 ;
    END
  END mprj_vcc_pwrgood
  PIN mprj_vdd_pwrgood
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1832.270 847.600 1832.550 850.000 ;
    END
  END mprj_vdd_pwrgood
  PIN mprj_we_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1835.030 847.600 1835.310 850.000 ;
    END
  END mprj_we_o
  PIN porb
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2147.600 810.600 2150.000 811.200 ;
    END
  END porb
  PIN pwr_ctrl_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2147.600 38.120 2150.000 38.720 ;
    END
  END pwr_ctrl_out[0]
  PIN pwr_ctrl_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2147.600 114.960 2150.000 115.560 ;
    END
  END pwr_ctrl_out[1]
  PIN pwr_ctrl_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2147.600 192.480 2150.000 193.080 ;
    END
  END pwr_ctrl_out[2]
  PIN pwr_ctrl_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2147.600 269.320 2150.000 269.920 ;
    END
  END pwr_ctrl_out[3]
  PIN resetb
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 2.400 ;
    END
  END resetb
  PIN sdo_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2147.600 656.240 2150.000 656.840 ;
    END
  END sdo_out
  PIN sdo_outenb
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2147.600 733.080 2150.000 733.680 ;
    END
  END sdo_outenb
  PIN user_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 2.400 5.400 ;
    END
  END user_addr[0]
  PIN user_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 2.400 15.600 ;
    END
  END user_addr[1]
  PIN user_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 2.400 26.480 ;
    END
  END user_addr[2]
  PIN user_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 2.400 37.360 ;
    END
  END user_addr[3]
  PIN user_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 2.400 47.560 ;
    END
  END user_addr[4]
  PIN user_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 2.400 58.440 ;
    END
  END user_addr[5]
  PIN user_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 2.400 69.320 ;
    END
  END user_addr[6]
  PIN user_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 2.400 76.120 ;
    END
  END user_addr[7]
  PIN user_clk
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 2.400 2.000 ;
    END
  END user_clk
  PIN user_ena[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 2.400 8.800 ;
    END
  END user_ena[0]
  PIN user_ena[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 2.400 19.680 ;
    END
  END user_ena[1]
  PIN user_ena[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 2.400 29.880 ;
    END
  END user_ena[2]
  PIN user_ena[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 2.400 40.760 ;
    END
  END user_ena[3]
  PIN user_ena[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 2.400 51.640 ;
    END
  END user_ena[4]
  PIN user_ena[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 2.400 61.840 ;
    END
  END user_ena[5]
  PIN user_rdata[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 2.400 12.200 ;
    END
  END user_rdata[0]
  PIN user_rdata[100]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.080 2.400 410.680 ;
    END
  END user_rdata[100]
  PIN user_rdata[101]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 2.400 414.080 ;
    END
  END user_rdata[101]
  PIN user_rdata[102]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.880 2.400 417.480 ;
    END
  END user_rdata[102]
  PIN user_rdata[103]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.960 2.400 421.560 ;
    END
  END user_rdata[103]
  PIN user_rdata[104]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 424.360 2.400 424.960 ;
    END
  END user_rdata[104]
  PIN user_rdata[105]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.760 2.400 428.360 ;
    END
  END user_rdata[105]
  PIN user_rdata[106]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.160 2.400 431.760 ;
    END
  END user_rdata[106]
  PIN user_rdata[107]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 2.400 435.840 ;
    END
  END user_rdata[107]
  PIN user_rdata[108]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 2.400 439.240 ;
    END
  END user_rdata[108]
  PIN user_rdata[109]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 2.400 442.640 ;
    END
  END user_rdata[109]
  PIN user_rdata[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 2.400 90.400 ;
    END
  END user_rdata[10]
  PIN user_rdata[110]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 2.400 446.040 ;
    END
  END user_rdata[110]
  PIN user_rdata[111]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 2.400 449.440 ;
    END
  END user_rdata[111]
  PIN user_rdata[112]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 2.400 453.520 ;
    END
  END user_rdata[112]
  PIN user_rdata[113]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 456.320 2.400 456.920 ;
    END
  END user_rdata[113]
  PIN user_rdata[114]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.720 2.400 460.320 ;
    END
  END user_rdata[114]
  PIN user_rdata[115]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.120 2.400 463.720 ;
    END
  END user_rdata[115]
  PIN user_rdata[116]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.200 2.400 467.800 ;
    END
  END user_rdata[116]
  PIN user_rdata[117]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 2.400 471.200 ;
    END
  END user_rdata[117]
  PIN user_rdata[118]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.000 2.400 474.600 ;
    END
  END user_rdata[118]
  PIN user_rdata[119]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 477.400 2.400 478.000 ;
    END
  END user_rdata[119]
  PIN user_rdata[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 2.400 93.800 ;
    END
  END user_rdata[11]
  PIN user_rdata[120]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 481.480 2.400 482.080 ;
    END
  END user_rdata[120]
  PIN user_rdata[121]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.880 2.400 485.480 ;
    END
  END user_rdata[121]
  PIN user_rdata[122]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.280 2.400 488.880 ;
    END
  END user_rdata[122]
  PIN user_rdata[123]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.680 2.400 492.280 ;
    END
  END user_rdata[123]
  PIN user_rdata[124]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.080 2.400 495.680 ;
    END
  END user_rdata[124]
  PIN user_rdata[125]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 2.400 499.760 ;
    END
  END user_rdata[125]
  PIN user_rdata[126]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 502.560 2.400 503.160 ;
    END
  END user_rdata[126]
  PIN user_rdata[127]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 505.960 2.400 506.560 ;
    END
  END user_rdata[127]
  PIN user_rdata[128]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 509.360 2.400 509.960 ;
    END
  END user_rdata[128]
  PIN user_rdata[129]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 513.440 2.400 514.040 ;
    END
  END user_rdata[129]
  PIN user_rdata[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 2.400 97.880 ;
    END
  END user_rdata[12]
  PIN user_rdata[130]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 2.400 517.440 ;
    END
  END user_rdata[130]
  PIN user_rdata[131]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 2.400 520.840 ;
    END
  END user_rdata[131]
  PIN user_rdata[132]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 2.400 524.240 ;
    END
  END user_rdata[132]
  PIN user_rdata[133]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.720 2.400 528.320 ;
    END
  END user_rdata[133]
  PIN user_rdata[134]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.120 2.400 531.720 ;
    END
  END user_rdata[134]
  PIN user_rdata[135]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 534.520 2.400 535.120 ;
    END
  END user_rdata[135]
  PIN user_rdata[136]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.920 2.400 538.520 ;
    END
  END user_rdata[136]
  PIN user_rdata[137]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 541.320 2.400 541.920 ;
    END
  END user_rdata[137]
  PIN user_rdata[138]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 545.400 2.400 546.000 ;
    END
  END user_rdata[138]
  PIN user_rdata[139]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.800 2.400 549.400 ;
    END
  END user_rdata[139]
  PIN user_rdata[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 2.400 101.280 ;
    END
  END user_rdata[13]
  PIN user_rdata[140]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.200 2.400 552.800 ;
    END
  END user_rdata[140]
  PIN user_rdata[141]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 555.600 2.400 556.200 ;
    END
  END user_rdata[141]
  PIN user_rdata[142]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.680 2.400 560.280 ;
    END
  END user_rdata[142]
  PIN user_rdata[143]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.080 2.400 563.680 ;
    END
  END user_rdata[143]
  PIN user_rdata[144]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 566.480 2.400 567.080 ;
    END
  END user_rdata[144]
  PIN user_rdata[145]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.880 2.400 570.480 ;
    END
  END user_rdata[145]
  PIN user_rdata[146]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.960 2.400 574.560 ;
    END
  END user_rdata[146]
  PIN user_rdata[147]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 577.360 2.400 577.960 ;
    END
  END user_rdata[147]
  PIN user_rdata[148]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 580.760 2.400 581.360 ;
    END
  END user_rdata[148]
  PIN user_rdata[149]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.160 2.400 584.760 ;
    END
  END user_rdata[149]
  PIN user_rdata[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.080 2.400 104.680 ;
    END
  END user_rdata[14]
  PIN user_rdata[150]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 587.560 2.400 588.160 ;
    END
  END user_rdata[150]
  PIN user_rdata[151]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 2.400 592.240 ;
    END
  END user_rdata[151]
  PIN user_rdata[152]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 2.400 595.640 ;
    END
  END user_rdata[152]
  PIN user_rdata[153]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 2.400 599.040 ;
    END
  END user_rdata[153]
  PIN user_rdata[154]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.840 2.400 602.440 ;
    END
  END user_rdata[154]
  PIN user_rdata[155]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.920 2.400 606.520 ;
    END
  END user_rdata[155]
  PIN user_rdata[156]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 609.320 2.400 609.920 ;
    END
  END user_rdata[156]
  PIN user_rdata[157]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.720 2.400 613.320 ;
    END
  END user_rdata[157]
  PIN user_rdata[158]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.120 2.400 616.720 ;
    END
  END user_rdata[158]
  PIN user_rdata[159]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.200 2.400 620.800 ;
    END
  END user_rdata[159]
  PIN user_rdata[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 2.400 108.080 ;
    END
  END user_rdata[15]
  PIN user_rdata[160]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 623.600 2.400 624.200 ;
    END
  END user_rdata[160]
  PIN user_rdata[161]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.000 2.400 627.600 ;
    END
  END user_rdata[161]
  PIN user_rdata[162]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 630.400 2.400 631.000 ;
    END
  END user_rdata[162]
  PIN user_rdata[163]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 633.800 2.400 634.400 ;
    END
  END user_rdata[163]
  PIN user_rdata[164]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 637.880 2.400 638.480 ;
    END
  END user_rdata[164]
  PIN user_rdata[165]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 641.280 2.400 641.880 ;
    END
  END user_rdata[165]
  PIN user_rdata[166]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 644.680 2.400 645.280 ;
    END
  END user_rdata[166]
  PIN user_rdata[167]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.080 2.400 648.680 ;
    END
  END user_rdata[167]
  PIN user_rdata[168]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.160 2.400 652.760 ;
    END
  END user_rdata[168]
  PIN user_rdata[169]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 655.560 2.400 656.160 ;
    END
  END user_rdata[169]
  PIN user_rdata[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 2.400 112.160 ;
    END
  END user_rdata[16]
  PIN user_rdata[170]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 658.960 2.400 659.560 ;
    END
  END user_rdata[170]
  PIN user_rdata[171]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 662.360 2.400 662.960 ;
    END
  END user_rdata[171]
  PIN user_rdata[172]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 2.400 667.040 ;
    END
  END user_rdata[172]
  PIN user_rdata[173]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.840 2.400 670.440 ;
    END
  END user_rdata[173]
  PIN user_rdata[174]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 2.400 673.840 ;
    END
  END user_rdata[174]
  PIN user_rdata[175]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 676.640 2.400 677.240 ;
    END
  END user_rdata[175]
  PIN user_rdata[176]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 2.400 680.640 ;
    END
  END user_rdata[176]
  PIN user_rdata[177]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.120 2.400 684.720 ;
    END
  END user_rdata[177]
  PIN user_rdata[178]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 687.520 2.400 688.120 ;
    END
  END user_rdata[178]
  PIN user_rdata[179]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.920 2.400 691.520 ;
    END
  END user_rdata[179]
  PIN user_rdata[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 2.400 115.560 ;
    END
  END user_rdata[17]
  PIN user_rdata[180]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 694.320 2.400 694.920 ;
    END
  END user_rdata[180]
  PIN user_rdata[181]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 698.400 2.400 699.000 ;
    END
  END user_rdata[181]
  PIN user_rdata[182]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 701.800 2.400 702.400 ;
    END
  END user_rdata[182]
  PIN user_rdata[183]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.200 2.400 705.800 ;
    END
  END user_rdata[183]
  PIN user_rdata[184]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 708.600 2.400 709.200 ;
    END
  END user_rdata[184]
  PIN user_rdata[185]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 712.680 2.400 713.280 ;
    END
  END user_rdata[185]
  PIN user_rdata[186]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.080 2.400 716.680 ;
    END
  END user_rdata[186]
  PIN user_rdata[187]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 719.480 2.400 720.080 ;
    END
  END user_rdata[187]
  PIN user_rdata[188]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.880 2.400 723.480 ;
    END
  END user_rdata[188]
  PIN user_rdata[189]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 726.280 2.400 726.880 ;
    END
  END user_rdata[189]
  PIN user_rdata[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 2.400 118.960 ;
    END
  END user_rdata[18]
  PIN user_rdata[190]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 730.360 2.400 730.960 ;
    END
  END user_rdata[190]
  PIN user_rdata[191]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 733.760 2.400 734.360 ;
    END
  END user_rdata[191]
  PIN user_rdata[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.760 2.400 122.360 ;
    END
  END user_rdata[19]
  PIN user_rdata[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 2.400 23.080 ;
    END
  END user_rdata[1]
  PIN user_rdata[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 2.400 126.440 ;
    END
  END user_rdata[20]
  PIN user_rdata[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 2.400 129.840 ;
    END
  END user_rdata[21]
  PIN user_rdata[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 2.400 133.240 ;
    END
  END user_rdata[22]
  PIN user_rdata[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 2.400 136.640 ;
    END
  END user_rdata[23]
  PIN user_rdata[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 2.400 140.040 ;
    END
  END user_rdata[24]
  PIN user_rdata[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 2.400 144.120 ;
    END
  END user_rdata[25]
  PIN user_rdata[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 2.400 147.520 ;
    END
  END user_rdata[26]
  PIN user_rdata[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.320 2.400 150.920 ;
    END
  END user_rdata[27]
  PIN user_rdata[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 2.400 154.320 ;
    END
  END user_rdata[28]
  PIN user_rdata[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 2.400 158.400 ;
    END
  END user_rdata[29]
  PIN user_rdata[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 2.400 33.960 ;
    END
  END user_rdata[2]
  PIN user_rdata[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.200 2.400 161.800 ;
    END
  END user_rdata[30]
  PIN user_rdata[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 2.400 165.200 ;
    END
  END user_rdata[31]
  PIN user_rdata[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 2.400 168.600 ;
    END
  END user_rdata[32]
  PIN user_rdata[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.080 2.400 172.680 ;
    END
  END user_rdata[33]
  PIN user_rdata[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 2.400 176.080 ;
    END
  END user_rdata[34]
  PIN user_rdata[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 2.400 179.480 ;
    END
  END user_rdata[35]
  PIN user_rdata[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 2.400 182.880 ;
    END
  END user_rdata[36]
  PIN user_rdata[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.680 2.400 186.280 ;
    END
  END user_rdata[37]
  PIN user_rdata[38]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.760 2.400 190.360 ;
    END
  END user_rdata[38]
  PIN user_rdata[39]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 2.400 193.760 ;
    END
  END user_rdata[39]
  PIN user_rdata[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 2.400 44.160 ;
    END
  END user_rdata[3]
  PIN user_rdata[40]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 2.400 197.160 ;
    END
  END user_rdata[40]
  PIN user_rdata[41]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 2.400 200.560 ;
    END
  END user_rdata[41]
  PIN user_rdata[42]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 2.400 204.640 ;
    END
  END user_rdata[42]
  PIN user_rdata[43]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 2.400 208.040 ;
    END
  END user_rdata[43]
  PIN user_rdata[44]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 2.400 211.440 ;
    END
  END user_rdata[44]
  PIN user_rdata[45]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 2.400 214.840 ;
    END
  END user_rdata[45]
  PIN user_rdata[46]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.320 2.400 218.920 ;
    END
  END user_rdata[46]
  PIN user_rdata[47]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 2.400 222.320 ;
    END
  END user_rdata[47]
  PIN user_rdata[48]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.120 2.400 225.720 ;
    END
  END user_rdata[48]
  PIN user_rdata[49]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 2.400 229.120 ;
    END
  END user_rdata[49]
  PIN user_rdata[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 2.400 55.040 ;
    END
  END user_rdata[4]
  PIN user_rdata[50]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.920 2.400 232.520 ;
    END
  END user_rdata[50]
  PIN user_rdata[51]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.000 2.400 236.600 ;
    END
  END user_rdata[51]
  PIN user_rdata[52]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 2.400 240.000 ;
    END
  END user_rdata[52]
  PIN user_rdata[53]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.800 2.400 243.400 ;
    END
  END user_rdata[53]
  PIN user_rdata[54]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 2.400 246.800 ;
    END
  END user_rdata[54]
  PIN user_rdata[55]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 2.400 250.880 ;
    END
  END user_rdata[55]
  PIN user_rdata[56]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.680 2.400 254.280 ;
    END
  END user_rdata[56]
  PIN user_rdata[57]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 2.400 257.680 ;
    END
  END user_rdata[57]
  PIN user_rdata[58]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 260.480 2.400 261.080 ;
    END
  END user_rdata[58]
  PIN user_rdata[59]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.560 2.400 265.160 ;
    END
  END user_rdata[59]
  PIN user_rdata[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 2.400 65.920 ;
    END
  END user_rdata[5]
  PIN user_rdata[60]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 2.400 268.560 ;
    END
  END user_rdata[60]
  PIN user_rdata[61]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 271.360 2.400 271.960 ;
    END
  END user_rdata[61]
  PIN user_rdata[62]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 2.400 275.360 ;
    END
  END user_rdata[62]
  PIN user_rdata[63]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.160 2.400 278.760 ;
    END
  END user_rdata[63]
  PIN user_rdata[64]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 2.400 282.840 ;
    END
  END user_rdata[64]
  PIN user_rdata[65]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 2.400 286.240 ;
    END
  END user_rdata[65]
  PIN user_rdata[66]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 2.400 289.640 ;
    END
  END user_rdata[66]
  PIN user_rdata[67]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 2.400 293.040 ;
    END
  END user_rdata[67]
  PIN user_rdata[68]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 2.400 297.120 ;
    END
  END user_rdata[68]
  PIN user_rdata[69]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.920 2.400 300.520 ;
    END
  END user_rdata[69]
  PIN user_rdata[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 2.400 72.720 ;
    END
  END user_rdata[6]
  PIN user_rdata[70]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 2.400 303.920 ;
    END
  END user_rdata[70]
  PIN user_rdata[71]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.720 2.400 307.320 ;
    END
  END user_rdata[71]
  PIN user_rdata[72]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.800 2.400 311.400 ;
    END
  END user_rdata[72]
  PIN user_rdata[73]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 2.400 314.800 ;
    END
  END user_rdata[73]
  PIN user_rdata[74]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 317.600 2.400 318.200 ;
    END
  END user_rdata[74]
  PIN user_rdata[75]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 2.400 321.600 ;
    END
  END user_rdata[75]
  PIN user_rdata[76]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 324.400 2.400 325.000 ;
    END
  END user_rdata[76]
  PIN user_rdata[77]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 328.480 2.400 329.080 ;
    END
  END user_rdata[77]
  PIN user_rdata[78]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 2.400 332.480 ;
    END
  END user_rdata[78]
  PIN user_rdata[79]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.280 2.400 335.880 ;
    END
  END user_rdata[79]
  PIN user_rdata[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 2.400 80.200 ;
    END
  END user_rdata[7]
  PIN user_rdata[80]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 2.400 339.280 ;
    END
  END user_rdata[80]
  PIN user_rdata[81]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 2.400 343.360 ;
    END
  END user_rdata[81]
  PIN user_rdata[82]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.160 2.400 346.760 ;
    END
  END user_rdata[82]
  PIN user_rdata[83]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 2.400 350.160 ;
    END
  END user_rdata[83]
  PIN user_rdata[84]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.960 2.400 353.560 ;
    END
  END user_rdata[84]
  PIN user_rdata[85]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 2.400 357.640 ;
    END
  END user_rdata[85]
  PIN user_rdata[86]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 2.400 361.040 ;
    END
  END user_rdata[86]
  PIN user_rdata[87]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 2.400 364.440 ;
    END
  END user_rdata[87]
  PIN user_rdata[88]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 2.400 367.840 ;
    END
  END user_rdata[88]
  PIN user_rdata[89]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 2.400 371.240 ;
    END
  END user_rdata[89]
  PIN user_rdata[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 2.400 83.600 ;
    END
  END user_rdata[8]
  PIN user_rdata[90]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.720 2.400 375.320 ;
    END
  END user_rdata[90]
  PIN user_rdata[91]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 2.400 378.720 ;
    END
  END user_rdata[91]
  PIN user_rdata[92]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 381.520 2.400 382.120 ;
    END
  END user_rdata[92]
  PIN user_rdata[93]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 2.400 385.520 ;
    END
  END user_rdata[93]
  PIN user_rdata[94]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 2.400 389.600 ;
    END
  END user_rdata[94]
  PIN user_rdata[95]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 392.400 2.400 393.000 ;
    END
  END user_rdata[95]
  PIN user_rdata[96]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 2.400 396.400 ;
    END
  END user_rdata[96]
  PIN user_rdata[97]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.200 2.400 399.800 ;
    END
  END user_rdata[97]
  PIN user_rdata[98]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.280 2.400 403.880 ;
    END
  END user_rdata[98]
  PIN user_rdata[99]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.680 2.400 407.280 ;
    END
  END user_rdata[99]
  PIN user_rdata[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 2.400 87.000 ;
    END
  END user_rdata[9]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 2144.060 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 2144.060 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 3.365 10.795 2144.060 847.875 ;
      LAYER met1 ;
        RECT 0.070 1.740 2148.590 849.620 ;
      LAYER met2 ;
        RECT 0.100 847.320 1.190 849.650 ;
        RECT 2.030 847.320 3.950 849.650 ;
        RECT 4.790 847.320 7.170 849.650 ;
        RECT 8.010 847.320 10.390 849.650 ;
        RECT 11.230 847.320 13.610 849.650 ;
        RECT 14.450 847.320 16.830 849.650 ;
        RECT 17.670 847.320 19.590 849.650 ;
        RECT 20.430 847.320 22.810 849.650 ;
        RECT 23.650 847.320 26.030 849.650 ;
        RECT 26.870 847.320 29.250 849.650 ;
        RECT 30.090 847.320 32.470 849.650 ;
        RECT 33.310 847.320 35.230 849.650 ;
        RECT 36.070 847.320 38.450 849.650 ;
        RECT 39.290 847.320 41.670 849.650 ;
        RECT 42.510 847.320 44.890 849.650 ;
        RECT 45.730 847.320 48.110 849.650 ;
        RECT 48.950 847.320 50.870 849.650 ;
        RECT 51.710 847.320 54.090 849.650 ;
        RECT 54.930 847.320 57.310 849.650 ;
        RECT 58.150 847.320 60.530 849.650 ;
        RECT 61.370 847.320 63.750 849.650 ;
        RECT 64.590 847.320 66.510 849.650 ;
        RECT 67.350 847.320 69.730 849.650 ;
        RECT 70.570 847.320 72.950 849.650 ;
        RECT 73.790 847.320 76.170 849.650 ;
        RECT 77.010 847.320 79.390 849.650 ;
        RECT 80.230 847.320 82.150 849.650 ;
        RECT 82.990 847.320 85.370 849.650 ;
        RECT 86.210 847.320 88.590 849.650 ;
        RECT 89.430 847.320 91.810 849.650 ;
        RECT 92.650 847.320 95.030 849.650 ;
        RECT 95.870 847.320 97.790 849.650 ;
        RECT 98.630 847.320 101.010 849.650 ;
        RECT 101.850 847.320 104.230 849.650 ;
        RECT 105.070 847.320 107.450 849.650 ;
        RECT 108.290 847.320 110.670 849.650 ;
        RECT 111.510 847.320 113.430 849.650 ;
        RECT 114.270 847.320 116.650 849.650 ;
        RECT 117.490 847.320 119.870 849.650 ;
        RECT 120.710 847.320 123.090 849.650 ;
        RECT 123.930 847.320 126.310 849.650 ;
        RECT 127.150 847.320 129.070 849.650 ;
        RECT 129.910 847.320 132.290 849.650 ;
        RECT 133.130 847.320 135.510 849.650 ;
        RECT 136.350 847.320 138.730 849.650 ;
        RECT 139.570 847.320 141.950 849.650 ;
        RECT 142.790 847.320 144.710 849.650 ;
        RECT 145.550 847.320 147.930 849.650 ;
        RECT 148.770 847.320 151.150 849.650 ;
        RECT 151.990 847.320 154.370 849.650 ;
        RECT 155.210 847.320 157.590 849.650 ;
        RECT 158.430 847.320 160.350 849.650 ;
        RECT 161.190 847.320 163.570 849.650 ;
        RECT 164.410 847.320 166.790 849.650 ;
        RECT 167.630 847.320 170.010 849.650 ;
        RECT 170.850 847.320 173.230 849.650 ;
        RECT 174.070 847.320 175.990 849.650 ;
        RECT 176.830 847.320 179.210 849.650 ;
        RECT 180.050 847.320 182.430 849.650 ;
        RECT 183.270 847.320 185.650 849.650 ;
        RECT 186.490 847.320 188.870 849.650 ;
        RECT 189.710 847.320 192.090 849.650 ;
        RECT 192.930 847.320 194.850 849.650 ;
        RECT 195.690 847.320 198.070 849.650 ;
        RECT 198.910 847.320 201.290 849.650 ;
        RECT 202.130 847.320 204.510 849.650 ;
        RECT 205.350 847.320 207.730 849.650 ;
        RECT 208.570 847.320 210.490 849.650 ;
        RECT 211.330 847.320 213.710 849.650 ;
        RECT 214.550 847.320 216.930 849.650 ;
        RECT 217.770 847.320 220.150 849.650 ;
        RECT 220.990 847.320 223.370 849.650 ;
        RECT 224.210 847.320 226.130 849.650 ;
        RECT 226.970 847.320 229.350 849.650 ;
        RECT 230.190 847.320 232.570 849.650 ;
        RECT 233.410 847.320 235.790 849.650 ;
        RECT 236.630 847.320 239.010 849.650 ;
        RECT 239.850 847.320 241.770 849.650 ;
        RECT 242.610 847.320 244.990 849.650 ;
        RECT 245.830 847.320 248.210 849.650 ;
        RECT 249.050 847.320 251.430 849.650 ;
        RECT 252.270 847.320 254.650 849.650 ;
        RECT 255.490 847.320 257.410 849.650 ;
        RECT 258.250 847.320 260.630 849.650 ;
        RECT 261.470 847.320 263.850 849.650 ;
        RECT 264.690 847.320 267.070 849.650 ;
        RECT 267.910 847.320 270.290 849.650 ;
        RECT 271.130 847.320 273.050 849.650 ;
        RECT 273.890 847.320 276.270 849.650 ;
        RECT 277.110 847.320 279.490 849.650 ;
        RECT 280.330 847.320 282.710 849.650 ;
        RECT 283.550 847.320 285.930 849.650 ;
        RECT 286.770 847.320 288.690 849.650 ;
        RECT 289.530 847.320 291.910 849.650 ;
        RECT 292.750 847.320 295.130 849.650 ;
        RECT 295.970 847.320 298.350 849.650 ;
        RECT 299.190 847.320 301.570 849.650 ;
        RECT 302.410 847.320 304.330 849.650 ;
        RECT 305.170 847.320 307.550 849.650 ;
        RECT 308.390 847.320 310.770 849.650 ;
        RECT 311.610 847.320 313.990 849.650 ;
        RECT 314.830 847.320 317.210 849.650 ;
        RECT 318.050 847.320 319.970 849.650 ;
        RECT 320.810 847.320 323.190 849.650 ;
        RECT 324.030 847.320 326.410 849.650 ;
        RECT 327.250 847.320 329.630 849.650 ;
        RECT 330.470 847.320 332.850 849.650 ;
        RECT 333.690 847.320 335.610 849.650 ;
        RECT 336.450 847.320 338.830 849.650 ;
        RECT 339.670 847.320 342.050 849.650 ;
        RECT 342.890 847.320 345.270 849.650 ;
        RECT 346.110 847.320 348.490 849.650 ;
        RECT 349.330 847.320 351.250 849.650 ;
        RECT 352.090 847.320 354.470 849.650 ;
        RECT 355.310 847.320 357.690 849.650 ;
        RECT 358.530 847.320 360.910 849.650 ;
        RECT 361.750 847.320 364.130 849.650 ;
        RECT 364.970 847.320 367.350 849.650 ;
        RECT 368.190 847.320 370.110 849.650 ;
        RECT 370.950 847.320 373.330 849.650 ;
        RECT 374.170 847.320 376.550 849.650 ;
        RECT 377.390 847.320 379.770 849.650 ;
        RECT 380.610 847.320 382.990 849.650 ;
        RECT 383.830 847.320 385.750 849.650 ;
        RECT 386.590 847.320 388.970 849.650 ;
        RECT 389.810 847.320 392.190 849.650 ;
        RECT 393.030 847.320 395.410 849.650 ;
        RECT 396.250 847.320 398.630 849.650 ;
        RECT 399.470 847.320 401.390 849.650 ;
        RECT 402.230 847.320 404.610 849.650 ;
        RECT 405.450 847.320 407.830 849.650 ;
        RECT 408.670 847.320 411.050 849.650 ;
        RECT 411.890 847.320 414.270 849.650 ;
        RECT 415.110 847.320 417.030 849.650 ;
        RECT 417.870 847.320 420.250 849.650 ;
        RECT 421.090 847.320 423.470 849.650 ;
        RECT 424.310 847.320 426.690 849.650 ;
        RECT 427.530 847.320 429.910 849.650 ;
        RECT 430.750 847.320 432.670 849.650 ;
        RECT 433.510 847.320 435.890 849.650 ;
        RECT 436.730 847.320 439.110 849.650 ;
        RECT 439.950 847.320 442.330 849.650 ;
        RECT 443.170 847.320 445.550 849.650 ;
        RECT 446.390 847.320 448.310 849.650 ;
        RECT 449.150 847.320 451.530 849.650 ;
        RECT 452.370 847.320 454.750 849.650 ;
        RECT 455.590 847.320 457.970 849.650 ;
        RECT 458.810 847.320 461.190 849.650 ;
        RECT 462.030 847.320 463.950 849.650 ;
        RECT 464.790 847.320 467.170 849.650 ;
        RECT 468.010 847.320 470.390 849.650 ;
        RECT 471.230 847.320 473.610 849.650 ;
        RECT 474.450 847.320 476.830 849.650 ;
        RECT 477.670 847.320 479.590 849.650 ;
        RECT 480.430 847.320 482.810 849.650 ;
        RECT 483.650 847.320 486.030 849.650 ;
        RECT 486.870 847.320 489.250 849.650 ;
        RECT 490.090 847.320 492.470 849.650 ;
        RECT 493.310 847.320 495.230 849.650 ;
        RECT 496.070 847.320 498.450 849.650 ;
        RECT 499.290 847.320 501.670 849.650 ;
        RECT 502.510 847.320 504.890 849.650 ;
        RECT 505.730 847.320 508.110 849.650 ;
        RECT 508.950 847.320 510.870 849.650 ;
        RECT 511.710 847.320 514.090 849.650 ;
        RECT 514.930 847.320 517.310 849.650 ;
        RECT 518.150 847.320 520.530 849.650 ;
        RECT 521.370 847.320 523.750 849.650 ;
        RECT 524.590 847.320 526.510 849.650 ;
        RECT 527.350 847.320 529.730 849.650 ;
        RECT 530.570 847.320 532.950 849.650 ;
        RECT 533.790 847.320 536.170 849.650 ;
        RECT 537.010 847.320 539.390 849.650 ;
        RECT 540.230 847.320 542.610 849.650 ;
        RECT 543.450 847.320 545.370 849.650 ;
        RECT 546.210 847.320 548.590 849.650 ;
        RECT 549.430 847.320 551.810 849.650 ;
        RECT 552.650 847.320 555.030 849.650 ;
        RECT 555.870 847.320 558.250 849.650 ;
        RECT 559.090 847.320 561.010 849.650 ;
        RECT 561.850 847.320 564.230 849.650 ;
        RECT 565.070 847.320 567.450 849.650 ;
        RECT 568.290 847.320 570.670 849.650 ;
        RECT 571.510 847.320 573.890 849.650 ;
        RECT 574.730 847.320 576.650 849.650 ;
        RECT 577.490 847.320 579.870 849.650 ;
        RECT 580.710 847.320 583.090 849.650 ;
        RECT 583.930 847.320 586.310 849.650 ;
        RECT 587.150 847.320 589.530 849.650 ;
        RECT 590.370 847.320 592.290 849.650 ;
        RECT 593.130 847.320 595.510 849.650 ;
        RECT 596.350 847.320 598.730 849.650 ;
        RECT 599.570 847.320 601.950 849.650 ;
        RECT 602.790 847.320 605.170 849.650 ;
        RECT 606.010 847.320 607.930 849.650 ;
        RECT 608.770 847.320 611.150 849.650 ;
        RECT 611.990 847.320 614.370 849.650 ;
        RECT 615.210 847.320 617.590 849.650 ;
        RECT 618.430 847.320 620.810 849.650 ;
        RECT 621.650 847.320 623.570 849.650 ;
        RECT 624.410 847.320 626.790 849.650 ;
        RECT 627.630 847.320 630.010 849.650 ;
        RECT 630.850 847.320 633.230 849.650 ;
        RECT 634.070 847.320 636.450 849.650 ;
        RECT 637.290 847.320 639.210 849.650 ;
        RECT 640.050 847.320 642.430 849.650 ;
        RECT 643.270 847.320 645.650 849.650 ;
        RECT 646.490 847.320 648.870 849.650 ;
        RECT 649.710 847.320 652.090 849.650 ;
        RECT 652.930 847.320 654.850 849.650 ;
        RECT 655.690 847.320 658.070 849.650 ;
        RECT 658.910 847.320 661.290 849.650 ;
        RECT 662.130 847.320 664.510 849.650 ;
        RECT 665.350 847.320 667.730 849.650 ;
        RECT 668.570 847.320 670.490 849.650 ;
        RECT 671.330 847.320 673.710 849.650 ;
        RECT 674.550 847.320 676.930 849.650 ;
        RECT 677.770 847.320 680.150 849.650 ;
        RECT 680.990 847.320 683.370 849.650 ;
        RECT 684.210 847.320 686.130 849.650 ;
        RECT 686.970 847.320 689.350 849.650 ;
        RECT 690.190 847.320 692.570 849.650 ;
        RECT 693.410 847.320 695.790 849.650 ;
        RECT 696.630 847.320 699.010 849.650 ;
        RECT 699.850 847.320 701.770 849.650 ;
        RECT 702.610 847.320 704.990 849.650 ;
        RECT 705.830 847.320 708.210 849.650 ;
        RECT 709.050 847.320 711.430 849.650 ;
        RECT 712.270 847.320 714.650 849.650 ;
        RECT 715.490 847.320 717.870 849.650 ;
        RECT 718.710 847.320 720.630 849.650 ;
        RECT 721.470 847.320 723.850 849.650 ;
        RECT 724.690 847.320 727.070 849.650 ;
        RECT 727.910 847.320 730.290 849.650 ;
        RECT 731.130 847.320 733.510 849.650 ;
        RECT 734.350 847.320 736.270 849.650 ;
        RECT 737.110 847.320 739.490 849.650 ;
        RECT 740.330 847.320 742.710 849.650 ;
        RECT 743.550 847.320 745.930 849.650 ;
        RECT 746.770 847.320 749.150 849.650 ;
        RECT 749.990 847.320 751.910 849.650 ;
        RECT 752.750 847.320 755.130 849.650 ;
        RECT 755.970 847.320 758.350 849.650 ;
        RECT 759.190 847.320 761.570 849.650 ;
        RECT 762.410 847.320 764.790 849.650 ;
        RECT 765.630 847.320 767.550 849.650 ;
        RECT 768.390 847.320 770.770 849.650 ;
        RECT 771.610 847.320 773.990 849.650 ;
        RECT 774.830 847.320 777.210 849.650 ;
        RECT 778.050 847.320 780.430 849.650 ;
        RECT 781.270 847.320 783.190 849.650 ;
        RECT 784.030 847.320 786.410 849.650 ;
        RECT 787.250 847.320 789.630 849.650 ;
        RECT 790.470 847.320 792.850 849.650 ;
        RECT 793.690 847.320 796.070 849.650 ;
        RECT 796.910 847.320 798.830 849.650 ;
        RECT 799.670 847.320 802.050 849.650 ;
        RECT 802.890 847.320 805.270 849.650 ;
        RECT 806.110 847.320 808.490 849.650 ;
        RECT 809.330 847.320 811.710 849.650 ;
        RECT 812.550 847.320 814.470 849.650 ;
        RECT 815.310 847.320 817.690 849.650 ;
        RECT 818.530 847.320 820.910 849.650 ;
        RECT 821.750 847.320 824.130 849.650 ;
        RECT 824.970 847.320 827.350 849.650 ;
        RECT 828.190 847.320 830.110 849.650 ;
        RECT 830.950 847.320 833.330 849.650 ;
        RECT 834.170 847.320 836.550 849.650 ;
        RECT 837.390 847.320 839.770 849.650 ;
        RECT 840.610 847.320 842.990 849.650 ;
        RECT 843.830 847.320 845.750 849.650 ;
        RECT 846.590 847.320 848.970 849.650 ;
        RECT 849.810 847.320 852.190 849.650 ;
        RECT 853.030 847.320 855.410 849.650 ;
        RECT 856.250 847.320 858.630 849.650 ;
        RECT 859.470 847.320 861.390 849.650 ;
        RECT 862.230 847.320 864.610 849.650 ;
        RECT 865.450 847.320 867.830 849.650 ;
        RECT 868.670 847.320 871.050 849.650 ;
        RECT 871.890 847.320 874.270 849.650 ;
        RECT 875.110 847.320 877.030 849.650 ;
        RECT 877.870 847.320 880.250 849.650 ;
        RECT 881.090 847.320 883.470 849.650 ;
        RECT 884.310 847.320 886.690 849.650 ;
        RECT 887.530 847.320 889.910 849.650 ;
        RECT 890.750 847.320 892.670 849.650 ;
        RECT 893.510 847.320 895.890 849.650 ;
        RECT 896.730 847.320 899.110 849.650 ;
        RECT 899.950 847.320 902.330 849.650 ;
        RECT 903.170 847.320 905.550 849.650 ;
        RECT 906.390 847.320 908.770 849.650 ;
        RECT 909.610 847.320 911.530 849.650 ;
        RECT 912.370 847.320 914.750 849.650 ;
        RECT 915.590 847.320 917.970 849.650 ;
        RECT 918.810 847.320 921.190 849.650 ;
        RECT 922.030 847.320 924.410 849.650 ;
        RECT 925.250 847.320 927.170 849.650 ;
        RECT 928.010 847.320 930.390 849.650 ;
        RECT 931.230 847.320 933.610 849.650 ;
        RECT 934.450 847.320 936.830 849.650 ;
        RECT 937.670 847.320 940.050 849.650 ;
        RECT 940.890 847.320 942.810 849.650 ;
        RECT 943.650 847.320 946.030 849.650 ;
        RECT 946.870 847.320 949.250 849.650 ;
        RECT 950.090 847.320 952.470 849.650 ;
        RECT 953.310 847.320 955.690 849.650 ;
        RECT 956.530 847.320 958.450 849.650 ;
        RECT 959.290 847.320 961.670 849.650 ;
        RECT 962.510 847.320 964.890 849.650 ;
        RECT 965.730 847.320 968.110 849.650 ;
        RECT 968.950 847.320 971.330 849.650 ;
        RECT 972.170 847.320 974.090 849.650 ;
        RECT 974.930 847.320 977.310 849.650 ;
        RECT 978.150 847.320 980.530 849.650 ;
        RECT 981.370 847.320 983.750 849.650 ;
        RECT 984.590 847.320 986.970 849.650 ;
        RECT 987.810 847.320 989.730 849.650 ;
        RECT 990.570 847.320 992.950 849.650 ;
        RECT 993.790 847.320 996.170 849.650 ;
        RECT 997.010 847.320 999.390 849.650 ;
        RECT 1000.230 847.320 1002.610 849.650 ;
        RECT 1003.450 847.320 1005.370 849.650 ;
        RECT 1006.210 847.320 1008.590 849.650 ;
        RECT 1009.430 847.320 1011.810 849.650 ;
        RECT 1012.650 847.320 1015.030 849.650 ;
        RECT 1015.870 847.320 1018.250 849.650 ;
        RECT 1019.090 847.320 1021.010 849.650 ;
        RECT 1021.850 847.320 1024.230 849.650 ;
        RECT 1025.070 847.320 1027.450 849.650 ;
        RECT 1028.290 847.320 1030.670 849.650 ;
        RECT 1031.510 847.320 1033.890 849.650 ;
        RECT 1034.730 847.320 1036.650 849.650 ;
        RECT 1037.490 847.320 1039.870 849.650 ;
        RECT 1040.710 847.320 1043.090 849.650 ;
        RECT 1043.930 847.320 1046.310 849.650 ;
        RECT 1047.150 847.320 1049.530 849.650 ;
        RECT 1050.370 847.320 1052.290 849.650 ;
        RECT 1053.130 847.320 1055.510 849.650 ;
        RECT 1056.350 847.320 1058.730 849.650 ;
        RECT 1059.570 847.320 1061.950 849.650 ;
        RECT 1062.790 847.320 1065.170 849.650 ;
        RECT 1066.010 847.320 1067.930 849.650 ;
        RECT 1068.770 847.320 1071.150 849.650 ;
        RECT 1071.990 847.320 1074.370 849.650 ;
        RECT 1075.210 847.320 1077.590 849.650 ;
        RECT 1078.430 847.320 1080.810 849.650 ;
        RECT 1081.650 847.320 1084.030 849.650 ;
        RECT 1084.870 847.320 1086.790 849.650 ;
        RECT 1087.630 847.320 1090.010 849.650 ;
        RECT 1090.850 847.320 1093.230 849.650 ;
        RECT 1094.070 847.320 1096.450 849.650 ;
        RECT 1097.290 847.320 1099.670 849.650 ;
        RECT 1100.510 847.320 1102.430 849.650 ;
        RECT 1103.270 847.320 1105.650 849.650 ;
        RECT 1106.490 847.320 1108.870 849.650 ;
        RECT 1109.710 847.320 1112.090 849.650 ;
        RECT 1112.930 847.320 1115.310 849.650 ;
        RECT 1116.150 847.320 1118.070 849.650 ;
        RECT 1118.910 847.320 1121.290 849.650 ;
        RECT 1122.130 847.320 1124.510 849.650 ;
        RECT 1125.350 847.320 1127.730 849.650 ;
        RECT 1128.570 847.320 1130.950 849.650 ;
        RECT 1131.790 847.320 1133.710 849.650 ;
        RECT 1134.550 847.320 1136.930 849.650 ;
        RECT 1137.770 847.320 1140.150 849.650 ;
        RECT 1140.990 847.320 1143.370 849.650 ;
        RECT 1144.210 847.320 1146.590 849.650 ;
        RECT 1147.430 847.320 1149.350 849.650 ;
        RECT 1150.190 847.320 1152.570 849.650 ;
        RECT 1153.410 847.320 1155.790 849.650 ;
        RECT 1156.630 847.320 1159.010 849.650 ;
        RECT 1159.850 847.320 1162.230 849.650 ;
        RECT 1163.070 847.320 1164.990 849.650 ;
        RECT 1165.830 847.320 1168.210 849.650 ;
        RECT 1169.050 847.320 1171.430 849.650 ;
        RECT 1172.270 847.320 1174.650 849.650 ;
        RECT 1175.490 847.320 1177.870 849.650 ;
        RECT 1178.710 847.320 1180.630 849.650 ;
        RECT 1181.470 847.320 1183.850 849.650 ;
        RECT 1184.690 847.320 1187.070 849.650 ;
        RECT 1187.910 847.320 1190.290 849.650 ;
        RECT 1191.130 847.320 1193.510 849.650 ;
        RECT 1194.350 847.320 1196.270 849.650 ;
        RECT 1197.110 847.320 1199.490 849.650 ;
        RECT 1200.330 847.320 1202.710 849.650 ;
        RECT 1203.550 847.320 1205.930 849.650 ;
        RECT 1206.770 847.320 1209.150 849.650 ;
        RECT 1209.990 847.320 1211.910 849.650 ;
        RECT 1212.750 847.320 1215.130 849.650 ;
        RECT 1215.970 847.320 1218.350 849.650 ;
        RECT 1219.190 847.320 1221.570 849.650 ;
        RECT 1222.410 847.320 1224.790 849.650 ;
        RECT 1225.630 847.320 1227.550 849.650 ;
        RECT 1228.390 847.320 1230.770 849.650 ;
        RECT 1231.610 847.320 1233.990 849.650 ;
        RECT 1234.830 847.320 1237.210 849.650 ;
        RECT 1238.050 847.320 1240.430 849.650 ;
        RECT 1241.270 847.320 1243.190 849.650 ;
        RECT 1244.030 847.320 1246.410 849.650 ;
        RECT 1247.250 847.320 1249.630 849.650 ;
        RECT 1250.470 847.320 1252.850 849.650 ;
        RECT 1253.690 847.320 1256.070 849.650 ;
        RECT 1256.910 847.320 1259.290 849.650 ;
        RECT 1260.130 847.320 1262.050 849.650 ;
        RECT 1262.890 847.320 1265.270 849.650 ;
        RECT 1266.110 847.320 1268.490 849.650 ;
        RECT 1269.330 847.320 1271.710 849.650 ;
        RECT 1272.550 847.320 1274.930 849.650 ;
        RECT 1275.770 847.320 1277.690 849.650 ;
        RECT 1278.530 847.320 1280.910 849.650 ;
        RECT 1281.750 847.320 1284.130 849.650 ;
        RECT 1284.970 847.320 1287.350 849.650 ;
        RECT 1288.190 847.320 1290.570 849.650 ;
        RECT 1291.410 847.320 1293.330 849.650 ;
        RECT 1294.170 847.320 1296.550 849.650 ;
        RECT 1297.390 847.320 1299.770 849.650 ;
        RECT 1300.610 847.320 1302.990 849.650 ;
        RECT 1303.830 847.320 1306.210 849.650 ;
        RECT 1307.050 847.320 1308.970 849.650 ;
        RECT 1309.810 847.320 1312.190 849.650 ;
        RECT 1313.030 847.320 1315.410 849.650 ;
        RECT 1316.250 847.320 1318.630 849.650 ;
        RECT 1319.470 847.320 1321.850 849.650 ;
        RECT 1322.690 847.320 1324.610 849.650 ;
        RECT 1325.450 847.320 1327.830 849.650 ;
        RECT 1328.670 847.320 1331.050 849.650 ;
        RECT 1331.890 847.320 1334.270 849.650 ;
        RECT 1335.110 847.320 1337.490 849.650 ;
        RECT 1338.330 847.320 1340.250 849.650 ;
        RECT 1341.090 847.320 1343.470 849.650 ;
        RECT 1344.310 847.320 1346.690 849.650 ;
        RECT 1347.530 847.320 1349.910 849.650 ;
        RECT 1350.750 847.320 1353.130 849.650 ;
        RECT 1353.970 847.320 1355.890 849.650 ;
        RECT 1356.730 847.320 1359.110 849.650 ;
        RECT 1359.950 847.320 1362.330 849.650 ;
        RECT 1363.170 847.320 1365.550 849.650 ;
        RECT 1366.390 847.320 1368.770 849.650 ;
        RECT 1369.610 847.320 1371.530 849.650 ;
        RECT 1372.370 847.320 1374.750 849.650 ;
        RECT 1375.590 847.320 1377.970 849.650 ;
        RECT 1378.810 847.320 1381.190 849.650 ;
        RECT 1382.030 847.320 1384.410 849.650 ;
        RECT 1385.250 847.320 1387.170 849.650 ;
        RECT 1388.010 847.320 1390.390 849.650 ;
        RECT 1391.230 847.320 1393.610 849.650 ;
        RECT 1394.450 847.320 1396.830 849.650 ;
        RECT 1397.670 847.320 1400.050 849.650 ;
        RECT 1400.890 847.320 1402.810 849.650 ;
        RECT 1403.650 847.320 1406.030 849.650 ;
        RECT 1406.870 847.320 1409.250 849.650 ;
        RECT 1410.090 847.320 1412.470 849.650 ;
        RECT 1413.310 847.320 1415.690 849.650 ;
        RECT 1416.530 847.320 1418.450 849.650 ;
        RECT 1419.290 847.320 1421.670 849.650 ;
        RECT 1422.510 847.320 1424.890 849.650 ;
        RECT 1425.730 847.320 1428.110 849.650 ;
        RECT 1428.950 847.320 1431.330 849.650 ;
        RECT 1432.170 847.320 1434.550 849.650 ;
        RECT 1435.390 847.320 1437.310 849.650 ;
        RECT 1438.150 847.320 1440.530 849.650 ;
        RECT 1441.370 847.320 1443.750 849.650 ;
        RECT 1444.590 847.320 1446.970 849.650 ;
        RECT 1447.810 847.320 1450.190 849.650 ;
        RECT 1451.030 847.320 1452.950 849.650 ;
        RECT 1453.790 847.320 1456.170 849.650 ;
        RECT 1457.010 847.320 1459.390 849.650 ;
        RECT 1460.230 847.320 1462.610 849.650 ;
        RECT 1463.450 847.320 1465.830 849.650 ;
        RECT 1466.670 847.320 1468.590 849.650 ;
        RECT 1469.430 847.320 1471.810 849.650 ;
        RECT 1472.650 847.320 1475.030 849.650 ;
        RECT 1475.870 847.320 1478.250 849.650 ;
        RECT 1479.090 847.320 1481.470 849.650 ;
        RECT 1482.310 847.320 1484.230 849.650 ;
        RECT 1485.070 847.320 1487.450 849.650 ;
        RECT 1488.290 847.320 1490.670 849.650 ;
        RECT 1491.510 847.320 1493.890 849.650 ;
        RECT 1494.730 847.320 1497.110 849.650 ;
        RECT 1497.950 847.320 1499.870 849.650 ;
        RECT 1500.710 847.320 1503.090 849.650 ;
        RECT 1503.930 847.320 1506.310 849.650 ;
        RECT 1507.150 847.320 1509.530 849.650 ;
        RECT 1510.370 847.320 1512.750 849.650 ;
        RECT 1513.590 847.320 1515.510 849.650 ;
        RECT 1516.350 847.320 1518.730 849.650 ;
        RECT 1519.570 847.320 1521.950 849.650 ;
        RECT 1522.790 847.320 1525.170 849.650 ;
        RECT 1526.010 847.320 1528.390 849.650 ;
        RECT 1529.230 847.320 1531.150 849.650 ;
        RECT 1531.990 847.320 1534.370 849.650 ;
        RECT 1535.210 847.320 1537.590 849.650 ;
        RECT 1538.430 847.320 1540.810 849.650 ;
        RECT 1541.650 847.320 1544.030 849.650 ;
        RECT 1544.870 847.320 1546.790 849.650 ;
        RECT 1547.630 847.320 1550.010 849.650 ;
        RECT 1550.850 847.320 1553.230 849.650 ;
        RECT 1554.070 847.320 1556.450 849.650 ;
        RECT 1557.290 847.320 1559.670 849.650 ;
        RECT 1560.510 847.320 1562.430 849.650 ;
        RECT 1563.270 847.320 1565.650 849.650 ;
        RECT 1566.490 847.320 1568.870 849.650 ;
        RECT 1569.710 847.320 1572.090 849.650 ;
        RECT 1572.930 847.320 1575.310 849.650 ;
        RECT 1576.150 847.320 1578.070 849.650 ;
        RECT 1578.910 847.320 1581.290 849.650 ;
        RECT 1582.130 847.320 1584.510 849.650 ;
        RECT 1585.350 847.320 1587.730 849.650 ;
        RECT 1588.570 847.320 1590.950 849.650 ;
        RECT 1591.790 847.320 1593.710 849.650 ;
        RECT 1594.550 847.320 1596.930 849.650 ;
        RECT 1597.770 847.320 1600.150 849.650 ;
        RECT 1600.990 847.320 1603.370 849.650 ;
        RECT 1604.210 847.320 1606.590 849.650 ;
        RECT 1607.430 847.320 1609.350 849.650 ;
        RECT 1610.190 847.320 1612.570 849.650 ;
        RECT 1613.410 847.320 1615.790 849.650 ;
        RECT 1616.630 847.320 1619.010 849.650 ;
        RECT 1619.850 847.320 1622.230 849.650 ;
        RECT 1623.070 847.320 1625.450 849.650 ;
        RECT 1626.290 847.320 1628.210 849.650 ;
        RECT 1629.050 847.320 1631.430 849.650 ;
        RECT 1632.270 847.320 1634.650 849.650 ;
        RECT 1635.490 847.320 1637.870 849.650 ;
        RECT 1638.710 847.320 1641.090 849.650 ;
        RECT 1641.930 847.320 1643.850 849.650 ;
        RECT 1644.690 847.320 1647.070 849.650 ;
        RECT 1647.910 847.320 1650.290 849.650 ;
        RECT 1651.130 847.320 1653.510 849.650 ;
        RECT 1654.350 847.320 1656.730 849.650 ;
        RECT 1657.570 847.320 1659.490 849.650 ;
        RECT 1660.330 847.320 1662.710 849.650 ;
        RECT 1663.550 847.320 1665.930 849.650 ;
        RECT 1666.770 847.320 1669.150 849.650 ;
        RECT 1669.990 847.320 1672.370 849.650 ;
        RECT 1673.210 847.320 1675.130 849.650 ;
        RECT 1675.970 847.320 1678.350 849.650 ;
        RECT 1679.190 847.320 1681.570 849.650 ;
        RECT 1682.410 847.320 1684.790 849.650 ;
        RECT 1685.630 847.320 1688.010 849.650 ;
        RECT 1688.850 847.320 1690.770 849.650 ;
        RECT 1691.610 847.320 1693.990 849.650 ;
        RECT 1694.830 847.320 1697.210 849.650 ;
        RECT 1698.050 847.320 1700.430 849.650 ;
        RECT 1701.270 847.320 1703.650 849.650 ;
        RECT 1704.490 847.320 1706.410 849.650 ;
        RECT 1707.250 847.320 1709.630 849.650 ;
        RECT 1710.470 847.320 1712.850 849.650 ;
        RECT 1713.690 847.320 1716.070 849.650 ;
        RECT 1716.910 847.320 1719.290 849.650 ;
        RECT 1720.130 847.320 1722.050 849.650 ;
        RECT 1722.890 847.320 1725.270 849.650 ;
        RECT 1726.110 847.320 1728.490 849.650 ;
        RECT 1729.330 847.320 1731.710 849.650 ;
        RECT 1732.550 847.320 1734.930 849.650 ;
        RECT 1735.770 847.320 1737.690 849.650 ;
        RECT 1738.530 847.320 1740.910 849.650 ;
        RECT 1741.750 847.320 1744.130 849.650 ;
        RECT 1744.970 847.320 1747.350 849.650 ;
        RECT 1748.190 847.320 1750.570 849.650 ;
        RECT 1751.410 847.320 1753.330 849.650 ;
        RECT 1754.170 847.320 1756.550 849.650 ;
        RECT 1757.390 847.320 1759.770 849.650 ;
        RECT 1760.610 847.320 1762.990 849.650 ;
        RECT 1763.830 847.320 1766.210 849.650 ;
        RECT 1767.050 847.320 1768.970 849.650 ;
        RECT 1769.810 847.320 1772.190 849.650 ;
        RECT 1773.030 847.320 1775.410 849.650 ;
        RECT 1776.250 847.320 1778.630 849.650 ;
        RECT 1779.470 847.320 1781.850 849.650 ;
        RECT 1782.690 847.320 1784.610 849.650 ;
        RECT 1785.450 847.320 1787.830 849.650 ;
        RECT 1788.670 847.320 1791.050 849.650 ;
        RECT 1791.890 847.320 1794.270 849.650 ;
        RECT 1795.110 847.320 1797.490 849.650 ;
        RECT 1798.330 847.320 1800.710 849.650 ;
        RECT 1801.550 847.320 1803.470 849.650 ;
        RECT 1804.310 847.320 1806.690 849.650 ;
        RECT 1807.530 847.320 1809.910 849.650 ;
        RECT 1810.750 847.320 1813.130 849.650 ;
        RECT 1813.970 847.320 1816.350 849.650 ;
        RECT 1817.190 847.320 1819.110 849.650 ;
        RECT 1819.950 847.320 1822.330 849.650 ;
        RECT 1823.170 847.320 1825.550 849.650 ;
        RECT 1826.390 847.320 1828.770 849.650 ;
        RECT 1829.610 847.320 1831.990 849.650 ;
        RECT 1832.830 847.320 1834.750 849.650 ;
        RECT 1835.590 847.320 1837.970 849.650 ;
        RECT 1838.810 847.320 1841.190 849.650 ;
        RECT 1842.030 847.320 1844.410 849.650 ;
        RECT 1845.250 847.320 1847.630 849.650 ;
        RECT 1848.470 847.320 1850.390 849.650 ;
        RECT 1851.230 847.320 1853.610 849.650 ;
        RECT 1854.450 847.320 1856.830 849.650 ;
        RECT 1857.670 847.320 1860.050 849.650 ;
        RECT 1860.890 847.320 1863.270 849.650 ;
        RECT 1864.110 847.320 1866.030 849.650 ;
        RECT 1866.870 847.320 1869.250 849.650 ;
        RECT 1870.090 847.320 1872.470 849.650 ;
        RECT 1873.310 847.320 1875.690 849.650 ;
        RECT 1876.530 847.320 1878.910 849.650 ;
        RECT 1879.750 847.320 1881.670 849.650 ;
        RECT 1882.510 847.320 1884.890 849.650 ;
        RECT 1885.730 847.320 1888.110 849.650 ;
        RECT 1888.950 847.320 1891.330 849.650 ;
        RECT 1892.170 847.320 1894.550 849.650 ;
        RECT 1895.390 847.320 1897.310 849.650 ;
        RECT 1898.150 847.320 1900.530 849.650 ;
        RECT 1901.370 847.320 1903.750 849.650 ;
        RECT 1904.590 847.320 1906.970 849.650 ;
        RECT 1907.810 847.320 1910.190 849.650 ;
        RECT 1911.030 847.320 1912.950 849.650 ;
        RECT 1913.790 847.320 1916.170 849.650 ;
        RECT 1917.010 847.320 1919.390 849.650 ;
        RECT 1920.230 847.320 1922.610 849.650 ;
        RECT 1923.450 847.320 1925.830 849.650 ;
        RECT 1926.670 847.320 1928.590 849.650 ;
        RECT 1929.430 847.320 1931.810 849.650 ;
        RECT 1932.650 847.320 1935.030 849.650 ;
        RECT 1935.870 847.320 1938.250 849.650 ;
        RECT 1939.090 847.320 1941.470 849.650 ;
        RECT 1942.310 847.320 1944.230 849.650 ;
        RECT 1945.070 847.320 1947.450 849.650 ;
        RECT 1948.290 847.320 1950.670 849.650 ;
        RECT 1951.510 847.320 1953.890 849.650 ;
        RECT 1954.730 847.320 1957.110 849.650 ;
        RECT 1957.950 847.320 1959.870 849.650 ;
        RECT 1960.710 847.320 1963.090 849.650 ;
        RECT 1963.930 847.320 1966.310 849.650 ;
        RECT 1967.150 847.320 1969.530 849.650 ;
        RECT 1970.370 847.320 1972.750 849.650 ;
        RECT 1973.590 847.320 1975.970 849.650 ;
        RECT 1976.810 847.320 1978.730 849.650 ;
        RECT 1979.570 847.320 1981.950 849.650 ;
        RECT 1982.790 847.320 1985.170 849.650 ;
        RECT 1986.010 847.320 1988.390 849.650 ;
        RECT 1989.230 847.320 1991.610 849.650 ;
        RECT 1992.450 847.320 1994.370 849.650 ;
        RECT 1995.210 847.320 1997.590 849.650 ;
        RECT 1998.430 847.320 2000.810 849.650 ;
        RECT 2001.650 847.320 2004.030 849.650 ;
        RECT 2004.870 847.320 2007.250 849.650 ;
        RECT 2008.090 847.320 2010.010 849.650 ;
        RECT 2010.850 847.320 2013.230 849.650 ;
        RECT 2014.070 847.320 2016.450 849.650 ;
        RECT 2017.290 847.320 2019.670 849.650 ;
        RECT 2020.510 847.320 2022.890 849.650 ;
        RECT 2023.730 847.320 2025.650 849.650 ;
        RECT 2026.490 847.320 2028.870 849.650 ;
        RECT 2029.710 847.320 2032.090 849.650 ;
        RECT 2032.930 847.320 2035.310 849.650 ;
        RECT 2036.150 847.320 2038.530 849.650 ;
        RECT 2039.370 847.320 2041.290 849.650 ;
        RECT 2042.130 847.320 2044.510 849.650 ;
        RECT 2045.350 847.320 2047.730 849.650 ;
        RECT 2048.570 847.320 2050.950 849.650 ;
        RECT 2051.790 847.320 2054.170 849.650 ;
        RECT 2055.010 847.320 2056.930 849.650 ;
        RECT 2057.770 847.320 2060.150 849.650 ;
        RECT 2060.990 847.320 2063.370 849.650 ;
        RECT 2064.210 847.320 2066.590 849.650 ;
        RECT 2067.430 847.320 2069.810 849.650 ;
        RECT 2070.650 847.320 2072.570 849.650 ;
        RECT 2073.410 847.320 2075.790 849.650 ;
        RECT 2076.630 847.320 2079.010 849.650 ;
        RECT 2079.850 847.320 2082.230 849.650 ;
        RECT 2083.070 847.320 2085.450 849.650 ;
        RECT 2086.290 847.320 2088.210 849.650 ;
        RECT 2089.050 847.320 2091.430 849.650 ;
        RECT 2092.270 847.320 2094.650 849.650 ;
        RECT 2095.490 847.320 2097.870 849.650 ;
        RECT 2098.710 847.320 2101.090 849.650 ;
        RECT 2101.930 847.320 2103.850 849.650 ;
        RECT 2104.690 847.320 2107.070 849.650 ;
        RECT 2107.910 847.320 2110.290 849.650 ;
        RECT 2111.130 847.320 2113.510 849.650 ;
        RECT 2114.350 847.320 2116.730 849.650 ;
        RECT 2117.570 847.320 2119.490 849.650 ;
        RECT 2120.330 847.320 2122.710 849.650 ;
        RECT 2123.550 847.320 2125.930 849.650 ;
        RECT 2126.770 847.320 2129.150 849.650 ;
        RECT 2129.990 847.320 2132.370 849.650 ;
        RECT 2133.210 847.320 2135.130 849.650 ;
        RECT 2135.970 847.320 2138.350 849.650 ;
        RECT 2139.190 847.320 2141.570 849.650 ;
        RECT 2142.410 847.320 2144.790 849.650 ;
        RECT 2145.630 847.320 2148.010 849.650 ;
        RECT 0.100 2.680 2148.560 847.320 ;
        RECT 0.100 1.515 48.570 2.680 ;
        RECT 49.410 1.515 146.090 2.680 ;
        RECT 146.930 1.515 243.610 2.680 ;
        RECT 244.450 1.515 341.590 2.680 ;
        RECT 342.430 1.515 439.110 2.680 ;
        RECT 439.950 1.515 537.090 2.680 ;
        RECT 537.930 1.515 634.610 2.680 ;
        RECT 635.450 1.515 732.590 2.680 ;
        RECT 733.430 1.515 830.110 2.680 ;
        RECT 830.950 1.515 928.090 2.680 ;
        RECT 928.930 1.515 1025.610 2.680 ;
        RECT 1026.450 1.515 1123.590 2.680 ;
        RECT 1124.430 1.515 1221.110 2.680 ;
        RECT 1221.950 1.515 1318.630 2.680 ;
        RECT 1319.470 1.515 1416.610 2.680 ;
        RECT 1417.450 1.515 1514.130 2.680 ;
        RECT 1514.970 1.515 1612.110 2.680 ;
        RECT 1612.950 1.515 1709.630 2.680 ;
        RECT 1710.470 1.515 1807.610 2.680 ;
        RECT 1808.450 1.515 1905.130 2.680 ;
        RECT 1905.970 1.515 2003.110 2.680 ;
        RECT 2003.950 1.515 2100.630 2.680 ;
        RECT 2101.470 1.515 2148.560 2.680 ;
      LAYER met3 ;
        RECT 2.800 846.920 2147.600 847.785 ;
        RECT 0.270 844.920 2147.600 846.920 ;
        RECT 2.800 843.520 2147.600 844.920 ;
        RECT 0.270 841.520 2147.600 843.520 ;
        RECT 2.800 840.120 2147.600 841.520 ;
        RECT 0.270 838.120 2147.600 840.120 ;
        RECT 2.800 836.720 2147.600 838.120 ;
        RECT 0.270 834.040 2147.600 836.720 ;
        RECT 2.800 832.640 2147.600 834.040 ;
        RECT 0.270 830.640 2147.600 832.640 ;
        RECT 2.800 829.240 2147.600 830.640 ;
        RECT 0.270 827.240 2147.600 829.240 ;
        RECT 2.800 825.840 2147.600 827.240 ;
        RECT 0.270 823.840 2147.600 825.840 ;
        RECT 2.800 822.440 2147.600 823.840 ;
        RECT 0.270 819.760 2147.600 822.440 ;
        RECT 2.800 818.360 2147.600 819.760 ;
        RECT 0.270 816.360 2147.600 818.360 ;
        RECT 2.800 814.960 2147.600 816.360 ;
        RECT 0.270 812.960 2147.600 814.960 ;
        RECT 2.800 811.600 2147.600 812.960 ;
        RECT 2.800 811.560 2147.200 811.600 ;
        RECT 0.270 810.200 2147.200 811.560 ;
        RECT 0.270 809.560 2147.600 810.200 ;
        RECT 2.800 808.160 2147.600 809.560 ;
        RECT 0.270 806.160 2147.600 808.160 ;
        RECT 2.800 804.760 2147.600 806.160 ;
        RECT 0.270 802.080 2147.600 804.760 ;
        RECT 2.800 800.680 2147.600 802.080 ;
        RECT 0.270 798.680 2147.600 800.680 ;
        RECT 2.800 797.280 2147.600 798.680 ;
        RECT 0.270 795.280 2147.600 797.280 ;
        RECT 2.800 793.880 2147.600 795.280 ;
        RECT 0.270 791.880 2147.600 793.880 ;
        RECT 2.800 790.480 2147.600 791.880 ;
        RECT 0.270 787.800 2147.600 790.480 ;
        RECT 2.800 786.400 2147.600 787.800 ;
        RECT 0.270 784.400 2147.600 786.400 ;
        RECT 2.800 783.000 2147.600 784.400 ;
        RECT 0.270 781.000 2147.600 783.000 ;
        RECT 2.800 779.600 2147.600 781.000 ;
        RECT 0.270 777.600 2147.600 779.600 ;
        RECT 2.800 776.200 2147.600 777.600 ;
        RECT 0.270 773.520 2147.600 776.200 ;
        RECT 2.800 772.120 2147.600 773.520 ;
        RECT 0.270 770.120 2147.600 772.120 ;
        RECT 2.800 768.720 2147.600 770.120 ;
        RECT 0.270 766.720 2147.600 768.720 ;
        RECT 2.800 765.320 2147.600 766.720 ;
        RECT 0.270 763.320 2147.600 765.320 ;
        RECT 2.800 761.920 2147.600 763.320 ;
        RECT 0.270 759.920 2147.600 761.920 ;
        RECT 2.800 758.520 2147.600 759.920 ;
        RECT 0.270 755.840 2147.600 758.520 ;
        RECT 2.800 754.440 2147.600 755.840 ;
        RECT 0.270 752.440 2147.600 754.440 ;
        RECT 2.800 751.040 2147.600 752.440 ;
        RECT 0.270 749.040 2147.600 751.040 ;
        RECT 2.800 747.640 2147.600 749.040 ;
        RECT 0.270 745.640 2147.600 747.640 ;
        RECT 2.800 744.240 2147.600 745.640 ;
        RECT 0.270 741.560 2147.600 744.240 ;
        RECT 2.800 740.160 2147.600 741.560 ;
        RECT 0.270 738.160 2147.600 740.160 ;
        RECT 2.800 736.760 2147.600 738.160 ;
        RECT 0.270 734.760 2147.600 736.760 ;
        RECT 2.800 734.080 2147.600 734.760 ;
        RECT 2.800 733.360 2147.200 734.080 ;
        RECT 0.270 732.680 2147.200 733.360 ;
        RECT 0.270 731.360 2147.600 732.680 ;
        RECT 2.800 729.960 2147.600 731.360 ;
        RECT 0.270 727.280 2147.600 729.960 ;
        RECT 2.800 725.880 2147.600 727.280 ;
        RECT 0.270 723.880 2147.600 725.880 ;
        RECT 2.800 722.480 2147.600 723.880 ;
        RECT 0.270 720.480 2147.600 722.480 ;
        RECT 2.800 719.080 2147.600 720.480 ;
        RECT 0.270 717.080 2147.600 719.080 ;
        RECT 2.800 715.680 2147.600 717.080 ;
        RECT 0.270 713.680 2147.600 715.680 ;
        RECT 2.800 712.280 2147.600 713.680 ;
        RECT 0.270 709.600 2147.600 712.280 ;
        RECT 2.800 708.200 2147.600 709.600 ;
        RECT 0.270 706.200 2147.600 708.200 ;
        RECT 2.800 704.800 2147.600 706.200 ;
        RECT 0.270 702.800 2147.600 704.800 ;
        RECT 2.800 701.400 2147.600 702.800 ;
        RECT 0.270 699.400 2147.600 701.400 ;
        RECT 2.800 698.000 2147.600 699.400 ;
        RECT 0.270 695.320 2147.600 698.000 ;
        RECT 2.800 693.920 2147.600 695.320 ;
        RECT 0.270 691.920 2147.600 693.920 ;
        RECT 2.800 690.520 2147.600 691.920 ;
        RECT 0.270 688.520 2147.600 690.520 ;
        RECT 2.800 687.120 2147.600 688.520 ;
        RECT 0.270 685.120 2147.600 687.120 ;
        RECT 2.800 683.720 2147.600 685.120 ;
        RECT 0.270 681.040 2147.600 683.720 ;
        RECT 2.800 679.640 2147.600 681.040 ;
        RECT 0.270 677.640 2147.600 679.640 ;
        RECT 2.800 676.240 2147.600 677.640 ;
        RECT 0.270 674.240 2147.600 676.240 ;
        RECT 2.800 672.840 2147.600 674.240 ;
        RECT 0.270 670.840 2147.600 672.840 ;
        RECT 2.800 669.440 2147.600 670.840 ;
        RECT 0.270 667.440 2147.600 669.440 ;
        RECT 2.800 666.040 2147.600 667.440 ;
        RECT 0.270 663.360 2147.600 666.040 ;
        RECT 2.800 661.960 2147.600 663.360 ;
        RECT 0.270 659.960 2147.600 661.960 ;
        RECT 2.800 658.560 2147.600 659.960 ;
        RECT 0.270 657.240 2147.600 658.560 ;
        RECT 0.270 656.560 2147.200 657.240 ;
        RECT 2.800 655.840 2147.200 656.560 ;
        RECT 2.800 655.160 2147.600 655.840 ;
        RECT 0.270 653.160 2147.600 655.160 ;
        RECT 2.800 651.760 2147.600 653.160 ;
        RECT 0.270 649.080 2147.600 651.760 ;
        RECT 2.800 647.680 2147.600 649.080 ;
        RECT 0.270 645.680 2147.600 647.680 ;
        RECT 2.800 644.280 2147.600 645.680 ;
        RECT 0.270 642.280 2147.600 644.280 ;
        RECT 2.800 640.880 2147.600 642.280 ;
        RECT 0.270 638.880 2147.600 640.880 ;
        RECT 2.800 637.480 2147.600 638.880 ;
        RECT 0.270 634.800 2147.600 637.480 ;
        RECT 2.800 633.400 2147.600 634.800 ;
        RECT 0.270 631.400 2147.600 633.400 ;
        RECT 2.800 630.000 2147.600 631.400 ;
        RECT 0.270 628.000 2147.600 630.000 ;
        RECT 2.800 626.600 2147.600 628.000 ;
        RECT 0.270 624.600 2147.600 626.600 ;
        RECT 2.800 623.200 2147.600 624.600 ;
        RECT 0.270 621.200 2147.600 623.200 ;
        RECT 2.800 619.800 2147.600 621.200 ;
        RECT 0.270 617.120 2147.600 619.800 ;
        RECT 2.800 615.720 2147.600 617.120 ;
        RECT 0.270 613.720 2147.600 615.720 ;
        RECT 2.800 612.320 2147.600 613.720 ;
        RECT 0.270 610.320 2147.600 612.320 ;
        RECT 2.800 608.920 2147.600 610.320 ;
        RECT 0.270 606.920 2147.600 608.920 ;
        RECT 2.800 605.520 2147.600 606.920 ;
        RECT 0.270 602.840 2147.600 605.520 ;
        RECT 2.800 601.440 2147.600 602.840 ;
        RECT 0.270 599.440 2147.600 601.440 ;
        RECT 2.800 598.040 2147.600 599.440 ;
        RECT 0.270 596.040 2147.600 598.040 ;
        RECT 2.800 594.640 2147.600 596.040 ;
        RECT 0.270 592.640 2147.600 594.640 ;
        RECT 2.800 591.240 2147.600 592.640 ;
        RECT 0.270 588.560 2147.600 591.240 ;
        RECT 2.800 587.160 2147.600 588.560 ;
        RECT 0.270 585.160 2147.600 587.160 ;
        RECT 2.800 583.760 2147.600 585.160 ;
        RECT 0.270 581.760 2147.600 583.760 ;
        RECT 2.800 580.360 2147.600 581.760 ;
        RECT 0.270 579.720 2147.600 580.360 ;
        RECT 0.270 578.360 2147.200 579.720 ;
        RECT 2.800 578.320 2147.200 578.360 ;
        RECT 2.800 576.960 2147.600 578.320 ;
        RECT 0.270 574.960 2147.600 576.960 ;
        RECT 2.800 573.560 2147.600 574.960 ;
        RECT 0.270 570.880 2147.600 573.560 ;
        RECT 2.800 569.480 2147.600 570.880 ;
        RECT 0.270 567.480 2147.600 569.480 ;
        RECT 2.800 566.080 2147.600 567.480 ;
        RECT 0.270 564.080 2147.600 566.080 ;
        RECT 2.800 562.680 2147.600 564.080 ;
        RECT 0.270 560.680 2147.600 562.680 ;
        RECT 2.800 559.280 2147.600 560.680 ;
        RECT 0.270 556.600 2147.600 559.280 ;
        RECT 2.800 555.200 2147.600 556.600 ;
        RECT 0.270 553.200 2147.600 555.200 ;
        RECT 2.800 551.800 2147.600 553.200 ;
        RECT 0.270 549.800 2147.600 551.800 ;
        RECT 2.800 548.400 2147.600 549.800 ;
        RECT 0.270 546.400 2147.600 548.400 ;
        RECT 2.800 545.000 2147.600 546.400 ;
        RECT 0.270 542.320 2147.600 545.000 ;
        RECT 2.800 540.920 2147.600 542.320 ;
        RECT 0.270 538.920 2147.600 540.920 ;
        RECT 2.800 537.520 2147.600 538.920 ;
        RECT 0.270 535.520 2147.600 537.520 ;
        RECT 2.800 534.120 2147.600 535.520 ;
        RECT 0.270 532.120 2147.600 534.120 ;
        RECT 2.800 530.720 2147.600 532.120 ;
        RECT 0.270 528.720 2147.600 530.720 ;
        RECT 2.800 527.320 2147.600 528.720 ;
        RECT 0.270 524.640 2147.600 527.320 ;
        RECT 2.800 523.240 2147.600 524.640 ;
        RECT 0.270 521.240 2147.600 523.240 ;
        RECT 2.800 519.840 2147.600 521.240 ;
        RECT 0.270 517.840 2147.600 519.840 ;
        RECT 2.800 516.440 2147.600 517.840 ;
        RECT 0.270 514.440 2147.600 516.440 ;
        RECT 2.800 513.040 2147.600 514.440 ;
        RECT 0.270 510.360 2147.600 513.040 ;
        RECT 2.800 508.960 2147.600 510.360 ;
        RECT 0.270 506.960 2147.600 508.960 ;
        RECT 2.800 505.560 2147.600 506.960 ;
        RECT 0.270 503.560 2147.600 505.560 ;
        RECT 2.800 502.200 2147.600 503.560 ;
        RECT 2.800 502.160 2147.200 502.200 ;
        RECT 0.270 500.800 2147.200 502.160 ;
        RECT 0.270 500.160 2147.600 500.800 ;
        RECT 2.800 498.760 2147.600 500.160 ;
        RECT 0.270 496.080 2147.600 498.760 ;
        RECT 2.800 494.680 2147.600 496.080 ;
        RECT 0.270 492.680 2147.600 494.680 ;
        RECT 2.800 491.280 2147.600 492.680 ;
        RECT 0.270 489.280 2147.600 491.280 ;
        RECT 2.800 487.880 2147.600 489.280 ;
        RECT 0.270 485.880 2147.600 487.880 ;
        RECT 2.800 484.480 2147.600 485.880 ;
        RECT 0.270 482.480 2147.600 484.480 ;
        RECT 2.800 481.080 2147.600 482.480 ;
        RECT 0.270 478.400 2147.600 481.080 ;
        RECT 2.800 477.000 2147.600 478.400 ;
        RECT 0.270 475.000 2147.600 477.000 ;
        RECT 2.800 473.600 2147.600 475.000 ;
        RECT 0.270 471.600 2147.600 473.600 ;
        RECT 2.800 470.200 2147.600 471.600 ;
        RECT 0.270 468.200 2147.600 470.200 ;
        RECT 2.800 466.800 2147.600 468.200 ;
        RECT 0.270 464.120 2147.600 466.800 ;
        RECT 2.800 462.720 2147.600 464.120 ;
        RECT 0.270 460.720 2147.600 462.720 ;
        RECT 2.800 459.320 2147.600 460.720 ;
        RECT 0.270 457.320 2147.600 459.320 ;
        RECT 2.800 455.920 2147.600 457.320 ;
        RECT 0.270 453.920 2147.600 455.920 ;
        RECT 2.800 452.520 2147.600 453.920 ;
        RECT 0.270 449.840 2147.600 452.520 ;
        RECT 2.800 448.440 2147.600 449.840 ;
        RECT 0.270 446.440 2147.600 448.440 ;
        RECT 2.800 445.040 2147.600 446.440 ;
        RECT 0.270 443.040 2147.600 445.040 ;
        RECT 2.800 441.640 2147.600 443.040 ;
        RECT 0.270 439.640 2147.600 441.640 ;
        RECT 2.800 438.240 2147.600 439.640 ;
        RECT 0.270 436.240 2147.600 438.240 ;
        RECT 2.800 434.840 2147.600 436.240 ;
        RECT 0.270 432.160 2147.600 434.840 ;
        RECT 2.800 430.760 2147.600 432.160 ;
        RECT 0.270 428.760 2147.600 430.760 ;
        RECT 2.800 427.360 2147.600 428.760 ;
        RECT 0.270 425.360 2147.600 427.360 ;
        RECT 2.800 423.960 2147.200 425.360 ;
        RECT 0.270 421.960 2147.600 423.960 ;
        RECT 2.800 420.560 2147.600 421.960 ;
        RECT 0.270 417.880 2147.600 420.560 ;
        RECT 2.800 416.480 2147.600 417.880 ;
        RECT 0.270 414.480 2147.600 416.480 ;
        RECT 2.800 413.080 2147.600 414.480 ;
        RECT 0.270 411.080 2147.600 413.080 ;
        RECT 2.800 409.680 2147.600 411.080 ;
        RECT 0.270 407.680 2147.600 409.680 ;
        RECT 2.800 406.280 2147.600 407.680 ;
        RECT 0.270 404.280 2147.600 406.280 ;
        RECT 2.800 402.880 2147.600 404.280 ;
        RECT 0.270 400.200 2147.600 402.880 ;
        RECT 2.800 398.800 2147.600 400.200 ;
        RECT 0.270 396.800 2147.600 398.800 ;
        RECT 2.800 395.400 2147.600 396.800 ;
        RECT 0.270 393.400 2147.600 395.400 ;
        RECT 2.800 392.000 2147.600 393.400 ;
        RECT 0.270 390.000 2147.600 392.000 ;
        RECT 2.800 388.600 2147.600 390.000 ;
        RECT 0.270 385.920 2147.600 388.600 ;
        RECT 2.800 384.520 2147.600 385.920 ;
        RECT 0.270 382.520 2147.600 384.520 ;
        RECT 2.800 381.120 2147.600 382.520 ;
        RECT 0.270 379.120 2147.600 381.120 ;
        RECT 2.800 377.720 2147.600 379.120 ;
        RECT 0.270 375.720 2147.600 377.720 ;
        RECT 2.800 374.320 2147.600 375.720 ;
        RECT 0.270 371.640 2147.600 374.320 ;
        RECT 2.800 370.240 2147.600 371.640 ;
        RECT 0.270 368.240 2147.600 370.240 ;
        RECT 2.800 366.840 2147.600 368.240 ;
        RECT 0.270 364.840 2147.600 366.840 ;
        RECT 2.800 363.440 2147.600 364.840 ;
        RECT 0.270 361.440 2147.600 363.440 ;
        RECT 2.800 360.040 2147.600 361.440 ;
        RECT 0.270 358.040 2147.600 360.040 ;
        RECT 2.800 356.640 2147.600 358.040 ;
        RECT 0.270 353.960 2147.600 356.640 ;
        RECT 2.800 352.560 2147.600 353.960 ;
        RECT 0.270 350.560 2147.600 352.560 ;
        RECT 2.800 349.160 2147.600 350.560 ;
        RECT 0.270 347.840 2147.600 349.160 ;
        RECT 0.270 347.160 2147.200 347.840 ;
        RECT 2.800 346.440 2147.200 347.160 ;
        RECT 2.800 345.760 2147.600 346.440 ;
        RECT 0.270 343.760 2147.600 345.760 ;
        RECT 2.800 342.360 2147.600 343.760 ;
        RECT 0.270 339.680 2147.600 342.360 ;
        RECT 2.800 338.280 2147.600 339.680 ;
        RECT 0.270 336.280 2147.600 338.280 ;
        RECT 2.800 334.880 2147.600 336.280 ;
        RECT 0.270 332.880 2147.600 334.880 ;
        RECT 2.800 331.480 2147.600 332.880 ;
        RECT 0.270 329.480 2147.600 331.480 ;
        RECT 2.800 328.080 2147.600 329.480 ;
        RECT 0.270 325.400 2147.600 328.080 ;
        RECT 2.800 324.000 2147.600 325.400 ;
        RECT 0.270 322.000 2147.600 324.000 ;
        RECT 2.800 320.600 2147.600 322.000 ;
        RECT 0.270 318.600 2147.600 320.600 ;
        RECT 2.800 317.200 2147.600 318.600 ;
        RECT 0.270 315.200 2147.600 317.200 ;
        RECT 2.800 313.800 2147.600 315.200 ;
        RECT 0.270 311.800 2147.600 313.800 ;
        RECT 2.800 310.400 2147.600 311.800 ;
        RECT 0.270 307.720 2147.600 310.400 ;
        RECT 2.800 306.320 2147.600 307.720 ;
        RECT 0.270 304.320 2147.600 306.320 ;
        RECT 2.800 302.920 2147.600 304.320 ;
        RECT 0.270 300.920 2147.600 302.920 ;
        RECT 2.800 299.520 2147.600 300.920 ;
        RECT 0.270 297.520 2147.600 299.520 ;
        RECT 2.800 296.120 2147.600 297.520 ;
        RECT 0.270 293.440 2147.600 296.120 ;
        RECT 2.800 292.040 2147.600 293.440 ;
        RECT 0.270 290.040 2147.600 292.040 ;
        RECT 2.800 288.640 2147.600 290.040 ;
        RECT 0.270 286.640 2147.600 288.640 ;
        RECT 2.800 285.240 2147.600 286.640 ;
        RECT 0.270 283.240 2147.600 285.240 ;
        RECT 2.800 281.840 2147.600 283.240 ;
        RECT 0.270 279.160 2147.600 281.840 ;
        RECT 2.800 277.760 2147.600 279.160 ;
        RECT 0.270 275.760 2147.600 277.760 ;
        RECT 2.800 274.360 2147.600 275.760 ;
        RECT 0.270 272.360 2147.600 274.360 ;
        RECT 2.800 270.960 2147.600 272.360 ;
        RECT 0.270 270.320 2147.600 270.960 ;
        RECT 0.270 268.960 2147.200 270.320 ;
        RECT 2.800 268.920 2147.200 268.960 ;
        RECT 2.800 267.560 2147.600 268.920 ;
        RECT 0.270 265.560 2147.600 267.560 ;
        RECT 2.800 264.160 2147.600 265.560 ;
        RECT 0.270 261.480 2147.600 264.160 ;
        RECT 2.800 260.080 2147.600 261.480 ;
        RECT 0.270 258.080 2147.600 260.080 ;
        RECT 2.800 256.680 2147.600 258.080 ;
        RECT 0.270 254.680 2147.600 256.680 ;
        RECT 2.800 253.280 2147.600 254.680 ;
        RECT 0.270 251.280 2147.600 253.280 ;
        RECT 2.800 249.880 2147.600 251.280 ;
        RECT 0.270 247.200 2147.600 249.880 ;
        RECT 2.800 245.800 2147.600 247.200 ;
        RECT 0.270 243.800 2147.600 245.800 ;
        RECT 2.800 242.400 2147.600 243.800 ;
        RECT 0.270 240.400 2147.600 242.400 ;
        RECT 2.800 239.000 2147.600 240.400 ;
        RECT 0.270 237.000 2147.600 239.000 ;
        RECT 2.800 235.600 2147.600 237.000 ;
        RECT 0.270 232.920 2147.600 235.600 ;
        RECT 2.800 231.520 2147.600 232.920 ;
        RECT 0.270 229.520 2147.600 231.520 ;
        RECT 2.800 228.120 2147.600 229.520 ;
        RECT 0.270 226.120 2147.600 228.120 ;
        RECT 2.800 224.720 2147.600 226.120 ;
        RECT 0.270 222.720 2147.600 224.720 ;
        RECT 2.800 221.320 2147.600 222.720 ;
        RECT 0.270 219.320 2147.600 221.320 ;
        RECT 2.800 217.920 2147.600 219.320 ;
        RECT 0.270 215.240 2147.600 217.920 ;
        RECT 2.800 213.840 2147.600 215.240 ;
        RECT 0.270 211.840 2147.600 213.840 ;
        RECT 2.800 210.440 2147.600 211.840 ;
        RECT 0.270 208.440 2147.600 210.440 ;
        RECT 2.800 207.040 2147.600 208.440 ;
        RECT 0.270 205.040 2147.600 207.040 ;
        RECT 2.800 203.640 2147.600 205.040 ;
        RECT 0.270 200.960 2147.600 203.640 ;
        RECT 2.800 199.560 2147.600 200.960 ;
        RECT 0.270 197.560 2147.600 199.560 ;
        RECT 2.800 196.160 2147.600 197.560 ;
        RECT 0.270 194.160 2147.600 196.160 ;
        RECT 2.800 193.480 2147.600 194.160 ;
        RECT 2.800 192.760 2147.200 193.480 ;
        RECT 0.270 192.080 2147.200 192.760 ;
        RECT 0.270 190.760 2147.600 192.080 ;
        RECT 2.800 189.360 2147.600 190.760 ;
        RECT 0.270 186.680 2147.600 189.360 ;
        RECT 2.800 185.280 2147.600 186.680 ;
        RECT 0.270 183.280 2147.600 185.280 ;
        RECT 2.800 181.880 2147.600 183.280 ;
        RECT 0.270 179.880 2147.600 181.880 ;
        RECT 2.800 178.480 2147.600 179.880 ;
        RECT 0.270 176.480 2147.600 178.480 ;
        RECT 2.800 175.080 2147.600 176.480 ;
        RECT 0.270 173.080 2147.600 175.080 ;
        RECT 2.800 171.680 2147.600 173.080 ;
        RECT 0.270 169.000 2147.600 171.680 ;
        RECT 2.800 167.600 2147.600 169.000 ;
        RECT 0.270 165.600 2147.600 167.600 ;
        RECT 2.800 164.200 2147.600 165.600 ;
        RECT 0.270 162.200 2147.600 164.200 ;
        RECT 2.800 160.800 2147.600 162.200 ;
        RECT 0.270 158.800 2147.600 160.800 ;
        RECT 2.800 157.400 2147.600 158.800 ;
        RECT 0.270 154.720 2147.600 157.400 ;
        RECT 2.800 153.320 2147.600 154.720 ;
        RECT 0.270 151.320 2147.600 153.320 ;
        RECT 2.800 149.920 2147.600 151.320 ;
        RECT 0.270 147.920 2147.600 149.920 ;
        RECT 2.800 146.520 2147.600 147.920 ;
        RECT 0.270 144.520 2147.600 146.520 ;
        RECT 2.800 143.120 2147.600 144.520 ;
        RECT 0.270 140.440 2147.600 143.120 ;
        RECT 2.800 139.040 2147.600 140.440 ;
        RECT 0.270 137.040 2147.600 139.040 ;
        RECT 2.800 135.640 2147.600 137.040 ;
        RECT 0.270 133.640 2147.600 135.640 ;
        RECT 2.800 132.240 2147.600 133.640 ;
        RECT 0.270 130.240 2147.600 132.240 ;
        RECT 2.800 128.840 2147.600 130.240 ;
        RECT 0.270 126.840 2147.600 128.840 ;
        RECT 2.800 125.440 2147.600 126.840 ;
        RECT 0.270 122.760 2147.600 125.440 ;
        RECT 2.800 121.360 2147.600 122.760 ;
        RECT 0.270 119.360 2147.600 121.360 ;
        RECT 2.800 117.960 2147.600 119.360 ;
        RECT 0.270 115.960 2147.600 117.960 ;
        RECT 2.800 114.560 2147.200 115.960 ;
        RECT 0.270 112.560 2147.600 114.560 ;
        RECT 2.800 111.160 2147.600 112.560 ;
        RECT 0.270 108.480 2147.600 111.160 ;
        RECT 2.800 107.080 2147.600 108.480 ;
        RECT 0.270 105.080 2147.600 107.080 ;
        RECT 2.800 103.680 2147.600 105.080 ;
        RECT 0.270 101.680 2147.600 103.680 ;
        RECT 2.800 100.280 2147.600 101.680 ;
        RECT 0.270 98.280 2147.600 100.280 ;
        RECT 2.800 96.880 2147.600 98.280 ;
        RECT 0.270 94.200 2147.600 96.880 ;
        RECT 2.800 92.800 2147.600 94.200 ;
        RECT 0.270 90.800 2147.600 92.800 ;
        RECT 2.800 89.400 2147.600 90.800 ;
        RECT 0.270 87.400 2147.600 89.400 ;
        RECT 2.800 86.000 2147.600 87.400 ;
        RECT 0.270 84.000 2147.600 86.000 ;
        RECT 2.800 82.600 2147.600 84.000 ;
        RECT 0.270 80.600 2147.600 82.600 ;
        RECT 2.800 79.200 2147.600 80.600 ;
        RECT 0.270 76.520 2147.600 79.200 ;
        RECT 2.800 75.120 2147.600 76.520 ;
        RECT 0.270 73.120 2147.600 75.120 ;
        RECT 2.800 71.720 2147.600 73.120 ;
        RECT 0.270 69.720 2147.600 71.720 ;
        RECT 2.800 68.320 2147.600 69.720 ;
        RECT 0.270 66.320 2147.600 68.320 ;
        RECT 2.800 64.920 2147.600 66.320 ;
        RECT 0.270 62.240 2147.600 64.920 ;
        RECT 2.800 60.840 2147.600 62.240 ;
        RECT 0.270 58.840 2147.600 60.840 ;
        RECT 2.800 57.440 2147.600 58.840 ;
        RECT 0.270 55.440 2147.600 57.440 ;
        RECT 2.800 54.040 2147.600 55.440 ;
        RECT 0.270 52.040 2147.600 54.040 ;
        RECT 2.800 50.640 2147.600 52.040 ;
        RECT 0.270 47.960 2147.600 50.640 ;
        RECT 2.800 46.560 2147.600 47.960 ;
        RECT 0.270 44.560 2147.600 46.560 ;
        RECT 2.800 43.160 2147.600 44.560 ;
        RECT 0.270 41.160 2147.600 43.160 ;
        RECT 2.800 39.760 2147.600 41.160 ;
        RECT 0.270 39.120 2147.600 39.760 ;
        RECT 0.270 37.760 2147.200 39.120 ;
        RECT 2.800 37.720 2147.200 37.760 ;
        RECT 2.800 36.360 2147.600 37.720 ;
        RECT 0.270 34.360 2147.600 36.360 ;
        RECT 2.800 32.960 2147.600 34.360 ;
        RECT 0.270 30.280 2147.600 32.960 ;
        RECT 2.800 28.880 2147.600 30.280 ;
        RECT 0.270 26.880 2147.600 28.880 ;
        RECT 2.800 25.480 2147.600 26.880 ;
        RECT 0.270 23.480 2147.600 25.480 ;
        RECT 2.800 22.080 2147.600 23.480 ;
        RECT 0.270 20.080 2147.600 22.080 ;
        RECT 2.800 18.680 2147.600 20.080 ;
        RECT 0.270 16.000 2147.600 18.680 ;
        RECT 2.800 14.600 2147.600 16.000 ;
        RECT 0.270 12.600 2147.600 14.600 ;
        RECT 2.800 11.200 2147.600 12.600 ;
        RECT 0.270 9.200 2147.600 11.200 ;
        RECT 2.800 7.800 2147.600 9.200 ;
        RECT 0.270 5.800 2147.600 7.800 ;
        RECT 2.800 4.400 2147.600 5.800 ;
        RECT 0.270 2.400 2147.600 4.400 ;
        RECT 2.800 1.535 2147.600 2.400 ;
      LAYER met4 ;
        RECT 0.295 10.640 2122.640 839.625 ;
      LAYER met5 ;
        RECT 5.520 179.670 2144.060 793.990 ;
  END
END mgmt_core
END LIBRARY

