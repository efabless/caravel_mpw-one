magic
tech sky130A
magscale 1 2
timestamp 1624038509
<< nwell >>
rect 335772 997737 347593 998041
rect 577972 997737 589793 998041
rect 39559 872172 39863 883993
rect 39559 829972 39863 841793
rect 677737 819207 678041 831028
rect 677737 504607 678041 516428
rect 39559 485372 39863 497193
rect 677737 416407 678041 428228
rect 39559 112572 39863 124393
rect 79607 39559 91428 39863
rect 569807 39559 581628 39863
rect 623607 39559 635428 39863
<< pwell >>
rect 35242 870499 39813 872057
rect 677787 831143 682358 832701
rect 677787 516543 682358 518101
rect 35242 483699 39813 485257
rect 35242 110899 39813 112457
rect 635543 35242 637101 39813
<< obsli1 >>
rect 76168 997646 92232 1037541
rect 127568 997646 143632 1037541
rect 178968 997646 195032 1037541
rect 230368 997646 246432 1037541
rect 281968 997646 298032 1037541
rect 333614 998007 347955 1037539
rect 335813 997978 336009 998007
rect 347352 997978 347530 998007
rect 335813 997800 347530 997978
rect 383768 997646 399832 1037541
rect 472768 997646 488832 1037541
rect 524168 997646 540232 1037541
rect 575814 998007 590155 1037539
rect 578013 997978 578209 998007
rect 589552 997978 589730 998007
rect 578013 997800 589730 997978
rect 625968 997646 642032 1037541
rect 59 954168 39954 970232
rect 677646 951568 717541 967632
rect 44 912048 39396 926951
rect 678204 907649 717556 922552
rect 61 883936 39593 884371
rect 61 883746 39806 883936
rect 61 872409 39593 883746
rect 39616 872409 39806 883746
rect 61 872207 39806 872409
rect 61 872031 39593 872207
rect 61 869922 39787 872031
rect 677646 862368 717541 878432
rect 61 841730 39593 842155
rect 61 841552 39800 841730
rect 61 830209 39593 841552
rect 39622 830209 39800 841552
rect 677813 831169 717539 833278
rect 678007 830993 717539 831169
rect 61 830013 39800 830209
rect 677794 830791 717539 830993
rect 61 827814 39593 830013
rect 677794 819454 677984 830791
rect 678007 819454 717539 830791
rect 677794 819264 717539 819454
rect 678007 818829 717539 819264
rect 59 784368 39954 800432
rect 677646 773168 717541 789232
rect 59 741168 39954 757232
rect 677646 728168 717541 744232
rect 59 697968 39954 714032
rect 677646 683168 717541 699232
rect 59 654768 39954 670832
rect 677646 637968 717541 654032
rect 59 611568 39954 627632
rect 677646 592968 717541 609032
rect 59 568368 39954 584432
rect 677646 547768 717541 563832
rect 59 525168 39954 541232
rect 677813 516569 717539 518678
rect 678007 516393 717539 516569
rect 677794 516191 717539 516393
rect 677794 504854 677984 516191
rect 678007 504854 717539 516191
rect 677794 504664 717539 504854
rect 678007 504229 717539 504664
rect 61 497136 39593 497571
rect 61 496946 39806 497136
rect 61 485609 39593 496946
rect 39616 485609 39806 496946
rect 61 485407 39806 485609
rect 61 485231 39593 485407
rect 61 483122 39787 485231
rect 678204 459849 717556 474752
rect 44 440848 39396 455751
rect 678007 428187 717539 430386
rect 677800 427991 717539 428187
rect 677800 416648 677978 427991
rect 678007 416648 717539 427991
rect 677800 416470 717539 416648
rect 678007 416045 717539 416470
rect 59 397568 39954 413632
rect 677646 370568 717541 386632
rect 59 354368 39954 370432
rect 59 311168 39954 327232
rect 677646 325368 717541 341432
rect 59 267968 39954 284032
rect 677646 280368 717541 296432
rect 59 224768 39954 240832
rect 677646 235368 717541 251432
rect 59 181568 39954 197632
rect 677646 190168 717541 206232
rect 677646 145168 717541 161232
rect 61 124336 39593 124771
rect 61 124146 39806 124336
rect 61 112809 39593 124146
rect 39616 112809 39806 124146
rect 61 112607 39806 112809
rect 61 112431 39593 112607
rect 61 110322 39787 112431
rect 677646 99968 717541 116032
rect 44 68048 39396 82951
rect 79670 39622 91387 39800
rect 79670 39593 79848 39622
rect 91191 39593 91387 39622
rect 79245 61 93586 39593
rect 132600 156 147600 39963
rect 186368 59 202432 39954
rect 241249 44 256152 39396
rect 294968 59 311032 39954
rect 349768 59 365832 39954
rect 404568 59 420632 39954
rect 459368 59 475432 39954
rect 514168 59 530232 39954
rect 569870 39622 581587 39800
rect 569870 39593 570048 39622
rect 581391 39593 581587 39622
rect 623664 39616 635393 39806
rect 623664 39593 623854 39616
rect 635191 39593 635393 39616
rect 635569 39593 637678 39787
rect 569445 61 583786 39593
rect 623229 61 637678 39593
<< metal1 >>
rect 78858 990564 78864 990616
rect 78916 990604 78922 990616
rect 83182 990604 83188 990616
rect 78916 990576 83188 990604
rect 78916 990564 78922 990576
rect 83182 990564 83188 990576
rect 83240 990604 83246 990616
rect 130286 990604 130292 990616
rect 83240 990576 130292 990604
rect 83240 990564 83246 990576
rect 130286 990564 130292 990576
rect 130344 990604 130350 990616
rect 134610 990604 134616 990616
rect 130344 990576 134616 990604
rect 130344 990564 130350 990576
rect 134610 990564 134616 990576
rect 134668 990604 134674 990616
rect 181714 990604 181720 990616
rect 134668 990576 181720 990604
rect 134668 990564 134674 990576
rect 181714 990564 181720 990576
rect 181772 990604 181778 990616
rect 186038 990604 186044 990616
rect 181772 990576 186044 990604
rect 181772 990564 181778 990576
rect 186038 990564 186044 990576
rect 186096 990604 186102 990616
rect 233050 990604 233056 990616
rect 186096 990576 233056 990604
rect 186096 990564 186102 990576
rect 233050 990564 233056 990576
rect 233108 990604 233114 990616
rect 237374 990604 237380 990616
rect 233108 990576 237380 990604
rect 233108 990564 233114 990576
rect 237374 990564 237380 990576
rect 237432 990604 237438 990616
rect 274450 990604 274456 990616
rect 237432 990576 274456 990604
rect 237432 990564 237438 990576
rect 274450 990564 274456 990576
rect 274508 990564 274514 990616
rect 274726 990632 274732 990684
rect 274784 990672 274790 990684
rect 284662 990672 284668 990684
rect 274784 990644 284668 990672
rect 274784 990632 274790 990644
rect 284662 990632 284668 990644
rect 284720 990672 284726 990684
rect 288986 990672 288992 990684
rect 284720 990644 288992 990672
rect 284720 990632 284726 990644
rect 288986 990632 288992 990644
rect 289044 990672 289050 990684
rect 289044 990644 386552 990672
rect 289044 990632 289050 990644
rect 386524 990616 386552 990644
rect 386506 990564 386512 990616
rect 386564 990604 386570 990616
rect 390830 990604 390836 990616
rect 386564 990576 390836 990604
rect 386564 990564 386570 990576
rect 390830 990564 390836 990576
rect 390888 990604 390894 990616
rect 475470 990604 475476 990616
rect 390888 990576 475476 990604
rect 390888 990564 390894 990576
rect 475470 990564 475476 990576
rect 475528 990604 475534 990616
rect 479794 990604 479800 990616
rect 475528 990576 479800 990604
rect 475528 990564 475534 990576
rect 479794 990564 479800 990576
rect 479852 990604 479858 990616
rect 526898 990604 526904 990616
rect 479852 990576 526904 990604
rect 479852 990564 479858 990576
rect 526898 990564 526904 990576
rect 526956 990604 526962 990616
rect 531222 990604 531228 990616
rect 526956 990576 531228 990604
rect 526956 990564 526962 990576
rect 531222 990564 531228 990576
rect 531280 990604 531286 990616
rect 628650 990604 628656 990616
rect 531280 990576 628656 990604
rect 531280 990564 531286 990576
rect 628650 990564 628656 990576
rect 628708 990604 628714 990616
rect 632974 990604 632980 990616
rect 628708 990576 632980 990604
rect 628708 990564 628714 990576
rect 632974 990564 632980 990576
rect 633032 990604 633038 990616
rect 634722 990604 634728 990616
rect 633032 990576 634728 990604
rect 633032 990564 633038 990576
rect 634722 990564 634728 990576
rect 634780 990564 634786 990616
rect 42334 990224 42340 990276
rect 42392 990264 42398 990276
rect 78858 990264 78864 990276
rect 42392 990236 78864 990264
rect 42392 990224 42398 990236
rect 78858 990224 78864 990236
rect 78916 990224 78922 990276
rect 634722 990088 634728 990140
rect 634780 990128 634786 990140
rect 673822 990128 673828 990140
rect 634780 990100 673828 990128
rect 634780 990088 634786 990100
rect 673822 990088 673828 990100
rect 673880 990088 673886 990140
rect 673822 965268 673828 965320
rect 673880 965308 673886 965320
rect 675386 965308 675392 965320
rect 673880 965280 675392 965308
rect 673880 965268 673886 965280
rect 675386 965268 675392 965280
rect 675444 965268 675450 965320
rect 41782 961120 41788 961172
rect 41840 961160 41846 961172
rect 42518 961160 42524 961172
rect 41840 961132 42524 961160
rect 41840 961120 41846 961132
rect 42518 961120 42524 961132
rect 42576 961120 42582 961172
rect 673638 960032 673644 960084
rect 673696 960072 673702 960084
rect 675386 960072 675392 960084
rect 673696 960044 675392 960072
rect 673696 960032 673702 960044
rect 675386 960032 675392 960044
rect 675444 960032 675450 960084
rect 673638 875780 673644 875832
rect 673696 875820 673702 875832
rect 675386 875820 675392 875832
rect 673696 875792 675392 875820
rect 673696 875780 673702 875792
rect 675386 875780 675392 875792
rect 675444 875780 675450 875832
rect 673822 871292 673828 871344
rect 673880 871332 673886 871344
rect 675294 871332 675300 871344
rect 673880 871304 675300 871332
rect 673880 871292 673886 871304
rect 675294 871292 675300 871304
rect 675352 871292 675358 871344
rect 41782 791936 41788 791988
rect 41840 791976 41846 791988
rect 42518 791976 42524 791988
rect 41840 791948 42524 791976
rect 41840 791936 41846 791948
rect 42518 791936 42524 791948
rect 42576 791936 42582 791988
rect 41782 786972 41788 787024
rect 41840 787012 41846 787024
rect 42426 787012 42432 787024
rect 41840 786984 42432 787012
rect 41840 786972 41846 786984
rect 42426 786972 42432 786984
rect 42484 786972 42490 787024
rect 673822 785952 673828 786004
rect 673880 785992 673886 786004
rect 675202 785992 675208 786004
rect 673880 785964 675208 785992
rect 673880 785952 673886 785964
rect 675202 785952 675208 785964
rect 675260 785992 675266 786004
rect 675386 785992 675392 786004
rect 675260 785964 675392 785992
rect 675260 785952 675266 785964
rect 675386 785952 675392 785964
rect 675444 785952 675450 786004
rect 673730 781600 673736 781652
rect 673788 781640 673794 781652
rect 675202 781640 675208 781652
rect 673788 781612 675208 781640
rect 673788 781600 673794 781612
rect 675202 781600 675208 781612
rect 675260 781640 675266 781652
rect 675386 781640 675392 781652
rect 675260 781612 675392 781640
rect 675260 781600 675266 781612
rect 675386 781600 675392 781612
rect 675444 781600 675450 781652
rect 42426 756576 42432 756628
rect 42484 756576 42490 756628
rect 42444 756424 42472 756576
rect 42426 756372 42432 756424
rect 42484 756372 42490 756424
rect 41966 747872 41972 747924
rect 42024 747912 42030 747924
rect 42334 747912 42340 747924
rect 42024 747884 42340 747912
rect 42024 747872 42030 747884
rect 42334 747872 42340 747884
rect 42392 747872 42398 747924
rect 41782 743452 41788 743504
rect 41840 743492 41846 743504
rect 42334 743492 42340 743504
rect 41840 743464 42340 743492
rect 41840 743452 41846 743464
rect 42334 743452 42340 743464
rect 42392 743452 42398 743504
rect 673730 740936 673736 740988
rect 673788 740976 673794 740988
rect 675202 740976 675208 740988
rect 673788 740948 675208 740976
rect 673788 740936 673794 740948
rect 675202 740936 675208 740948
rect 675260 740976 675266 740988
rect 675386 740976 675392 740988
rect 675260 740948 675392 740976
rect 675260 740936 675266 740948
rect 675386 740936 675392 740948
rect 675444 740936 675450 740988
rect 673730 736992 673736 737044
rect 673788 737032 673794 737044
rect 675202 737032 675208 737044
rect 673788 737004 675208 737032
rect 673788 736992 673794 737004
rect 675202 736992 675208 737004
rect 675260 737032 675266 737044
rect 675386 737032 675392 737044
rect 675260 737004 675392 737032
rect 675260 736992 675266 737004
rect 675386 736992 675392 737004
rect 675444 736992 675450 737044
rect 42334 719040 42340 719092
rect 42392 719040 42398 719092
rect 42352 718888 42380 719040
rect 42334 718836 42340 718888
rect 42392 718836 42398 718888
rect 673730 695920 673736 695972
rect 673788 695960 673794 695972
rect 675202 695960 675208 695972
rect 673788 695932 675208 695960
rect 673788 695920 673794 695932
rect 675202 695920 675208 695932
rect 675260 695960 675266 695972
rect 675386 695960 675392 695972
rect 675260 695932 675392 695960
rect 675260 695920 675266 695932
rect 675386 695920 675392 695932
rect 675444 695920 675450 695972
rect 673730 692044 673736 692096
rect 673788 692084 673794 692096
rect 675202 692084 675208 692096
rect 673788 692056 675208 692084
rect 673788 692044 673794 692056
rect 675202 692044 675208 692056
rect 675260 692084 675266 692096
rect 675386 692084 675392 692096
rect 675260 692056 675392 692084
rect 675260 692044 675266 692056
rect 675386 692044 675392 692056
rect 675444 692044 675450 692096
rect 673730 651108 673736 651160
rect 673788 651148 673794 651160
rect 675386 651148 675392 651160
rect 673788 651120 675392 651148
rect 673788 651108 673794 651120
rect 675386 651108 675392 651120
rect 675444 651108 675450 651160
rect 673730 646416 673736 646468
rect 673788 646456 673794 646468
rect 675386 646456 675392 646468
rect 673788 646428 675392 646456
rect 673788 646416 673794 646428
rect 675386 646416 675392 646428
rect 675444 646416 675450 646468
rect 673730 605752 673736 605804
rect 673788 605792 673794 605804
rect 675202 605792 675208 605804
rect 673788 605764 675208 605792
rect 673788 605752 673794 605764
rect 675202 605752 675208 605764
rect 675260 605792 675266 605804
rect 675386 605792 675392 605804
rect 675260 605764 675392 605792
rect 675260 605752 675266 605764
rect 675386 605752 675392 605764
rect 675444 605752 675450 605804
rect 673730 601808 673736 601860
rect 673788 601848 673794 601860
rect 675202 601848 675208 601860
rect 673788 601820 675208 601848
rect 673788 601808 673794 601820
rect 675202 601808 675208 601820
rect 675260 601848 675266 601860
rect 675386 601848 675392 601860
rect 675260 601820 675392 601848
rect 675260 601808 675266 601820
rect 675386 601808 675392 601820
rect 675444 601808 675450 601860
rect 673730 561212 673736 561264
rect 673788 561252 673794 561264
rect 675202 561252 675208 561264
rect 673788 561224 675208 561252
rect 673788 561212 673794 561224
rect 675202 561212 675208 561224
rect 675260 561252 675266 561264
rect 675386 561252 675392 561264
rect 675260 561224 675392 561252
rect 675260 561212 675266 561224
rect 675386 561212 675392 561224
rect 675444 561212 675450 561264
rect 675202 557268 675208 557320
rect 675260 557308 675266 557320
rect 675386 557308 675392 557320
rect 675260 557280 675392 557308
rect 675260 557268 675266 557280
rect 675386 557268 675392 557280
rect 675444 557268 675450 557320
rect 673638 379040 673644 379092
rect 673696 379080 673702 379092
rect 675386 379080 675392 379092
rect 673696 379052 675392 379080
rect 673696 379040 673702 379052
rect 675386 379040 675392 379052
rect 675444 379040 675450 379092
rect 673638 338784 673644 338836
rect 673696 338824 673702 338836
rect 675386 338824 675392 338836
rect 673696 338796 675392 338824
rect 673696 338784 673702 338796
rect 675386 338784 675392 338796
rect 675444 338784 675450 338836
rect 673822 334228 673828 334280
rect 673880 334268 673886 334280
rect 675386 334268 675392 334280
rect 673880 334240 675392 334268
rect 673880 334228 673886 334240
rect 675386 334228 675392 334240
rect 675444 334228 675450 334280
rect 673822 293700 673828 293752
rect 673880 293740 673886 293752
rect 675294 293740 675300 293752
rect 673880 293712 675300 293740
rect 673880 293700 673886 293712
rect 675294 293700 675300 293712
rect 675352 293700 675358 293752
rect 673730 288804 673736 288856
rect 673788 288844 673794 288856
rect 675386 288844 675392 288856
rect 673788 288816 675392 288844
rect 673788 288804 673794 288816
rect 675386 288804 675392 288816
rect 675444 288804 675450 288856
rect 673730 249092 673736 249144
rect 673788 249132 673794 249144
rect 675386 249132 675392 249144
rect 673788 249104 675392 249132
rect 673788 249092 673794 249104
rect 675386 249092 675392 249104
rect 675444 249092 675450 249144
rect 673730 243788 673736 243840
rect 673788 243828 673794 243840
rect 675386 243828 675392 243840
rect 673788 243800 675392 243828
rect 673788 243788 673794 243800
rect 675386 243788 675392 243800
rect 675444 243788 675450 243840
rect 673730 203464 673736 203516
rect 673788 203504 673794 203516
rect 675294 203504 675300 203516
rect 673788 203476 675300 203504
rect 673788 203464 673794 203476
rect 675294 203464 675300 203476
rect 675352 203464 675358 203516
rect 673730 199044 673736 199096
rect 673788 199084 673794 199096
rect 675386 199084 675392 199096
rect 673788 199056 675392 199084
rect 673788 199044 673794 199056
rect 675386 199044 675392 199056
rect 675444 199044 675450 199096
rect 42334 197480 42340 197532
rect 42392 197480 42398 197532
rect 42352 197328 42380 197480
rect 42334 197276 42340 197328
rect 42392 197276 42398 197328
rect 673730 158584 673736 158636
rect 673788 158624 673794 158636
rect 675386 158624 675392 158636
rect 673788 158596 675392 158624
rect 673788 158584 673794 158596
rect 675386 158584 675392 158596
rect 675444 158584 675450 158636
rect 673730 154096 673736 154148
rect 673788 154136 673794 154148
rect 675294 154136 675300 154148
rect 673788 154108 675300 154136
rect 673788 154096 673794 154108
rect 675294 154096 675300 154108
rect 675352 154096 675358 154148
rect 673638 113704 673644 113756
rect 673696 113744 673702 113756
rect 675386 113744 675392 113756
rect 673696 113716 675392 113744
rect 673696 113704 673702 113716
rect 675386 113704 675392 113716
rect 675444 113704 675450 113756
rect 673638 108400 673644 108452
rect 673696 108440 673702 108452
rect 675386 108440 675392 108452
rect 673696 108412 675392 108440
rect 673696 108400 673702 108412
rect 675386 108400 675392 108412
rect 675444 108400 675450 108452
rect 673638 46968 673644 46980
rect 527468 46940 673644 46968
rect 527468 46912 527496 46940
rect 673638 46928 673644 46940
rect 673696 46928 673702 46980
rect 527450 46860 527456 46912
rect 527508 46860 527514 46912
rect 42334 45568 42340 45620
rect 42392 45608 42398 45620
rect 143626 45608 143632 45620
rect 42392 45580 143632 45608
rect 42392 45568 42398 45580
rect 143626 45568 143632 45580
rect 143684 45568 143690 45620
rect 199654 44412 199660 44464
rect 199712 44452 199718 44464
rect 199712 44424 207014 44452
rect 199712 44412 199718 44424
rect 143626 44140 143632 44192
rect 143684 44180 143690 44192
rect 145098 44180 145104 44192
rect 143684 44152 145104 44180
rect 143684 44140 143690 44152
rect 145098 44140 145104 44152
rect 145156 44180 145162 44192
rect 195330 44180 195336 44192
rect 145156 44152 195336 44180
rect 145156 44140 145162 44152
rect 195330 44140 195336 44152
rect 195388 44180 195394 44192
rect 199654 44180 199660 44192
rect 195388 44152 199660 44180
rect 195388 44140 195394 44152
rect 199654 44140 199660 44152
rect 199712 44140 199718 44192
rect 206986 44248 207014 44424
rect 363046 44316 363052 44328
rect 284266 44288 303936 44316
rect 284266 44248 284294 44288
rect 303908 44260 303936 44288
rect 361546 44288 363052 44316
rect 206986 44220 284294 44248
rect 303890 44208 303896 44260
rect 303948 44248 303954 44260
rect 308214 44248 308220 44260
rect 303948 44220 308220 44248
rect 303948 44208 303954 44220
rect 308214 44208 308220 44220
rect 308272 44248 308278 44260
rect 358722 44248 358728 44260
rect 308272 44220 358728 44248
rect 308272 44208 308278 44220
rect 358722 44208 358728 44220
rect 358780 44248 358786 44260
rect 361546 44248 361574 44288
rect 363046 44276 363052 44288
rect 363104 44316 363110 44328
rect 413554 44316 413560 44328
rect 363104 44288 413560 44316
rect 363104 44276 363110 44288
rect 413554 44276 413560 44288
rect 413612 44316 413618 44328
rect 417878 44316 417884 44328
rect 413612 44288 417884 44316
rect 413612 44276 413618 44288
rect 417878 44276 417884 44288
rect 417936 44316 417942 44328
rect 468294 44316 468300 44328
rect 417936 44288 468300 44316
rect 417936 44276 417942 44288
rect 468294 44276 468300 44288
rect 468352 44316 468358 44328
rect 472618 44316 472624 44328
rect 468352 44288 472624 44316
rect 468352 44276 468358 44288
rect 472618 44276 472624 44288
rect 472676 44316 472682 44328
rect 472676 44288 523172 44316
rect 472676 44276 472682 44288
rect 358780 44220 361574 44248
rect 358780 44208 358786 44220
rect 523144 44192 523172 44288
rect 523126 44140 523132 44192
rect 523184 44180 523190 44192
rect 527450 44180 527456 44192
rect 523184 44152 527456 44180
rect 523184 44140 523190 44152
rect 527450 44140 527456 44152
rect 527508 44140 527514 44192
rect 409322 41760 409328 41812
rect 409380 41800 409386 41812
rect 412358 41800 412364 41812
rect 409380 41772 412364 41800
rect 409380 41760 409386 41772
rect 412358 41760 412364 41772
rect 412416 41800 412422 41812
rect 415210 41800 415216 41812
rect 412416 41772 415216 41800
rect 412416 41760 412422 41772
rect 415210 41760 415216 41772
rect 415268 41760 415274 41812
rect 464154 41760 464160 41812
rect 464212 41800 464218 41812
rect 467190 41800 467196 41812
rect 464212 41772 467196 41800
rect 464212 41760 464218 41772
rect 467190 41760 467196 41772
rect 467248 41800 467254 41812
rect 470042 41800 470048 41812
rect 467248 41772 470048 41800
rect 467248 41760 467254 41772
rect 470042 41760 470048 41772
rect 470100 41760 470106 41812
<< via1 >>
rect 78864 990564 78916 990616
rect 83188 990564 83240 990616
rect 130292 990564 130344 990616
rect 134616 990564 134668 990616
rect 181720 990564 181772 990616
rect 186044 990564 186096 990616
rect 233056 990564 233108 990616
rect 237380 990564 237432 990616
rect 274456 990564 274508 990616
rect 274732 990632 274784 990684
rect 284668 990632 284720 990684
rect 288992 990632 289044 990684
rect 386512 990564 386564 990616
rect 390836 990564 390888 990616
rect 475476 990564 475528 990616
rect 479800 990564 479852 990616
rect 526904 990564 526956 990616
rect 531228 990564 531280 990616
rect 628656 990564 628708 990616
rect 632980 990564 633032 990616
rect 634728 990564 634780 990616
rect 42340 990224 42392 990276
rect 78864 990224 78916 990276
rect 634728 990088 634780 990140
rect 673828 990088 673880 990140
rect 673828 965268 673880 965320
rect 675392 965268 675444 965320
rect 41788 961120 41840 961172
rect 42524 961120 42576 961172
rect 673644 960032 673696 960084
rect 675392 960032 675444 960084
rect 673644 875780 673696 875832
rect 675392 875780 675444 875832
rect 673828 871292 673880 871344
rect 675300 871292 675352 871344
rect 41788 791936 41840 791988
rect 42524 791936 42576 791988
rect 41788 786972 41840 787024
rect 42432 786972 42484 787024
rect 673828 785952 673880 786004
rect 675208 785952 675260 786004
rect 675392 785952 675444 786004
rect 673736 781600 673788 781652
rect 675208 781600 675260 781652
rect 675392 781600 675444 781652
rect 42432 756576 42484 756628
rect 42432 756372 42484 756424
rect 41972 747872 42024 747924
rect 42340 747872 42392 747924
rect 41788 743452 41840 743504
rect 42340 743452 42392 743504
rect 673736 740936 673788 740988
rect 675208 740936 675260 740988
rect 675392 740936 675444 740988
rect 673736 736992 673788 737044
rect 675208 736992 675260 737044
rect 675392 736992 675444 737044
rect 42340 719040 42392 719092
rect 42340 718836 42392 718888
rect 673736 695920 673788 695972
rect 675208 695920 675260 695972
rect 675392 695920 675444 695972
rect 673736 692044 673788 692096
rect 675208 692044 675260 692096
rect 675392 692044 675444 692096
rect 673736 651108 673788 651160
rect 675392 651108 675444 651160
rect 673736 646416 673788 646468
rect 675392 646416 675444 646468
rect 673736 605752 673788 605804
rect 675208 605752 675260 605804
rect 675392 605752 675444 605804
rect 673736 601808 673788 601860
rect 675208 601808 675260 601860
rect 675392 601808 675444 601860
rect 673736 561212 673788 561264
rect 675208 561212 675260 561264
rect 675392 561212 675444 561264
rect 675208 557268 675260 557320
rect 675392 557268 675444 557320
rect 673644 379040 673696 379092
rect 675392 379040 675444 379092
rect 673644 338784 673696 338836
rect 675392 338784 675444 338836
rect 673828 334228 673880 334280
rect 675392 334228 675444 334280
rect 673828 293700 673880 293752
rect 675300 293700 675352 293752
rect 673736 288804 673788 288856
rect 675392 288804 675444 288856
rect 673736 249092 673788 249144
rect 675392 249092 675444 249144
rect 673736 243788 673788 243840
rect 675392 243788 675444 243840
rect 673736 203464 673788 203516
rect 675300 203464 675352 203516
rect 673736 199044 673788 199096
rect 675392 199044 675444 199096
rect 42340 197480 42392 197532
rect 42340 197276 42392 197328
rect 673736 158584 673788 158636
rect 675392 158584 675444 158636
rect 673736 154096 673788 154148
rect 675300 154096 675352 154148
rect 673644 113704 673696 113756
rect 675392 113704 675444 113756
rect 673644 108400 673696 108452
rect 675392 108400 675444 108452
rect 673644 46928 673696 46980
rect 527456 46860 527508 46912
rect 42340 45568 42392 45620
rect 143632 45568 143684 45620
rect 199660 44412 199712 44464
rect 143632 44140 143684 44192
rect 145104 44140 145156 44192
rect 195336 44140 195388 44192
rect 199660 44140 199712 44192
rect 303896 44208 303948 44260
rect 308220 44208 308272 44260
rect 358728 44208 358780 44260
rect 363052 44276 363104 44328
rect 413560 44276 413612 44328
rect 417884 44276 417936 44328
rect 468300 44276 468352 44328
rect 472624 44276 472676 44328
rect 523132 44140 523184 44192
rect 527456 44140 527508 44192
rect 409328 41760 409380 41812
rect 412364 41760 412416 41812
rect 415216 41760 415268 41812
rect 464160 41760 464212 41812
rect 467196 41760 467248 41812
rect 470048 41760 470100 41812
<< obsm1 >>
rect 76171 996231 92229 1037600
rect 127571 996231 143629 1037600
rect 178971 996231 195029 1037600
rect 230371 996231 246429 1037600
rect 281971 996231 298029 1037600
rect 333437 998007 348124 1037545
rect 335807 997984 336070 998007
tri 336070 997984 336093 998007 sw
tri 347285 997984 347308 998007 se
rect 347308 997984 347536 998007
rect 335807 997794 347536 997984
rect 383771 996231 399829 1037600
rect 472771 996231 488829 1037600
rect 524171 996231 540229 1037600
rect 575637 998007 590324 1037545
rect 578007 997984 578270 998007
tri 578270 997984 578293 998007 sw
tri 589485 997984 589508 998007 se
rect 589508 997984 589736 998007
rect 578007 997794 589736 997984
rect 625971 996231 642029 1037600
rect 84010 995636 84074 995648
rect 91738 995636 91802 995648
rect 84010 995608 91802 995636
rect 84010 995596 84074 995608
rect 91738 995596 91802 995608
rect 238202 995636 238266 995648
rect 245930 995636 245994 995648
rect 238202 995608 245994 995636
rect 238202 995596 238266 995608
rect 245930 995596 245994 995608
rect 531958 995636 532022 995648
rect 539686 995636 539750 995648
rect 531958 995608 539750 995636
rect 531958 995596 532022 995608
rect 539686 995596 539750 995608
rect 135346 995500 135410 995512
rect 143166 995500 143230 995512
rect 135346 995472 143230 995500
rect 135346 995460 135410 995472
rect 143166 995460 143230 995472
rect 633802 995500 633866 995512
rect 641530 995500 641594 995512
rect 633802 995472 641594 995500
rect 633802 995460 633866 995472
rect 641530 995460 641594 995472
rect 289630 995296 289694 995308
rect 297634 995296 297698 995308
rect 289630 995268 297698 995296
rect 289630 995256 289694 995268
rect 297634 995256 297698 995268
rect 391474 995296 391538 995308
rect 399478 995296 399542 995308
rect 391474 995268 399542 995296
rect 391474 995256 391538 995268
rect 399478 995256 399542 995268
rect 480438 995296 480502 995308
rect 488442 995296 488506 995308
rect 480438 995268 488506 995296
rect 480438 995256 480502 995268
rect 488442 995256 488506 995268
rect 585042 992236 585106 992248
rect 674742 992236 674806 992248
rect 585042 992208 674806 992236
rect 585042 992196 585106 992208
rect 674742 992196 674806 992208
rect 82538 990808 82602 990820
rect 133966 990808 134030 990820
rect 135162 990808 135226 990820
rect 82538 990780 135226 990808
rect 82538 990768 82602 990780
rect 133966 990768 134030 990780
rect 135162 990768 135226 990780
rect 184934 990808 184998 990820
rect 185394 990808 185458 990820
rect 236730 990808 236794 990820
rect 184934 990780 236794 990808
rect 184934 990768 184998 990780
rect 185394 990768 185458 990780
rect 236730 990768 236794 990780
rect 88334 990740 88398 990752
rect 89990 990740 90054 990752
rect 141418 990740 141482 990752
rect 192846 990740 192910 990752
rect 244182 990740 244246 990752
rect 295794 990740 295858 990752
rect 397638 990740 397702 990752
rect 486602 990740 486666 990752
rect 538030 990740 538094 990752
rect 639782 990740 639846 990752
rect 88334 990712 639846 990740
rect 88334 990700 88398 990712
rect 89990 990700 90054 990712
rect 141418 990700 141482 990712
rect 192846 990700 192910 990712
rect 244182 990700 244246 990712
rect 295794 990700 295858 990712
rect 397638 990700 397702 990712
rect 486602 990700 486666 990712
rect 538030 990700 538094 990712
rect 639782 990700 639846 990712
rect 79502 990672 79566 990684
rect 130930 990672 130994 990684
rect 182358 990672 182422 990684
rect 233694 990672 233758 990684
rect 79502 990644 274680 990672
rect 79502 990632 79566 990644
rect 130930 990632 130994 990644
rect 182358 990632 182422 990644
rect 233694 990632 233758 990644
rect 274652 990604 274680 990644
rect 390186 990672 390250 990684
rect 479150 990672 479214 990684
rect 480162 990672 480226 990684
rect 390186 990644 480226 990672
rect 390186 990632 390250 990644
rect 479150 990632 479214 990644
rect 480162 990632 480226 990644
rect 527542 990672 527606 990684
rect 629294 990672 629358 990684
rect 631778 990672 631842 990684
rect 527542 990644 631842 990672
rect 527542 990632 527606 990644
rect 629294 990632 629358 990644
rect 631778 990632 631842 990644
rect 285306 990604 285370 990616
rect 342162 990604 342226 990616
rect 386414 990604 386478 990616
rect 274652 990576 386478 990604
rect 285306 990564 285370 990576
rect 342162 990564 342226 990576
rect 386414 990564 386478 990576
rect 186682 990536 186746 990548
rect 194686 990536 194750 990548
rect 186682 990508 194750 990536
rect 186682 990496 186746 990508
rect 194686 990496 194750 990508
rect 236730 990536 236794 990548
rect 288342 990536 288406 990548
rect 390186 990536 390250 990548
rect 476114 990536 476178 990548
rect 527542 990536 527606 990548
rect 632330 990536 632394 990548
rect 236730 990508 390250 990536
rect 236730 990496 236794 990508
rect 288342 990496 288406 990508
rect 390186 990496 390250 990508
rect 438826 990508 527606 990536
rect 135162 990468 135226 990480
rect 184934 990468 184998 990480
rect 135162 990440 184998 990468
rect 135162 990428 135226 990440
rect 184934 990428 184998 990440
rect 386414 990468 386478 990480
rect 387150 990468 387214 990480
rect 438826 990468 438854 990508
rect 476114 990496 476178 990508
rect 527542 990496 527606 990508
rect 535426 990508 632394 990536
rect 386414 990440 438854 990468
rect 480162 990468 480226 990480
rect 530578 990468 530642 990480
rect 535426 990468 535454 990508
rect 480162 990440 535454 990468
rect 386414 990428 386478 990440
rect 387150 990428 387214 990440
rect 480162 990428 480226 990440
rect 530578 990428 530642 990440
rect 42242 990196 42306 990208
rect 79502 990196 79566 990208
rect 42242 990168 79566 990196
rect 632026 990196 632054 990508
rect 632330 990496 632394 990508
rect 639782 990264 639846 990276
rect 673730 990264 673794 990276
rect 639782 990236 673794 990264
rect 639782 990224 639846 990236
rect 673730 990224 673794 990236
rect 673454 990196 673518 990208
rect 632026 990168 673518 990196
rect 42242 990156 42306 990168
rect 79502 990156 79566 990168
rect 673454 990156 673518 990168
rect 44910 990128 44974 990140
rect 82538 990128 82602 990140
rect 44910 990100 82602 990128
rect 44910 990088 44974 990100
rect 82538 990088 82602 990100
rect 88334 990088 88398 990140
rect 631778 990128 631842 990140
rect 631778 990100 632054 990128
rect 631778 990088 631842 990100
rect 42610 990060 42674 990072
rect 88352 990060 88380 990088
rect 42610 990032 88380 990060
rect 632026 990060 632054 990100
rect 673638 990060 673702 990072
rect 632026 990032 673702 990060
rect 42610 990020 42674 990032
rect 673638 990020 673702 990032
rect 0 954171 41369 970229
rect 41782 969388 41846 969400
rect 42334 969388 42398 969400
rect 41782 969360 42398 969388
rect 41782 969348 41846 969360
rect 42334 969348 42398 969360
rect 41782 968504 41846 968516
rect 42610 968504 42674 968516
rect 41782 968476 42674 968504
rect 41782 968464 41846 968476
rect 42610 968464 42674 968476
rect 673638 964764 673702 964776
rect 675386 964764 675450 964776
rect 673638 964736 675450 964764
rect 673638 964724 673702 964736
rect 675386 964724 675450 964736
rect 41782 962452 41846 962464
rect 42334 962452 42398 962464
rect 41782 962424 42398 962452
rect 41782 962412 41846 962424
rect 42334 962412 42398 962424
rect 673454 961364 673518 961376
rect 675386 961364 675450 961376
rect 673454 961336 675450 961364
rect 673454 961324 673518 961336
rect 675386 961324 675450 961336
rect 41966 960480 42030 960492
rect 44818 960480 44882 960492
rect 41966 960452 44882 960480
rect 41966 960440 42030 960452
rect 44818 960440 44882 960452
rect 44174 955040 44238 955052
rect 44818 955040 44882 955052
rect 44174 955012 44882 955040
rect 44174 955000 44238 955012
rect 44818 955000 44882 955012
rect 673730 953340 673794 953352
rect 675386 953340 675450 953352
rect 673730 953312 675450 953340
rect 673730 953300 673794 953312
rect 675386 953300 675450 953312
rect 676231 951571 717600 967629
rect 24523 928387 40977 929187
tri 40977 928387 41777 929187 sw
rect 24523 927240 41777 928387
rect 32 923313 39593 927000
rect 39756 923313 41777 927240
rect 32 916185 41777 923313
rect 678007 919269 717568 922576
rect 678000 918415 717568 919269
rect 32 915331 39600 916185
rect 32 912024 39593 915331
rect 675823 911287 717568 918415
rect 675823 907360 677844 911287
rect 678007 907600 717568 911287
rect 675823 906213 693077 907360
tri 675823 905413 676623 906213 ne
rect 676623 905413 693077 906213
rect 55 883936 39593 884383
rect 55 883708 39806 883936
rect 55 872470 39593 883708
tri 39593 883685 39616 883708 ne
tri 39593 872470 39616 872493 se
rect 39616 872470 39806 883708
rect 673546 874528 673610 874540
rect 675386 874528 675450 874540
rect 673546 874500 675450 874528
rect 673546 874488 673610 874500
rect 675386 874488 675450 874500
rect 55 872207 39806 872470
rect 673454 872420 673518 872432
rect 674006 872420 674070 872432
rect 675386 872420 675450 872432
rect 673454 872392 675450 872420
rect 673454 872380 673518 872392
rect 674006 872380 674070 872392
rect 675386 872380 675450 872392
rect 55 871571 39593 872207
rect 55 870525 39774 871571
rect 673454 870584 673518 870596
rect 673730 870584 673794 870596
rect 673454 870556 673794 870584
rect 673454 870544 673518 870556
rect 673730 870544 673794 870556
rect 55 869837 39593 870525
rect 673914 870176 673978 870188
rect 675386 870176 675450 870188
rect 673914 870148 675450 870176
rect 673914 870136 673978 870148
rect 675386 870136 675450 870148
rect 673454 864464 673518 864476
rect 675386 864464 675450 864476
rect 673454 864436 675450 864464
rect 673454 864424 673518 864436
rect 675386 864424 675450 864436
rect 673914 863240 673978 863252
rect 675386 863240 675450 863252
rect 673914 863212 675450 863240
rect 673914 863200 673978 863212
rect 675386 863200 675450 863212
rect 676231 862371 717600 878429
rect 55 841736 39593 842324
rect 55 841508 39806 841736
rect 55 830270 39593 841508
tri 39593 841485 39616 841508 ne
tri 39593 830270 39616 830293 se
rect 39616 830270 39806 841508
rect 678007 832675 717545 833363
rect 677826 831629 717545 832675
rect 678007 830993 717545 831629
rect 55 830007 39806 830270
rect 677794 830730 717545 830993
rect 55 827637 39593 830007
rect 677794 819492 677984 830730
tri 677984 830707 678007 830730 nw
tri 677984 819492 678007 819515 sw
rect 678007 819492 717545 830730
rect 677794 819264 717545 819492
rect 678007 818817 717545 819264
rect 675294 818360 675358 818372
rect 677594 818360 677658 818372
rect 675294 818332 677658 818360
rect 675294 818320 675358 818332
rect 677594 818320 677658 818332
rect 0 784371 41369 800429
rect 41782 797756 41846 797768
rect 42334 797756 42398 797768
rect 41782 797728 42398 797756
rect 41782 797716 41846 797728
rect 42334 797716 42398 797728
rect 41782 791364 41846 791376
rect 42242 791364 42306 791376
rect 42426 791364 42490 791376
rect 41782 791336 42490 791364
rect 41782 791324 41846 791336
rect 42242 791324 42306 791336
rect 42426 791324 42490 791336
rect 41782 787284 41846 787296
rect 42610 787284 42674 787296
rect 41782 787256 42674 787284
rect 41782 787244 41846 787256
rect 42610 787244 42674 787256
rect 673546 785720 673610 785732
rect 675386 785720 675450 785732
rect 673546 785692 675450 785720
rect 673546 785680 673610 785692
rect 675386 785680 675450 785692
rect 673638 782320 673702 782332
rect 674006 782320 674070 782332
rect 675386 782320 675450 782332
rect 673638 782292 675450 782320
rect 673638 782280 673702 782292
rect 674006 782280 674070 782292
rect 675386 782280 675450 782292
rect 675202 781028 675266 781040
rect 675386 781028 675450 781040
rect 675202 781000 675450 781028
rect 675202 780988 675266 781000
rect 675386 780988 675450 781000
rect 673454 775860 673518 775872
rect 675386 775860 675450 775872
rect 673454 775832 675450 775860
rect 673454 775820 673518 775832
rect 675386 775820 675450 775832
rect 676231 773171 717600 789229
rect 0 741171 41369 757229
rect 41782 756412 41846 756424
rect 42334 756412 42398 756424
rect 41782 756384 42398 756412
rect 41782 756372 41846 756384
rect 42334 756372 42398 756384
rect 41782 755460 41846 755472
rect 42518 755460 42582 755472
rect 41782 755432 42582 755460
rect 41782 755420 41846 755432
rect 42518 755420 42582 755432
rect 41782 749408 41846 749420
rect 42334 749408 42398 749420
rect 41782 749380 42398 749408
rect 41782 749368 41846 749380
rect 42334 749368 42398 749380
rect 41782 744036 41846 744048
rect 42610 744036 42674 744048
rect 41782 744008 42674 744036
rect 41782 743996 41846 744008
rect 42610 743996 42674 744008
rect 673546 740364 673610 740376
rect 673822 740364 673886 740376
rect 675386 740364 675450 740376
rect 673546 740336 675450 740364
rect 673546 740324 673610 740336
rect 673822 740324 673886 740336
rect 675386 740324 675450 740336
rect 673638 738120 673702 738132
rect 675386 738120 675450 738132
rect 673638 738092 675450 738120
rect 673638 738080 673702 738092
rect 675386 738080 675450 738092
rect 673454 730912 673518 730924
rect 673914 730912 673978 730924
rect 675386 730912 675450 730924
rect 673454 730884 675450 730912
rect 673454 730872 673518 730884
rect 673914 730872 673978 730884
rect 675386 730872 675450 730884
rect 676231 728171 717600 744229
rect 0 697971 41369 714029
rect 41782 712280 41846 712292
rect 42518 712280 42582 712292
rect 41782 712252 42582 712280
rect 41782 712240 41846 712252
rect 42518 712240 42582 712252
rect 41782 703984 41846 703996
rect 42426 703984 42490 703996
rect 41782 703956 42490 703984
rect 41782 703944 41846 703956
rect 42426 703944 42490 703956
rect 41782 700856 41846 700868
rect 42610 700856 42674 700868
rect 41782 700828 42674 700856
rect 41782 700816 41846 700828
rect 42610 700816 42674 700828
rect 673454 695348 673518 695360
rect 673822 695348 673886 695360
rect 675386 695348 675450 695360
rect 673454 695320 675450 695348
rect 673454 695308 673518 695320
rect 673822 695308 673886 695320
rect 675386 695308 675450 695320
rect 673638 692288 673702 692300
rect 675386 692288 675450 692300
rect 673638 692260 675450 692288
rect 673638 692248 673702 692260
rect 675386 692248 675450 692260
rect 673546 685216 673610 685228
rect 673914 685216 673978 685228
rect 675386 685216 675450 685228
rect 673546 685188 675450 685216
rect 673546 685176 673610 685188
rect 673914 685176 673978 685188
rect 675386 685176 675450 685188
rect 676231 683171 717600 699229
rect 0 654771 41369 670829
rect 41782 668148 41846 668160
rect 42518 668148 42582 668160
rect 41782 668120 42582 668148
rect 41782 668108 41846 668120
rect 42518 668108 42582 668120
rect 41782 661076 41846 661088
rect 42426 661076 42490 661088
rect 41782 661048 42490 661076
rect 41782 661036 41846 661048
rect 42426 661036 42490 661048
rect 41782 658696 41846 658708
rect 42610 658696 42674 658708
rect 41782 658668 42674 658696
rect 41782 658656 41846 658668
rect 42610 658656 42674 658668
rect 673454 650536 673518 650548
rect 675386 650536 675450 650548
rect 673454 650508 675450 650536
rect 673454 650496 673518 650508
rect 675386 650496 675450 650508
rect 673638 647068 673702 647080
rect 675386 647068 675450 647080
rect 673638 647040 675450 647068
rect 673638 647028 673702 647040
rect 675386 647028 675450 647040
rect 675202 645776 675266 645788
rect 675386 645776 675450 645788
rect 675202 645748 675450 645776
rect 675202 645736 675266 645748
rect 675386 645736 675450 645748
rect 673546 640676 673610 640688
rect 675386 640676 675450 640688
rect 673546 640648 675450 640676
rect 673546 640636 673610 640648
rect 675386 640636 675450 640648
rect 676231 637971 717600 654029
rect 0 611571 41369 627629
rect 41782 624968 41846 624980
rect 42518 624968 42582 624980
rect 41782 624940 42582 624968
rect 41782 624928 41846 624940
rect 42518 624928 42582 624940
rect 41782 618508 41846 618520
rect 42426 618508 42490 618520
rect 41782 618480 42490 618508
rect 41782 618468 41846 618480
rect 42426 618468 42490 618480
rect 41782 615516 41846 615528
rect 42610 615516 42674 615528
rect 41782 615488 42674 615516
rect 41782 615476 41846 615488
rect 42610 615476 42674 615488
rect 673454 605112 673518 605124
rect 675386 605112 675450 605124
rect 673454 605084 675450 605112
rect 673454 605072 673518 605084
rect 675386 605072 675450 605084
rect 42518 603168 42582 603220
rect 42536 603016 42564 603168
rect 42518 602964 42582 603016
rect 673638 602936 673702 602948
rect 673822 602936 673886 602948
rect 675386 602936 675450 602948
rect 673638 602908 675450 602936
rect 673638 602896 673702 602908
rect 673822 602896 673886 602908
rect 675386 602896 675450 602908
rect 673546 595660 673610 595672
rect 673914 595660 673978 595672
rect 675386 595660 675450 595672
rect 673546 595632 675450 595660
rect 673546 595620 673610 595632
rect 673914 595620 673978 595632
rect 675386 595620 675450 595632
rect 676231 592971 717600 609029
rect 0 568371 41369 584429
rect 41782 581720 41846 581732
rect 42426 581720 42490 581732
rect 41782 581692 42490 581720
rect 41782 581680 41846 581692
rect 42426 581680 42490 581692
rect 41782 575260 41846 575272
rect 42702 575260 42766 575272
rect 41782 575232 42766 575260
rect 41782 575220 41846 575232
rect 42702 575220 42766 575232
rect 41782 572268 41846 572280
rect 42518 572268 42582 572280
rect 42794 572268 42858 572280
rect 41782 572240 42858 572268
rect 41782 572228 41846 572240
rect 42518 572228 42582 572240
rect 42794 572228 42858 572240
rect 42242 571180 42306 571192
rect 42426 571180 42490 571192
rect 42242 571152 42490 571180
rect 42242 571140 42306 571152
rect 42426 571140 42490 571152
rect 673454 559960 673518 559972
rect 675386 559960 675450 559972
rect 673454 559932 675450 559960
rect 673454 559920 673518 559932
rect 675386 559920 675450 559932
rect 673822 557852 673886 557864
rect 675386 557852 675450 557864
rect 673822 557824 675450 557852
rect 673822 557812 673886 557824
rect 675386 557812 675450 557824
rect 675202 555608 675266 555620
rect 675386 555608 675450 555620
rect 675202 555580 675450 555608
rect 675202 555568 675266 555580
rect 675386 555568 675450 555580
rect 673914 550508 673978 550520
rect 675386 550508 675450 550520
rect 673914 550480 675450 550508
rect 673914 550468 673978 550480
rect 675386 550468 675450 550480
rect 676231 547771 717600 563829
rect 42242 543096 42306 543108
rect 42426 543096 42490 543108
rect 42242 543068 42490 543096
rect 42242 543056 42306 543068
rect 42426 543056 42490 543068
rect 0 525171 41369 541229
rect 41782 539492 41846 539504
rect 42426 539492 42490 539504
rect 42702 539492 42766 539504
rect 41782 539464 42766 539492
rect 41782 539452 41846 539464
rect 42426 539452 42490 539464
rect 42702 539452 42766 539464
rect 41782 531196 41846 531208
rect 42610 531196 42674 531208
rect 41782 531168 42674 531196
rect 41782 531156 41846 531168
rect 42610 531156 42674 531168
rect 41782 528068 41846 528080
rect 42518 528068 42582 528080
rect 41782 528040 42582 528068
rect 41782 528028 41846 528040
rect 42518 528028 42582 528040
rect 678007 518075 717545 518763
rect 677826 517029 717545 518075
rect 678007 516393 717545 517029
rect 677794 516130 717545 516393
rect 675294 513788 675358 513800
rect 677686 513788 677750 513800
rect 675294 513760 677750 513788
rect 675294 513748 675358 513760
rect 677686 513748 677750 513760
rect 677794 504892 677984 516130
tri 677984 516107 678007 516130 nw
tri 677984 504892 678007 504915 sw
rect 678007 504892 717545 516130
rect 677794 504664 717545 504892
rect 678007 504217 717545 504664
rect 55 497136 39593 497583
rect 55 496908 39806 497136
rect 55 485670 39593 496908
tri 39593 496885 39616 496908 ne
tri 39593 485670 39616 485693 se
rect 39616 485670 39806 496908
rect 55 485407 39806 485670
rect 55 484771 39593 485407
rect 55 483725 39774 484771
rect 55 483037 39593 483725
rect 678007 471469 717568 474776
rect 678000 470615 717568 471469
rect 675823 463487 717568 470615
rect 675823 459560 677844 463487
rect 678007 459800 717568 463487
rect 675823 458413 693077 459560
tri 675823 457987 676249 458413 ne
rect 676249 457987 693077 458413
rect 24523 457187 40977 457987
tri 40977 457187 41777 457987 sw
tri 676249 457613 676623 457987 ne
rect 676623 457613 693077 457987
rect 24523 456040 41777 457187
rect 32 452113 39593 455800
rect 39756 452113 41777 456040
rect 32 444985 41777 452113
rect 32 444131 39600 444985
rect 32 440824 39593 444131
rect 678007 428193 717545 430563
rect 677794 427930 717545 428193
rect 674742 427836 674806 427848
rect 677502 427836 677566 427848
rect 674742 427808 677566 427836
rect 674742 427796 674806 427808
rect 677502 427796 677566 427808
rect 677794 416692 677984 427930
tri 677984 427907 678007 427930 nw
tri 677984 416692 678007 416715 sw
rect 678007 416692 717545 427930
rect 677794 416464 717545 416692
rect 678007 415876 717545 416464
rect 0 397571 41369 413629
rect 41782 410972 41846 410984
rect 42426 410972 42490 410984
rect 42702 410972 42766 410984
rect 41782 410944 42766 410972
rect 41782 410932 41846 410944
rect 42426 410932 42490 410944
rect 42702 410932 42766 410944
rect 41782 404512 41846 404524
rect 42610 404512 42674 404524
rect 41782 404484 42674 404512
rect 41782 404472 41846 404484
rect 42610 404472 42674 404484
rect 41782 401520 41846 401532
rect 42518 401520 42582 401532
rect 42702 401520 42766 401532
rect 41782 401492 42766 401520
rect 41782 401480 41846 401492
rect 42518 401480 42582 401492
rect 42702 401480 42766 401492
rect 673454 383568 673518 383580
rect 675386 383568 675450 383580
rect 673454 383540 675450 383568
rect 673454 383528 673518 383540
rect 675386 383528 675450 383540
rect 673730 379692 673794 379704
rect 675386 379692 675450 379704
rect 673730 379664 675450 379692
rect 673730 379652 673794 379664
rect 675386 379652 675450 379664
rect 673454 372348 673518 372360
rect 673822 372348 673886 372360
rect 675386 372348 675450 372360
rect 673454 372320 675450 372348
rect 673454 372308 673518 372320
rect 673822 372308 673886 372320
rect 675386 372308 675450 372320
rect 676231 370571 717600 386629
rect 0 354371 41369 370429
rect 41782 369560 41846 369572
rect 42334 369560 42398 369572
rect 41782 369532 42398 369560
rect 41782 369520 41846 369532
rect 42334 369520 42398 369532
rect 41782 368676 41846 368688
rect 42426 368676 42490 368688
rect 41782 368648 42490 368676
rect 41782 368636 41846 368648
rect 42426 368636 42490 368648
rect 41782 362624 41846 362636
rect 42334 362624 42398 362636
rect 41782 362596 42398 362624
rect 41782 362584 41846 362596
rect 42334 362584 42398 362596
rect 41782 360720 41846 360732
rect 42610 360720 42674 360732
rect 41782 360692 42674 360720
rect 41782 360680 41846 360692
rect 42610 360680 42674 360692
rect 41782 357252 41846 357264
rect 42334 357252 42398 357264
rect 42702 357252 42766 357264
rect 41782 357224 42766 357252
rect 41782 357212 41846 357224
rect 42334 357212 42398 357224
rect 42702 357212 42766 357224
rect 673546 337532 673610 337544
rect 675386 337532 675450 337544
rect 673546 337504 675450 337532
rect 673546 337492 673610 337504
rect 675386 337492 675450 337504
rect 673730 334472 673794 334484
rect 675386 334472 675450 334484
rect 673730 334444 675450 334472
rect 673730 334432 673794 334444
rect 675386 334432 675450 334444
rect 673454 328080 673518 328092
rect 675386 328080 675450 328092
rect 673454 328052 675450 328080
rect 673454 328040 673518 328052
rect 675386 328040 675450 328052
rect 0 311171 41369 327229
rect 41782 325496 41846 325508
rect 42518 325496 42582 325508
rect 42702 325496 42766 325508
rect 41782 325468 42766 325496
rect 41782 325456 41846 325468
rect 42518 325456 42582 325468
rect 42702 325456 42766 325468
rect 676231 325371 717600 341429
rect 41782 317200 41846 317212
rect 42518 317200 42582 317212
rect 41782 317172 42582 317200
rect 41782 317160 41846 317172
rect 42518 317160 42582 317172
rect 41782 314072 41846 314084
rect 42426 314072 42490 314084
rect 42610 314072 42674 314084
rect 41782 314044 42674 314072
rect 41782 314032 41846 314044
rect 42426 314032 42490 314044
rect 42610 314032 42674 314044
rect 673454 313256 673518 313268
rect 673638 313256 673702 313268
rect 673454 313228 673702 313256
rect 673454 313216 673518 313228
rect 673638 313216 673702 313228
rect 673454 293196 673518 293208
rect 675386 293196 675450 293208
rect 673454 293168 675450 293196
rect 673454 293156 673518 293168
rect 675386 293156 675450 293168
rect 673546 289524 673610 289536
rect 673730 289524 673794 289536
rect 675386 289524 675450 289536
rect 673546 289496 675450 289524
rect 673546 289484 673610 289496
rect 673730 289484 673794 289496
rect 675386 289484 675450 289496
rect 0 267971 41369 284029
rect 673638 283064 673702 283076
rect 673914 283064 673978 283076
rect 675386 283064 675450 283076
rect 673638 283036 675450 283064
rect 673638 283024 673702 283036
rect 673914 283024 673978 283036
rect 675386 283024 675450 283036
rect 41782 281364 41846 281376
rect 42426 281364 42490 281376
rect 42702 281364 42766 281376
rect 41782 281336 42766 281364
rect 41782 281324 41846 281336
rect 42426 281324 42490 281336
rect 42702 281324 42766 281336
rect 676231 280371 717600 296429
rect 41782 274564 41846 274576
rect 42518 274564 42582 274576
rect 41782 274536 42582 274564
rect 41782 274524 41846 274536
rect 42518 274524 42582 274536
rect 41782 271912 41846 271924
rect 42610 271912 42674 271924
rect 41782 271884 42674 271912
rect 41782 271872 41846 271884
rect 42610 271872 42674 271884
rect 673454 248588 673518 248600
rect 674006 248588 674070 248600
rect 675386 248588 675450 248600
rect 673454 248560 675450 248588
rect 673454 248548 673518 248560
rect 674006 248548 674070 248560
rect 675386 248548 675450 248560
rect 673638 244916 673702 244928
rect 675386 244916 675450 244928
rect 673638 244888 675450 244916
rect 673638 244876 673702 244888
rect 675386 244876 675450 244888
rect 0 224771 41369 240829
rect 41782 238116 41846 238128
rect 42426 238116 42490 238128
rect 41782 238088 42490 238116
rect 41782 238076 41846 238088
rect 42426 238076 42490 238088
rect 673822 237708 673886 237720
rect 675386 237708 675450 237720
rect 673822 237680 675450 237708
rect 673822 237668 673886 237680
rect 675386 237668 675450 237680
rect 676231 235371 717600 251429
rect 41782 231724 41846 231736
rect 42518 231724 42582 231736
rect 41782 231696 42582 231724
rect 41782 231684 41846 231696
rect 42518 231684 42582 231696
rect 41782 228664 41846 228676
rect 42610 228664 42674 228676
rect 41782 228636 42674 228664
rect 41782 228624 41846 228636
rect 42610 228624 42674 228636
rect 42242 227508 42306 227520
rect 42518 227508 42582 227520
rect 42242 227480 42582 227508
rect 42242 227468 42306 227480
rect 42518 227468 42582 227480
rect 673546 202348 673610 202360
rect 674006 202348 674070 202360
rect 675386 202348 675450 202360
rect 673546 202320 675450 202348
rect 673546 202308 673610 202320
rect 674006 202308 674070 202320
rect 675386 202308 675450 202320
rect 673638 199288 673702 199300
rect 675386 199288 675450 199300
rect 673638 199260 675450 199288
rect 673638 199248 673702 199260
rect 675386 199248 675450 199260
rect 0 181571 41369 197629
rect 42426 197520 42490 197532
rect 42610 197520 42674 197532
rect 42426 197492 42674 197520
rect 42426 197480 42490 197492
rect 42610 197480 42674 197492
rect 41782 195888 41846 195900
rect 42610 195888 42674 195900
rect 41782 195860 42674 195888
rect 41782 195848 41846 195860
rect 42610 195848 42674 195860
rect 673914 191944 673978 191956
rect 675386 191944 675450 191956
rect 673914 191916 675450 191944
rect 673914 191904 673978 191916
rect 675386 191904 675450 191916
rect 676231 190171 717600 206229
rect 41782 187660 41846 187672
rect 42426 187660 42490 187672
rect 41782 187632 42490 187660
rect 41782 187620 41846 187632
rect 42426 187620 42490 187632
rect 41782 184464 41846 184476
rect 42518 184464 42582 184476
rect 41782 184436 42582 184464
rect 41782 184424 41846 184436
rect 42260 184204 42288 184436
rect 42518 184424 42582 184436
rect 42242 184152 42306 184204
rect 673546 158352 673610 158364
rect 675386 158352 675450 158364
rect 673546 158324 675450 158352
rect 673546 158312 673610 158324
rect 675386 158312 675450 158324
rect 673638 155224 673702 155236
rect 675386 155224 675450 155236
rect 673638 155196 675450 155224
rect 673638 155184 673702 155196
rect 675386 155184 675450 155196
rect 673822 146928 673886 146940
rect 675386 146928 675450 146940
rect 673822 146900 675450 146928
rect 673822 146888 673886 146900
rect 675386 146888 675450 146900
rect 676231 145171 717600 161229
rect 55 124336 39593 124783
rect 55 124108 39806 124336
rect 55 112870 39593 124108
tri 39593 124085 39616 124108 ne
tri 39593 112870 39616 112893 se
rect 39616 112870 39806 124108
rect 42426 121496 42490 121508
rect 44174 121496 44238 121508
rect 42426 121468 44238 121496
rect 42426 121456 42490 121468
rect 44174 121456 44238 121468
rect 673454 113200 673518 113212
rect 675386 113200 675450 113212
rect 673454 113172 675450 113200
rect 673454 113160 673518 113172
rect 675386 113160 675450 113172
rect 55 112607 39806 112870
rect 55 111971 39593 112607
rect 55 110925 39774 111971
rect 55 110237 39593 110925
rect 673546 109528 673610 109540
rect 675386 109528 675450 109540
rect 673546 109500 675450 109528
rect 673546 109488 673610 109500
rect 675386 109488 675450 109500
rect 673730 101708 673794 101720
rect 675386 101708 675450 101720
rect 673730 101680 675450 101708
rect 673730 101668 673794 101680
rect 675386 101668 675450 101680
rect 676231 99971 717600 116029
rect 31928 85187 32702 85239
rect 31928 84387 40900 85187
tri 40900 84387 41700 85187 sw
rect 31928 83240 41700 84387
rect 31928 83049 32702 83240
rect 32 79313 39593 83000
rect 39756 79313 41700 83240
rect 42610 80356 42674 80368
rect 44174 80356 44238 80368
rect 42610 80328 44238 80356
rect 42610 80316 42674 80328
rect 44174 80316 44238 80328
rect 32 72099 41700 79313
rect 32 71331 39600 72099
rect 39796 71731 41700 72099
tri 39796 71331 40196 71731 ne
rect 40196 71331 41300 71731
tri 41300 71331 41700 71731 nw
rect 32 68024 39593 71331
rect 44818 46928 44882 46980
rect 200868 46940 297772 46968
rect 44836 46900 44864 46928
rect 200868 46912 200896 46940
rect 248432 46912 248460 46940
rect 297744 46912 297772 46940
rect 309428 46940 352604 46968
rect 309428 46912 309456 46940
rect 352576 46912 352604 46940
rect 364260 46940 407436 46968
rect 364260 46912 364288 46940
rect 407408 46912 407436 46940
rect 419092 46940 462176 46968
rect 419092 46912 419120 46940
rect 462148 46912 462176 46940
rect 473832 46940 517008 46968
rect 473832 46912 473860 46940
rect 516980 46912 517008 46940
rect 143534 46900 143598 46912
rect 44836 46872 143598 46900
rect 143534 46860 143598 46872
rect 200850 46860 200914 46912
rect 248414 46860 248478 46912
rect 297726 46860 297790 46912
rect 309410 46860 309474 46912
rect 352558 46860 352622 46912
rect 364242 46860 364306 46912
rect 407390 46860 407454 46912
rect 419074 46860 419138 46912
rect 462130 46860 462194 46912
rect 473814 46860 473878 46912
rect 516962 46860 517026 46912
rect 42242 45676 42306 45688
rect 140958 45676 141022 45688
rect 42242 45648 141022 45676
rect 42242 45636 42306 45648
rect 140958 45636 141022 45648
rect 186682 45676 186746 45688
rect 194686 45676 194750 45688
rect 186682 45648 194750 45676
rect 186682 45636 186746 45648
rect 194686 45636 194750 45648
rect 523770 45608 523834 45620
rect 673546 45608 673610 45620
rect 523770 45580 673610 45608
rect 523770 45568 523834 45580
rect 673546 45568 673610 45580
rect 44910 45540 44974 45552
rect 195974 45540 196038 45552
rect 44910 45512 196038 45540
rect 44910 45500 44974 45512
rect 195974 45500 196038 45512
rect 518710 45540 518774 45552
rect 673730 45540 673794 45552
rect 518710 45512 673794 45540
rect 518710 45500 518774 45512
rect 673730 45500 673794 45512
rect 349982 44452 350046 44464
rect 359366 44452 359430 44464
rect 414198 44452 414262 44464
rect 188522 44384 188586 44396
rect 192846 44384 192910 44396
rect 201494 44384 201558 44396
rect 188522 44356 201558 44384
rect 188522 44344 188586 44356
rect 192846 44344 192910 44356
rect 201494 44344 201558 44356
rect 195974 44316 196038 44328
rect 195974 44288 204392 44316
rect 195974 44276 196038 44288
rect 201494 44180 201558 44192
rect 204162 44180 204226 44192
rect 201494 44152 204226 44180
rect 204364 44180 204392 44288
rect 349982 44424 414262 44452
rect 349982 44412 350046 44424
rect 359366 44412 359430 44424
rect 414198 44412 414262 44424
rect 360470 44384 360534 44396
rect 406746 44384 406810 44396
rect 360470 44356 406810 44384
rect 360470 44344 360534 44356
rect 406746 44344 406810 44356
rect 468938 44384 469002 44396
rect 523770 44384 523834 44396
rect 468938 44356 523834 44384
rect 468938 44344 469002 44356
rect 523770 44344 523834 44356
rect 305730 44316 305794 44328
rect 351914 44316 351978 44328
rect 305730 44288 351978 44316
rect 305730 44276 305794 44288
rect 351914 44276 351978 44288
rect 295242 44248 295306 44260
rect 303246 44248 303310 44260
rect 295242 44220 303310 44248
rect 295242 44208 295306 44220
rect 303246 44208 303310 44220
rect 406746 44248 406810 44260
rect 461486 44248 461550 44260
rect 516318 44248 516382 44260
rect 518710 44248 518774 44260
rect 406746 44220 518774 44248
rect 406746 44208 406810 44220
rect 461486 44208 461550 44220
rect 516318 44208 516382 44220
rect 518710 44208 518774 44220
rect 304534 44180 304598 44192
rect 349982 44180 350046 44192
rect 204364 44152 350046 44180
rect 201494 44140 201558 44152
rect 204162 44140 204226 44152
rect 304534 44140 304598 44152
rect 349982 44140 350046 44152
rect 350074 44180 350138 44192
rect 358078 44180 358142 44192
rect 350074 44152 358142 44180
rect 350074 44140 350138 44152
rect 358078 44140 358142 44152
rect 414198 44180 414262 44192
rect 468938 44180 469002 44192
rect 414198 44152 469002 44180
rect 414198 44140 414262 44152
rect 468938 44140 469002 44152
rect 576762 42752 576826 42764
rect 673454 42752 673518 42764
rect 576762 42724 673518 42752
rect 576762 42712 576826 42724
rect 673454 42712 673518 42724
rect 297726 42276 297790 42288
rect 300762 42276 300826 42288
rect 297726 42248 300826 42276
rect 297726 42236 297790 42248
rect 300762 42236 300826 42248
rect 305638 42004 305702 42016
rect 299492 41976 305702 42004
rect 299492 41948 299520 41976
rect 305638 41964 305702 41976
rect 352650 42004 352714 42016
rect 355502 42004 355566 42016
rect 352650 41976 355566 42004
rect 352650 41964 352714 41976
rect 355502 41964 355566 41976
rect 356974 42004 357038 42016
rect 359826 42004 359890 42016
rect 361114 42004 361178 42016
rect 356974 41976 361178 42004
rect 356974 41964 357038 41976
rect 359826 41964 359890 41976
rect 361114 41964 361178 41976
rect 189258 41936 189322 41948
rect 191098 41936 191162 41948
rect 192294 41936 192358 41948
rect 193582 41936 193646 41948
rect 196434 41936 196498 41948
rect 189258 41908 196498 41936
rect 189258 41896 189322 41908
rect 191098 41896 191162 41908
rect 192294 41896 192358 41908
rect 193582 41896 193646 41908
rect 196434 41896 196498 41908
rect 198458 41936 198522 41948
rect 200114 41936 200178 41948
rect 198458 41908 200178 41936
rect 198458 41896 198522 41908
rect 200114 41896 200178 41908
rect 297266 41936 297330 41948
rect 299474 41936 299538 41948
rect 297266 41908 299538 41936
rect 297266 41896 297330 41908
rect 299474 41896 299538 41908
rect 302234 41936 302298 41948
rect 305270 41936 305334 41948
rect 306558 41936 306622 41948
rect 308674 41936 308738 41948
rect 302234 41908 308738 41936
rect 302234 41896 302298 41908
rect 305270 41896 305334 41908
rect 306558 41896 306622 41908
rect 308674 41896 308738 41908
rect 352006 41936 352070 41948
rect 354306 41936 354370 41948
rect 360470 41936 360534 41948
rect 352006 41908 360534 41936
rect 361132 41936 361160 41964
rect 363506 41936 363570 41948
rect 361132 41908 363570 41936
rect 352006 41896 352070 41908
rect 354306 41896 354370 41908
rect 360470 41896 360534 41908
rect 363506 41896 363570 41908
rect 407482 41936 407546 41948
rect 410242 41936 410306 41948
rect 411530 41936 411594 41948
rect 414566 41936 414630 41948
rect 415854 41936 415918 41948
rect 418246 41936 418310 41948
rect 407482 41908 418310 41936
rect 407482 41896 407546 41908
rect 410242 41896 410306 41908
rect 411530 41896 411594 41908
rect 414566 41896 414630 41908
rect 415854 41896 415918 41908
rect 418246 41896 418310 41908
rect 462314 41936 462378 41948
rect 465074 41936 465138 41948
rect 466362 41936 466426 41948
rect 469398 41936 469462 41948
rect 470686 41936 470750 41948
rect 473078 41936 473142 41948
rect 462314 41908 473142 41936
rect 462314 41896 462378 41908
rect 465074 41896 465138 41908
rect 466362 41896 466426 41908
rect 469398 41896 469462 41908
rect 470686 41896 470750 41908
rect 473078 41896 473142 41908
rect 517054 41936 517118 41948
rect 519906 41936 519970 41948
rect 521194 41936 521258 41948
rect 524230 41936 524294 41948
rect 525518 41936 525582 41948
rect 527910 41936 527974 41948
rect 517054 41908 527974 41936
rect 517054 41896 517118 41908
rect 519906 41896 519970 41908
rect 521194 41896 521258 41908
rect 524230 41896 524294 41908
rect 525518 41896 525582 41908
rect 527910 41896 527974 41908
rect 146294 41868 146358 41880
rect 569126 41868 569190 41880
rect 576762 41868 576826 41880
rect 146294 41840 576826 41868
rect 146294 41828 146358 41840
rect 569126 41828 569190 41840
rect 576762 41828 576826 41840
rect 198918 41800 198982 41812
rect 307754 41800 307818 41812
rect 362494 41800 362558 41812
rect 168346 41772 380894 41800
rect 93762 41528 93826 41540
rect 168346 41528 168374 41772
rect 198918 41760 198982 41772
rect 307754 41760 307818 41772
rect 362494 41760 362558 41772
rect 93762 41500 168374 41528
rect 93762 41488 93826 41500
tri 239482 41369 239813 41700 se
rect 239813 41369 252469 41700
rect 135162 40236 135226 40248
rect 143534 40236 143598 40248
rect 135162 40208 143598 40236
rect 135162 40196 135226 40208
rect 143534 40196 143598 40208
rect 140990 40100 141054 40112
rect 143066 40100 143130 40112
rect 144546 40100 144610 40112
rect 146294 40100 146358 40112
rect 140990 40072 146358 40100
rect 140990 40060 141054 40072
rect 142586 40000 142614 40072
rect 143066 40060 143130 40072
rect 144546 40060 144610 40072
rect 146294 40060 146358 40072
rect 79664 39616 91393 39806
rect 79664 39593 79892 39616
tri 79892 39593 79915 39616 nw
tri 91107 39593 91130 39616 ne
rect 91130 39593 91393 39616
rect 79076 55 93763 39593
rect 132600 37949 142517 40000
rect 142573 38005 142619 40000
rect 142675 37949 147600 40000
rect 132600 158 147600 37949
rect 186371 0 202429 41369
tri 239013 40900 239482 41369 se
rect 239482 41300 252469 41369
tri 252469 41300 252869 41700 sw
rect 380866 41528 380894 41772
rect 417326 41800 417390 41812
rect 417252 41772 417390 41800
rect 417252 41528 417280 41772
rect 417326 41760 417390 41772
rect 472158 41800 472222 41812
rect 526714 41800 526778 41812
rect 472084 41772 472222 41800
rect 472084 41528 472112 41772
rect 472158 41760 472222 41772
rect 516106 41772 526778 41800
rect 516106 41528 516134 41772
rect 526714 41760 526778 41772
rect 380866 41500 516134 41528
rect 239482 40900 252869 41300
rect 239013 40196 252869 40900
rect 239013 39796 252469 40196
tri 252469 39796 252869 40196 nw
rect 239013 39756 252101 39796
rect 239013 32702 240960 39756
rect 244887 39600 252101 39756
rect 244887 39593 252869 39600
rect 238961 31928 241151 32702
rect 241200 32 256176 39593
rect 294971 0 311029 41369
rect 349771 0 365829 41369
rect 404571 0 420629 41369
rect 459371 0 475429 41369
rect 514171 0 530229 41369
rect 569864 39616 581593 39806
rect 569864 39593 570092 39616
tri 570092 39593 570115 39616 nw
tri 581307 39593 581330 39616 ne
rect 581330 39593 581593 39616
rect 623664 39616 635393 39806
rect 623664 39593 623892 39616
tri 623892 39593 623915 39616 nw
tri 635107 39593 635130 39616 ne
rect 635130 39593 635393 39616
rect 636029 39593 637075 39774
rect 569276 55 583963 39593
rect 623217 55 637763 39593
<< metal2 >>
rect 77049 995407 77105 995887
rect 77693 995407 77749 995887
rect 78337 995407 78393 995887
rect 78889 995452 78945 995887
rect 78876 995407 78945 995452
rect 80177 995407 80233 995887
rect 80729 995407 80785 995887
rect 81373 995407 81429 995887
rect 82017 995407 82073 995887
rect 83213 995452 83269 995887
rect 83200 995407 83269 995452
rect 84501 995407 84557 995887
rect 85053 995407 85109 995887
rect 85697 995407 85753 995887
rect 86341 995407 86397 995887
rect 87537 995407 87593 995887
rect 88733 995407 88789 995887
rect 89377 995407 89433 995887
rect 91217 995407 91273 995887
rect 128449 995407 128505 995887
rect 129093 995407 129149 995887
rect 129737 995407 129793 995887
rect 130289 995407 130345 995887
rect 131577 995407 131633 995887
rect 132129 995407 132185 995887
rect 132773 995407 132829 995887
rect 133417 995407 133473 995887
rect 134613 995407 134669 995887
rect 135901 995407 135957 995887
rect 136453 995407 136509 995887
rect 137097 995407 137153 995887
rect 137741 995407 137797 995887
rect 138937 995407 138993 995887
rect 140133 995407 140189 995887
rect 140777 995407 140833 995887
rect 142617 995407 142673 995887
rect 179849 995407 179905 995887
rect 180493 995407 180549 995887
rect 181137 995407 181193 995887
rect 181689 995466 181745 995887
rect 181689 995407 181760 995466
rect 182977 995407 183033 995887
rect 183529 995407 183585 995887
rect 184173 995407 184229 995887
rect 184817 995407 184873 995887
rect 186013 995466 186069 995887
rect 186013 995407 186084 995466
rect 187301 995407 187357 995887
rect 187853 995407 187909 995887
rect 188497 995407 188553 995887
rect 189141 995407 189197 995887
rect 190337 995407 190393 995887
rect 191533 995407 191589 995887
rect 192177 995407 192233 995887
rect 194017 995407 194073 995887
rect 231249 995407 231305 995887
rect 231893 995407 231949 995887
rect 232537 995407 232593 995887
rect 233089 995466 233145 995887
rect 233068 995407 233145 995466
rect 234377 995407 234433 995887
rect 234929 995407 234985 995887
rect 235573 995407 235629 995887
rect 236217 995407 236273 995887
rect 237413 995466 237469 995887
rect 237392 995407 237469 995466
rect 238701 995407 238757 995887
rect 239253 995407 239309 995887
rect 239897 995407 239953 995887
rect 240541 995407 240597 995887
rect 241737 995407 241793 995887
rect 242933 995407 242989 995887
rect 243577 995407 243633 995887
rect 245417 995407 245473 995887
rect 282849 995407 282905 995887
rect 283493 995407 283549 995887
rect 284137 995407 284193 995887
rect 284689 995452 284745 995887
rect 284680 995407 284745 995452
rect 285977 995407 286033 995887
rect 286529 995407 286585 995887
rect 287173 995407 287229 995887
rect 287817 995407 287873 995887
rect 289013 995452 289069 995887
rect 289004 995407 289069 995452
rect 290301 995407 290357 995887
rect 290853 995407 290909 995887
rect 291497 995407 291553 995887
rect 292141 995407 292197 995887
rect 293337 995407 293393 995887
rect 294533 995407 294589 995887
rect 295177 995407 295233 995887
rect 297017 995407 297073 995887
rect 78876 990622 78904 995407
rect 78864 990616 78916 990622
rect 78864 990558 78916 990564
rect 78876 990282 78904 990558
rect 42340 990276 42392 990282
rect 42340 990218 42392 990224
rect 78864 990276 78916 990282
rect 78864 990218 78916 990224
rect 41713 969217 42193 969273
rect 41713 967377 42193 967433
rect 41713 966733 42193 966789
rect 41713 965537 42193 965593
rect 41713 964341 42193 964397
rect 41713 963697 42193 963753
rect 41713 963053 42193 963109
rect 41713 962501 42193 962557
rect 41713 961213 42193 961269
rect 41800 961178 41828 961213
rect 41788 961172 41840 961178
rect 41788 961114 41840 961120
rect 41713 960017 42193 960073
rect 41713 959373 42193 959429
rect 41713 958729 42193 958785
rect 41713 958177 42193 958233
rect 42352 969626 42380 990218
rect 83200 990622 83228 995407
rect 83188 990616 83240 990622
rect 83188 990558 83240 990564
rect 130304 990622 130332 995407
rect 134628 990622 134656 995407
rect 130292 990616 130344 990622
rect 130292 990558 130344 990564
rect 134616 990616 134668 990622
rect 134616 990558 134668 990564
rect 181732 990622 181760 995407
rect 181720 990616 181772 990622
rect 181720 990558 181772 990564
rect 186056 990622 186084 995407
rect 186044 990616 186096 990622
rect 186044 990558 186096 990564
rect 233068 990622 233096 995407
rect 233056 990616 233108 990622
rect 233056 990558 233108 990564
rect 237392 990622 237420 995407
rect 284680 990690 284708 995407
rect 274732 990684 274784 990690
rect 274652 990644 274732 990672
rect 237380 990616 237432 990622
rect 237380 990558 237432 990564
rect 274456 990616 274508 990622
rect 274652 990570 274680 990644
rect 274732 990626 274784 990632
rect 284668 990684 284720 990690
rect 284668 990626 284720 990632
rect 274508 990564 274680 990570
rect 274456 990558 274680 990564
rect 274468 990542 274680 990558
rect 289004 990690 289032 995407
rect 288992 990684 289044 990690
rect 288992 990626 289044 990632
rect 384649 995407 384705 995887
rect 385293 995407 385349 995887
rect 385937 995407 385993 995887
rect 386489 995452 386545 995887
rect 386489 995407 386552 995452
rect 387777 995407 387833 995887
rect 388329 995407 388385 995887
rect 388973 995407 389029 995887
rect 389617 995407 389673 995887
rect 390813 995452 390869 995887
rect 390813 995407 390876 995452
rect 392101 995407 392157 995887
rect 392653 995407 392709 995887
rect 393297 995407 393353 995887
rect 393941 995407 393997 995887
rect 395137 995407 395193 995887
rect 396333 995407 396389 995887
rect 396977 995407 397033 995887
rect 398817 995407 398873 995887
rect 473649 995407 473705 995887
rect 474293 995407 474349 995887
rect 474937 995407 474993 995887
rect 475489 995452 475545 995887
rect 475488 995407 475545 995452
rect 476777 995407 476833 995887
rect 477329 995407 477385 995887
rect 477973 995407 478029 995887
rect 478617 995407 478673 995887
rect 479813 995452 479869 995887
rect 479812 995407 479869 995452
rect 481101 995407 481157 995887
rect 481653 995407 481709 995887
rect 482297 995407 482353 995887
rect 482941 995407 482997 995887
rect 484137 995407 484193 995887
rect 485333 995407 485389 995887
rect 485977 995407 486033 995887
rect 487817 995407 487873 995887
rect 525049 995407 525105 995887
rect 525693 995407 525749 995887
rect 526337 995407 526393 995887
rect 526889 995407 526945 995887
rect 528177 995407 528233 995887
rect 528729 995407 528785 995887
rect 529373 995407 529429 995887
rect 530017 995407 530073 995887
rect 531213 995407 531269 995887
rect 532501 995407 532557 995887
rect 533053 995407 533109 995887
rect 533697 995407 533753 995887
rect 534341 995407 534397 995887
rect 535537 995407 535593 995887
rect 536733 995407 536789 995887
rect 537377 995407 537433 995887
rect 539217 995407 539273 995887
rect 386524 990622 386552 995407
rect 386512 990616 386564 990622
rect 386512 990558 386564 990564
rect 390848 990622 390876 995407
rect 475488 990622 475516 995407
rect 390836 990616 390888 990622
rect 390836 990558 390888 990564
rect 475476 990616 475528 990622
rect 475476 990558 475528 990564
rect 479812 990622 479840 995407
rect 479800 990616 479852 990622
rect 479800 990558 479852 990564
rect 526916 990622 526944 995407
rect 526904 990616 526956 990622
rect 526904 990558 526956 990564
rect 531240 990622 531268 995407
rect 626849 995407 626905 995887
rect 627493 995407 627549 995887
rect 628137 995407 628193 995887
rect 628689 995466 628745 995887
rect 628668 995407 628745 995466
rect 629977 995407 630033 995887
rect 630529 995407 630585 995887
rect 631173 995407 631229 995887
rect 631817 995407 631873 995887
rect 633013 995466 633069 995887
rect 632992 995407 633069 995466
rect 634301 995407 634357 995887
rect 634853 995407 634909 995887
rect 635497 995407 635553 995887
rect 636141 995407 636197 995887
rect 637337 995407 637393 995887
rect 638533 995407 638589 995887
rect 639177 995407 639233 995887
rect 641017 995407 641073 995887
rect 628668 990622 628696 995407
rect 531228 990616 531280 990622
rect 531228 990558 531280 990564
rect 628656 990616 628708 990622
rect 628656 990558 628708 990564
rect 632992 990622 633020 995407
rect 632980 990616 633032 990622
rect 632980 990558 633032 990564
rect 634728 990616 634780 990622
rect 634728 990558 634780 990564
rect 634740 990146 634768 990558
rect 634728 990140 634780 990146
rect 634728 990082 634780 990088
rect 42352 969598 42564 969626
rect 42536 961178 42564 969598
rect 42524 961172 42576 961178
rect 42524 961114 42576 961120
rect 41713 956889 42193 956945
rect 41800 956842 41828 956889
rect 42536 956842 42564 961114
rect 41800 956814 42564 956842
rect 41713 956337 42193 956393
rect 41713 955693 42193 955749
rect 41713 955049 42193 955105
rect 42260 941174 42288 956814
rect 42260 941146 42564 941174
rect 41713 799417 42193 799473
rect 41713 797577 42193 797633
rect 41713 796933 42193 796989
rect 41713 795737 42193 795793
rect 41713 794541 42193 794597
rect 41713 793897 42193 793953
rect 41713 793253 42193 793309
rect 41713 792701 42193 792757
rect 41788 791988 41840 791994
rect 41788 791930 41840 791936
rect 41800 791469 41828 791930
rect 41713 791413 42193 791469
rect 41713 790217 42193 790273
rect 41713 789573 42193 789629
rect 41713 788929 42193 788985
rect 41713 788377 42193 788433
rect 41713 787089 42193 787145
rect 41722 787086 41828 787089
rect 41800 787030 41828 787086
rect 41788 787024 41840 787030
rect 41788 786966 41840 786972
rect 41713 786537 42193 786593
rect 41713 785893 42193 785949
rect 41713 785249 42193 785305
rect 41713 756217 42193 756273
rect 41713 754377 42193 754433
rect 41713 753733 42193 753789
rect 41713 752537 42193 752593
rect 41713 751341 42193 751397
rect 41713 750697 42193 750753
rect 41713 750053 42193 750109
rect 41713 749501 42193 749557
rect 41713 748213 42193 748269
rect 41984 747930 42012 748213
rect 41972 747924 42024 747930
rect 41972 747866 42024 747872
rect 42536 791994 42564 941146
rect 673644 960084 673696 960090
rect 673644 960026 673696 960032
rect 673656 875838 673684 960026
rect 673828 990140 673880 990146
rect 673828 990082 673880 990088
rect 673840 965326 673868 990082
rect 673828 965320 673880 965326
rect 673828 965262 673880 965268
rect 673644 875832 673696 875838
rect 673644 875774 673696 875780
rect 42524 791988 42576 791994
rect 42524 791930 42576 791936
rect 42536 787658 42564 791930
rect 42444 787630 42564 787658
rect 42444 787030 42472 787630
rect 42432 787024 42484 787030
rect 42432 786966 42484 786972
rect 42444 756634 42472 786966
rect 42432 756628 42484 756634
rect 42432 756570 42484 756576
rect 42432 756424 42484 756430
rect 42432 756366 42484 756372
rect 42444 749306 42472 756366
rect 42352 749278 42472 749306
rect 42352 747930 42380 749278
rect 42340 747924 42392 747930
rect 42340 747866 42392 747872
rect 41713 747017 42193 747073
rect 41713 746373 42193 746429
rect 41713 745729 42193 745785
rect 41713 745177 42193 745233
rect 41713 743889 42193 743945
rect 41800 743510 41828 743889
rect 41788 743504 41840 743510
rect 41788 743446 41840 743452
rect 41713 743337 42193 743393
rect 41713 742693 42193 742749
rect 41713 742049 42193 742105
rect 42352 743510 42380 747866
rect 42340 743504 42392 743510
rect 42340 743446 42392 743452
rect 42352 719098 42380 743446
rect 42340 719092 42392 719098
rect 42340 719034 42392 719040
rect 42340 718888 42392 718894
rect 42340 718830 42392 718836
rect 41713 713017 42193 713073
rect 41713 711177 42193 711233
rect 41713 710533 42193 710589
rect 41713 709337 42193 709393
rect 41713 708141 42193 708197
rect 41713 707497 42193 707553
rect 41713 706853 42193 706909
rect 41713 706301 42193 706357
rect 41713 705013 42193 705069
rect 41892 704970 41920 705013
rect 42352 704970 42380 718830
rect 41892 704942 42380 704970
rect 41713 703817 42193 703873
rect 41713 703173 42193 703229
rect 41713 702529 42193 702585
rect 41713 701977 42193 702033
rect 41722 700745 41920 700754
rect 41713 700689 42193 700745
rect 41892 700618 41920 700689
rect 42260 700618 42288 704942
rect 673828 871344 673880 871350
rect 673828 871286 673880 871292
rect 673840 786010 673868 871286
rect 673828 786004 673880 786010
rect 673828 785946 673880 785952
rect 41892 700590 42288 700618
rect 41713 700137 42193 700193
rect 41713 699493 42193 699549
rect 41713 698849 42193 698905
rect 42260 690014 42288 700590
rect 42260 689986 42380 690014
rect 41713 669817 42193 669873
rect 41713 667977 42193 668033
rect 41713 667333 42193 667389
rect 41713 666137 42193 666193
rect 41713 664941 42193 664997
rect 41713 664297 42193 664353
rect 41713 663653 42193 663709
rect 41713 663101 42193 663157
rect 42352 661994 42380 689986
rect 41800 661966 42380 661994
rect 41800 661869 41828 661966
rect 41713 661813 42193 661869
rect 41713 660617 42193 660673
rect 41713 659973 42193 660029
rect 41713 659329 42193 659385
rect 41713 658777 42193 658833
rect 42260 657642 42288 661966
rect 673736 781652 673788 781658
rect 673736 781594 673788 781600
rect 673748 740994 673776 781594
rect 673736 740988 673788 740994
rect 673736 740930 673788 740936
rect 41892 657614 42288 657642
rect 41892 657545 41920 657614
rect 41713 657489 42193 657545
rect 41722 657478 41920 657489
rect 41713 656937 42193 656993
rect 41713 656293 42193 656349
rect 41713 655649 42193 655705
rect 42260 651374 42288 657614
rect 42260 651346 42380 651374
rect 41713 626617 42193 626673
rect 41713 624777 42193 624833
rect 41713 624133 42193 624189
rect 41713 622937 42193 622993
rect 41713 621741 42193 621797
rect 41713 621097 42193 621153
rect 41713 620453 42193 620509
rect 41713 619901 42193 619957
rect 42352 618746 42380 651346
rect 41800 618718 42380 618746
rect 41800 618669 41828 618718
rect 41713 618613 42193 618669
rect 41713 617417 42193 617473
rect 41713 616773 42193 616829
rect 41713 616129 42193 616185
rect 41713 615577 42193 615633
rect 41713 614331 42193 614345
rect 42260 614331 42288 618718
rect 41713 614303 42288 614331
rect 41713 614289 42193 614303
rect 41713 613737 42193 613793
rect 41713 613093 42193 613149
rect 42260 612734 42288 614303
rect 42260 612706 42380 612734
rect 41713 612449 42193 612505
rect 41713 583417 42193 583473
rect 41713 581577 42193 581633
rect 41713 580933 42193 580989
rect 41713 579737 42193 579793
rect 41713 578541 42193 578597
rect 41713 577897 42193 577953
rect 41713 577253 42193 577309
rect 41713 576701 42193 576757
rect 41713 575455 42193 575469
rect 42352 575455 42380 612706
rect 673736 737044 673788 737050
rect 673736 736986 673788 736992
rect 673748 695978 673776 736986
rect 673736 695972 673788 695978
rect 673736 695914 673788 695920
rect 41713 575427 42380 575455
rect 41713 575413 42193 575427
rect 41713 574217 42193 574273
rect 41713 573573 42193 573629
rect 41713 572929 42193 572985
rect 41713 572377 42193 572433
rect 42260 571282 42288 575427
rect 41800 571254 42380 571282
rect 41800 571146 41828 571254
rect 41722 571145 41828 571146
rect 41713 571089 42193 571145
rect 41713 570537 42193 570593
rect 41713 569893 42193 569949
rect 41713 569249 42193 569305
rect 41713 540217 42193 540273
rect 41713 538377 42193 538433
rect 41713 537733 42193 537789
rect 41713 536537 42193 536593
rect 41713 535341 42193 535397
rect 41713 534697 42193 534753
rect 41713 534053 42193 534109
rect 41713 533501 42193 533557
rect 41713 532213 42193 532269
rect 41892 532114 41920 532213
rect 42352 532114 42380 571254
rect 41892 532086 42380 532114
rect 41713 531017 42193 531073
rect 41713 530373 42193 530429
rect 41713 529729 42193 529785
rect 41713 529177 42193 529233
rect 41713 527917 42193 527945
rect 41708 527898 42193 527917
rect 42260 527898 42288 532086
rect 673736 692096 673788 692102
rect 673736 692038 673788 692044
rect 673748 651166 673776 692038
rect 673736 651160 673788 651166
rect 673736 651102 673788 651108
rect 673748 646474 673776 651102
rect 673736 646468 673788 646474
rect 673736 646410 673788 646416
rect 673748 605810 673776 646410
rect 673736 605804 673788 605810
rect 673736 605746 673788 605752
rect 673736 601860 673788 601866
rect 673736 601802 673788 601808
rect 673748 561270 673776 601802
rect 673736 561264 673788 561270
rect 673736 561206 673788 561212
rect 41708 527870 42288 527898
rect 41713 527337 42193 527393
rect 41713 526693 42193 526749
rect 41713 526049 42193 526105
rect 42260 419534 42288 527870
rect 42260 419506 42380 419534
rect 41713 412617 42193 412673
rect 41713 410777 42193 410833
rect 41713 410133 42193 410189
rect 41713 408937 42193 408993
rect 41713 407741 42193 407797
rect 41713 407097 42193 407153
rect 41713 406453 42193 406509
rect 41713 405901 42193 405957
rect 42352 405226 42380 419506
rect 41800 405198 42380 405226
rect 41800 404682 41828 405198
rect 41722 404669 41828 404682
rect 41713 404613 42193 404669
rect 41713 403417 42193 403473
rect 41713 402773 42193 402829
rect 41713 402129 42193 402185
rect 41713 401577 42193 401633
rect 41713 400330 42193 400345
rect 42260 400330 42288 405198
rect 41713 400302 42288 400330
rect 41713 400289 42193 400302
rect 41713 399737 42193 399793
rect 41713 399093 42193 399149
rect 41713 398449 42193 398505
rect 41713 369417 42193 369473
rect 41713 367577 42193 367633
rect 41713 366933 42193 366989
rect 41713 365737 42193 365793
rect 41713 364541 42193 364597
rect 41713 363897 42193 363953
rect 41713 363253 42193 363309
rect 41713 362701 42193 362757
rect 41713 361434 42193 361469
rect 42260 361434 42288 400302
rect 41713 361413 42288 361434
rect 41722 361406 42288 361413
rect 41713 360217 42193 360273
rect 41713 359573 42193 359629
rect 41713 358929 42193 358985
rect 41713 358377 42193 358433
rect 41713 357089 42193 357145
rect 41984 356674 42012 357089
rect 42260 356674 42288 361406
rect 41984 356646 42288 356674
rect 41713 356537 42193 356593
rect 41713 355893 42193 355949
rect 41713 355249 42193 355305
rect 42260 332602 42288 356646
rect 42260 332574 42380 332602
rect 41713 326217 42193 326273
rect 41713 324377 42193 324433
rect 41713 323733 42193 323789
rect 41713 322537 42193 322593
rect 41713 321341 42193 321397
rect 41713 320697 42193 320753
rect 41713 320053 42193 320109
rect 41713 319501 42193 319557
rect 41713 318255 42193 318269
rect 42352 318255 42380 332574
rect 41713 318227 42380 318255
rect 41713 318213 42193 318227
rect 41713 317017 42193 317073
rect 41713 316373 42193 316429
rect 41713 315729 42193 315785
rect 41713 315177 42193 315233
rect 41713 313889 42193 313945
rect 41800 313834 41828 313889
rect 42260 313834 42288 318227
rect 673644 379092 673696 379098
rect 673644 379034 673696 379040
rect 673656 338842 673684 379034
rect 673644 338836 673696 338842
rect 673644 338778 673696 338784
rect 41800 313806 42288 313834
rect 41713 313337 42193 313393
rect 41713 312693 42193 312749
rect 41713 312049 42193 312105
rect 42260 303614 42288 313806
rect 42260 303586 42380 303614
rect 41713 283017 42193 283073
rect 41713 281177 42193 281233
rect 41713 280533 42193 280589
rect 41713 279337 42193 279393
rect 41713 278141 42193 278197
rect 41713 277497 42193 277553
rect 41713 276853 42193 276909
rect 41713 276301 42193 276357
rect 42352 275210 42380 303586
rect 41800 275182 42380 275210
rect 41800 275074 41828 275182
rect 41722 275069 41828 275074
rect 41713 275013 42193 275069
rect 41713 273817 42193 273873
rect 41713 273173 42193 273229
rect 41713 272529 42193 272585
rect 41713 271977 42193 272033
rect 42260 270858 42288 275182
rect 41892 270830 42288 270858
rect 41892 270745 41920 270830
rect 41713 270689 42193 270745
rect 41713 270137 42193 270193
rect 41713 269493 42193 269549
rect 41713 268849 42193 268905
rect 42260 264974 42288 270830
rect 42260 264946 42380 264974
rect 41713 239817 42193 239873
rect 41713 237977 42193 238033
rect 41713 236137 42193 236193
rect 41713 234941 42193 234997
rect 41713 234297 42193 234353
rect 41713 233653 42193 233709
rect 41713 233101 42193 233157
rect 41713 231855 42193 231869
rect 42352 231855 42380 264946
rect 41713 231827 42380 231855
rect 41713 231813 42193 231827
rect 41713 230617 42193 230673
rect 41713 229973 42193 230029
rect 41713 229329 42193 229385
rect 41713 228777 42193 228833
rect 42260 227610 42288 231827
rect 41800 227582 42380 227610
rect 41800 227545 41828 227582
rect 41713 227489 42193 227545
rect 41713 226937 42193 226993
rect 41713 226293 42193 226349
rect 41713 225649 42193 225705
rect 42352 197538 42380 227582
rect 675407 966695 675887 966751
rect 675407 966051 675887 966107
rect 675407 965407 675887 965463
rect 675392 965320 675444 965326
rect 675392 965262 675444 965268
rect 675404 964911 675432 965262
rect 675404 964897 675887 964911
rect 675312 964869 675887 964897
rect 675312 960573 675340 964869
rect 675407 964855 675887 964869
rect 675407 963567 675887 963623
rect 675407 963015 675887 963071
rect 675407 962371 675887 962427
rect 675407 961727 675887 961783
rect 675407 960573 675887 960587
rect 675312 960545 675887 960573
rect 675404 960531 675887 960545
rect 675404 960090 675432 960531
rect 675392 960084 675444 960090
rect 675392 960026 675444 960032
rect 675407 959243 675887 959299
rect 675407 958691 675887 958747
rect 675407 958047 675887 958103
rect 675407 957403 675887 957459
rect 675407 956207 675887 956263
rect 675407 955011 675887 955067
rect 675407 954367 675887 954423
rect 675407 952527 675887 952583
rect 675407 877495 675887 877551
rect 675407 876851 675887 876907
rect 675407 876207 675887 876263
rect 675392 875832 675444 875838
rect 675392 875774 675444 875780
rect 675404 875711 675432 875774
rect 675404 875697 675887 875711
rect 675312 875669 675887 875697
rect 675312 871373 675340 875669
rect 675407 875655 675887 875669
rect 675407 874367 675887 874423
rect 675407 873815 675887 873871
rect 675407 873171 675887 873227
rect 675407 872527 675887 872583
rect 675407 871373 675887 871387
rect 675312 871350 675887 871373
rect 675300 871345 675887 871350
rect 675300 871344 675352 871345
rect 675407 871331 675887 871345
rect 675300 871286 675352 871292
rect 675407 870043 675887 870099
rect 675407 869491 675887 869547
rect 675407 868847 675887 868903
rect 675407 868203 675887 868259
rect 675407 867007 675887 867063
rect 675407 865811 675887 865867
rect 675407 865167 675887 865223
rect 675407 863327 675887 863383
rect 675407 788295 675887 788351
rect 675407 787651 675887 787707
rect 675407 787007 675887 787063
rect 675407 786483 675887 786511
rect 675404 786455 675887 786483
rect 675404 786010 675432 786455
rect 675208 786004 675260 786010
rect 675208 785946 675260 785952
rect 675392 786004 675444 786010
rect 675392 785946 675444 785952
rect 675220 781658 675248 785946
rect 675407 785167 675887 785223
rect 675407 784615 675887 784671
rect 675407 783971 675887 784027
rect 675407 783327 675887 783383
rect 675407 782159 675887 782187
rect 675404 782131 675887 782159
rect 675404 781658 675432 782131
rect 675208 781652 675260 781658
rect 675208 781594 675260 781600
rect 675392 781652 675444 781658
rect 675392 781594 675444 781600
rect 675407 780843 675887 780899
rect 675407 780291 675887 780347
rect 675407 779647 675887 779703
rect 675407 779003 675887 779059
rect 675407 777807 675887 777863
rect 675407 776611 675887 776667
rect 675407 775967 675887 776023
rect 675407 774127 675887 774183
rect 675407 743295 675887 743351
rect 675407 742651 675887 742707
rect 675407 742007 675887 742063
rect 675407 741483 675887 741511
rect 675404 741455 675887 741483
rect 675404 740994 675432 741455
rect 675208 740988 675260 740994
rect 675208 740930 675260 740936
rect 675392 740988 675444 740994
rect 675392 740930 675444 740936
rect 675220 737050 675248 740930
rect 675407 740167 675887 740223
rect 675407 739615 675887 739671
rect 675407 738971 675887 739027
rect 675407 738327 675887 738383
rect 675407 737159 675887 737187
rect 675404 737131 675887 737159
rect 675404 737050 675432 737131
rect 675208 737044 675260 737050
rect 675208 736986 675260 736992
rect 675392 737044 675444 737050
rect 675392 736986 675444 736992
rect 675407 735843 675887 735899
rect 675407 735291 675887 735347
rect 675407 734647 675887 734703
rect 675407 734003 675887 734059
rect 675407 732807 675887 732863
rect 675407 731611 675887 731667
rect 675407 730967 675887 731023
rect 675407 729127 675887 729183
rect 675407 698295 675887 698351
rect 675407 697651 675887 697707
rect 675407 697007 675887 697063
rect 675407 696483 675887 696511
rect 675404 696455 675887 696483
rect 675404 695978 675432 696455
rect 675208 695972 675260 695978
rect 675208 695914 675260 695920
rect 675392 695972 675444 695978
rect 675392 695914 675444 695920
rect 675220 692102 675248 695914
rect 675407 695167 675887 695223
rect 675407 694615 675887 694671
rect 675407 693971 675887 694027
rect 675407 693327 675887 693383
rect 675407 692172 675887 692187
rect 675404 692131 675887 692172
rect 675404 692102 675432 692131
rect 675208 692096 675260 692102
rect 675208 692038 675260 692044
rect 675392 692096 675444 692102
rect 675392 692038 675444 692044
rect 675407 690843 675887 690899
rect 675407 690291 675887 690347
rect 675407 689647 675887 689703
rect 675407 689003 675887 689059
rect 675407 687807 675887 687863
rect 675407 686611 675887 686667
rect 675407 685967 675887 686023
rect 675407 684127 675887 684183
rect 675407 653095 675887 653151
rect 675407 652451 675887 652507
rect 675407 651807 675887 651863
rect 675407 651283 675887 651311
rect 675404 651255 675887 651283
rect 675404 651166 675432 651255
rect 675392 651160 675444 651166
rect 675392 651102 675444 651108
rect 675407 649967 675887 650023
rect 675407 649415 675887 649471
rect 675407 648771 675887 648827
rect 675407 648127 675887 648183
rect 675407 646959 675887 646987
rect 675404 646931 675887 646959
rect 675404 646474 675432 646931
rect 675392 646468 675444 646474
rect 675392 646410 675444 646416
rect 675407 645643 675887 645699
rect 675407 645091 675887 645147
rect 675407 644447 675887 644503
rect 675407 643803 675887 643859
rect 675407 642607 675887 642663
rect 675407 641411 675887 641467
rect 675407 640767 675887 640823
rect 675407 638927 675887 638983
rect 675407 608095 675887 608151
rect 675407 607451 675887 607507
rect 675407 606807 675887 606863
rect 675407 606283 675887 606311
rect 675404 606255 675887 606283
rect 675404 605810 675432 606255
rect 675208 605804 675260 605810
rect 675208 605746 675260 605752
rect 675392 605804 675444 605810
rect 675392 605746 675444 605752
rect 675220 601866 675248 605746
rect 675407 604967 675887 605023
rect 675407 604415 675887 604471
rect 675407 603771 675887 603827
rect 675407 603127 675887 603183
rect 675407 601959 675887 601987
rect 675404 601931 675887 601959
rect 675404 601866 675432 601931
rect 675208 601860 675260 601866
rect 675208 601802 675260 601808
rect 675392 601860 675444 601866
rect 675392 601802 675444 601808
rect 675407 600643 675887 600699
rect 675407 600091 675887 600147
rect 675407 599447 675887 599503
rect 675407 598803 675887 598859
rect 675407 597607 675887 597663
rect 675407 596411 675887 596467
rect 675407 595767 675887 595823
rect 675407 593927 675887 593983
rect 675407 562895 675887 562951
rect 675407 562251 675887 562307
rect 675407 561607 675887 561663
rect 675208 561264 675260 561270
rect 675208 561206 675260 561212
rect 675392 561264 675444 561270
rect 675392 561206 675444 561212
rect 675220 557326 675248 561206
rect 675404 561111 675432 561206
rect 675404 561068 675887 561111
rect 675407 561055 675887 561068
rect 675407 559767 675887 559823
rect 675407 559215 675887 559271
rect 675407 558571 675887 558627
rect 675407 557927 675887 557983
rect 675208 557320 675260 557326
rect 675208 557262 675260 557268
rect 675392 557320 675444 557326
rect 675392 557262 675444 557268
rect 675404 556787 675432 557262
rect 675404 556759 675887 556787
rect 675407 556731 675887 556759
rect 675407 555443 675887 555499
rect 675407 554891 675887 554947
rect 675407 554247 675887 554303
rect 675407 553603 675887 553659
rect 675407 552407 675887 552463
rect 675407 551211 675887 551267
rect 675407 550567 675887 550623
rect 675407 548727 675887 548783
rect 675407 385695 675887 385751
rect 675407 385051 675887 385107
rect 675407 384407 675887 384463
rect 675312 383982 675432 384010
rect 675312 379573 675340 383982
rect 675404 383911 675432 383982
rect 675404 383860 675887 383911
rect 675407 383855 675887 383860
rect 675407 382567 675887 382623
rect 675407 382015 675887 382071
rect 675407 381371 675887 381427
rect 675407 380727 675887 380783
rect 675407 379573 675887 379587
rect 675312 379545 675887 379573
rect 675404 379531 675887 379545
rect 675404 379098 675432 379531
rect 675392 379092 675444 379098
rect 675392 379034 675444 379040
rect 675407 378243 675887 378299
rect 675407 377691 675887 377747
rect 675407 377047 675887 377103
rect 675407 376403 675887 376459
rect 675407 375207 675887 375263
rect 675407 373367 675887 373423
rect 675407 371527 675887 371583
rect 675407 340495 675887 340551
rect 675407 339851 675887 339907
rect 675407 339207 675887 339263
rect 675392 338836 675444 338842
rect 675392 338778 675444 338784
rect 675404 338711 675432 338778
rect 675404 338655 675887 338711
rect 675404 338178 675432 338655
rect 675312 338150 675432 338178
rect 675312 334370 675340 338150
rect 675407 337367 675887 337423
rect 675407 336815 675887 336871
rect 675407 336171 675887 336227
rect 675407 335527 675887 335583
rect 675407 334370 675887 334387
rect 675312 334342 675887 334370
rect 675404 334331 675887 334342
rect 675404 334286 675432 334331
rect 673828 334280 673880 334286
rect 673828 334222 673880 334228
rect 675392 334280 675444 334286
rect 675392 334222 675444 334228
rect 673840 293758 673868 334222
rect 675407 333043 675887 333099
rect 675407 332491 675887 332547
rect 675407 331847 675887 331903
rect 675407 331203 675887 331259
rect 675407 330007 675887 330063
rect 675407 328167 675887 328223
rect 675407 326327 675887 326383
rect 675407 295495 675887 295551
rect 675407 294851 675887 294907
rect 675407 294207 675887 294263
rect 675312 293758 675340 293789
rect 673828 293752 673880 293758
rect 673828 293694 673880 293700
rect 675300 293752 675352 293758
rect 675407 293706 675887 293711
rect 675352 293700 675887 293706
rect 675300 293694 675887 293700
rect 675312 293678 675887 293694
rect 675312 289354 675340 293678
rect 675407 293655 675887 293678
rect 675407 292367 675887 292423
rect 675407 291815 675887 291871
rect 675407 291171 675887 291227
rect 675407 290527 675887 290583
rect 675407 289354 675887 289387
rect 675312 289331 675887 289354
rect 675312 289326 675432 289331
rect 675404 288862 675432 289326
rect 673736 288856 673788 288862
rect 673736 288798 673788 288804
rect 675392 288856 675444 288862
rect 675392 288798 675444 288804
rect 673748 249150 673776 288798
rect 673736 249144 673788 249150
rect 673736 249086 673788 249092
rect 675407 288043 675887 288099
rect 675407 287491 675887 287547
rect 675407 286847 675887 286903
rect 675407 286203 675887 286259
rect 675407 285007 675887 285063
rect 675407 283167 675887 283223
rect 675407 281327 675887 281383
rect 675407 250495 675887 250551
rect 675407 249851 675887 249907
rect 675407 249207 675887 249263
rect 675392 249144 675444 249150
rect 675392 249086 675444 249092
rect 675404 248711 675432 249086
rect 675404 248690 675887 248711
rect 675312 248662 675887 248690
rect 42340 197532 42392 197538
rect 42340 197474 42392 197480
rect 42340 197328 42392 197334
rect 42340 197270 42392 197276
rect 41713 196617 42193 196673
rect 41713 194777 42193 194833
rect 41713 192937 42193 192993
rect 41713 191741 42193 191797
rect 41713 191097 42193 191153
rect 41713 190453 42193 190509
rect 41713 189901 42193 189957
rect 42352 188850 42380 197270
rect 41800 188822 42380 188850
rect 41800 188669 41828 188822
rect 41713 188613 42193 188669
rect 41713 187417 42193 187473
rect 41713 186773 42193 186829
rect 41713 186129 42193 186185
rect 41713 185577 42193 185633
rect 41713 184331 42193 184345
rect 42260 184331 42288 188822
rect 41713 184303 42380 184331
rect 41713 184289 42193 184303
rect 41713 183737 42193 183793
rect 41713 183093 42193 183149
rect 41713 182449 42193 182505
rect 42352 45626 42380 184303
rect 673736 243840 673788 243846
rect 673736 243782 673788 243788
rect 673748 203522 673776 243782
rect 673736 203516 673788 203522
rect 673736 203458 673788 203464
rect 673736 199096 673788 199102
rect 673736 199038 673788 199044
rect 673748 158642 673776 199038
rect 675312 244373 675340 248662
rect 675407 248655 675887 248662
rect 675407 247367 675887 247423
rect 675407 246815 675887 246871
rect 675407 246171 675887 246227
rect 675407 245527 675887 245583
rect 675407 244373 675887 244387
rect 675312 244345 675887 244373
rect 675404 244331 675887 244345
rect 675404 243846 675432 244331
rect 675392 243840 675444 243846
rect 675392 243782 675444 243788
rect 675407 243043 675887 243099
rect 675407 242491 675887 242547
rect 675407 241847 675887 241903
rect 675407 241203 675887 241259
rect 675407 240007 675887 240063
rect 675407 238167 675887 238223
rect 675407 236327 675887 236383
rect 675407 205295 675887 205351
rect 675407 204651 675887 204707
rect 675407 204007 675887 204063
rect 675312 203522 675340 203580
rect 675300 203516 675352 203522
rect 675407 203497 675887 203511
rect 675352 203469 675887 203497
rect 675300 203458 675352 203464
rect 675312 199186 675340 203458
rect 675407 203455 675887 203469
rect 675407 202167 675887 202223
rect 675407 201615 675887 201671
rect 675407 200971 675887 201027
rect 675407 200327 675887 200383
rect 675407 199186 675887 199187
rect 675312 199158 675887 199186
rect 675404 199131 675887 199158
rect 675404 199102 675432 199131
rect 675392 199096 675444 199102
rect 675392 199038 675444 199044
rect 673736 158636 673788 158642
rect 673736 158578 673788 158584
rect 673736 154148 673788 154154
rect 673736 154090 673788 154096
rect 42340 45620 42392 45626
rect 42340 45562 42392 45568
rect 143632 45620 143684 45626
rect 143632 45562 143684 45568
rect 143644 44198 143672 45562
rect 143632 44192 143684 44198
rect 143632 44134 143684 44140
rect 145104 44192 145156 44198
rect 145104 44134 145156 44140
rect 145116 40202 145144 44134
rect 145103 40174 145144 40202
rect 145103 40000 145131 40174
rect 199660 44464 199712 44470
rect 199660 44406 199712 44412
rect 195336 44192 195388 44198
rect 195336 44134 195388 44140
rect 195348 42193 195376 44134
rect 199672 44198 199700 44406
rect 199660 44192 199712 44198
rect 199660 44134 199712 44140
rect 199672 42193 199700 44134
rect 187327 41713 187383 42193
rect 194043 41713 194099 42193
rect 195331 41713 195387 42193
rect 199655 41713 199711 42193
rect 145091 39706 145143 40000
rect 527456 46912 527508 46918
rect 527456 46854 527508 46860
rect 303896 44260 303948 44266
rect 303896 44202 303948 44208
rect 303908 42193 303936 44202
rect 308220 44260 308272 44266
rect 308220 44202 308272 44208
rect 308232 42193 308260 44202
rect 358728 44260 358780 44266
rect 358728 44202 358780 44208
rect 358740 42193 358768 44202
rect 302643 41713 302699 42193
rect 303908 41806 303987 42193
rect 303931 41713 303987 41806
rect 306967 41713 307023 42193
rect 308232 41806 308311 42193
rect 308255 41713 308311 41806
rect 310095 41713 310151 42193
rect 357443 41713 357499 42193
rect 358731 41713 358787 42193
rect 363052 44328 363104 44334
rect 363052 44270 363104 44276
rect 363064 42193 363092 44270
rect 411074 44432 411130 44441
rect 411074 44367 411130 44376
rect 411088 42193 411116 44367
rect 413560 44328 413612 44334
rect 413560 44270 413612 44276
rect 413572 42193 413600 44270
rect 417884 44328 417936 44334
rect 417884 44270 417936 44276
rect 417896 42193 417924 44270
rect 419722 44296 419778 44305
rect 419722 44231 419778 44240
rect 419736 42193 419764 44231
rect 465814 44432 465870 44441
rect 465814 44367 465870 44376
rect 465828 42193 465856 44367
rect 468300 44328 468352 44334
rect 468300 44270 468352 44276
rect 468312 42193 468340 44270
rect 472624 44328 472676 44334
rect 472624 44270 472676 44276
rect 472636 42193 472664 44270
rect 474462 44432 474518 44441
rect 474462 44367 474518 44376
rect 474476 42193 474504 44367
rect 518806 44296 518862 44305
rect 518806 44231 518862 44240
rect 518820 42193 518848 44231
rect 523132 44192 523184 44198
rect 523132 44134 523184 44140
rect 523144 42193 523172 44134
rect 524970 44296 525026 44305
rect 524970 44231 525026 44240
rect 524984 42193 525012 44231
rect 527468 44198 527496 46854
rect 527456 44192 527508 44198
rect 527456 44134 527508 44140
rect 527468 42193 527496 44134
rect 673748 139346 673776 154090
rect 675407 197843 675887 197899
rect 675407 197291 675887 197347
rect 675407 196647 675887 196703
rect 675407 196003 675887 196059
rect 675407 194807 675887 194863
rect 675407 192967 675887 193023
rect 675407 191127 675887 191183
rect 675407 160295 675887 160351
rect 675407 159651 675887 159707
rect 675407 159007 675887 159063
rect 675392 158636 675444 158642
rect 675392 158578 675444 158584
rect 675404 158522 675432 158578
rect 675312 158511 675432 158522
rect 675312 158494 675887 158511
rect 675312 154170 675340 158494
rect 675407 158455 675887 158494
rect 675407 157167 675887 157223
rect 675407 156615 675887 156671
rect 675407 155971 675887 156027
rect 675407 155327 675887 155383
rect 675407 154170 675887 154187
rect 675312 154154 675887 154170
rect 675300 154148 675887 154154
rect 675352 154142 675887 154148
rect 675407 154131 675887 154142
rect 675300 154090 675352 154096
rect 675312 154059 675340 154090
rect 673656 139318 673776 139346
rect 673656 113762 673684 139318
rect 675407 152843 675887 152899
rect 675407 152291 675887 152347
rect 675407 151647 675887 151703
rect 675407 151003 675887 151059
rect 675407 149807 675887 149863
rect 675407 147967 675887 148023
rect 675407 146127 675887 146183
rect 673644 113756 673696 113762
rect 673644 113698 673696 113704
rect 673644 108452 673696 108458
rect 673644 108394 673696 108400
rect 673656 46986 673684 108394
rect 675407 115095 675887 115151
rect 675407 114451 675887 114507
rect 675407 113807 675887 113863
rect 675392 113756 675444 113762
rect 675392 113698 675444 113704
rect 675404 113311 675432 113698
rect 675404 113297 675887 113311
rect 675312 113269 675887 113297
rect 675312 108973 675340 113269
rect 675407 113255 675887 113269
rect 675407 111967 675887 112023
rect 675407 111415 675887 111471
rect 675407 110771 675887 110827
rect 675407 110127 675887 110183
rect 675407 108973 675887 108987
rect 675312 108945 675887 108973
rect 675404 108931 675887 108945
rect 675404 108458 675432 108931
rect 675392 108452 675444 108458
rect 675392 108394 675444 108400
rect 673644 46980 673696 46986
rect 673644 46922 673696 46928
rect 675407 107643 675887 107699
rect 675407 107091 675887 107147
rect 675407 106447 675887 106503
rect 675407 105803 675887 105859
rect 675407 104607 675887 104663
rect 675407 102767 675887 102823
rect 675407 100927 675887 100983
rect 361767 41713 361823 42193
rect 363055 41713 363111 42193
rect 364895 41713 364951 42193
rect 405527 41713 405583 42193
rect 409207 41834 409263 42193
rect 409207 41818 409368 41834
rect 409207 41812 409380 41818
rect 409207 41806 409328 41812
rect 409207 41713 409263 41806
rect 409328 41754 409380 41760
rect 411047 41820 411116 42193
rect 411047 41713 411103 41820
rect 412243 41834 412299 42193
rect 412243 41818 412404 41834
rect 413531 41820 413600 42193
rect 415371 41834 415427 42193
rect 412243 41812 412416 41818
rect 412243 41806 412364 41812
rect 412243 41713 412299 41806
rect 412364 41754 412416 41760
rect 413531 41713 413587 41820
rect 415228 41818 415427 41834
rect 415216 41812 415427 41818
rect 415268 41806 415427 41812
rect 415216 41754 415268 41760
rect 415371 41713 415427 41806
rect 416567 41713 416623 42193
rect 417855 41820 417924 42193
rect 419695 41820 419764 42193
rect 417855 41713 417911 41820
rect 419695 41713 419751 41820
rect 460327 41713 460383 42193
rect 464007 41834 464063 42193
rect 464007 41818 464200 41834
rect 464007 41812 464212 41818
rect 464007 41806 464160 41812
rect 464007 41713 464063 41806
rect 464160 41754 464212 41760
rect 465828 41806 465903 42193
rect 465847 41713 465903 41806
rect 467043 41834 467099 42193
rect 467043 41818 467236 41834
rect 467043 41812 467248 41818
rect 467043 41806 467196 41812
rect 467043 41713 467099 41806
rect 468312 41806 468387 42193
rect 470171 41834 470227 42193
rect 470060 41818 470227 41834
rect 467196 41754 467248 41760
rect 468331 41713 468387 41806
rect 470048 41812 470227 41818
rect 470100 41806 470227 41812
rect 470048 41754 470100 41760
rect 470171 41713 470227 41806
rect 471367 41713 471423 42193
rect 472636 41806 472711 42193
rect 474476 41806 474551 42193
rect 472655 41713 472711 41806
rect 474495 41713 474551 41806
rect 515127 41713 515183 42193
rect 518807 41713 518863 42193
rect 520647 41713 520703 42193
rect 521843 41713 521899 42193
rect 523131 41713 523187 42193
rect 524971 41713 525027 42193
rect 526167 41713 526223 42193
rect 527455 41713 527511 42193
rect 529295 41713 529351 42193
<< via2 >>
rect 411074 44376 411130 44432
rect 419722 44240 419778 44296
rect 465814 44376 465870 44432
rect 474462 44376 474518 44432
rect 518806 44240 518862 44296
rect 524970 44240 525026 44296
<< obsm2 >>
rect 76242 995943 92183 1037600
rect 76242 995887 76441 995943
rect 76609 995887 76993 995943
rect 77161 995887 77637 995943
rect 77805 995887 78281 995943
rect 78449 995887 78833 995943
rect 79001 995887 79477 995943
rect 79645 995887 80121 995943
rect 80289 995887 80673 995943
rect 80841 995887 81317 995943
rect 81485 995887 81961 995943
rect 82129 995887 82513 995943
rect 82681 995887 83157 995943
rect 83325 995887 83801 995943
rect 83969 995887 84445 995943
rect 84613 995887 84997 995943
rect 85165 995887 85641 995943
rect 85809 995887 86285 995943
rect 86453 995887 86837 995943
rect 87005 995887 87481 995943
rect 87649 995887 88125 995943
rect 88293 995887 88677 995943
rect 88845 995887 89321 995943
rect 89489 995887 89965 995943
rect 90133 995887 90517 995943
rect 90685 995887 91161 995943
rect 91329 995887 91805 995943
rect 91973 995887 92183 995943
rect 127642 995943 143583 1037600
rect 127642 995887 127841 995943
rect 128009 995887 128393 995943
rect 128561 995887 129037 995943
rect 129205 995887 129681 995943
rect 129849 995887 130233 995943
rect 130401 995887 130877 995943
rect 131045 995887 131521 995943
rect 131689 995887 132073 995943
rect 132241 995887 132717 995943
rect 132885 995887 133361 995943
rect 133529 995887 133913 995943
rect 134081 995887 134557 995943
rect 134725 995887 135201 995943
rect 135369 995887 135845 995943
rect 136013 995887 136397 995943
rect 136565 995887 137041 995943
rect 137209 995887 137685 995943
rect 137853 995887 138237 995943
rect 138405 995887 138881 995943
rect 139049 995887 139525 995943
rect 139693 995887 140077 995943
rect 140245 995887 140721 995943
rect 140889 995887 141365 995943
rect 141533 995887 141917 995943
rect 142085 995887 142561 995943
rect 142729 995887 143205 995943
rect 143373 995887 143583 995943
rect 179042 995943 194983 1037600
rect 179042 995887 179241 995943
rect 179409 995887 179793 995943
rect 179961 995887 180437 995943
rect 180605 995887 181081 995943
rect 181249 995887 181633 995943
rect 181801 995887 182277 995943
rect 182445 995887 182921 995943
rect 183089 995887 183473 995943
rect 183641 995887 184117 995943
rect 184285 995887 184761 995943
rect 184929 995887 185313 995943
rect 185481 995887 185957 995943
rect 186125 995887 186601 995943
rect 186769 995887 187245 995943
rect 187413 995887 187797 995943
rect 187965 995887 188441 995943
rect 188609 995887 189085 995943
rect 189253 995887 189637 995943
rect 189805 995887 190281 995943
rect 190449 995887 190925 995943
rect 191093 995887 191477 995943
rect 191645 995887 192121 995943
rect 192289 995887 192765 995943
rect 192933 995887 193317 995943
rect 193485 995887 193961 995943
rect 194129 995887 194605 995943
rect 194773 995887 194983 995943
rect 230442 995943 246383 1037600
rect 230442 995887 230641 995943
rect 230809 995887 231193 995943
rect 231361 995887 231837 995943
rect 232005 995887 232481 995943
rect 232649 995887 233033 995943
rect 233201 995887 233677 995943
rect 233845 995887 234321 995943
rect 234489 995887 234873 995943
rect 235041 995887 235517 995943
rect 235685 995887 236161 995943
rect 236329 995887 236713 995943
rect 236881 995887 237357 995943
rect 237525 995887 238001 995943
rect 238169 995887 238645 995943
rect 238813 995887 239197 995943
rect 239365 995887 239841 995943
rect 240009 995887 240485 995943
rect 240653 995887 241037 995943
rect 241205 995887 241681 995943
rect 241849 995887 242325 995943
rect 242493 995887 242877 995943
rect 243045 995887 243521 995943
rect 243689 995887 244165 995943
rect 244333 995887 244717 995943
rect 244885 995887 245361 995943
rect 245529 995887 246005 995943
rect 246173 995887 246383 995943
rect 282042 995943 297983 1037600
rect 333453 998007 348258 1036615
rect 333499 997600 338279 998007
rect 338579 997600 338979 997984
rect 343478 997600 348258 998007
rect 342166 997455 342222 997529
rect 282042 995887 282241 995943
rect 282409 995887 282793 995943
rect 282961 995887 283437 995943
rect 283605 995887 284081 995943
rect 284249 995887 284633 995943
rect 284801 995887 285277 995943
rect 285445 995887 285921 995943
rect 286089 995887 286473 995943
rect 286641 995887 287117 995943
rect 287285 995887 287761 995943
rect 287929 995887 288313 995943
rect 288481 995887 288957 995943
rect 289125 995887 289601 995943
rect 289769 995887 290245 995943
rect 290413 995887 290797 995943
rect 290965 995887 291441 995943
rect 291609 995887 292085 995943
rect 292253 995887 292637 995943
rect 292805 995887 293281 995943
rect 293449 995887 293925 995943
rect 294093 995887 294477 995943
rect 294645 995887 295121 995943
rect 295289 995887 295765 995943
rect 295933 995887 296317 995943
rect 296485 995887 296961 995943
rect 297129 995887 297605 995943
rect 297773 995887 297983 995943
rect 76497 995407 76553 995887
rect 79533 995452 79589 995887
rect 79520 995407 79589 995452
rect 82569 995452 82625 995887
rect 82556 995407 82625 995452
rect 83857 995466 83913 995887
rect 84016 995590 84068 995654
rect 84028 995466 84056 995590
rect 83857 995438 84056 995466
rect 83857 995407 83913 995438
rect 86893 995407 86949 995887
rect 88181 995407 88237 995887
rect 90021 995452 90077 995887
rect 90008 995407 90077 995452
rect 90573 995407 90629 995887
rect 91744 995590 91796 995654
rect 91756 995466 91784 995590
rect 91861 995466 91917 995887
rect 91756 995438 91917 995466
rect 91861 995407 91917 995438
rect 127897 995407 127953 995887
rect 130933 995407 130989 995887
rect 133969 995407 134025 995887
rect 135257 995466 135313 995887
rect 135352 995466 135404 995518
rect 135257 995454 135404 995466
rect 135257 995438 135392 995454
rect 135257 995407 135313 995438
rect 138293 995407 138349 995887
rect 139581 995407 139637 995887
rect 141421 995407 141477 995887
rect 141973 995407 142029 995887
rect 143172 995466 143224 995518
rect 143261 995466 143317 995887
rect 143172 995454 143317 995466
rect 143184 995438 143317 995454
rect 143261 995407 143317 995438
rect 179297 995407 179353 995887
rect 182333 995466 182389 995887
rect 182333 995407 182404 995466
rect 185369 995466 185425 995887
rect 186657 995466 186713 995887
rect 185369 995407 185440 995466
rect 186657 995407 186728 995466
rect 189693 995407 189749 995887
rect 190981 995407 191037 995887
rect 192821 995466 192877 995887
rect 192821 995407 192892 995466
rect 193373 995407 193429 995887
rect 194661 995466 194717 995887
rect 194661 995407 194732 995466
rect 230697 995407 230753 995887
rect 233733 995466 233789 995887
rect 233712 995407 233789 995466
rect 236769 995466 236825 995887
rect 236748 995407 236825 995466
rect 238057 995466 238113 995887
rect 238208 995590 238260 995654
rect 238220 995466 238248 995590
rect 238057 995438 238248 995466
rect 238057 995407 238113 995438
rect 241093 995407 241149 995887
rect 242381 995407 242437 995887
rect 244221 995466 244277 995887
rect 244200 995407 244277 995466
rect 244773 995407 244829 995887
rect 245936 995590 245988 995654
rect 245948 995466 245976 995590
rect 246061 995466 246117 995887
rect 245948 995438 246117 995466
rect 246061 995407 246117 995438
rect 282297 995407 282353 995887
rect 285333 995452 285389 995887
rect 285324 995407 285389 995452
rect 288369 995452 288425 995887
rect 289657 995452 289713 995887
rect 288360 995407 288425 995452
rect 289648 995407 289713 995452
rect 292693 995407 292749 995887
rect 293981 995407 294037 995887
rect 295821 995452 295877 995887
rect 295812 995407 295877 995452
rect 296373 995407 296429 995887
rect 297661 995452 297717 995887
rect 297652 995407 297717 995452
rect 79520 990690 79548 995407
rect 82556 990826 82584 995407
rect 82544 990762 82596 990826
rect 79508 990626 79560 990690
rect 42248 990150 42300 990214
rect 0 969973 41713 970183
rect 0 969805 41657 969973
rect 41713 969861 42193 969917
rect 0 969329 41713 969805
rect 41800 969406 41828 969861
rect 41788 969342 41840 969406
rect 0 969161 41657 969329
rect 0 968685 41713 969161
rect 0 968517 41657 968685
rect 41713 968573 42193 968629
rect 0 968133 41713 968517
rect 41788 968458 41840 968522
rect 0 967965 41657 968133
rect 41800 968077 41828 968458
rect 41713 968021 42193 968077
rect 0 967489 41713 967965
rect 0 967321 41657 967489
rect 0 966845 41713 967321
rect 0 966677 41657 966845
rect 0 966293 41713 966677
rect 0 966125 41657 966293
rect 41713 966181 42193 966237
rect 0 965649 41713 966125
rect 0 965481 41657 965649
rect 0 965005 41713 965481
rect 0 964837 41657 965005
rect 41713 964893 42193 964949
rect 0 964453 41713 964837
rect 0 964285 41657 964453
rect 0 963809 41713 964285
rect 0 963641 41657 963809
rect 0 963165 41713 963641
rect 0 962997 41657 963165
rect 0 962613 41713 962997
rect 0 962445 41657 962613
rect 0 961969 41713 962445
rect 41788 962406 41840 962470
rect 0 961801 41657 961969
rect 41800 961913 41828 962406
rect 41713 961857 42193 961913
rect 41722 961846 41828 961857
rect 0 961325 41713 961801
rect 0 961157 41657 961325
rect 0 960681 41713 961157
rect 0 960513 41657 960681
rect 41713 960569 42193 960625
rect 0 960129 41713 960513
rect 41984 960498 42012 960569
rect 41972 960434 42024 960498
rect 0 959961 41657 960129
rect 0 959485 41713 959961
rect 0 959317 41657 959485
rect 0 958841 41713 959317
rect 0 958673 41657 958841
rect 0 958289 41713 958673
rect 0 958121 41657 958289
rect 0 957645 41713 958121
rect 42260 957658 42288 990150
rect 79520 990214 79548 990626
rect 79508 990150 79560 990214
rect 82556 990146 82584 990762
rect 90008 990758 90036 995407
rect 88340 990694 88392 990758
rect 89996 990694 90048 990758
rect 88352 990146 88380 990694
rect 130948 990690 130976 995407
rect 133984 990826 134012 995407
rect 133972 990762 134024 990826
rect 130936 990626 130988 990690
rect 135168 990762 135220 990826
rect 135180 990486 135208 990762
rect 141436 990758 141464 995407
rect 141424 990694 141476 990758
rect 182376 990690 182404 995407
rect 185412 990826 185440 995407
rect 184940 990762 184992 990826
rect 185400 990762 185452 990826
rect 182364 990626 182416 990690
rect 184952 990486 184980 990762
rect 186700 990554 186728 995407
rect 192864 990758 192892 995407
rect 192852 990694 192904 990758
rect 194704 990554 194732 995407
rect 233712 990690 233740 995407
rect 236748 990826 236776 995407
rect 236736 990762 236788 990826
rect 233700 990626 233752 990690
rect 236748 990554 236776 990762
rect 244200 990758 244228 995407
rect 244188 990694 244240 990758
rect 285324 990622 285352 995407
rect 285312 990558 285364 990622
rect 186688 990490 186740 990554
rect 194692 990490 194744 990554
rect 236736 990490 236788 990554
rect 288360 990554 288388 995407
rect 289648 995314 289676 995407
rect 289636 995250 289688 995314
rect 295812 990758 295840 995407
rect 297652 995314 297680 995407
rect 297640 995250 297692 995314
rect 295800 990694 295852 990758
rect 342180 990622 342208 997455
rect 383842 995943 399783 1037600
rect 383842 995887 384041 995943
rect 384209 995887 384593 995943
rect 384761 995887 385237 995943
rect 385405 995887 385881 995943
rect 386049 995887 386433 995943
rect 386601 995887 387077 995943
rect 387245 995887 387721 995943
rect 387889 995887 388273 995943
rect 388441 995887 388917 995943
rect 389085 995887 389561 995943
rect 389729 995887 390113 995943
rect 390281 995887 390757 995943
rect 390925 995887 391401 995943
rect 391569 995887 392045 995943
rect 392213 995887 392597 995943
rect 392765 995887 393241 995943
rect 393409 995887 393885 995943
rect 394053 995887 394437 995943
rect 394605 995887 395081 995943
rect 395249 995887 395725 995943
rect 395893 995887 396277 995943
rect 396445 995887 396921 995943
rect 397089 995887 397565 995943
rect 397733 995887 398117 995943
rect 398285 995887 398761 995943
rect 398929 995887 399405 995943
rect 399573 995887 399783 995943
rect 472842 995943 488783 1037600
rect 472842 995887 473041 995943
rect 473209 995887 473593 995943
rect 473761 995887 474237 995943
rect 474405 995887 474881 995943
rect 475049 995887 475433 995943
rect 475601 995887 476077 995943
rect 476245 995887 476721 995943
rect 476889 995887 477273 995943
rect 477441 995887 477917 995943
rect 478085 995887 478561 995943
rect 478729 995887 479113 995943
rect 479281 995887 479757 995943
rect 479925 995887 480401 995943
rect 480569 995887 481045 995943
rect 481213 995887 481597 995943
rect 481765 995887 482241 995943
rect 482409 995887 482885 995943
rect 483053 995887 483437 995943
rect 483605 995887 484081 995943
rect 484249 995887 484725 995943
rect 484893 995887 485277 995943
rect 485445 995887 485921 995943
rect 486089 995887 486565 995943
rect 486733 995887 487117 995943
rect 487285 995887 487761 995943
rect 487929 995887 488405 995943
rect 488573 995887 488783 995943
rect 524242 995943 540183 1037600
rect 575653 998007 590458 1036615
rect 575699 997600 580479 998007
rect 580779 997600 581179 997984
rect 585678 997600 590458 998007
rect 585046 997455 585102 997529
rect 524242 995887 524441 995943
rect 524609 995887 524993 995943
rect 525161 995887 525637 995943
rect 525805 995887 526281 995943
rect 526449 995887 526833 995943
rect 527001 995887 527477 995943
rect 527645 995887 528121 995943
rect 528289 995887 528673 995943
rect 528841 995887 529317 995943
rect 529485 995887 529961 995943
rect 530129 995887 530513 995943
rect 530681 995887 531157 995943
rect 531325 995887 531801 995943
rect 531969 995887 532445 995943
rect 532613 995887 532997 995943
rect 533165 995887 533641 995943
rect 533809 995887 534285 995943
rect 534453 995887 534837 995943
rect 535005 995887 535481 995943
rect 535649 995887 536125 995943
rect 536293 995887 536677 995943
rect 536845 995887 537321 995943
rect 537489 995887 537965 995943
rect 538133 995887 538517 995943
rect 538685 995887 539161 995943
rect 539329 995887 539805 995943
rect 539973 995887 540183 995943
rect 384097 995407 384153 995887
rect 387133 995452 387189 995887
rect 387133 995407 387196 995452
rect 390169 995452 390225 995887
rect 391457 995452 391513 995887
rect 390169 995407 390232 995452
rect 391457 995407 391520 995452
rect 394493 995407 394549 995887
rect 395781 995407 395837 995887
rect 397621 995452 397677 995887
rect 397621 995407 397684 995452
rect 398173 995407 398229 995887
rect 399461 995452 399517 995887
rect 399461 995407 399524 995452
rect 473097 995407 473153 995887
rect 476133 995452 476189 995887
rect 476132 995407 476189 995452
rect 479169 995452 479225 995887
rect 480457 995452 480513 995887
rect 479168 995407 479225 995452
rect 480456 995407 480513 995452
rect 483493 995407 483549 995887
rect 484781 995407 484837 995887
rect 486621 995452 486677 995887
rect 486620 995407 486677 995452
rect 487173 995407 487229 995887
rect 488461 995452 488517 995887
rect 488460 995407 488517 995452
rect 524497 995407 524553 995887
rect 527533 995407 527589 995887
rect 530569 995407 530625 995887
rect 531857 995466 531913 995887
rect 531964 995590 532016 995654
rect 531976 995466 532004 995590
rect 531857 995438 532004 995466
rect 531857 995407 531913 995438
rect 534893 995407 534949 995887
rect 536181 995407 536237 995887
rect 538021 995407 538077 995887
rect 538573 995407 538629 995887
rect 539692 995590 539744 995654
rect 539704 995466 539732 995590
rect 539861 995466 539917 995887
rect 539704 995438 539917 995466
rect 539861 995407 539917 995438
rect 342168 990558 342220 990622
rect 386420 990558 386472 990622
rect 288348 990490 288400 990554
rect 386432 990486 386460 990558
rect 387168 990486 387196 995407
rect 390204 990690 390232 995407
rect 390192 990626 390244 990690
rect 390204 990554 390232 990626
rect 391492 995314 391520 995407
rect 391480 995250 391532 995314
rect 397656 990758 397684 995407
rect 399496 995314 399524 995407
rect 399484 995250 399536 995314
rect 397644 990694 397696 990758
rect 476132 990554 476160 995407
rect 479168 990690 479196 995407
rect 479156 990626 479208 990690
rect 480456 995314 480484 995407
rect 480444 995250 480496 995314
rect 486620 990758 486648 995407
rect 488460 995314 488488 995407
rect 488448 995250 488500 995314
rect 486608 990694 486660 990758
rect 480168 990626 480220 990690
rect 390192 990490 390244 990554
rect 476120 990490 476172 990554
rect 480180 990486 480208 990626
rect 527560 990690 527588 995407
rect 527548 990626 527600 990690
rect 527560 990554 527588 990626
rect 527548 990490 527600 990554
rect 530596 990486 530624 995407
rect 538048 990758 538076 995407
rect 585060 992254 585088 997455
rect 626042 995943 641983 1037600
rect 626042 995887 626241 995943
rect 626409 995887 626793 995943
rect 626961 995887 627437 995943
rect 627605 995887 628081 995943
rect 628249 995887 628633 995943
rect 628801 995887 629277 995943
rect 629445 995887 629921 995943
rect 630089 995887 630473 995943
rect 630641 995887 631117 995943
rect 631285 995887 631761 995943
rect 631929 995887 632313 995943
rect 632481 995887 632957 995943
rect 633125 995887 633601 995943
rect 633769 995887 634245 995943
rect 634413 995887 634797 995943
rect 634965 995887 635441 995943
rect 635609 995887 636085 995943
rect 636253 995887 636637 995943
rect 636805 995887 637281 995943
rect 637449 995887 637925 995943
rect 638093 995887 638477 995943
rect 638645 995887 639121 995943
rect 639289 995887 639765 995943
rect 639933 995887 640317 995943
rect 640485 995887 640961 995943
rect 641129 995887 641605 995943
rect 641773 995887 641983 995943
rect 626297 995407 626353 995887
rect 629333 995466 629389 995887
rect 629312 995407 629389 995466
rect 632369 995466 632425 995887
rect 632348 995407 632425 995466
rect 633657 995466 633713 995887
rect 633808 995466 633860 995518
rect 633657 995454 633860 995466
rect 633657 995438 633848 995454
rect 633657 995407 633713 995438
rect 636693 995407 636749 995887
rect 637981 995407 638037 995887
rect 639821 995466 639877 995887
rect 639800 995407 639877 995466
rect 640373 995407 640429 995887
rect 641536 995466 641588 995518
rect 641661 995466 641717 995887
rect 641536 995454 641717 995466
rect 641548 995438 641717 995454
rect 641661 995407 641717 995438
rect 585048 992190 585100 992254
rect 538036 990694 538088 990758
rect 629312 990690 629340 995407
rect 629300 990626 629352 990690
rect 631784 990626 631836 990690
rect 135168 990422 135220 990486
rect 184940 990422 184992 990486
rect 386420 990422 386472 990486
rect 387156 990422 387208 990486
rect 480168 990422 480220 990486
rect 530584 990422 530636 990486
rect 631796 990146 631824 990626
rect 632348 990554 632376 995407
rect 639800 990758 639828 995407
rect 674748 992190 674800 992254
rect 639788 990694 639840 990758
rect 632336 990490 632388 990554
rect 639800 990282 639828 990694
rect 639788 990218 639840 990282
rect 673736 990218 673788 990282
rect 673460 990150 673512 990214
rect 44916 990082 44968 990146
rect 82544 990082 82596 990146
rect 88340 990082 88392 990146
rect 631784 990082 631836 990146
rect 42616 990014 42668 990078
rect 42340 969342 42392 969406
rect 42352 962470 42380 969342
rect 42340 962406 42392 962470
rect 42628 968522 42656 990014
rect 42616 968458 42668 968522
rect 0 957477 41657 957645
rect 41800 957630 42288 957658
rect 41800 957589 41828 957630
rect 41713 957533 42193 957589
rect 0 957001 41713 957477
rect 0 956833 41657 957001
rect 44824 960494 44876 960498
rect 44928 960494 44956 990082
rect 673472 961382 673500 990150
rect 673644 990014 673696 990078
rect 673656 964782 673684 990014
rect 673644 964718 673696 964782
rect 673460 961318 673512 961382
rect 44824 960466 44956 960494
rect 44824 960434 44876 960466
rect 0 956449 41713 956833
rect 0 956281 41657 956449
rect 0 955805 41713 956281
rect 0 955637 41657 955805
rect 0 955161 41713 955637
rect 0 954993 41657 955161
rect 0 954609 41713 954993
rect 0 954441 41657 954609
rect 41713 954497 42193 954553
rect 0 954242 41713 954441
rect 44836 955058 44864 960434
rect 44180 954994 44232 955058
rect 44824 954994 44876 955058
rect 7 927240 30281 929187
rect 30753 927000 31683 929228
rect 32033 927240 34915 929187
rect 7 926940 39593 927000
rect 7 922819 39600 926940
rect 7 922707 39593 922819
rect 7 916185 39600 922707
rect 7 916099 39593 916185
rect 7 912100 39600 916099
rect 7 912000 39593 912100
rect 30760 909805 31690 912000
rect 985 879878 40000 884658
rect 985 874679 39593 879878
rect 39616 874979 40000 875379
rect 985 869899 40000 874679
rect 42246 870023 42302 870097
rect 985 869853 39593 869899
rect 985 837678 40000 842458
rect 985 832479 39593 837678
rect 39616 832779 40000 833179
rect 985 827699 40000 832479
rect 985 827653 39593 827699
rect 42260 805934 42288 870023
rect 42260 805906 42472 805934
rect 0 800173 41713 800383
rect 0 800005 41657 800173
rect 41713 800103 42193 800117
rect 41713 800075 42288 800103
rect 41713 800061 42193 800075
rect 0 799529 41713 800005
rect 0 799361 41657 799529
rect 0 798885 41713 799361
rect 0 798717 41657 798885
rect 41713 798773 42193 798829
rect 0 798333 41713 798717
rect 0 798165 41657 798333
rect 41713 798221 42193 798277
rect 0 797689 41713 798165
rect 41800 797774 41828 798221
rect 41788 797710 41840 797774
rect 0 797521 41657 797689
rect 0 797045 41713 797521
rect 0 796877 41657 797045
rect 0 796493 41713 796877
rect 0 796325 41657 796493
rect 41713 796381 42193 796437
rect 0 795849 41713 796325
rect 0 795681 41657 795849
rect 0 795205 41713 795681
rect 0 795037 41657 795205
rect 41713 795093 42193 795149
rect 0 794653 41713 795037
rect 0 794485 41657 794653
rect 0 794009 41713 794485
rect 0 793841 41657 794009
rect 0 793365 41713 793841
rect 0 793197 41657 793365
rect 0 792813 41713 793197
rect 0 792645 41657 792813
rect 0 792169 41713 792645
rect 42260 792282 42288 800075
rect 42340 797710 42392 797774
rect 41800 792254 42288 792282
rect 0 792001 41657 792169
rect 41800 792113 41828 792254
rect 41713 792057 42193 792113
rect 0 791525 41713 792001
rect 0 791357 41657 791525
rect 0 790881 41713 791357
rect 41788 791318 41840 791382
rect 42248 791318 42300 791382
rect 0 790713 41657 790881
rect 41800 790825 41828 791318
rect 41713 790769 42193 790825
rect 41722 790758 41828 790769
rect 0 790329 41713 790713
rect 0 790161 41657 790329
rect 0 789685 41713 790161
rect 0 789517 41657 789685
rect 0 789041 41713 789517
rect 0 788873 41657 789041
rect 0 788489 41713 788873
rect 0 788321 41657 788489
rect 0 787845 41713 788321
rect 0 787677 41657 787845
rect 41722 787789 41828 787794
rect 41713 787733 42193 787789
rect 0 787201 41713 787677
rect 41800 787302 41828 787733
rect 41788 787238 41840 787302
rect 0 787033 41657 787201
rect 0 786649 41713 787033
rect 0 786481 41657 786649
rect 0 786005 41713 786481
rect 0 785837 41657 786005
rect 0 785361 41713 785837
rect 0 785193 41657 785361
rect 0 784809 41713 785193
rect 0 784641 41657 784809
rect 41713 784697 42193 784753
rect 0 784442 41713 784641
rect 0 756973 41713 757183
rect 0 756805 41657 756973
rect 41722 756917 41828 756922
rect 41713 756861 42193 756917
rect 0 756329 41713 756805
rect 41800 756430 41828 756861
rect 41788 756366 41840 756430
rect 0 756161 41657 756329
rect 0 755685 41713 756161
rect 0 755517 41657 755685
rect 41713 755573 42193 755629
rect 0 755133 41713 755517
rect 41788 755414 41840 755478
rect 0 754965 41657 755133
rect 41800 755077 41828 755414
rect 41713 755021 42193 755077
rect 0 754489 41713 754965
rect 0 754321 41657 754489
rect 0 753845 41713 754321
rect 0 753677 41657 753845
rect 0 753293 41713 753677
rect 0 753125 41657 753293
rect 41713 753181 42193 753237
rect 0 752649 41713 753125
rect 0 752481 41657 752649
rect 0 752005 41713 752481
rect 0 751837 41657 752005
rect 41713 751893 42193 751949
rect 0 751453 41713 751837
rect 0 751285 41657 751453
rect 0 750809 41713 751285
rect 0 750641 41657 750809
rect 0 750165 41713 750641
rect 0 749997 41657 750165
rect 0 749613 41713 749997
rect 0 749445 41657 749613
rect 0 748969 41713 749445
rect 41788 749362 41840 749426
rect 0 748801 41657 748969
rect 41800 748913 41828 749362
rect 41713 748857 42193 748913
rect 0 748325 41713 748801
rect 0 748157 41657 748325
rect 0 747681 41713 748157
rect 0 747513 41657 747681
rect 41713 747611 42193 747625
rect 42260 747611 42288 791318
rect 42352 756514 42380 797710
rect 42444 791382 42472 805906
rect 44192 870097 44220 954994
rect 673472 872438 673500 961318
rect 673656 960494 673684 964718
rect 673564 960466 673684 960494
rect 673564 874546 673592 960466
rect 673748 953358 673776 990218
rect 673736 953294 673788 953358
rect 673552 874482 673604 874546
rect 673460 872374 673512 872438
rect 673460 870538 673512 870602
rect 44178 870023 44234 870097
rect 673472 864482 673500 870538
rect 673460 864418 673512 864482
rect 42432 791318 42484 791382
rect 42616 787238 42668 787302
rect 42352 756486 42564 756514
rect 42340 756366 42392 756430
rect 42352 749426 42380 756366
rect 42340 749362 42392 749426
rect 42536 755478 42564 756486
rect 42524 755414 42576 755478
rect 41713 747583 42288 747611
rect 41713 747569 42193 747583
rect 0 747129 41713 747513
rect 0 746961 41657 747129
rect 0 746485 41713 746961
rect 0 746317 41657 746485
rect 0 745841 41713 746317
rect 0 745673 41657 745841
rect 0 745289 41713 745673
rect 0 745121 41657 745289
rect 0 744645 41713 745121
rect 0 744477 41657 744645
rect 41713 744533 42193 744589
rect 0 744001 41713 744477
rect 41800 744054 41828 744533
rect 0 743833 41657 744001
rect 41788 743990 41840 744054
rect 0 743449 41713 743833
rect 0 743281 41657 743449
rect 0 742805 41713 743281
rect 0 742637 41657 742805
rect 0 742161 41713 742637
rect 0 741993 41657 742161
rect 0 741609 41713 741993
rect 0 741441 41657 741609
rect 41713 741497 42193 741553
rect 0 741242 41713 741441
rect 42260 718978 42288 747583
rect 42260 718950 42472 718978
rect 0 713773 41713 713983
rect 0 713605 41657 713773
rect 41713 713703 42193 713717
rect 41713 713675 42288 713703
rect 41713 713661 42193 713675
rect 0 713129 41713 713605
rect 0 712961 41657 713129
rect 0 712485 41713 712961
rect 0 712317 41657 712485
rect 41713 712373 42193 712429
rect 0 711933 41713 712317
rect 41788 712234 41840 712298
rect 0 711765 41657 711933
rect 41800 711877 41828 712234
rect 41713 711821 42193 711877
rect 0 711289 41713 711765
rect 0 711121 41657 711289
rect 0 710645 41713 711121
rect 0 710477 41657 710645
rect 0 710093 41713 710477
rect 0 709925 41657 710093
rect 41713 709981 42193 710037
rect 0 709449 41713 709925
rect 0 709281 41657 709449
rect 0 708805 41713 709281
rect 0 708637 41657 708805
rect 41713 708693 42193 708749
rect 0 708253 41713 708637
rect 0 708085 41657 708253
rect 0 707609 41713 708085
rect 0 707441 41657 707609
rect 0 706965 41713 707441
rect 0 706797 41657 706965
rect 0 706413 41713 706797
rect 0 706245 41657 706413
rect 0 705769 41713 706245
rect 42260 706194 42288 713675
rect 41892 706166 42288 706194
rect 0 705601 41657 705769
rect 41892 705713 41920 706166
rect 41713 705657 42193 705713
rect 0 705125 41713 705601
rect 0 704957 41657 705125
rect 0 704481 41713 704957
rect 0 704313 41657 704481
rect 41722 704425 41828 704426
rect 41713 704369 42193 704425
rect 0 703929 41713 704313
rect 41800 704002 41828 704369
rect 41788 703938 41840 704002
rect 0 703761 41657 703929
rect 0 703285 41713 703761
rect 0 703117 41657 703285
rect 0 702641 41713 703117
rect 0 702473 41657 702641
rect 0 702089 41713 702473
rect 0 701921 41657 702089
rect 0 701445 41713 701921
rect 0 701277 41657 701445
rect 41713 701333 42193 701389
rect 0 700801 41713 701277
rect 41800 700874 41828 701333
rect 41788 700810 41840 700874
rect 0 700633 41657 700801
rect 0 700249 41713 700633
rect 42444 704002 42472 718950
rect 42536 712298 42564 755414
rect 42628 744054 42656 787238
rect 673472 775878 673500 864418
rect 673564 785738 673592 874482
rect 673748 870602 673776 953294
rect 674012 872374 674064 872438
rect 673736 870538 673788 870602
rect 673920 870130 673972 870194
rect 673932 863258 673960 870130
rect 673920 863194 673972 863258
rect 673552 785674 673604 785738
rect 673460 775814 673512 775878
rect 42616 743990 42668 744054
rect 42524 712234 42576 712298
rect 42432 703938 42484 704002
rect 0 700081 41657 700249
rect 0 699605 41713 700081
rect 0 699437 41657 699605
rect 0 698961 41713 699437
rect 0 698793 41657 698961
rect 0 698409 41713 698793
rect 0 698241 41657 698409
rect 41713 698297 42193 698353
rect 0 698042 41713 698241
rect 0 670573 41713 670783
rect 0 670405 41657 670573
rect 41713 670503 42193 670517
rect 41713 670475 42288 670503
rect 41713 670461 42193 670475
rect 0 669929 41713 670405
rect 0 669761 41657 669929
rect 0 669285 41713 669761
rect 0 669117 41657 669285
rect 41713 669173 42193 669229
rect 0 668733 41713 669117
rect 0 668565 41657 668733
rect 41713 668621 42193 668677
rect 0 668089 41713 668565
rect 41800 668166 41828 668621
rect 41788 668102 41840 668166
rect 0 667921 41657 668089
rect 0 667445 41713 667921
rect 0 667277 41657 667445
rect 0 666893 41713 667277
rect 0 666725 41657 666893
rect 41713 666781 42193 666837
rect 0 666249 41713 666725
rect 0 666081 41657 666249
rect 0 665605 41713 666081
rect 0 665437 41657 665605
rect 41713 665493 42193 665549
rect 0 665053 41713 665437
rect 0 664885 41657 665053
rect 0 664409 41713 664885
rect 0 664241 41657 664409
rect 0 663765 41713 664241
rect 0 663597 41657 663765
rect 0 663213 41713 663597
rect 0 663045 41657 663213
rect 0 662569 41713 663045
rect 0 662401 41657 662569
rect 42260 662538 42288 670475
rect 41708 662510 42288 662538
rect 41708 662485 42193 662510
rect 41713 662457 42193 662485
rect 0 661925 41713 662401
rect 0 661757 41657 661925
rect 0 661281 41713 661757
rect 0 661113 41657 661281
rect 41713 661169 42193 661225
rect 0 660729 41713 661113
rect 41800 661094 41828 661169
rect 41788 661030 41840 661094
rect 0 660561 41657 660729
rect 0 660085 41713 660561
rect 0 659917 41657 660085
rect 0 659441 41713 659917
rect 0 659273 41657 659441
rect 0 658889 41713 659273
rect 0 658721 41657 658889
rect 0 658245 41713 658721
rect 41788 658650 41840 658714
rect 0 658077 41657 658245
rect 41800 658189 41828 658650
rect 41713 658133 42193 658189
rect 0 657601 41713 658077
rect 42444 661094 42472 703938
rect 42536 668166 42564 712234
rect 42628 700874 42656 743990
rect 673472 730930 673500 775814
rect 673564 740382 673592 785674
rect 674024 782338 674052 872374
rect 673644 782274 673696 782338
rect 674012 782274 674064 782338
rect 673552 740318 673604 740382
rect 673656 738138 673684 782274
rect 673828 740318 673880 740382
rect 673644 738074 673696 738138
rect 673460 730866 673512 730930
rect 42616 700810 42668 700874
rect 42524 668102 42576 668166
rect 42432 661030 42484 661094
rect 0 657433 41657 657601
rect 0 657049 41713 657433
rect 0 656881 41657 657049
rect 0 656405 41713 656881
rect 0 656237 41657 656405
rect 0 655761 41713 656237
rect 0 655593 41657 655761
rect 0 655209 41713 655593
rect 0 655041 41657 655209
rect 41713 655097 42193 655153
rect 0 654842 41713 655041
rect 0 627373 41713 627583
rect 0 627205 41657 627373
rect 41713 627314 42193 627317
rect 41713 627286 42288 627314
rect 41713 627261 42193 627286
rect 0 626729 41713 627205
rect 0 626561 41657 626729
rect 0 626085 41713 626561
rect 0 625917 41657 626085
rect 41713 625973 42193 626029
rect 0 625533 41713 625917
rect 0 625365 41657 625533
rect 41713 625421 42193 625477
rect 0 624889 41713 625365
rect 41800 624986 41828 625421
rect 41788 624922 41840 624986
rect 0 624721 41657 624889
rect 0 624245 41713 624721
rect 0 624077 41657 624245
rect 0 623693 41713 624077
rect 0 623525 41657 623693
rect 41713 623581 42193 623637
rect 0 623049 41713 623525
rect 0 622881 41657 623049
rect 0 622405 41713 622881
rect 0 622237 41657 622405
rect 41713 622293 42193 622349
rect 0 621853 41713 622237
rect 0 621685 41657 621853
rect 0 621209 41713 621685
rect 0 621041 41657 621209
rect 0 620565 41713 621041
rect 0 620397 41657 620565
rect 0 620013 41713 620397
rect 0 619845 41657 620013
rect 0 619369 41713 619845
rect 42260 619426 42288 627286
rect 41800 619398 42288 619426
rect 0 619201 41657 619369
rect 41800 619313 41828 619398
rect 41713 619257 42193 619313
rect 0 618725 41713 619201
rect 0 618557 41657 618725
rect 0 618081 41713 618557
rect 41788 618462 41840 618526
rect 0 617913 41657 618081
rect 41800 618025 41828 618462
rect 41713 617969 42193 618025
rect 0 617529 41713 617913
rect 0 617361 41657 617529
rect 0 616885 41713 617361
rect 0 616717 41657 616885
rect 0 616241 41713 616717
rect 0 616073 41657 616241
rect 0 615689 41713 616073
rect 0 615521 41657 615689
rect 0 615045 41713 615521
rect 41788 615470 41840 615534
rect 0 614877 41657 615045
rect 41800 614989 41828 615470
rect 41713 614933 42193 614989
rect 0 614401 41713 614877
rect 0 614233 41657 614401
rect 42444 618526 42472 661030
rect 42536 624986 42564 668102
rect 42628 658714 42656 700810
rect 673460 695302 673512 695366
rect 42616 658650 42668 658714
rect 42524 624922 42576 624986
rect 42432 618462 42484 618526
rect 0 613849 41713 614233
rect 0 613681 41657 613849
rect 0 613205 41713 613681
rect 0 613037 41657 613205
rect 0 612561 41713 613037
rect 0 612393 41657 612561
rect 0 612009 41713 612393
rect 0 611841 41657 612009
rect 41713 611897 42193 611953
rect 0 611642 41713 611841
rect 0 584173 41713 584383
rect 0 584005 41657 584173
rect 41713 584103 42193 584117
rect 41713 584075 42288 584103
rect 41713 584061 42193 584075
rect 0 583529 41713 584005
rect 0 583361 41657 583529
rect 0 582885 41713 583361
rect 0 582717 41657 582885
rect 41713 582773 42193 582829
rect 0 582333 41713 582717
rect 0 582165 41657 582333
rect 41713 582221 42193 582277
rect 0 581689 41713 582165
rect 41800 581738 41828 582221
rect 0 581521 41657 581689
rect 41788 581674 41840 581738
rect 0 581045 41713 581521
rect 0 580877 41657 581045
rect 0 580493 41713 580877
rect 0 580325 41657 580493
rect 41713 580381 42193 580437
rect 0 579849 41713 580325
rect 0 579681 41657 579849
rect 0 579205 41713 579681
rect 0 579037 41657 579205
rect 41713 579093 42193 579149
rect 0 578653 41713 579037
rect 0 578485 41657 578653
rect 0 578009 41713 578485
rect 0 577841 41657 578009
rect 0 577365 41713 577841
rect 0 577197 41657 577365
rect 0 576813 41713 577197
rect 0 576645 41657 576813
rect 0 576169 41713 576645
rect 42260 576178 42288 584075
rect 0 576001 41657 576169
rect 41800 576150 42288 576178
rect 41800 576113 41828 576150
rect 41713 576057 42193 576113
rect 0 575525 41713 576001
rect 0 575357 41657 575525
rect 42444 603106 42472 618462
rect 42536 603226 42564 624922
rect 42628 615534 42656 658650
rect 673472 650554 673500 695302
rect 673656 692306 673684 738074
rect 673840 695366 673868 740318
rect 673920 730866 673972 730930
rect 673828 695302 673880 695366
rect 673644 692242 673696 692306
rect 673552 685170 673604 685234
rect 673460 650490 673512 650554
rect 42616 615470 42668 615534
rect 42628 612734 42656 615470
rect 42628 612706 42840 612734
rect 42524 603162 42576 603226
rect 42444 603078 42656 603106
rect 42524 602958 42576 603022
rect 42536 585134 42564 602958
rect 42628 593414 42656 603078
rect 42628 593386 42748 593414
rect 42444 585106 42564 585134
rect 42444 581738 42472 585106
rect 42432 581674 42484 581738
rect 0 574881 41713 575357
rect 41788 575214 41840 575278
rect 0 574713 41657 574881
rect 41800 574825 41828 575214
rect 41713 574769 42193 574825
rect 0 574329 41713 574713
rect 0 574161 41657 574329
rect 0 573685 41713 574161
rect 0 573517 41657 573685
rect 0 573041 41713 573517
rect 0 572873 41657 573041
rect 0 572489 41713 572873
rect 0 572321 41657 572489
rect 0 571845 41713 572321
rect 41788 572222 41840 572286
rect 0 571677 41657 571845
rect 41800 571789 41828 572222
rect 41713 571733 42193 571789
rect 0 571201 41713 571677
rect 0 571033 41657 571201
rect 42248 571134 42300 571198
rect 0 570649 41713 571033
rect 0 570481 41657 570649
rect 0 570005 41713 570481
rect 0 569837 41657 570005
rect 0 569361 41713 569837
rect 0 569193 41657 569361
rect 0 568809 41713 569193
rect 0 568641 41657 568809
rect 41713 568697 42193 568753
rect 0 568442 41713 568641
rect 42260 543114 42288 571134
rect 42248 543050 42300 543114
rect 0 540973 41713 541183
rect 0 540805 41657 540973
rect 41713 540903 42193 540917
rect 41713 540875 42288 540903
rect 41713 540861 42193 540875
rect 0 540329 41713 540805
rect 0 540161 41657 540329
rect 0 539685 41713 540161
rect 0 539517 41657 539685
rect 41713 539573 42193 539629
rect 0 539133 41713 539517
rect 41788 539446 41840 539510
rect 0 538965 41657 539133
rect 41800 539077 41828 539446
rect 41713 539021 42193 539077
rect 0 538489 41713 538965
rect 0 538321 41657 538489
rect 0 537845 41713 538321
rect 0 537677 41657 537845
rect 0 537293 41713 537677
rect 0 537125 41657 537293
rect 41713 537181 42193 537237
rect 0 536649 41713 537125
rect 0 536481 41657 536649
rect 0 536005 41713 536481
rect 0 535837 41657 536005
rect 41713 535893 42193 535949
rect 0 535453 41713 535837
rect 0 535285 41657 535453
rect 0 534809 41713 535285
rect 0 534641 41657 534809
rect 0 534165 41713 534641
rect 0 533997 41657 534165
rect 0 533613 41713 533997
rect 0 533445 41657 533613
rect 0 532969 41713 533445
rect 42260 533066 42288 540875
rect 41800 533038 42288 533066
rect 0 532801 41657 532969
rect 41800 532913 41828 533038
rect 41713 532857 42193 532913
rect 0 532325 41713 532801
rect 0 532157 41657 532325
rect 0 531681 41713 532157
rect 42444 571198 42472 581674
rect 42720 575278 42748 593386
rect 42708 575214 42760 575278
rect 42524 572222 42576 572286
rect 42432 571134 42484 571198
rect 42432 543050 42484 543114
rect 42444 539510 42472 543050
rect 42432 539446 42484 539510
rect 0 531513 41657 531681
rect 41713 531569 42193 531625
rect 0 531129 41713 531513
rect 41800 531214 41828 531569
rect 41788 531150 41840 531214
rect 0 530961 41657 531129
rect 0 530485 41713 530961
rect 0 530317 41657 530485
rect 0 529841 41713 530317
rect 0 529673 41657 529841
rect 0 529289 41713 529673
rect 0 529121 41657 529289
rect 0 528645 41713 529121
rect 0 528477 41657 528645
rect 41713 528533 42193 528589
rect 0 528001 41713 528477
rect 41800 528086 41828 528533
rect 41788 528022 41840 528086
rect 0 527833 41657 528001
rect 42536 528086 42564 572222
rect 42720 554774 42748 575214
rect 42812 572286 42840 612706
rect 673472 605130 673500 650490
rect 673564 640694 673592 685170
rect 673656 647086 673684 692242
rect 673932 685234 673960 730866
rect 673920 685170 673972 685234
rect 673644 647022 673696 647086
rect 673552 640630 673604 640694
rect 673460 605066 673512 605130
rect 42800 572222 42852 572286
rect 673472 559978 673500 605066
rect 673564 595678 673592 640630
rect 673656 602954 673684 647022
rect 673644 602890 673696 602954
rect 673828 602890 673880 602954
rect 673552 595614 673604 595678
rect 673460 559914 673512 559978
rect 42628 554746 42748 554774
rect 42628 531214 42656 554746
rect 42708 539446 42760 539510
rect 42616 531150 42668 531214
rect 42524 528022 42576 528086
rect 0 527449 41713 527833
rect 0 527281 41657 527449
rect 0 526805 41713 527281
rect 0 526637 41657 526805
rect 0 526161 41713 526637
rect 0 525993 41657 526161
rect 0 525609 41713 525993
rect 0 525441 41657 525609
rect 41713 525497 42193 525553
rect 0 525242 41713 525441
rect 985 493078 40000 497858
rect 985 487879 39593 493078
rect 39616 488179 40000 488579
rect 985 483099 40000 487879
rect 985 483053 39593 483099
rect 7 456040 30281 457987
rect 30753 455800 31683 458028
rect 32033 456040 34915 457987
rect 7 455740 39593 455800
rect 7 451619 39600 455740
rect 7 451507 39593 451619
rect 7 444985 39600 451507
rect 7 444899 39593 444985
rect 7 440900 39600 444899
rect 7 440800 39593 440900
rect 30760 438605 31690 440800
rect 0 413373 41713 413583
rect 0 413205 41657 413373
rect 41713 413303 42193 413317
rect 41713 413275 42288 413303
rect 41713 413261 42193 413275
rect 0 412729 41713 413205
rect 0 412561 41657 412729
rect 0 412085 41713 412561
rect 0 411917 41657 412085
rect 41713 411973 42193 412029
rect 0 411533 41713 411917
rect 0 411365 41657 411533
rect 41722 411477 41828 411482
rect 41713 411421 42193 411477
rect 0 410889 41713 411365
rect 41800 410990 41828 411421
rect 41788 410926 41840 410990
rect 0 410721 41657 410889
rect 0 410245 41713 410721
rect 0 410077 41657 410245
rect 0 409693 41713 410077
rect 0 409525 41657 409693
rect 41713 409581 42193 409637
rect 0 409049 41713 409525
rect 0 408881 41657 409049
rect 0 408405 41713 408881
rect 0 408237 41657 408405
rect 41713 408293 42193 408349
rect 0 407853 41713 408237
rect 0 407685 41657 407853
rect 0 407209 41713 407685
rect 0 407041 41657 407209
rect 0 406565 41713 407041
rect 0 406397 41657 406565
rect 0 406013 41713 406397
rect 0 405845 41657 406013
rect 0 405369 41713 405845
rect 42260 405498 42288 413275
rect 41800 405470 42288 405498
rect 0 405201 41657 405369
rect 41800 405313 41828 405470
rect 41713 405257 42193 405313
rect 42432 410926 42484 410990
rect 0 404725 41713 405201
rect 0 404557 41657 404725
rect 0 404081 41713 404557
rect 41788 404466 41840 404530
rect 0 403913 41657 404081
rect 41800 404025 41828 404466
rect 41713 403969 42193 404025
rect 0 403529 41713 403913
rect 0 403361 41657 403529
rect 0 402885 41713 403361
rect 0 402717 41657 402885
rect 0 402241 41713 402717
rect 0 402073 41657 402241
rect 0 401689 41713 402073
rect 0 401521 41657 401689
rect 0 401045 41713 401521
rect 41788 401474 41840 401538
rect 0 400877 41657 401045
rect 41800 400989 41828 401474
rect 41713 400933 42193 400989
rect 0 400401 41713 400877
rect 0 400233 41657 400401
rect 0 399849 41713 400233
rect 0 399681 41657 399849
rect 0 399205 41713 399681
rect 0 399037 41657 399205
rect 0 398561 41713 399037
rect 0 398393 41657 398561
rect 0 398009 41713 398393
rect 0 397841 41657 398009
rect 41713 397897 42193 397953
rect 0 397642 41713 397841
rect 0 370173 41713 370383
rect 0 370005 41657 370173
rect 41713 370061 42193 370117
rect 0 369529 41713 370005
rect 41800 369578 41828 370061
rect 0 369361 41657 369529
rect 41788 369514 41840 369578
rect 0 368885 41713 369361
rect 0 368717 41657 368885
rect 41713 368773 42193 368829
rect 0 368333 41713 368717
rect 41788 368630 41840 368694
rect 0 368165 41657 368333
rect 41800 368277 41828 368630
rect 41713 368221 42193 368277
rect 0 367689 41713 368165
rect 0 367521 41657 367689
rect 0 367045 41713 367521
rect 0 366877 41657 367045
rect 0 366493 41713 366877
rect 0 366325 41657 366493
rect 41713 366381 42193 366437
rect 0 365849 41713 366325
rect 0 365681 41657 365849
rect 0 365205 41713 365681
rect 0 365037 41657 365205
rect 41713 365093 42193 365149
rect 0 364653 41713 365037
rect 0 364485 41657 364653
rect 0 364009 41713 364485
rect 0 363841 41657 364009
rect 0 363365 41713 363841
rect 0 363197 41657 363365
rect 0 362813 41713 363197
rect 0 362645 41657 362813
rect 0 362169 41713 362645
rect 41788 362578 41840 362642
rect 0 362001 41657 362169
rect 41800 362114 41828 362578
rect 41722 362113 41828 362114
rect 41713 362057 42193 362113
rect 0 361525 41713 362001
rect 0 361357 41657 361525
rect 42340 369514 42392 369578
rect 42352 362642 42380 369514
rect 42444 368694 42472 410926
rect 42536 401538 42564 528022
rect 42628 404530 42656 531150
rect 42720 410990 42748 539446
rect 42708 410926 42760 410990
rect 42616 404466 42668 404530
rect 42524 401474 42576 401538
rect 42432 368630 42484 368694
rect 42340 362578 42392 362642
rect 42444 361574 42472 368630
rect 42444 361546 42564 361574
rect 0 360881 41713 361357
rect 0 360713 41657 360881
rect 41713 360769 42193 360825
rect 41800 360738 41828 360769
rect 0 360329 41713 360713
rect 41788 360674 41840 360738
rect 0 360161 41657 360329
rect 0 359685 41713 360161
rect 0 359517 41657 359685
rect 0 359041 41713 359517
rect 0 358873 41657 359041
rect 0 358489 41713 358873
rect 0 358321 41657 358489
rect 0 357845 41713 358321
rect 0 357677 41657 357845
rect 41713 357733 42193 357789
rect 0 357201 41713 357677
rect 41800 357270 41828 357733
rect 41788 357206 41840 357270
rect 0 357033 41657 357201
rect 0 356649 41713 357033
rect 42340 357206 42392 357270
rect 0 356481 41657 356649
rect 0 356005 41713 356481
rect 0 355837 41657 356005
rect 0 355361 41713 355837
rect 0 355193 41657 355361
rect 0 354809 41713 355193
rect 0 354641 41657 354809
rect 41713 354697 42193 354753
rect 0 354442 41713 354641
rect 42352 342254 42380 357206
rect 42352 342226 42472 342254
rect 0 326973 41713 327183
rect 0 326805 41657 326973
rect 41713 326861 42193 326917
rect 0 326329 41713 326805
rect 41800 326754 41828 326861
rect 41800 326726 42288 326754
rect 0 326161 41657 326329
rect 0 325685 41713 326161
rect 0 325517 41657 325685
rect 41713 325573 42193 325629
rect 0 325133 41713 325517
rect 41788 325450 41840 325514
rect 0 324965 41657 325133
rect 41800 325077 41828 325450
rect 41713 325021 42193 325077
rect 0 324489 41713 324965
rect 0 324321 41657 324489
rect 0 323845 41713 324321
rect 0 323677 41657 323845
rect 0 323293 41713 323677
rect 0 323125 41657 323293
rect 41713 323181 42193 323237
rect 0 322649 41713 323125
rect 0 322481 41657 322649
rect 0 322005 41713 322481
rect 0 321837 41657 322005
rect 41713 321893 42193 321949
rect 0 321453 41713 321837
rect 0 321285 41657 321453
rect 0 320809 41713 321285
rect 0 320641 41657 320809
rect 0 320165 41713 320641
rect 0 319997 41657 320165
rect 0 319613 41713 319997
rect 0 319445 41657 319613
rect 0 318969 41713 319445
rect 0 318801 41657 318969
rect 41713 318899 42193 318913
rect 42260 318899 42288 326726
rect 41713 318871 42288 318899
rect 41713 318857 42193 318871
rect 0 318325 41713 318801
rect 0 318157 41657 318325
rect 0 317681 41713 318157
rect 0 317513 41657 317681
rect 41713 317569 42193 317625
rect 0 317129 41713 317513
rect 41800 317218 41828 317569
rect 41788 317154 41840 317218
rect 0 316961 41657 317129
rect 0 316485 41713 316961
rect 0 316317 41657 316485
rect 0 315841 41713 316317
rect 0 315673 41657 315841
rect 0 315289 41713 315673
rect 0 315121 41657 315289
rect 0 314645 41713 315121
rect 0 314477 41657 314645
rect 41713 314533 42193 314589
rect 0 314001 41713 314477
rect 41800 314090 41828 314533
rect 41788 314026 41840 314090
rect 0 313833 41657 314001
rect 42444 314090 42472 342226
rect 42536 325514 42564 361546
rect 42628 360738 42656 404466
rect 42708 401474 42760 401538
rect 42616 360674 42668 360738
rect 42524 325450 42576 325514
rect 42628 322934 42656 360674
rect 42720 357270 42748 401474
rect 673472 383586 673500 559914
rect 673840 557870 673868 602890
rect 673920 595614 673972 595678
rect 673828 557806 673880 557870
rect 673932 550526 673960 595614
rect 673920 550462 673972 550526
rect 673932 546494 673960 550462
rect 673840 546466 673960 546494
rect 673460 383522 673512 383586
rect 673472 380894 673500 383522
rect 673472 380866 673592 380894
rect 673460 372302 673512 372366
rect 42708 357206 42760 357270
rect 673472 328098 673500 372302
rect 673564 337550 673592 380866
rect 673736 379646 673788 379710
rect 673552 337486 673604 337550
rect 673460 328034 673512 328098
rect 42708 325450 42760 325514
rect 42536 322906 42656 322934
rect 42536 317218 42564 322906
rect 42524 317154 42576 317218
rect 42432 314026 42484 314090
rect 0 313449 41713 313833
rect 0 313281 41657 313449
rect 0 312805 41713 313281
rect 0 312637 41657 312805
rect 0 312161 41713 312637
rect 0 311993 41657 312161
rect 0 311609 41713 311993
rect 0 311441 41657 311609
rect 41713 311497 42193 311553
rect 0 311242 41713 311441
rect 0 283773 41713 283983
rect 0 283605 41657 283773
rect 41713 283703 42193 283717
rect 41713 283675 42288 283703
rect 41713 283661 42193 283675
rect 0 283129 41713 283605
rect 0 282961 41657 283129
rect 0 282485 41713 282961
rect 0 282317 41657 282485
rect 41713 282373 42193 282429
rect 0 281933 41713 282317
rect 0 281765 41657 281933
rect 41713 281821 42193 281877
rect 0 281289 41713 281765
rect 41800 281382 41828 281821
rect 41788 281318 41840 281382
rect 0 281121 41657 281289
rect 0 280645 41713 281121
rect 0 280477 41657 280645
rect 0 280093 41713 280477
rect 0 279925 41657 280093
rect 41713 279981 42193 280037
rect 0 279449 41713 279925
rect 0 279281 41657 279449
rect 0 278805 41713 279281
rect 0 278637 41657 278805
rect 41713 278693 42193 278749
rect 0 278253 41713 278637
rect 0 278085 41657 278253
rect 0 277609 41713 278085
rect 0 277441 41657 277609
rect 0 276965 41713 277441
rect 0 276797 41657 276965
rect 0 276413 41713 276797
rect 0 276245 41657 276413
rect 0 275769 41713 276245
rect 0 275601 41657 275769
rect 41713 275699 42193 275713
rect 42260 275699 42288 283675
rect 41713 275671 42288 275699
rect 41713 275657 42193 275671
rect 0 275125 41713 275601
rect 42432 281318 42484 281382
rect 0 274957 41657 275125
rect 0 274481 41713 274957
rect 41788 274518 41840 274582
rect 0 274313 41657 274481
rect 41800 274425 41828 274518
rect 41713 274369 42193 274425
rect 41722 274366 41828 274369
rect 0 273929 41713 274313
rect 0 273761 41657 273929
rect 0 273285 41713 273761
rect 0 273117 41657 273285
rect 0 272641 41713 273117
rect 0 272473 41657 272641
rect 0 272089 41713 272473
rect 0 271921 41657 272089
rect 0 271445 41713 271921
rect 41788 271866 41840 271930
rect 0 271277 41657 271445
rect 41800 271402 41828 271866
rect 41722 271389 41828 271402
rect 41713 271333 42193 271389
rect 0 270801 41713 271277
rect 0 270633 41657 270801
rect 0 270249 41713 270633
rect 0 270081 41657 270249
rect 0 269605 41713 270081
rect 0 269437 41657 269605
rect 0 268961 41713 269437
rect 0 268793 41657 268961
rect 0 268409 41713 268793
rect 0 268241 41657 268409
rect 41713 268297 42193 268353
rect 0 268042 41713 268241
rect 0 240573 41713 240783
rect 0 240405 41657 240573
rect 41722 240517 42288 240530
rect 41713 240502 42288 240517
rect 41713 240461 42193 240502
rect 0 239929 41713 240405
rect 0 239761 41657 239929
rect 0 239285 41713 239761
rect 0 239117 41657 239285
rect 41713 239173 42193 239229
rect 0 238733 41713 239117
rect 0 238565 41657 238733
rect 41713 238621 42193 238677
rect 0 238089 41713 238565
rect 41800 238134 41828 238621
rect 0 237921 41657 238089
rect 41788 238070 41840 238134
rect 0 237445 41713 237921
rect 0 237277 41657 237445
rect 41713 237333 42193 237389
rect 0 236893 41713 237277
rect 0 236725 41657 236893
rect 41713 236781 42193 236837
rect 0 236249 41713 236725
rect 0 236081 41657 236249
rect 0 235605 41713 236081
rect 0 235437 41657 235605
rect 41713 235493 42193 235549
rect 0 235053 41713 235437
rect 0 234885 41657 235053
rect 0 234409 41713 234885
rect 0 234241 41657 234409
rect 0 233765 41713 234241
rect 0 233597 41657 233765
rect 0 233213 41713 233597
rect 0 233045 41657 233213
rect 0 232569 41713 233045
rect 42260 232642 42288 240502
rect 41800 232614 42288 232642
rect 0 232401 41657 232569
rect 41800 232513 41828 232614
rect 41713 232457 42193 232513
rect 0 231925 41713 232401
rect 0 231757 41657 231925
rect 42444 238134 42472 281318
rect 42536 274582 42564 317154
rect 42616 314026 42668 314090
rect 42524 274518 42576 274582
rect 42432 238070 42484 238134
rect 0 231281 41713 231757
rect 41788 231678 41840 231742
rect 0 231113 41657 231281
rect 41800 231225 41828 231678
rect 41713 231169 42193 231225
rect 0 230729 41713 231113
rect 0 230561 41657 230729
rect 0 230085 41713 230561
rect 0 229917 41657 230085
rect 0 229441 41713 229917
rect 0 229273 41657 229441
rect 0 228889 41713 229273
rect 0 228721 41657 228889
rect 0 228245 41713 228721
rect 41788 228618 41840 228682
rect 0 228077 41657 228245
rect 41800 228189 41828 228618
rect 41713 228133 42193 228189
rect 41722 228126 41828 228133
rect 0 227601 41713 228077
rect 0 227433 41657 227601
rect 42248 227462 42300 227526
rect 0 227049 41713 227433
rect 0 226881 41657 227049
rect 0 226405 41713 226881
rect 0 226237 41657 226405
rect 0 225761 41713 226237
rect 0 225593 41657 225761
rect 0 225209 41713 225593
rect 0 225041 41657 225209
rect 41713 225097 42193 225153
rect 0 224842 41713 225041
rect 0 197373 41713 197583
rect 42260 197418 42288 227462
rect 42444 197538 42472 238070
rect 42536 231742 42564 274518
rect 42628 271930 42656 314026
rect 42720 281382 42748 325450
rect 673472 313274 673500 328034
rect 673460 313210 673512 313274
rect 673564 295334 673592 337486
rect 673748 334490 673776 379646
rect 673840 372366 673868 546466
rect 674760 427854 674788 992190
rect 675887 967359 717600 967558
rect 675407 967247 675887 967303
rect 675943 967191 717600 967359
rect 675887 966807 717600 967191
rect 675943 966639 717600 966807
rect 675887 966163 717600 966639
rect 675943 965995 717600 966163
rect 675887 965519 717600 965995
rect 675943 965351 717600 965519
rect 675887 964967 717600 965351
rect 675943 964799 717600 964967
rect 675392 964718 675444 964782
rect 675404 964267 675432 964718
rect 675887 964323 717600 964799
rect 675404 964239 675887 964267
rect 675407 964211 675887 964239
rect 675943 964155 717600 964323
rect 675887 963679 717600 964155
rect 675943 963511 717600 963679
rect 675887 963127 717600 963511
rect 675943 962959 717600 963127
rect 675887 962483 717600 962959
rect 675943 962315 717600 962483
rect 675887 961839 717600 962315
rect 675943 961671 717600 961839
rect 675392 961318 675444 961382
rect 675404 961231 675432 961318
rect 675887 961287 717600 961671
rect 675404 961180 675887 961231
rect 675407 961175 675887 961180
rect 675943 961119 717600 961287
rect 675887 960643 717600 961119
rect 675943 960475 717600 960643
rect 675887 959999 717600 960475
rect 675407 959929 675887 959943
rect 675312 959901 675887 959929
rect 675312 951810 675340 959901
rect 675407 959887 675887 959901
rect 675943 959831 717600 959999
rect 675887 959355 717600 959831
rect 675943 959187 717600 959355
rect 675887 958803 717600 959187
rect 675943 958635 717600 958803
rect 675887 958159 717600 958635
rect 675943 957991 717600 958159
rect 675887 957515 717600 957991
rect 675943 957347 717600 957515
rect 675887 956963 717600 957347
rect 675407 956851 675887 956907
rect 675943 956795 717600 956963
rect 675887 956319 717600 956795
rect 675943 956151 717600 956319
rect 675887 955675 717600 956151
rect 675407 955563 675887 955619
rect 675943 955507 717600 955675
rect 675887 955123 717600 955507
rect 675943 954955 717600 955123
rect 675887 954479 717600 954955
rect 675943 954311 717600 954479
rect 675887 953835 717600 954311
rect 675407 953751 675887 953779
rect 675404 953723 675887 953751
rect 675404 953358 675432 953723
rect 675943 953667 717600 953835
rect 675392 953294 675444 953358
rect 675887 953283 717600 953667
rect 675407 953171 675887 953227
rect 675943 953115 717600 953283
rect 675887 952639 717600 953115
rect 675943 952471 717600 952639
rect 675887 951995 717600 952471
rect 675407 951932 675887 951939
rect 675404 951883 675887 951932
rect 675404 951810 675432 951883
rect 675943 951827 717600 951995
rect 675312 951782 675432 951810
rect 675887 951617 717600 951827
rect 685910 922600 686840 924795
rect 678007 922500 717593 922600
rect 678000 918501 717593 922500
rect 678007 918415 717593 918501
rect 678000 911893 717593 918415
rect 678007 911781 717593 911893
rect 678000 907660 717593 911781
rect 678007 907600 717593 907660
rect 682685 905413 685567 907360
rect 685917 905372 686847 907600
rect 687319 905413 717593 907360
rect 675887 878159 717600 878358
rect 675407 878047 675887 878103
rect 675943 877991 717600 878159
rect 675887 877607 717600 877991
rect 675943 877439 717600 877607
rect 675887 876963 717600 877439
rect 675943 876795 717600 876963
rect 675887 876319 717600 876795
rect 675943 876151 717600 876319
rect 675887 875767 717600 876151
rect 675943 875599 717600 875767
rect 675887 875123 717600 875599
rect 675407 875039 675887 875067
rect 675404 875011 675887 875039
rect 675404 874546 675432 875011
rect 675943 874955 717600 875123
rect 675392 874482 675444 874546
rect 675887 874479 717600 874955
rect 675943 874311 717600 874479
rect 675887 873927 717600 874311
rect 675943 873759 717600 873927
rect 675887 873283 717600 873759
rect 675943 873115 717600 873283
rect 675887 872639 717600 873115
rect 675943 872471 717600 872639
rect 675392 872374 675444 872438
rect 675404 872031 675432 872374
rect 675887 872087 717600 872471
rect 675404 872003 675887 872031
rect 675407 871975 675887 872003
rect 675943 871919 717600 872087
rect 675887 871443 717600 871919
rect 675943 871275 717600 871443
rect 675887 870799 717600 871275
rect 675407 870740 675887 870743
rect 675404 870687 675887 870740
rect 675404 870194 675432 870687
rect 675943 870631 717600 870799
rect 675392 870130 675444 870194
rect 675887 870155 717600 870631
rect 675943 869987 717600 870155
rect 675887 869603 717600 869987
rect 675943 869435 717600 869603
rect 675887 868959 717600 869435
rect 675943 868791 717600 868959
rect 675887 868315 717600 868791
rect 675943 868147 717600 868315
rect 675887 867763 717600 868147
rect 675407 867651 675887 867707
rect 675943 867595 717600 867763
rect 675887 867119 717600 867595
rect 675943 866951 717600 867119
rect 675887 866475 717600 866951
rect 675407 866363 675887 866419
rect 675943 866307 717600 866475
rect 675887 865923 717600 866307
rect 675943 865755 717600 865923
rect 675887 865279 717600 865755
rect 675943 865111 717600 865279
rect 675887 864635 717600 865111
rect 675407 864551 675887 864579
rect 675404 864523 675887 864551
rect 675404 864482 675432 864523
rect 675392 864418 675444 864482
rect 675943 864467 717600 864635
rect 675887 864083 717600 864467
rect 675407 863971 675887 864027
rect 675943 863915 717600 864083
rect 675887 863439 717600 863915
rect 675943 863271 717600 863439
rect 675392 863194 675444 863258
rect 675404 862739 675432 863194
rect 675887 862795 717600 863271
rect 675404 862716 675887 862739
rect 675407 862683 675887 862716
rect 675943 862627 717600 862795
rect 675887 862417 717600 862627
rect 678007 833301 716615 833347
rect 677600 828521 716615 833301
rect 677600 827821 677984 828221
rect 678007 823322 716615 828521
rect 677600 818542 716615 823322
rect 675300 818314 675352 818378
rect 677598 818343 677654 818417
rect 677600 818314 677652 818343
rect 675312 786614 675340 818314
rect 675887 788959 717600 789158
rect 675407 788847 675887 788903
rect 675943 788791 717600 788959
rect 675887 788407 717600 788791
rect 675943 788239 717600 788407
rect 675887 787763 717600 788239
rect 675943 787595 717600 787763
rect 675887 787119 717600 787595
rect 675943 786951 717600 787119
rect 675128 786586 675340 786614
rect 675128 728906 675156 786586
rect 675887 786567 717600 786951
rect 675943 786399 717600 786567
rect 675887 785923 717600 786399
rect 675407 785839 675887 785867
rect 675404 785811 675887 785839
rect 675404 785738 675432 785811
rect 675943 785755 717600 785923
rect 675392 785674 675444 785738
rect 675887 785279 717600 785755
rect 675943 785111 717600 785279
rect 675887 784727 717600 785111
rect 675943 784559 717600 784727
rect 675887 784083 717600 784559
rect 675943 783915 717600 784083
rect 675887 783439 717600 783915
rect 675943 783271 717600 783439
rect 675887 782887 717600 783271
rect 675407 782803 675887 782831
rect 675404 782775 675887 782803
rect 675404 782338 675432 782775
rect 675943 782719 717600 782887
rect 675392 782274 675444 782338
rect 675887 782243 717600 782719
rect 675943 782075 717600 782243
rect 675887 781599 717600 782075
rect 675407 781524 675887 781543
rect 675404 781487 675887 781524
rect 675404 781046 675432 781487
rect 675943 781431 717600 781599
rect 675208 780982 675260 781046
rect 675392 780982 675444 781046
rect 675220 773514 675248 780982
rect 675887 780955 717600 781431
rect 675943 780787 717600 780955
rect 675887 780403 717600 780787
rect 675943 780235 717600 780403
rect 675887 779759 717600 780235
rect 675943 779591 717600 779759
rect 675887 779115 717600 779591
rect 675943 778947 717600 779115
rect 675887 778563 717600 778947
rect 675407 778451 675887 778507
rect 675943 778395 717600 778563
rect 675887 777919 717600 778395
rect 675943 777751 717600 777919
rect 675887 777275 717600 777751
rect 675407 777163 675887 777219
rect 675943 777107 717600 777275
rect 675887 776723 717600 777107
rect 675943 776555 717600 776723
rect 675887 776079 717600 776555
rect 675943 775911 717600 776079
rect 675392 775814 675444 775878
rect 675404 775379 675432 775814
rect 675887 775435 717600 775911
rect 675404 775351 675887 775379
rect 675407 775323 675887 775351
rect 675943 775267 717600 775435
rect 675887 774883 717600 775267
rect 675407 774771 675887 774827
rect 675943 774715 717600 774883
rect 675887 774239 717600 774715
rect 675943 774071 717600 774239
rect 675887 773595 717600 774071
rect 675407 773514 675887 773539
rect 675220 773486 675887 773514
rect 675407 773483 675887 773486
rect 675943 773427 717600 773595
rect 675887 773217 717600 773427
rect 675887 743959 717600 744158
rect 675407 743847 675887 743903
rect 675943 743791 717600 743959
rect 675887 743407 717600 743791
rect 675943 743239 717600 743407
rect 675887 742763 717600 743239
rect 675943 742595 717600 742763
rect 675887 742119 717600 742595
rect 675943 741951 717600 742119
rect 675887 741567 717600 741951
rect 675943 741399 717600 741567
rect 675887 740923 717600 741399
rect 675407 740860 675887 740867
rect 675404 740811 675887 740860
rect 675404 740382 675432 740811
rect 675943 740755 717600 740923
rect 675392 740318 675444 740382
rect 675887 740279 717600 740755
rect 675943 740111 717600 740279
rect 675887 739727 717600 740111
rect 675943 739559 717600 739727
rect 675887 739083 717600 739559
rect 675943 738915 717600 739083
rect 675887 738439 717600 738915
rect 675943 738271 717600 738439
rect 675392 738074 675444 738138
rect 675404 737831 675432 738074
rect 675887 737887 717600 738271
rect 675404 737803 675887 737831
rect 675407 737775 675887 737803
rect 675943 737719 717600 737887
rect 675887 737243 717600 737719
rect 675943 737075 717600 737243
rect 675887 736599 717600 737075
rect 675407 736522 675887 736543
rect 675312 736494 675887 736522
rect 675312 729042 675340 736494
rect 675407 736487 675887 736494
rect 675943 736431 717600 736599
rect 675887 735955 717600 736431
rect 675943 735787 717600 735955
rect 675887 735403 717600 735787
rect 675943 735235 717600 735403
rect 675887 734759 717600 735235
rect 675943 734591 717600 734759
rect 675887 734115 717600 734591
rect 675943 733947 717600 734115
rect 675887 733563 717600 733947
rect 675407 733451 675887 733507
rect 675943 733395 717600 733563
rect 675887 732919 717600 733395
rect 675943 732751 717600 732919
rect 675887 732275 717600 732751
rect 675407 732163 675887 732219
rect 675943 732107 717600 732275
rect 675887 731723 717600 732107
rect 675943 731555 717600 731723
rect 675887 731079 717600 731555
rect 675392 730866 675444 730930
rect 675943 730911 717600 731079
rect 675404 730379 675432 730866
rect 675887 730435 717600 730911
rect 675404 730351 675887 730379
rect 675407 730323 675887 730351
rect 675943 730267 717600 730435
rect 675887 729883 717600 730267
rect 675407 729771 675887 729827
rect 675943 729715 717600 729883
rect 675887 729239 717600 729715
rect 675943 729071 717600 729239
rect 675312 729014 675432 729042
rect 675128 728878 675340 728906
rect 675312 701054 675340 728878
rect 675404 728539 675432 729014
rect 675887 728595 717600 729071
rect 675404 728484 675887 728539
rect 675407 728483 675887 728484
rect 675943 728427 717600 728595
rect 675887 728217 717600 728427
rect 675128 701026 675340 701054
rect 675128 681734 675156 701026
rect 675887 698959 717600 699158
rect 675407 698847 675887 698903
rect 675943 698791 717600 698959
rect 675887 698407 717600 698791
rect 675943 698239 717600 698407
rect 675887 697763 717600 698239
rect 675943 697595 717600 697763
rect 675887 697119 717600 697595
rect 675943 696951 717600 697119
rect 675887 696567 717600 696951
rect 675943 696399 717600 696567
rect 675887 695923 717600 696399
rect 675407 695844 675887 695867
rect 675404 695811 675887 695844
rect 675404 695366 675432 695811
rect 675943 695755 717600 695923
rect 675392 695302 675444 695366
rect 675887 695279 717600 695755
rect 675943 695111 717600 695279
rect 675887 694727 717600 695111
rect 675943 694559 717600 694727
rect 675887 694083 717600 694559
rect 675943 693915 717600 694083
rect 675887 693439 717600 693915
rect 675943 693271 717600 693439
rect 675887 692887 717600 693271
rect 675407 692803 675887 692831
rect 675404 692775 675887 692803
rect 675404 692306 675432 692775
rect 675943 692719 717600 692887
rect 675392 692242 675444 692306
rect 675887 692243 717600 692719
rect 675943 692075 717600 692243
rect 675312 691614 675432 691642
rect 675312 683525 675340 691614
rect 675404 691543 675432 691614
rect 675887 691599 717600 692075
rect 675404 691492 675887 691543
rect 675407 691487 675887 691492
rect 675943 691431 717600 691599
rect 675887 690955 717600 691431
rect 675943 690787 717600 690955
rect 675887 690403 717600 690787
rect 675943 690235 717600 690403
rect 675887 689759 717600 690235
rect 675943 689591 717600 689759
rect 675887 689115 717600 689591
rect 675943 688947 717600 689115
rect 675887 688563 717600 688947
rect 675407 688451 675887 688507
rect 675943 688395 717600 688563
rect 675887 687919 717600 688395
rect 675943 687751 717600 687919
rect 675887 687275 717600 687751
rect 675407 687163 675887 687219
rect 675943 687107 717600 687275
rect 675887 686723 717600 687107
rect 675943 686555 717600 686723
rect 675887 686079 717600 686555
rect 675943 685911 717600 686079
rect 675887 685435 717600 685911
rect 675407 685372 675887 685379
rect 675404 685323 675887 685372
rect 675404 685234 675432 685323
rect 675943 685267 717600 685435
rect 675392 685170 675444 685234
rect 675887 684883 717600 685267
rect 675407 684771 675887 684827
rect 675943 684715 717600 684883
rect 675887 684239 717600 684715
rect 675943 684071 717600 684239
rect 675887 683595 717600 684071
rect 675407 683525 675887 683539
rect 675312 683497 675887 683525
rect 675407 683483 675887 683497
rect 675943 683427 717600 683595
rect 675887 683217 717600 683427
rect 675128 681706 675340 681734
rect 675312 651374 675340 681706
rect 675887 653759 717600 653958
rect 675407 653647 675887 653703
rect 675943 653591 717600 653759
rect 675887 653207 717600 653591
rect 675943 653039 717600 653207
rect 675887 652563 717600 653039
rect 675943 652395 717600 652563
rect 675887 651919 717600 652395
rect 675943 651751 717600 651919
rect 675128 651346 675340 651374
rect 675887 651367 717600 651751
rect 675128 632054 675156 651346
rect 675943 651199 717600 651367
rect 675887 650723 717600 651199
rect 675407 650639 675887 650667
rect 675404 650611 675887 650639
rect 675404 650554 675432 650611
rect 675943 650555 717600 650723
rect 675392 650490 675444 650554
rect 675887 650079 717600 650555
rect 675943 649911 717600 650079
rect 675887 649527 717600 649911
rect 675943 649359 717600 649527
rect 675887 648883 717600 649359
rect 675943 648715 717600 648883
rect 675887 648239 717600 648715
rect 675943 648071 717600 648239
rect 675887 647687 717600 648071
rect 675407 647603 675887 647631
rect 675404 647575 675887 647603
rect 675404 647086 675432 647575
rect 675943 647519 717600 647687
rect 675392 647022 675444 647086
rect 675887 647043 717600 647519
rect 675943 646875 717600 647043
rect 675887 646399 717600 646875
rect 675407 646340 675887 646343
rect 675404 646287 675887 646340
rect 675404 645794 675432 646287
rect 675943 646231 717600 646399
rect 675208 645730 675260 645794
rect 675392 645730 675444 645794
rect 675887 645755 717600 646231
rect 675220 638330 675248 645730
rect 675943 645587 717600 645755
rect 675887 645203 717600 645587
rect 675943 645035 717600 645203
rect 675887 644559 717600 645035
rect 675943 644391 717600 644559
rect 675887 643915 717600 644391
rect 675943 643747 717600 643915
rect 675887 643363 717600 643747
rect 675407 643251 675887 643307
rect 675943 643195 717600 643363
rect 675887 642719 717600 643195
rect 675943 642551 717600 642719
rect 675887 642075 717600 642551
rect 675407 641963 675887 642019
rect 675943 641907 717600 642075
rect 675887 641523 717600 641907
rect 675943 641355 717600 641523
rect 675887 640879 717600 641355
rect 675943 640711 717600 640879
rect 675392 640630 675444 640694
rect 675404 640179 675432 640630
rect 675887 640235 717600 640711
rect 675404 640151 675887 640179
rect 675407 640123 675887 640151
rect 675943 640067 717600 640235
rect 675887 639683 717600 640067
rect 675407 639571 675887 639627
rect 675943 639515 717600 639683
rect 675887 639039 717600 639515
rect 675943 638871 717600 639039
rect 675887 638395 717600 638871
rect 675407 638330 675887 638339
rect 675220 638302 675887 638330
rect 675407 638283 675887 638302
rect 675943 638227 717600 638395
rect 675887 638017 717600 638227
rect 675128 632026 675340 632054
rect 675312 612734 675340 632026
rect 675128 612706 675340 612734
rect 675128 593722 675156 612706
rect 675887 608759 717600 608958
rect 675407 608647 675887 608703
rect 675943 608591 717600 608759
rect 675887 608207 717600 608591
rect 675943 608039 717600 608207
rect 675887 607563 717600 608039
rect 675943 607395 717600 607563
rect 675887 606919 717600 607395
rect 675943 606751 717600 606919
rect 675887 606367 717600 606751
rect 675943 606199 717600 606367
rect 675887 605723 717600 606199
rect 675407 605639 675887 605667
rect 675404 605611 675887 605639
rect 675404 605130 675432 605611
rect 675943 605555 717600 605723
rect 675392 605066 675444 605130
rect 675887 605079 717600 605555
rect 675943 604911 717600 605079
rect 675887 604527 717600 604911
rect 675943 604359 717600 604527
rect 675887 603883 717600 604359
rect 675943 603715 717600 603883
rect 675887 603239 717600 603715
rect 675943 603071 717600 603239
rect 675392 602890 675444 602954
rect 675404 602631 675432 602890
rect 675887 602687 717600 603071
rect 675404 602603 675887 602631
rect 675407 602575 675887 602603
rect 675943 602519 717600 602687
rect 675887 602043 717600 602519
rect 675943 601875 717600 602043
rect 675887 601399 717600 601875
rect 675407 601338 675887 601343
rect 675312 601310 675887 601338
rect 675312 593858 675340 601310
rect 675407 601287 675887 601310
rect 675943 601231 717600 601399
rect 675887 600755 717600 601231
rect 675943 600587 717600 600755
rect 675887 600203 717600 600587
rect 675943 600035 717600 600203
rect 675887 599559 717600 600035
rect 675943 599391 717600 599559
rect 675887 598915 717600 599391
rect 675943 598747 717600 598915
rect 675887 598363 717600 598747
rect 675407 598251 675887 598307
rect 675943 598195 717600 598363
rect 675887 597719 717600 598195
rect 675943 597551 717600 597719
rect 675887 597075 717600 597551
rect 675407 596963 675887 597019
rect 675943 596907 717600 597075
rect 675887 596523 717600 596907
rect 675943 596355 717600 596523
rect 675887 595879 717600 596355
rect 675943 595711 717600 595879
rect 675392 595614 675444 595678
rect 675404 595179 675432 595614
rect 675887 595235 717600 595711
rect 675404 595151 675887 595179
rect 675407 595123 675887 595151
rect 675943 595067 717600 595235
rect 675887 594683 717600 595067
rect 675407 594571 675887 594627
rect 675943 594515 717600 594683
rect 675887 594039 717600 594515
rect 675943 593871 717600 594039
rect 675312 593830 675432 593858
rect 675128 593694 675340 593722
rect 675312 574094 675340 593694
rect 675404 593339 675432 593830
rect 675887 593395 717600 593871
rect 675404 593300 675887 593339
rect 675407 593283 675887 593300
rect 675943 593227 717600 593395
rect 675887 593017 717600 593227
rect 675128 574066 675340 574094
rect 675128 546494 675156 574066
rect 675887 563559 717600 563758
rect 675407 563447 675887 563503
rect 675943 563391 717600 563559
rect 675887 563007 717600 563391
rect 675943 562839 717600 563007
rect 675887 562363 717600 562839
rect 675943 562195 717600 562363
rect 675887 561719 717600 562195
rect 675943 561551 717600 561719
rect 675887 561167 717600 561551
rect 675943 560999 717600 561167
rect 675887 560523 717600 560999
rect 675407 560439 675887 560467
rect 675404 560411 675887 560439
rect 675404 559978 675432 560411
rect 675943 560355 717600 560523
rect 675392 559914 675444 559978
rect 675887 559879 717600 560355
rect 675943 559711 717600 559879
rect 675887 559327 717600 559711
rect 675943 559159 717600 559327
rect 675887 558683 717600 559159
rect 675943 558515 717600 558683
rect 675887 558039 717600 558515
rect 675943 557871 717600 558039
rect 675392 557806 675444 557870
rect 675404 557431 675432 557806
rect 675887 557487 717600 557871
rect 675404 557396 675887 557431
rect 675407 557375 675887 557396
rect 675943 557319 717600 557487
rect 675887 556843 717600 557319
rect 675943 556675 717600 556843
rect 675887 556199 717600 556675
rect 675407 556115 675887 556143
rect 675404 556087 675887 556115
rect 675404 555626 675432 556087
rect 675943 556031 717600 556199
rect 675208 555562 675260 555626
rect 675392 555562 675444 555626
rect 675220 548125 675248 555562
rect 675887 555555 717600 556031
rect 675943 555387 717600 555555
rect 675887 555003 717600 555387
rect 675943 554835 717600 555003
rect 675887 554359 717600 554835
rect 675943 554191 717600 554359
rect 675887 553715 717600 554191
rect 675943 553547 717600 553715
rect 675887 553163 717600 553547
rect 675407 553051 675887 553107
rect 675943 552995 717600 553163
rect 675887 552519 717600 552995
rect 675943 552351 717600 552519
rect 675887 551875 717600 552351
rect 675407 551763 675887 551819
rect 675943 551707 717600 551875
rect 675887 551323 717600 551707
rect 675943 551155 717600 551323
rect 675887 550679 717600 551155
rect 675392 550462 675444 550526
rect 675943 550511 717600 550679
rect 675404 549979 675432 550462
rect 675887 550035 717600 550511
rect 675404 549951 675887 549979
rect 675407 549923 675887 549951
rect 675943 549867 717600 550035
rect 675887 549483 717600 549867
rect 675407 549371 675887 549427
rect 675943 549315 717600 549483
rect 675887 548839 717600 549315
rect 675943 548671 717600 548839
rect 675887 548195 717600 548671
rect 675407 548125 675887 548139
rect 675220 548097 675887 548125
rect 675407 548083 675887 548097
rect 675943 548027 717600 548195
rect 675887 547817 717600 548027
rect 675128 546466 675340 546494
rect 675312 513806 675340 546466
rect 678007 518701 716615 518747
rect 677600 513921 716615 518701
rect 675300 513742 675352 513806
rect 677692 513777 677744 513806
rect 677690 513703 677746 513777
rect 677600 513221 677984 513621
rect 678007 508722 716615 513921
rect 677600 503942 716615 508722
rect 685910 474800 686840 476995
rect 678007 474700 717593 474800
rect 678000 470701 717593 474700
rect 678007 470615 717593 470701
rect 678000 464093 717593 470615
rect 678007 463981 717593 464093
rect 678000 459860 717593 463981
rect 678007 459800 717593 459860
rect 682685 457613 685567 459560
rect 685917 457572 686847 459800
rect 687319 457613 717593 459560
rect 678007 430501 716615 430547
rect 674748 427790 674800 427854
rect 677508 427790 677560 427854
rect 677520 425649 677548 427790
rect 677600 425721 716615 430501
rect 677506 425575 677562 425649
rect 677600 425021 677984 425421
rect 678007 420522 716615 425721
rect 677600 415742 716615 420522
rect 675887 386359 717600 386558
rect 675407 386247 675887 386303
rect 675943 386191 717600 386359
rect 675887 385807 717600 386191
rect 675943 385639 717600 385807
rect 675887 385163 717600 385639
rect 675943 384995 717600 385163
rect 675887 384519 717600 384995
rect 675943 384351 717600 384519
rect 675887 383967 717600 384351
rect 675943 383799 717600 383967
rect 675392 383522 675444 383586
rect 675404 383267 675432 383522
rect 675887 383323 717600 383799
rect 675404 383239 675887 383267
rect 675407 383211 675887 383239
rect 675943 383155 717600 383323
rect 675887 382679 717600 383155
rect 675943 382511 717600 382679
rect 675887 382127 717600 382511
rect 675943 381959 717600 382127
rect 675887 381483 717600 381959
rect 675943 381315 717600 381483
rect 675887 380839 717600 381315
rect 675943 380671 717600 380839
rect 675887 380287 717600 380671
rect 675407 380188 675887 380231
rect 675404 380175 675887 380188
rect 675404 379710 675432 380175
rect 675943 380119 717600 380287
rect 675392 379646 675444 379710
rect 675887 379643 717600 380119
rect 675943 379475 717600 379643
rect 675887 378999 717600 379475
rect 675407 378929 675887 378943
rect 675312 378901 675887 378929
rect 673828 372302 673880 372366
rect 675312 370925 675340 378901
rect 675407 378887 675887 378901
rect 675943 378831 717600 378999
rect 675887 378355 717600 378831
rect 675943 378187 717600 378355
rect 675887 377803 717600 378187
rect 675943 377635 717600 377803
rect 675887 377159 717600 377635
rect 675943 376991 717600 377159
rect 675887 376515 717600 376991
rect 675943 376347 717600 376515
rect 675887 375963 717600 376347
rect 675407 375851 675887 375907
rect 675943 375795 717600 375963
rect 675887 375319 717600 375795
rect 675943 375151 717600 375319
rect 675887 374675 717600 375151
rect 675407 374563 675887 374619
rect 675943 374507 717600 374675
rect 675887 374123 717600 374507
rect 675407 374011 675887 374067
rect 675943 373955 717600 374123
rect 675887 373479 717600 373955
rect 675943 373311 717600 373479
rect 675887 372835 717600 373311
rect 675407 372751 675887 372779
rect 675404 372723 675887 372751
rect 675404 372366 675432 372723
rect 675943 372667 717600 372835
rect 675392 372302 675444 372366
rect 675887 372283 717600 372667
rect 675407 372171 675887 372227
rect 675943 372115 717600 372283
rect 675887 371639 717600 372115
rect 675943 371471 717600 371639
rect 675887 370995 717600 371471
rect 675407 370925 675887 370939
rect 675312 370897 675887 370925
rect 675407 370883 675887 370897
rect 675943 370827 717600 370995
rect 675887 370617 717600 370827
rect 675887 341159 717600 341358
rect 675407 341047 675887 341103
rect 675943 340991 717600 341159
rect 675887 340607 717600 340991
rect 675943 340439 717600 340607
rect 675887 339963 717600 340439
rect 675943 339795 717600 339963
rect 675887 339319 717600 339795
rect 675943 339151 717600 339319
rect 675887 338767 717600 339151
rect 675943 338599 717600 338767
rect 673736 334426 673788 334490
rect 673644 313210 673696 313274
rect 673472 295306 673592 295334
rect 673472 293214 673500 295306
rect 673460 293150 673512 293214
rect 42708 281318 42760 281382
rect 42616 271866 42668 271930
rect 42524 231678 42576 231742
rect 42536 227526 42564 231678
rect 42628 228682 42656 271866
rect 673472 248606 673500 293150
rect 673552 289478 673604 289542
rect 673564 264974 673592 289478
rect 673656 283082 673684 313210
rect 673748 289542 673776 334426
rect 675887 338123 717600 338599
rect 675407 338028 675887 338067
rect 675404 338011 675887 338028
rect 675404 337550 675432 338011
rect 675943 337955 717600 338123
rect 675392 337486 675444 337550
rect 675887 337479 717600 337955
rect 675943 337311 717600 337479
rect 675887 336927 717600 337311
rect 675943 336759 717600 336927
rect 675887 336283 717600 336759
rect 675943 336115 717600 336283
rect 675887 335639 717600 336115
rect 675943 335471 717600 335639
rect 675887 335087 717600 335471
rect 675407 335003 675887 335031
rect 675404 334975 675887 335003
rect 675404 334490 675432 334975
rect 675943 334919 717600 335087
rect 675392 334426 675444 334490
rect 675887 334443 717600 334919
rect 675943 334275 717600 334443
rect 675887 333799 717600 334275
rect 675407 333729 675887 333743
rect 675312 333701 675887 333729
rect 675312 325725 675340 333701
rect 675407 333687 675887 333701
rect 675943 333631 717600 333799
rect 675887 333155 717600 333631
rect 675943 332987 717600 333155
rect 675887 332603 717600 332987
rect 675943 332435 717600 332603
rect 675887 331959 717600 332435
rect 675943 331791 717600 331959
rect 675887 331315 717600 331791
rect 675943 331147 717600 331315
rect 675887 330763 717600 331147
rect 675407 330651 675887 330707
rect 675943 330595 717600 330763
rect 675887 330119 717600 330595
rect 675943 329951 717600 330119
rect 675887 329475 717600 329951
rect 675407 329363 675887 329419
rect 675943 329307 717600 329475
rect 675887 328923 717600 329307
rect 675407 328811 675887 328867
rect 675943 328755 717600 328923
rect 675887 328279 717600 328755
rect 675943 328111 717600 328279
rect 675392 328034 675444 328098
rect 675404 327579 675432 328034
rect 675887 327635 717600 328111
rect 675404 327556 675887 327579
rect 675407 327523 675887 327556
rect 675943 327467 717600 327635
rect 675887 327083 717600 327467
rect 675407 326971 675887 327027
rect 675943 326915 717600 327083
rect 675887 326439 717600 326915
rect 675943 326271 717600 326439
rect 675887 325795 717600 326271
rect 675407 325725 675887 325739
rect 675312 325697 675887 325725
rect 675407 325683 675887 325697
rect 675943 325627 717600 325795
rect 675887 325417 717600 325627
rect 675887 296159 717600 296358
rect 675407 296047 675887 296103
rect 675943 295991 717600 296159
rect 675887 295607 717600 295991
rect 675943 295439 717600 295607
rect 675887 294963 717600 295439
rect 675943 294795 717600 294963
rect 675887 294319 717600 294795
rect 675943 294151 717600 294319
rect 675887 293767 717600 294151
rect 673736 289478 673788 289542
rect 675943 293599 717600 293767
rect 675392 293150 675444 293214
rect 675404 293067 675432 293150
rect 675887 293123 717600 293599
rect 675404 293012 675887 293067
rect 675407 293011 675887 293012
rect 675943 292955 717600 293123
rect 675887 292479 717600 292955
rect 675943 292311 717600 292479
rect 675887 291927 717600 292311
rect 675943 291759 717600 291927
rect 675887 291283 717600 291759
rect 675943 291115 717600 291283
rect 675887 290639 717600 291115
rect 675943 290471 717600 290639
rect 675887 290087 717600 290471
rect 675407 290020 675887 290031
rect 675404 289975 675887 290020
rect 675404 289542 675432 289975
rect 675943 289919 717600 290087
rect 675392 289478 675444 289542
rect 675887 289443 717600 289919
rect 675943 289275 717600 289443
rect 675887 288799 717600 289275
rect 673644 283018 673696 283082
rect 673564 264946 673684 264974
rect 673460 248542 673512 248606
rect 673656 244934 673684 264946
rect 675407 288729 675887 288743
rect 675312 288701 675887 288729
rect 673920 283018 673972 283082
rect 673932 245654 673960 283018
rect 675312 280725 675340 288701
rect 675407 288687 675887 288701
rect 675943 288631 717600 288799
rect 675887 288155 717600 288631
rect 675943 287987 717600 288155
rect 675887 287603 717600 287987
rect 675943 287435 717600 287603
rect 675887 286959 717600 287435
rect 675943 286791 717600 286959
rect 675887 286315 717600 286791
rect 675943 286147 717600 286315
rect 675887 285763 717600 286147
rect 675407 285651 675887 285707
rect 675943 285595 717600 285763
rect 675887 285119 717600 285595
rect 675943 284951 717600 285119
rect 675887 284475 717600 284951
rect 675407 284363 675887 284419
rect 675943 284307 717600 284475
rect 675887 283923 717600 284307
rect 675407 283811 675887 283867
rect 675943 283755 717600 283923
rect 675887 283279 717600 283755
rect 675943 283111 717600 283279
rect 675392 283018 675444 283082
rect 675404 282579 675432 283018
rect 675887 282635 717600 283111
rect 675404 282540 675887 282579
rect 675407 282523 675887 282540
rect 675943 282467 717600 282635
rect 675887 282083 717600 282467
rect 675407 281971 675887 282027
rect 675943 281915 717600 282083
rect 675887 281439 717600 281915
rect 675943 281271 717600 281439
rect 675887 280795 717600 281271
rect 675407 280725 675887 280739
rect 675312 280697 675887 280725
rect 675407 280683 675887 280697
rect 675943 280627 717600 280795
rect 675887 280417 717600 280627
rect 675887 251159 717600 251358
rect 675407 251047 675887 251103
rect 675943 250991 717600 251159
rect 675887 250607 717600 250991
rect 675943 250439 717600 250607
rect 675887 249963 717600 250439
rect 675943 249795 717600 249963
rect 675887 249319 717600 249795
rect 675943 249151 717600 249319
rect 675887 248767 717600 249151
rect 674012 248542 674064 248606
rect 673840 245626 673960 245654
rect 673644 244870 673696 244934
rect 42616 228618 42668 228682
rect 42524 227462 42576 227526
rect 42628 207014 42656 228618
rect 42536 206986 42656 207014
rect 42432 197474 42484 197538
rect 42260 197390 42472 197418
rect 0 197205 41657 197373
rect 41713 197282 42193 197317
rect 41713 197261 42288 197282
rect 41722 197254 42288 197261
rect 0 196729 41713 197205
rect 0 196561 41657 196729
rect 0 196085 41713 196561
rect 0 195917 41657 196085
rect 41713 195973 42193 196029
rect 0 195533 41713 195917
rect 41788 195842 41840 195906
rect 0 195365 41657 195533
rect 41800 195477 41828 195842
rect 41713 195421 42193 195477
rect 0 194889 41713 195365
rect 0 194721 41657 194889
rect 0 194245 41713 194721
rect 0 194077 41657 194245
rect 41713 194133 42193 194189
rect 0 193693 41713 194077
rect 0 193525 41657 193693
rect 41713 193581 42193 193637
rect 0 193049 41713 193525
rect 0 192881 41657 193049
rect 0 192405 41713 192881
rect 0 192237 41657 192405
rect 41713 192293 42193 192349
rect 0 191853 41713 192237
rect 0 191685 41657 191853
rect 0 191209 41713 191685
rect 0 191041 41657 191209
rect 0 190565 41713 191041
rect 0 190397 41657 190565
rect 0 190013 41713 190397
rect 0 189845 41657 190013
rect 0 189369 41713 189845
rect 42260 189394 42288 197254
rect 0 189201 41657 189369
rect 41892 189366 42288 189394
rect 41892 189313 41920 189366
rect 41713 189257 42193 189313
rect 0 188725 41713 189201
rect 0 188557 41657 188725
rect 0 188081 41713 188557
rect 0 187913 41657 188081
rect 41722 188025 41828 188034
rect 41713 187969 42193 188025
rect 0 187529 41713 187913
rect 41800 187678 41828 187969
rect 41788 187614 41840 187678
rect 0 187361 41657 187529
rect 0 186885 41713 187361
rect 0 186717 41657 186885
rect 0 186241 41713 186717
rect 0 186073 41657 186241
rect 0 185689 41713 186073
rect 0 185521 41657 185689
rect 0 185045 41713 185521
rect 0 184877 41657 185045
rect 41713 184933 42193 184989
rect 0 184401 41713 184877
rect 41800 184482 41828 184933
rect 41788 184418 41840 184482
rect 0 184233 41657 184401
rect 42444 187678 42472 197390
rect 42432 187614 42484 187678
rect 0 183849 41713 184233
rect 42248 184146 42300 184210
rect 0 183681 41657 183849
rect 0 183205 41713 183681
rect 0 183037 41657 183205
rect 0 182561 41713 183037
rect 0 182393 41657 182561
rect 0 182009 41713 182393
rect 0 181841 41657 182009
rect 41713 181897 42193 181953
rect 0 181642 41713 181841
rect 985 120278 40000 125058
rect 985 115079 39593 120278
rect 39616 115379 40000 115779
rect 985 110299 40000 115079
rect 985 110253 39593 110299
rect 30753 83000 31683 85228
rect 31928 83049 32702 85239
rect 714 82940 39593 83000
rect 714 78819 39600 82940
rect 714 78707 39593 78819
rect 714 72185 39600 78707
rect 714 72099 39593 72185
rect 714 68100 39600 72099
rect 714 68098 39593 68100
rect 42260 45694 42288 184146
rect 42248 45630 42300 45694
rect 42444 121514 42472 187614
rect 42536 184482 42564 206986
rect 673552 202302 673604 202366
rect 42616 197474 42668 197538
rect 42628 195906 42656 197474
rect 42616 195842 42668 195906
rect 42524 184418 42576 184482
rect 42432 121450 42484 121514
rect 42628 80374 42656 195842
rect 673564 158370 673592 202302
rect 673656 199306 673684 244870
rect 673840 237726 673868 245626
rect 673828 237662 673880 237726
rect 673644 199242 673696 199306
rect 673552 158306 673604 158370
rect 673564 158250 673592 158306
rect 673472 158222 673592 158250
rect 44180 121450 44232 121514
rect 44192 110537 44220 121450
rect 673472 113218 673500 158222
rect 673656 155242 673684 199242
rect 673840 198734 673868 237662
rect 674024 202366 674052 248542
rect 675392 248542 675444 248606
rect 675943 248599 717600 248767
rect 675404 248067 675432 248542
rect 675887 248123 717600 248599
rect 675404 248039 675887 248067
rect 675407 248011 675887 248039
rect 675943 247955 717600 248123
rect 675887 247479 717600 247955
rect 675943 247311 717600 247479
rect 675887 246927 717600 247311
rect 675943 246759 717600 246927
rect 675887 246283 717600 246759
rect 675943 246115 717600 246283
rect 675887 245639 717600 246115
rect 675943 245471 717600 245639
rect 675887 245087 717600 245471
rect 675407 245004 675887 245031
rect 675404 244975 675887 245004
rect 675404 244934 675432 244975
rect 675392 244870 675444 244934
rect 675943 244919 717600 245087
rect 675887 244443 717600 244919
rect 675943 244275 717600 244443
rect 675887 243799 717600 244275
rect 675407 243729 675887 243743
rect 675312 243701 675887 243729
rect 675312 235725 675340 243701
rect 675407 243687 675887 243701
rect 675943 243631 717600 243799
rect 675887 243155 717600 243631
rect 675943 242987 717600 243155
rect 675887 242603 717600 242987
rect 675943 242435 717600 242603
rect 675887 241959 717600 242435
rect 675943 241791 717600 241959
rect 675887 241315 717600 241791
rect 675943 241147 717600 241315
rect 675887 240763 717600 241147
rect 675407 240651 675887 240707
rect 675943 240595 717600 240763
rect 675887 240119 717600 240595
rect 675943 239951 717600 240119
rect 675887 239475 717600 239951
rect 675407 239363 675887 239419
rect 675943 239307 717600 239475
rect 675887 238923 717600 239307
rect 675407 238811 675887 238867
rect 675943 238755 717600 238923
rect 675887 238279 717600 238755
rect 675943 238111 717600 238279
rect 675392 237662 675444 237726
rect 675404 237579 675432 237662
rect 675887 237635 717600 238111
rect 675404 237524 675887 237579
rect 675407 237523 675887 237524
rect 675943 237467 717600 237635
rect 675887 237083 717600 237467
rect 675407 236971 675887 237027
rect 675943 236915 717600 237083
rect 675887 236439 717600 236915
rect 675943 236271 717600 236439
rect 675887 235795 717600 236271
rect 675407 235725 675887 235739
rect 675312 235697 675887 235725
rect 675407 235683 675887 235697
rect 675943 235627 717600 235795
rect 675887 235417 717600 235627
rect 675887 205959 717600 206158
rect 675407 205847 675887 205903
rect 675943 205791 717600 205959
rect 675887 205407 717600 205791
rect 675943 205239 717600 205407
rect 675887 204763 717600 205239
rect 675943 204595 717600 204763
rect 675887 204119 717600 204595
rect 675943 203951 717600 204119
rect 675887 203567 717600 203951
rect 674012 202302 674064 202366
rect 675943 203399 717600 203567
rect 675887 202923 717600 203399
rect 675407 202844 675887 202867
rect 675404 202811 675887 202844
rect 675404 202366 675432 202811
rect 675943 202755 717600 202923
rect 675392 202302 675444 202366
rect 675887 202279 717600 202755
rect 675943 202111 717600 202279
rect 675887 201727 717600 202111
rect 675943 201559 717600 201727
rect 675887 201083 717600 201559
rect 675943 200915 717600 201083
rect 675887 200439 717600 200915
rect 675943 200271 717600 200439
rect 675887 199887 717600 200271
rect 675407 199803 675887 199831
rect 675404 199775 675887 199803
rect 675404 199306 675432 199775
rect 675943 199719 717600 199887
rect 675392 199242 675444 199306
rect 675887 199243 717600 199719
rect 675943 199075 717600 199243
rect 673840 198706 673960 198734
rect 673932 191962 673960 198706
rect 675312 198614 675432 198642
rect 673920 191898 673972 191962
rect 673644 155178 673696 155242
rect 673656 149054 673684 155178
rect 673564 149026 673684 149054
rect 673460 113154 673512 113218
rect 44178 110463 44234 110537
rect 44822 110463 44878 110537
rect 44836 110414 44864 110463
rect 44836 110386 44956 110414
rect 42616 80310 42668 80374
rect 44180 80310 44232 80374
rect 44192 71913 44220 80310
rect 44178 71839 44234 71913
rect 44822 71839 44878 71913
rect 44836 46986 44864 71839
rect 44824 46922 44876 46986
rect 44928 45558 44956 110386
rect 143540 46854 143592 46918
rect 140964 45630 141016 45694
rect 44916 45494 44968 45558
rect 93768 41482 93820 41546
rect 93780 40225 93808 41482
rect 135168 40225 135220 40254
rect 93766 40151 93822 40225
rect 135166 40151 135222 40225
rect 140976 40202 141004 45630
rect 143552 40497 143580 46854
rect 151726 46815 151782 46889
rect 188526 46815 188582 46889
rect 200856 46854 200908 46918
rect 143538 40423 143594 40497
rect 143540 40225 143592 40254
rect 140976 40174 141036 40202
rect 141008 40118 141036 40174
rect 143078 40151 143134 40225
rect 143538 40151 143594 40225
rect 146300 41822 146352 41886
rect 143084 40118 143112 40151
rect 140996 40054 141048 40118
rect 143072 40054 143124 40118
rect 144552 40054 144604 40118
rect 141008 40000 141036 40054
rect 143084 40000 143112 40054
rect 144564 40000 144592 40054
rect 146312 40118 146340 41822
rect 151740 40497 151768 46815
rect 186688 45630 186740 45694
rect 186700 42193 186728 45630
rect 188540 44402 188568 46815
rect 194692 45630 194744 45694
rect 188528 44338 188580 44402
rect 192852 44338 192904 44402
rect 188540 42193 188568 44338
rect 192864 42193 192892 44338
rect 194704 42193 194732 45630
rect 195980 45494 196032 45558
rect 195992 44334 196020 45494
rect 195980 44270 196032 44334
rect 195992 42193 196020 44270
rect 200868 42193 200896 46854
rect 204166 46815 204222 46889
rect 248420 46854 248472 46918
rect 201500 44338 201552 44402
rect 201512 44198 201540 44338
rect 204180 44198 204208 46815
rect 201500 44134 201552 44198
rect 204168 44134 204220 44198
rect 201512 42193 201540 44134
rect 186683 41713 186739 42193
rect 187971 41713 188027 42193
rect 188523 41713 188579 42193
rect 189167 41834 189223 42193
rect 189264 41890 189316 41954
rect 189276 41834 189304 41890
rect 189167 41806 189304 41834
rect 189167 41713 189223 41806
rect 189811 41713 189867 42193
rect 190363 41713 190419 42193
rect 191007 41834 191063 42193
rect 191104 41890 191156 41954
rect 191116 41834 191144 41890
rect 191007 41806 191144 41834
rect 191007 41713 191063 41806
rect 191651 41713 191707 42193
rect 192203 41834 192259 42193
rect 192300 41890 192352 41954
rect 192312 41834 192340 41890
rect 192203 41806 192340 41834
rect 192203 41713 192259 41806
rect 192847 41713 192903 42193
rect 193491 41834 193547 42193
rect 193588 41890 193640 41954
rect 193600 41834 193628 41890
rect 193491 41806 193628 41834
rect 193491 41713 193547 41806
rect 194687 41713 194743 42193
rect 195975 41713 196031 42193
rect 196440 41890 196492 41954
rect 196452 41834 196480 41890
rect 196527 41834 196583 42193
rect 197171 41834 197227 42193
rect 197815 41834 197871 42193
rect 198367 41834 198423 42193
rect 198464 41890 198516 41954
rect 198476 41834 198504 41890
rect 199011 41834 199067 42193
rect 196452 41806 198504 41834
rect 198936 41818 199067 41834
rect 198924 41806 199067 41818
rect 196527 41713 196583 41806
rect 197171 41713 197227 41806
rect 197815 41713 197871 41806
rect 198367 41713 198423 41806
rect 198924 41754 198976 41806
rect 199011 41713 199067 41806
rect 200120 41890 200172 41954
rect 200132 41834 200160 41890
rect 200207 41834 200263 42193
rect 200851 41834 200907 42193
rect 200132 41806 200907 41834
rect 200207 41713 200263 41806
rect 200851 41713 200907 41806
rect 201495 41713 201551 42193
rect 202047 41713 202103 42193
rect 186417 41657 186627 41713
rect 186795 41657 187271 41713
rect 187439 41657 187915 41713
rect 188083 41657 188467 41713
rect 188635 41657 189111 41713
rect 189279 41657 189755 41713
rect 189923 41657 190307 41713
rect 190475 41657 190951 41713
rect 191119 41657 191595 41713
rect 191763 41657 192147 41713
rect 192315 41657 192791 41713
rect 192959 41657 193435 41713
rect 193603 41657 193987 41713
rect 194155 41657 194631 41713
rect 194799 41657 195275 41713
rect 195443 41657 195919 41713
rect 196087 41657 196471 41713
rect 196639 41657 197115 41713
rect 197283 41657 197759 41713
rect 197927 41657 198311 41713
rect 198479 41657 198955 41713
rect 199123 41657 199599 41713
rect 199767 41657 200151 41713
rect 200319 41657 200795 41713
rect 200963 41657 201439 41713
rect 201607 41657 201991 41713
rect 202159 41657 202358 41713
rect 151726 40423 151782 40497
rect 146300 40054 146352 40118
rect 78942 39593 83722 40000
rect 88221 39616 88621 40000
rect 88921 39593 93701 40000
rect 132617 39816 140940 40000
rect 140996 39872 141048 40000
rect 141104 39878 141313 40000
rect 141369 39934 141499 40000
rect 141555 39878 141898 40000
rect 141954 39934 142084 40000
rect 142140 39878 143012 40000
rect 141104 39816 143012 39878
rect 78942 985 93747 39593
rect 132617 39204 143012 39816
rect 132617 39147 142955 39204
rect 143068 39151 143128 40000
rect 143184 39747 144517 40000
rect 144564 39916 144689 40000
rect 144573 39803 144689 39916
rect 144745 39747 145035 40000
rect 143184 39650 145035 39747
rect 145199 39650 147532 40000
rect 143184 39369 147532 39650
rect 143184 39297 144495 39369
rect 145520 39341 147532 39369
rect 143184 39243 144441 39297
rect 144551 39285 145464 39313
rect 144551 39271 145530 39285
rect 145586 39275 147532 39341
rect 144551 39261 145436 39271
rect 143184 39207 144367 39243
rect 144551 39241 144623 39261
rect 144625 39241 144645 39261
rect 145414 39247 145461 39261
rect 145464 39247 145530 39271
rect 143244 39169 144367 39207
rect 144497 39233 144551 39241
rect 144571 39233 144625 39241
rect 144497 39205 144625 39233
rect 145414 39219 145530 39247
rect 145414 39214 145461 39219
rect 144497 39187 144551 39205
rect 144571 39187 144625 39205
rect 143068 39148 143188 39151
rect 132617 39076 141720 39147
rect 143011 39091 143188 39148
rect 143244 39147 144345 39169
rect 144423 39113 144571 39187
rect 144701 39185 145358 39205
rect 144681 39158 145358 39185
rect 145461 39191 145525 39214
rect 145530 39191 145599 39219
rect 145655 39206 147532 39275
rect 145461 39163 145599 39191
rect 144681 39131 145405 39158
rect 145461 39150 145525 39163
rect 145530 39150 145599 39163
rect 144401 39091 144497 39113
rect 132617 39010 141654 39076
rect 141776 39063 144497 39091
rect 141776 39049 141847 39063
rect 143068 39049 143128 39063
rect 144423 39049 144497 39063
rect 144627 39094 145405 39131
rect 145525 39135 145591 39150
rect 145599 39135 145653 39150
rect 144627 39057 145469 39094
rect 145525 39085 145653 39135
rect 145525 39084 145591 39085
rect 141776 39039 144497 39049
rect 141776 39020 141847 39039
rect 141850 39020 141869 39039
rect 144553 39028 145469 39057
rect 141710 39011 141776 39020
rect 141784 39011 141850 39020
rect 132617 37861 141628 39010
rect 141710 38969 141850 39011
rect 144553 38983 145545 39028
rect 141710 38954 141776 38969
rect 141784 38954 141850 38969
rect 141925 38964 145545 38983
rect 141684 38928 141710 38954
rect 141736 38928 141784 38954
rect 141684 38906 141784 38928
rect 132617 37823 141590 37861
rect 132617 36927 141538 37823
rect 141684 37805 141736 38906
rect 141906 38898 145545 38964
rect 141840 38850 145545 38898
rect 141646 37783 141736 37805
rect 141646 37767 141684 37783
rect 141720 37767 141736 37783
rect 141792 38284 145545 38850
rect 141792 38216 145477 38284
rect 145601 38228 145653 39085
rect 141792 38176 145437 38216
rect 145533 38178 145653 38228
rect 141792 38110 145371 38176
rect 145533 38160 145601 38178
rect 145607 38160 145653 38178
rect 145493 38150 145533 38160
rect 145567 38150 145607 38160
rect 145493 38136 145607 38150
rect 145493 38120 145533 38136
rect 145567 38120 145607 38136
rect 141594 37693 141720 37767
rect 141792 37711 145319 38110
rect 145427 38108 145493 38120
rect 145501 38108 145567 38120
rect 145427 38080 145567 38108
rect 145709 38104 147532 39206
rect 145427 38054 145493 38080
rect 145501 38054 145567 38080
rect 145663 38064 147532 38104
rect 132617 36860 141471 36927
rect 141594 36871 141646 37693
rect 141776 37637 145319 37711
rect 132617 35845 141419 36860
rect 141527 36821 141646 36871
rect 141527 36804 141594 36821
rect 141601 36804 141646 36821
rect 141475 36730 141601 36804
rect 141702 36748 145319 37637
rect 141475 35901 141527 36730
rect 141657 36674 145319 36748
rect 141583 35845 145319 36674
rect 132617 34484 145319 35845
rect 145375 37980 145501 38054
rect 145623 37998 147532 38064
rect 145375 34678 145427 37980
rect 145557 37924 147532 37998
rect 145483 34734 147532 37924
rect 145375 34540 145470 34678
rect 132617 34469 145362 34484
rect 132617 33839 145319 34469
rect 145418 34413 145470 34540
rect 145375 34371 145470 34413
rect 145375 34370 145418 34371
rect 145375 34275 145470 34370
rect 132617 33810 145290 33839
rect 132617 33765 145245 33810
rect 145375 33783 145427 34275
rect 145526 34219 147532 34734
rect 132617 32852 145240 33765
rect 145346 33754 145427 33783
rect 145301 33747 145346 33754
rect 145375 33747 145427 33754
rect 145301 33733 145427 33747
rect 145301 33709 145346 33733
rect 145375 33709 145427 33733
rect 145296 33704 145301 33709
rect 145348 33704 145375 33709
rect 145296 33682 145375 33704
rect 132617 32688 145114 32852
rect 145296 32796 145348 33682
rect 145483 33653 147532 34219
rect 145431 33626 147532 33653
rect 145170 32744 145348 32796
rect 145404 32688 147532 33626
rect 132617 158 147532 32688
rect 186417 0 202358 41657
rect 248432 39953 248460 46854
rect 297086 46815 297142 46889
rect 297732 46854 297784 46918
rect 309416 46854 309468 46918
rect 352564 46854 352616 46918
rect 364248 46854 364300 46918
rect 407396 46854 407448 46918
rect 419080 46854 419132 46918
rect 462136 46854 462188 46918
rect 473820 46854 473872 46918
rect 516968 46854 517020 46918
rect 295248 44202 295300 44266
rect 295260 42193 295288 44202
rect 297100 42193 297128 46815
rect 297744 42294 297772 46854
rect 305736 44270 305788 44334
rect 303252 44202 303304 44266
rect 297732 42230 297784 42294
rect 300768 42230 300820 42294
rect 297744 42193 297772 42230
rect 300780 42193 300808 42230
rect 303264 42193 303292 44202
rect 304540 44134 304592 44198
rect 304552 42193 304580 44134
rect 305748 42193 305776 44270
rect 309428 42193 309456 46854
rect 349988 44406 350040 44470
rect 350000 44198 350028 44406
rect 351920 44270 351972 44334
rect 349988 44134 350040 44198
rect 350080 44134 350132 44198
rect 350092 42193 350120 44134
rect 351932 42193 351960 44270
rect 352576 42193 352604 46854
rect 359372 44406 359424 44470
rect 358084 44134 358136 44198
rect 358096 42193 358124 44134
rect 359384 42193 359412 44406
rect 360476 44338 360528 44402
rect 295260 41806 295339 42193
rect 295283 41713 295339 41806
rect 295927 41713 295983 42193
rect 296571 41713 296627 42193
rect 297100 41834 297179 42193
rect 297272 41890 297324 41954
rect 297284 41834 297312 41890
rect 297100 41806 297312 41834
rect 297744 41806 297823 42193
rect 297123 41713 297179 41806
rect 297767 41713 297823 41806
rect 298411 41713 298467 42193
rect 298963 41713 299019 42193
rect 299480 41890 299532 41954
rect 299492 41834 299520 41890
rect 299607 41834 299663 42193
rect 299492 41806 299663 41834
rect 299607 41713 299663 41806
rect 300251 41713 300307 42193
rect 300780 41834 300859 42193
rect 301447 41834 301503 42193
rect 302091 41834 302147 42193
rect 302240 41890 302292 41954
rect 302252 41834 302280 41890
rect 300780 41806 302280 41834
rect 300803 41713 300859 41806
rect 301447 41713 301503 41806
rect 302091 41713 302147 41806
rect 303264 41806 303343 42193
rect 304552 41806 304631 42193
rect 303287 41713 303343 41806
rect 304575 41713 304631 41806
rect 305127 41834 305183 42193
rect 305644 41970 305696 42022
rect 305748 41970 305827 42193
rect 305644 41958 305827 41970
rect 305276 41890 305328 41954
rect 305656 41942 305827 41958
rect 305288 41834 305316 41890
rect 305127 41806 305316 41834
rect 305748 41806 305827 41942
rect 305127 41713 305183 41806
rect 305771 41713 305827 41806
rect 306415 41834 306471 42193
rect 306564 41890 306616 41954
rect 306576 41834 306604 41890
rect 306415 41806 306604 41834
rect 306415 41713 306471 41806
rect 307611 41834 307667 42193
rect 307611 41818 307800 41834
rect 307611 41806 307812 41818
rect 308680 41890 308732 41954
rect 308692 41834 308720 41890
rect 308807 41834 308863 42193
rect 309428 41834 309507 42193
rect 308692 41806 309507 41834
rect 307611 41713 307667 41806
rect 307760 41754 307812 41806
rect 308807 41713 308863 41806
rect 309451 41713 309507 41806
rect 310647 41713 310703 42193
rect 350083 41713 350139 42193
rect 350727 41713 350783 42193
rect 351371 41713 351427 42193
rect 351923 41970 351979 42193
rect 352567 41970 352623 42193
rect 352656 41970 352708 42022
rect 351923 41954 352052 41970
rect 352567 41958 352708 41970
rect 351923 41942 352064 41954
rect 351923 41713 351979 41942
rect 352012 41890 352064 41942
rect 352567 41942 352696 41958
rect 352567 41713 352623 41942
rect 353211 41713 353267 42193
rect 353763 41713 353819 42193
rect 354312 41890 354364 41954
rect 354324 41834 354352 41890
rect 354407 41834 354463 42193
rect 354324 41806 354463 41834
rect 354407 41713 354463 41806
rect 355051 41713 355107 42193
rect 355508 41958 355560 42022
rect 355520 41834 355548 41958
rect 355603 41834 355659 42193
rect 356247 41834 356303 42193
rect 356891 41834 356947 42193
rect 356980 41958 357032 42022
rect 356992 41834 357020 41958
rect 355520 41806 357020 41834
rect 355603 41713 355659 41806
rect 356247 41713 356303 41806
rect 356891 41713 356947 41806
rect 358087 41713 358143 42193
rect 359375 41713 359431 42193
rect 359832 41958 359884 42022
rect 359844 41834 359872 41958
rect 359927 41834 359983 42193
rect 360488 41954 360516 44338
rect 364260 42193 364288 46854
rect 406752 44338 406804 44402
rect 404910 44231 404966 44305
rect 406764 44266 406792 44338
rect 404924 42193 404952 44231
rect 406752 44202 406804 44266
rect 406764 42193 406792 44202
rect 407408 42193 407436 46854
rect 414204 44406 414256 44470
rect 412914 44231 412970 44305
rect 412928 42193 412956 44231
rect 414216 44198 414244 44406
rect 414204 44134 414256 44198
rect 414216 42193 414244 44134
rect 419092 42193 419120 46854
rect 459650 44231 459706 44305
rect 459664 42193 459692 44231
rect 461492 44202 461544 44266
rect 461504 42193 461532 44202
rect 462148 42193 462176 46854
rect 468944 44338 468996 44402
rect 467654 44231 467710 44305
rect 467668 42193 467696 44231
rect 468956 44198 468984 44338
rect 468944 44134 468996 44198
rect 468956 42193 468984 44134
rect 473832 42193 473860 46854
rect 514482 44231 514538 44305
rect 514496 42193 514524 44231
rect 516324 44202 516376 44266
rect 516336 42193 516364 44202
rect 516980 42193 517008 46854
rect 523776 45562 523828 45626
rect 518716 45494 518768 45558
rect 518728 44266 518756 45494
rect 522486 44367 522542 44441
rect 523788 44402 523816 45562
rect 518716 44202 518768 44266
rect 522500 42193 522528 44367
rect 523776 44338 523828 44402
rect 523788 42193 523816 44338
rect 673472 42770 673500 113154
rect 673564 109546 673592 149026
rect 673932 149054 673960 191898
rect 675312 190525 675340 198614
rect 675404 198543 675432 198614
rect 675887 198599 717600 199075
rect 675404 198492 675887 198543
rect 675407 198487 675887 198492
rect 675943 198431 717600 198599
rect 675887 197955 717600 198431
rect 675943 197787 717600 197955
rect 675887 197403 717600 197787
rect 675943 197235 717600 197403
rect 675887 196759 717600 197235
rect 675943 196591 717600 196759
rect 675887 196115 717600 196591
rect 675943 195947 717600 196115
rect 675887 195563 717600 195947
rect 675407 195451 675887 195507
rect 675943 195395 717600 195563
rect 675887 194919 717600 195395
rect 675943 194751 717600 194919
rect 675887 194275 717600 194751
rect 675407 194163 675887 194219
rect 675943 194107 717600 194275
rect 675887 193723 717600 194107
rect 675407 193611 675887 193667
rect 675943 193555 717600 193723
rect 675887 193079 717600 193555
rect 675943 192911 717600 193079
rect 675887 192435 717600 192911
rect 675407 192372 675887 192379
rect 675404 192323 675887 192372
rect 675404 191962 675432 192323
rect 675943 192267 717600 192435
rect 675392 191898 675444 191962
rect 675887 191883 717600 192267
rect 675407 191771 675887 191827
rect 675943 191715 717600 191883
rect 675887 191239 717600 191715
rect 675943 191071 717600 191239
rect 675887 190595 717600 191071
rect 675407 190525 675887 190539
rect 675312 190497 675887 190525
rect 675407 190483 675887 190497
rect 675943 190427 717600 190595
rect 675887 190217 717600 190427
rect 675887 160959 717600 161158
rect 675407 160847 675887 160903
rect 675943 160791 717600 160959
rect 675887 160407 717600 160791
rect 675943 160239 717600 160407
rect 675887 159763 717600 160239
rect 675943 159595 717600 159763
rect 675887 159119 717600 159595
rect 675943 158951 717600 159119
rect 675887 158567 717600 158951
rect 675943 158399 717600 158567
rect 675392 158306 675444 158370
rect 675404 157867 675432 158306
rect 675887 157923 717600 158399
rect 675404 157828 675887 157867
rect 675407 157811 675887 157828
rect 675943 157755 717600 157923
rect 675887 157279 717600 157755
rect 675943 157111 717600 157279
rect 675887 156727 717600 157111
rect 675943 156559 717600 156727
rect 675887 156083 717600 156559
rect 675943 155915 717600 156083
rect 675887 155439 717600 155915
rect 675943 155271 717600 155439
rect 675392 155178 675444 155242
rect 675404 154831 675432 155178
rect 675887 154887 717600 155271
rect 675404 154803 675887 154831
rect 675407 154775 675887 154803
rect 675943 154719 717600 154887
rect 675887 154243 717600 154719
rect 675943 154075 717600 154243
rect 675887 153599 717600 154075
rect 675407 153529 675887 153543
rect 673840 149026 673960 149054
rect 675312 153501 675887 153529
rect 673840 146946 673868 149026
rect 673828 146882 673880 146946
rect 673840 129734 673868 146882
rect 675312 145525 675340 153501
rect 675407 153487 675887 153501
rect 675943 153431 717600 153599
rect 675887 152955 717600 153431
rect 675943 152787 717600 152955
rect 675887 152403 717600 152787
rect 675943 152235 717600 152403
rect 675887 151759 717600 152235
rect 675943 151591 717600 151759
rect 675887 151115 717600 151591
rect 675943 150947 717600 151115
rect 675887 150563 717600 150947
rect 675407 150451 675887 150507
rect 675943 150395 717600 150563
rect 675887 149919 717600 150395
rect 675943 149751 717600 149919
rect 675887 149275 717600 149751
rect 675407 149163 675887 149219
rect 675943 149107 717600 149275
rect 675887 148723 717600 149107
rect 675407 148611 675887 148667
rect 675943 148555 717600 148723
rect 675887 148079 717600 148555
rect 675943 147911 717600 148079
rect 675887 147435 717600 147911
rect 675407 147356 675887 147379
rect 675404 147323 675887 147356
rect 675404 146946 675432 147323
rect 675943 147267 717600 147435
rect 675392 146882 675444 146946
rect 675887 146883 717600 147267
rect 675407 146771 675887 146827
rect 675943 146715 717600 146883
rect 675887 146239 717600 146715
rect 675943 146071 717600 146239
rect 675887 145595 717600 146071
rect 675407 145525 675887 145539
rect 675312 145497 675887 145525
rect 675407 145483 675887 145497
rect 675943 145427 717600 145595
rect 675887 145217 717600 145427
rect 673748 129706 673868 129734
rect 673552 109482 673604 109546
rect 673564 45626 673592 109482
rect 673748 101726 673776 129706
rect 675887 115759 717600 115958
rect 675407 115647 675887 115703
rect 675943 115591 717600 115759
rect 675887 115207 717600 115591
rect 675943 115039 717600 115207
rect 675887 114563 717600 115039
rect 675943 114395 717600 114563
rect 675887 113919 717600 114395
rect 675943 113751 717600 113919
rect 675887 113367 717600 113751
rect 675392 113154 675444 113218
rect 675943 113199 717600 113367
rect 675404 112667 675432 113154
rect 675887 112723 717600 113199
rect 675404 112639 675887 112667
rect 675407 112611 675887 112639
rect 675943 112555 717600 112723
rect 675887 112079 717600 112555
rect 675943 111911 717600 112079
rect 675887 111527 717600 111911
rect 675943 111359 717600 111527
rect 675887 110883 717600 111359
rect 675943 110715 717600 110883
rect 675887 110239 717600 110715
rect 675943 110071 717600 110239
rect 675887 109687 717600 110071
rect 675407 109603 675887 109631
rect 675404 109575 675887 109603
rect 675404 109546 675432 109575
rect 675392 109482 675444 109546
rect 675943 109519 717600 109687
rect 675887 109043 717600 109519
rect 675943 108875 717600 109043
rect 675887 108399 717600 108875
rect 675407 108338 675887 108343
rect 675312 108310 675887 108338
rect 673736 101662 673788 101726
rect 673552 45562 673604 45626
rect 673748 45558 673776 101662
rect 675312 100314 675340 108310
rect 675407 108287 675887 108310
rect 675943 108231 717600 108399
rect 675887 107755 717600 108231
rect 675943 107587 717600 107755
rect 675887 107203 717600 107587
rect 675943 107035 717600 107203
rect 675887 106559 717600 107035
rect 675943 106391 717600 106559
rect 675887 105915 717600 106391
rect 675943 105747 717600 105915
rect 675887 105363 717600 105747
rect 675407 105251 675887 105307
rect 675943 105195 717600 105363
rect 675887 104719 717600 105195
rect 675943 104551 717600 104719
rect 675887 104075 717600 104551
rect 675407 103963 675887 104019
rect 675943 103907 717600 104075
rect 675887 103523 717600 103907
rect 675407 103411 675887 103467
rect 675943 103355 717600 103523
rect 675887 102879 717600 103355
rect 675943 102711 717600 102879
rect 675887 102235 717600 102711
rect 675407 102151 675887 102179
rect 675404 102123 675887 102151
rect 675404 101726 675432 102123
rect 675943 102067 717600 102235
rect 675392 101662 675444 101726
rect 675887 101683 717600 102067
rect 675407 101571 675887 101627
rect 675943 101515 717600 101683
rect 675887 101039 717600 101515
rect 675943 100871 717600 101039
rect 675887 100395 717600 100871
rect 675407 100314 675887 100339
rect 675312 100286 675887 100314
rect 675407 100283 675887 100286
rect 675943 100227 717600 100395
rect 675887 100017 717600 100227
rect 673736 45494 673788 45558
rect 576768 42706 576820 42770
rect 673460 42706 673512 42770
rect 360476 41890 360528 41954
rect 359844 41806 359983 41834
rect 360488 41834 360516 41890
rect 360571 41834 360627 42193
rect 361120 41958 361172 42022
rect 360488 41806 360627 41834
rect 361132 41834 361160 41958
rect 361215 41834 361271 42193
rect 361132 41806 361271 41834
rect 359927 41713 359983 41806
rect 360571 41713 360627 41806
rect 361215 41713 361271 41806
rect 362411 41834 362467 42193
rect 362411 41818 362540 41834
rect 362411 41806 362552 41818
rect 362411 41713 362467 41806
rect 362500 41754 362552 41806
rect 363512 41890 363564 41954
rect 363524 41834 363552 41890
rect 363607 41834 363663 42193
rect 364251 41834 364307 42193
rect 363524 41806 364307 41834
rect 363607 41713 363663 41806
rect 364251 41713 364307 41806
rect 365447 41713 365503 42193
rect 404883 41820 404952 42193
rect 404883 41713 404939 41820
rect 406171 41713 406227 42193
rect 406723 41820 406792 42193
rect 407367 41970 407436 42193
rect 407367 41954 407528 41970
rect 407367 41942 407540 41954
rect 407367 41820 407436 41942
rect 407488 41890 407540 41942
rect 406723 41713 406779 41820
rect 407367 41713 407423 41820
rect 408011 41713 408067 42193
rect 408563 41713 408619 42193
rect 409851 41713 409907 42193
rect 410248 41890 410300 41954
rect 410260 41834 410288 41890
rect 410403 41834 410459 42193
rect 410260 41806 410459 41834
rect 410403 41713 410459 41806
rect 411536 41890 411588 41954
rect 411548 41834 411576 41890
rect 411691 41834 411747 42193
rect 411548 41806 411747 41834
rect 411691 41713 411747 41806
rect 412887 41820 412956 42193
rect 414175 41820 414244 42193
rect 414572 41890 414624 41954
rect 414584 41834 414612 41890
rect 414727 41834 414783 42193
rect 415860 41890 415912 41954
rect 412887 41713 412943 41820
rect 414175 41713 414231 41820
rect 414584 41806 414783 41834
rect 414727 41713 414783 41806
rect 415872 41834 415900 41890
rect 416015 41834 416071 42193
rect 415872 41806 416071 41834
rect 416015 41713 416071 41806
rect 417211 41834 417267 42193
rect 417211 41818 417372 41834
rect 418252 41890 418304 41954
rect 418264 41834 418292 41890
rect 418407 41834 418463 42193
rect 419051 41834 419120 42193
rect 418264 41820 419120 41834
rect 417211 41806 417384 41818
rect 417211 41713 417267 41806
rect 417332 41754 417384 41806
rect 418264 41806 419107 41820
rect 418407 41713 418463 41806
rect 419051 41713 419107 41806
rect 420247 41713 420303 42193
rect 459664 41806 459739 42193
rect 459683 41713 459739 41806
rect 460971 41713 461027 42193
rect 461504 41806 461579 42193
rect 462148 41834 462223 42193
rect 462320 41890 462372 41954
rect 462332 41834 462360 41890
rect 462148 41806 462360 41834
rect 461523 41713 461579 41806
rect 462167 41713 462223 41806
rect 462811 41713 462867 42193
rect 463363 41713 463419 42193
rect 464651 41713 464707 42193
rect 465080 41890 465132 41954
rect 465092 41834 465120 41890
rect 465203 41834 465259 42193
rect 465092 41806 465259 41834
rect 466368 41890 466420 41954
rect 466380 41834 466408 41890
rect 466491 41834 466547 42193
rect 466380 41806 466547 41834
rect 465203 41713 465259 41806
rect 466491 41713 466547 41806
rect 467668 41806 467743 42193
rect 468956 41806 469031 42193
rect 469404 41890 469456 41954
rect 469416 41834 469444 41890
rect 469527 41834 469583 42193
rect 470692 41890 470744 41954
rect 469416 41806 469583 41834
rect 467687 41713 467743 41806
rect 468975 41713 469031 41806
rect 469527 41713 469583 41806
rect 470704 41834 470732 41890
rect 470815 41834 470871 42193
rect 470704 41806 470871 41834
rect 470815 41713 470871 41806
rect 472011 41834 472067 42193
rect 472011 41818 472204 41834
rect 472011 41806 472216 41818
rect 473084 41890 473136 41954
rect 473096 41834 473124 41890
rect 473207 41834 473263 42193
rect 473832 41834 473907 42193
rect 473096 41806 473907 41834
rect 472011 41713 472067 41806
rect 472164 41754 472216 41806
rect 473207 41713 473263 41806
rect 473851 41713 473907 41806
rect 475047 41713 475103 42193
rect 514483 41713 514539 42193
rect 515771 41713 515827 42193
rect 516323 41713 516379 42193
rect 516967 41970 517023 42193
rect 516967 41954 517100 41970
rect 516967 41942 517112 41954
rect 516967 41713 517023 41942
rect 517060 41890 517112 41942
rect 517611 41713 517667 42193
rect 518163 41713 518219 42193
rect 519451 41713 519507 42193
rect 519912 41890 519964 41954
rect 519924 41834 519952 41890
rect 520003 41834 520059 42193
rect 519924 41806 520059 41834
rect 520003 41713 520059 41806
rect 521200 41890 521252 41954
rect 521212 41834 521240 41890
rect 521291 41834 521347 42193
rect 521212 41806 521347 41834
rect 521291 41713 521347 41806
rect 522487 41713 522543 42193
rect 523775 41713 523831 42193
rect 524236 41890 524288 41954
rect 524248 41834 524276 41890
rect 524327 41834 524383 42193
rect 524248 41806 524383 41834
rect 524327 41713 524383 41806
rect 525524 41890 525576 41954
rect 525536 41834 525564 41890
rect 525615 41834 525671 42193
rect 525536 41806 525671 41834
rect 525615 41713 525671 41806
rect 526811 41834 526867 42193
rect 526732 41818 526867 41834
rect 526720 41806 526867 41818
rect 526720 41754 526772 41806
rect 526811 41713 526867 41806
rect 527916 41890 527968 41954
rect 527928 41834 527956 41890
rect 528007 41834 528063 42193
rect 528651 41834 528707 42193
rect 527928 41806 528707 41834
rect 528007 41713 528063 41806
rect 528651 41713 528707 41806
rect 529847 41713 529903 42193
rect 576780 41886 576808 42706
rect 569132 41822 569184 41886
rect 576768 41822 576820 41886
rect 295017 41657 295227 41713
rect 295395 41657 295871 41713
rect 296039 41657 296515 41713
rect 296683 41657 297067 41713
rect 297235 41657 297711 41713
rect 297879 41657 298355 41713
rect 298523 41657 298907 41713
rect 299075 41657 299551 41713
rect 299719 41657 300195 41713
rect 300363 41657 300747 41713
rect 300915 41657 301391 41713
rect 301559 41657 302035 41713
rect 302203 41657 302587 41713
rect 302755 41657 303231 41713
rect 303399 41657 303875 41713
rect 304043 41657 304519 41713
rect 304687 41657 305071 41713
rect 305239 41657 305715 41713
rect 305883 41657 306359 41713
rect 306527 41657 306911 41713
rect 307079 41657 307555 41713
rect 307723 41657 308199 41713
rect 308367 41657 308751 41713
rect 308919 41657 309395 41713
rect 309563 41657 310039 41713
rect 310207 41657 310591 41713
rect 310759 41657 310958 41713
rect 248418 39879 248474 39953
rect 241260 39593 245381 39600
rect 245493 39593 252015 39600
rect 252101 39593 256100 39600
rect 238961 31928 241151 32702
rect 241200 31683 256100 39593
rect 238972 30753 256100 31683
rect 241200 714 256100 30753
rect 295017 0 310958 41657
rect 349817 41657 350027 41713
rect 350195 41657 350671 41713
rect 350839 41657 351315 41713
rect 351483 41657 351867 41713
rect 352035 41657 352511 41713
rect 352679 41657 353155 41713
rect 353323 41657 353707 41713
rect 353875 41657 354351 41713
rect 354519 41657 354995 41713
rect 355163 41657 355547 41713
rect 355715 41657 356191 41713
rect 356359 41657 356835 41713
rect 357003 41657 357387 41713
rect 357555 41657 358031 41713
rect 358199 41657 358675 41713
rect 358843 41657 359319 41713
rect 359487 41657 359871 41713
rect 360039 41657 360515 41713
rect 360683 41657 361159 41713
rect 361327 41657 361711 41713
rect 361879 41657 362355 41713
rect 362523 41657 362999 41713
rect 363167 41657 363551 41713
rect 363719 41657 364195 41713
rect 364363 41657 364839 41713
rect 365007 41657 365391 41713
rect 365559 41657 365758 41713
rect 349817 0 365758 41657
rect 404617 41657 404827 41713
rect 404995 41657 405471 41713
rect 405639 41657 406115 41713
rect 406283 41657 406667 41713
rect 406835 41657 407311 41713
rect 407479 41657 407955 41713
rect 408123 41657 408507 41713
rect 408675 41657 409151 41713
rect 409319 41657 409795 41713
rect 409963 41657 410347 41713
rect 410515 41657 410991 41713
rect 411159 41657 411635 41713
rect 411803 41657 412187 41713
rect 412355 41657 412831 41713
rect 412999 41657 413475 41713
rect 413643 41657 414119 41713
rect 414287 41657 414671 41713
rect 414839 41657 415315 41713
rect 415483 41657 415959 41713
rect 416127 41657 416511 41713
rect 416679 41657 417155 41713
rect 417323 41657 417799 41713
rect 417967 41657 418351 41713
rect 418519 41657 418995 41713
rect 419163 41657 419639 41713
rect 419807 41657 420191 41713
rect 420359 41657 420558 41713
rect 404617 0 420558 41657
rect 459417 41657 459627 41713
rect 459795 41657 460271 41713
rect 460439 41657 460915 41713
rect 461083 41657 461467 41713
rect 461635 41657 462111 41713
rect 462279 41657 462755 41713
rect 462923 41657 463307 41713
rect 463475 41657 463951 41713
rect 464119 41657 464595 41713
rect 464763 41657 465147 41713
rect 465315 41657 465791 41713
rect 465959 41657 466435 41713
rect 466603 41657 466987 41713
rect 467155 41657 467631 41713
rect 467799 41657 468275 41713
rect 468443 41657 468919 41713
rect 469087 41657 469471 41713
rect 469639 41657 470115 41713
rect 470283 41657 470759 41713
rect 470927 41657 471311 41713
rect 471479 41657 471955 41713
rect 472123 41657 472599 41713
rect 472767 41657 473151 41713
rect 473319 41657 473795 41713
rect 473963 41657 474439 41713
rect 474607 41657 474991 41713
rect 475159 41657 475358 41713
rect 459417 0 475358 41657
rect 514217 41657 514427 41713
rect 514595 41657 515071 41713
rect 515239 41657 515715 41713
rect 515883 41657 516267 41713
rect 516435 41657 516911 41713
rect 517079 41657 517555 41713
rect 517723 41657 518107 41713
rect 518275 41657 518751 41713
rect 518919 41657 519395 41713
rect 519563 41657 519947 41713
rect 520115 41657 520591 41713
rect 520759 41657 521235 41713
rect 521403 41657 521787 41713
rect 521955 41657 522431 41713
rect 522599 41657 523075 41713
rect 523243 41657 523719 41713
rect 523887 41657 524271 41713
rect 524439 41657 524915 41713
rect 525083 41657 525559 41713
rect 525727 41657 526111 41713
rect 526279 41657 526755 41713
rect 526923 41657 527399 41713
rect 527567 41657 527951 41713
rect 528119 41657 528595 41713
rect 528763 41657 529239 41713
rect 529407 41657 529791 41713
rect 529959 41657 530158 41713
rect 514217 0 530158 41657
rect 569144 40225 569172 41822
rect 569130 40151 569186 40225
rect 569142 39593 573922 40000
rect 578421 39616 578821 40000
rect 579121 39593 583901 40000
rect 622942 39593 627722 40000
rect 632221 39616 632621 40000
rect 632921 39593 637701 40000
rect 569142 985 583947 39593
rect 622942 985 637747 39593
<< metal3 >>
rect 678000 469900 685920 474700
rect 31680 440900 39600 445700
rect 411069 44434 411135 44437
rect 465809 44434 465875 44437
rect 474457 44434 474523 44437
rect 411069 44432 419550 44434
rect 411069 44376 411074 44432
rect 411130 44376 419550 44432
rect 411069 44374 419550 44376
rect 411069 44371 411135 44374
rect 419490 44298 419550 44374
rect 465809 44432 474523 44434
rect 465809 44376 465814 44432
rect 465870 44376 474462 44432
rect 474518 44376 474523 44432
rect 465809 44374 474523 44376
rect 465809 44371 465875 44374
rect 474457 44371 474523 44374
rect 419717 44298 419783 44301
rect 419490 44296 419783 44298
rect 419490 44240 419722 44296
rect 419778 44240 419783 44296
rect 419490 44238 419783 44240
rect 419717 44235 419783 44238
rect 518801 44298 518867 44301
rect 524965 44298 525031 44301
rect 518801 44296 525031 44298
rect 518801 44240 518806 44296
rect 518862 44240 524970 44296
rect 525026 44240 525031 44296
rect 518801 44238 525031 44240
rect 518801 44235 518867 44238
rect 524965 44235 525031 44238
rect 141667 38031 141813 40000
rect 141667 37971 141873 38031
rect 141667 37911 141820 37971
rect 141873 37911 141966 37971
rect 141667 37818 141966 37911
rect 141820 37046 141966 37818
<< obsm3 >>
rect 76262 997338 92114 1037600
rect 127662 997338 143514 1037600
rect 179062 997338 194914 1037600
rect 230462 997338 246314 1037600
rect 282062 997338 297914 1037600
rect 333448 1002850 348258 1037600
rect 333499 997600 338279 1002770
rect 338359 998007 343398 1002850
rect 338579 997600 340779 998007
rect 340978 997600 343178 998007
rect 343478 997600 348258 1002770
rect 342161 997522 342227 997525
rect 343590 997522 343650 997600
rect 342161 997462 343650 997522
rect 342161 997459 342227 997462
rect 383862 997338 399714 1037600
rect 472862 997338 488714 1037600
rect 524262 997338 540114 1037600
rect 575648 1005032 590458 1036620
rect 575648 1004183 585598 1005032
rect 575699 997600 580479 1004103
rect 580559 998007 585598 1004183
rect 580779 997600 582979 998007
rect 583178 997600 585378 998007
rect 585678 997600 590458 1004952
rect 585041 997522 585107 997525
rect 585734 997522 585794 997600
rect 585041 997462 585794 997522
rect 585041 997459 585107 997462
rect 626062 997338 641914 1037600
rect 0 954262 40262 970114
rect 677338 951686 717600 967538
rect 7 927240 4850 929187
rect 30753 927121 31683 929228
rect 33910 927240 34840 929187
rect 7 922071 38140 927000
rect 38220 922151 39600 926940
rect 685910 922779 686840 924795
rect 678007 922580 717593 922600
rect 7 921851 39593 922071
rect 7 919676 39600 921851
rect 7 919376 39593 919676
rect 7 917200 39600 919376
rect 678000 917700 679380 922500
rect 679460 917620 717593 922580
rect 678007 917400 717593 917620
rect 7 916980 39593 917200
rect 7 912020 38140 916980
rect 38220 912100 39600 916900
rect 678000 915224 717593 917400
rect 678007 914924 717593 915224
rect 678000 912749 717593 914924
rect 678007 912529 717593 912749
rect 7 912000 39593 912020
rect 30760 909805 31690 911821
rect 678000 907660 679380 912449
rect 679460 907600 717593 912529
rect 682760 905413 683690 907360
rect 685917 905372 686847 907479
rect 712750 905413 717593 907360
rect 0 879798 35960 884658
rect 36040 879878 40000 884658
rect 0 879578 39593 879798
rect 0 877378 40000 879578
rect 0 877179 39593 877378
rect 0 874979 40000 877179
rect 0 874759 39593 874979
rect 0 869848 35960 874759
rect 36040 870090 40000 874679
rect 42241 870090 42307 870093
rect 44173 870090 44239 870093
rect 36040 870030 44239 870090
rect 36040 869899 40000 870030
rect 42241 870027 42307 870030
rect 44173 870027 44239 870030
rect 677338 862486 717600 878338
rect 980 837598 32568 842458
rect 32648 837678 40000 842458
rect 980 837378 39593 837598
rect 980 835178 40000 837378
rect 980 834979 39593 835178
rect 980 832779 40000 834979
rect 980 832559 39593 832779
rect 980 827648 33417 832559
rect 33497 827699 40000 832479
rect 677600 828521 680592 833301
rect 680672 828441 717600 833352
rect 678007 828221 717600 828441
rect 677600 826021 717600 828221
rect 678007 825822 717600 826021
rect 677600 823622 717600 825822
rect 678007 823402 717600 823622
rect 677600 818542 680592 823322
rect 680672 818542 717600 823402
rect 677593 818410 677659 818413
rect 677734 818410 677794 818542
rect 677593 818350 677794 818410
rect 677593 818347 677659 818350
rect 0 784462 40262 800314
rect 677338 773286 717600 789138
rect 0 741262 40262 757114
rect 677338 728286 717600 744138
rect 0 698062 40262 713914
rect 677338 683286 717600 699138
rect 0 654862 40262 670714
rect 677338 638086 717600 653938
rect 0 611662 40262 627514
rect 677338 593086 717600 608938
rect 0 568462 40262 584314
rect 677338 547886 717600 563738
rect 0 525262 40262 541114
rect 677600 513921 680592 518701
rect 677734 513773 677794 513921
rect 680672 513841 717600 518752
rect 677685 513710 677794 513773
rect 677685 513707 677751 513710
rect 678007 513621 717600 513841
rect 677600 511421 717600 513621
rect 678007 511222 717600 511421
rect 677600 509022 717600 511222
rect 678007 508802 717600 509022
rect 677600 503942 680592 508722
rect 680672 503942 717600 508802
rect 0 492998 36928 497858
rect 37008 493078 40000 497858
rect 0 492778 39593 492998
rect 0 490578 40000 492778
rect 0 490379 39593 490578
rect 0 488179 40000 490379
rect 0 487959 39593 488179
rect 0 483048 36928 487959
rect 37008 483099 40000 487879
rect 685910 474979 686840 476995
rect 678007 474780 717593 474800
rect 686000 469820 717593 474780
rect 678007 469600 717593 469820
rect 678000 467424 717593 469600
rect 678007 467124 717593 467424
rect 678000 464949 717593 467124
rect 678007 464729 717593 464949
rect 678000 459860 685920 464649
rect 686000 459800 717593 464729
rect 7 456040 4850 457987
rect 30753 455921 31683 458028
rect 33910 456040 34840 457987
rect 682760 457613 683690 459560
rect 685917 457572 686847 459679
rect 712750 457613 717593 459560
rect 7 450871 31600 455800
rect 31680 450951 39600 455740
rect 7 450651 39593 450871
rect 7 448476 39600 450651
rect 7 448176 39593 448476
rect 7 446000 39600 448176
rect 7 445780 39593 446000
rect 7 440820 31600 445780
rect 7 440800 39593 440820
rect 30760 438605 31690 440621
rect 677600 425721 684103 430501
rect 677501 425642 677567 425645
rect 677734 425642 677794 425721
rect 677501 425582 677794 425642
rect 684183 425641 716620 430552
rect 677501 425579 677567 425582
rect 678007 425421 716620 425641
rect 677600 423221 716620 425421
rect 678007 423022 716620 423221
rect 677600 420822 716620 423022
rect 678007 420602 716620 420822
rect 677600 415742 684952 420522
rect 685032 415742 716620 420602
rect 0 397662 40262 413514
rect 677338 370686 717600 386538
rect 0 354462 40262 370314
rect 0 311262 40262 327114
rect 677338 325486 717600 341338
rect 0 268062 40262 283914
rect 677338 280486 717600 296338
rect 0 224862 40262 240714
rect 677338 235486 717600 251338
rect 0 181662 40262 197514
rect 677338 190286 717600 206138
rect 677338 145286 717600 161138
rect 0 120198 35960 125058
rect 36040 120278 40000 125058
rect 0 119978 39593 120198
rect 0 117778 40000 119978
rect 0 117579 39593 117778
rect 0 115379 40000 117579
rect 0 115159 39593 115379
rect 0 110248 35960 115159
rect 36040 110530 40000 115079
rect 44173 110530 44239 110533
rect 44817 110530 44883 110533
rect 36040 110470 44883 110530
rect 36040 110299 40000 110470
rect 44173 110467 44239 110470
rect 44817 110467 44883 110470
rect 677338 100086 717600 115938
rect 30753 83121 31683 85228
rect 31961 83088 32654 85228
rect 879 78071 38140 83000
rect 38220 78151 39600 82940
rect 879 77851 39593 78071
rect 879 75676 39600 77851
rect 879 75376 39593 75676
rect 879 73200 39600 75376
rect 879 72980 39593 73200
rect 879 68098 38140 72980
rect 38220 71906 39600 72900
rect 44173 71906 44239 71909
rect 44817 71906 44883 71909
rect 38220 71846 44883 71906
rect 38220 68100 39600 71846
rect 44173 71843 44239 71846
rect 44817 71843 44883 71846
rect 151721 46882 151787 46885
rect 188521 46882 188587 46885
rect 151721 46822 188587 46882
rect 151721 46819 151787 46822
rect 188521 46819 188587 46822
rect 204161 46882 204227 46885
rect 297081 46882 297147 46885
rect 204161 46822 297147 46882
rect 204161 46819 204227 46822
rect 297081 46819 297147 46822
rect 522481 44434 522547 44437
rect 404905 44298 404971 44301
rect 412909 44298 412975 44301
rect 404905 44238 412975 44298
rect 516090 44374 522547 44434
rect 404905 44235 404971 44238
rect 412909 44235 412975 44238
rect 459645 44298 459711 44301
rect 467649 44298 467715 44301
rect 459645 44238 467715 44298
rect 459645 44235 459711 44238
rect 467649 44235 467715 44238
rect 514477 44298 514543 44301
rect 516090 44298 516150 44374
rect 522481 44371 522547 44374
rect 514477 44238 516150 44298
rect 514477 44235 514543 44238
rect 143533 40490 143599 40493
rect 151721 40490 151787 40493
rect 143533 40430 151787 40490
rect 143533 40427 143599 40430
rect 145790 40354 145850 40430
rect 151721 40427 151787 40430
rect 145790 40294 145898 40354
rect 93761 40218 93827 40221
rect 135161 40218 135227 40221
rect 91142 40158 93827 40218
rect 91142 40000 91202 40158
rect 93761 40155 93827 40158
rect 133094 40158 135227 40218
rect 133094 40000 133154 40158
rect 135161 40155 135227 40158
rect 143073 40218 143139 40221
rect 143533 40218 143599 40221
rect 143073 40158 143458 40218
rect 143073 40155 143139 40158
rect 143398 40000 143458 40158
rect 143533 40158 144010 40218
rect 143533 40155 143599 40158
rect 143950 40000 144010 40158
rect 145838 40014 145898 40294
rect 145820 40000 145898 40014
rect 47600 32953 51202 36017
rect 51600 32953 55202 36017
rect 55600 32953 59202 36017
rect 59600 32953 63202 36017
rect 63600 32953 67202 36017
rect 67600 32953 71202 36017
rect 78942 32648 83722 40000
rect 84022 39593 86222 40000
rect 86421 39593 88621 40000
rect 83802 33417 88841 39593
rect 88921 33497 93701 40000
rect 83802 32568 93752 33417
rect 101400 32953 105002 36017
rect 105400 32953 109002 36017
rect 109400 32953 113002 36017
rect 113400 32953 117002 36017
rect 117400 32953 121002 36017
rect 121400 32953 125002 36017
rect 78942 980 93752 32568
rect 132660 30216 132868 39875
rect 132660 26680 132735 30216
rect 132948 30136 133162 40000
rect 132815 30016 133162 30136
rect 133242 37738 141587 39875
rect 141893 38746 143275 39875
rect 141893 38453 142982 38746
rect 143355 38666 143585 40000
rect 141893 38397 142926 38453
rect 143062 38420 143585 38666
rect 141893 38111 142710 38397
rect 143062 38373 143355 38420
rect 143388 38373 143585 38420
rect 143665 39293 143738 39875
rect 143818 39373 144151 40000
rect 144231 39293 145736 39875
rect 143006 38317 143062 38373
rect 143332 38317 143388 38373
rect 141953 38051 142710 38111
rect 133242 36966 141740 37738
rect 142046 37467 142710 38051
rect 142790 38300 143006 38317
rect 143019 38300 143332 38317
rect 142790 38120 143332 38300
rect 143665 38293 145736 39293
rect 143468 38237 145736 38293
rect 142790 38101 143006 38120
rect 143019 38101 143332 38120
rect 142790 38004 143332 38101
rect 142790 37547 143019 38004
rect 143412 37924 145736 38237
rect 143099 37467 145736 37924
rect 142046 36966 145736 37467
rect 133242 36603 145736 36966
rect 145816 36843 145920 40000
rect 146000 36923 147407 39875
rect 146042 36881 147407 36923
rect 145816 36801 145962 36843
rect 145816 36741 145934 36801
rect 145962 36741 146052 36801
rect 146132 36791 147407 36881
rect 145816 36711 146052 36741
rect 145816 36683 145934 36711
rect 145934 36651 146026 36683
rect 146052 36651 146142 36711
rect 146222 36701 147407 36791
rect 145934 36621 146142 36651
rect 133242 36511 145854 36603
rect 145934 36591 146245 36621
rect 146026 36531 146141 36591
rect 146142 36531 146245 36591
rect 133242 36396 145946 36511
rect 146026 36476 146245 36531
rect 133242 33821 146061 36396
rect 133242 33704 145944 33821
rect 146141 33741 146245 36476
rect 133242 33561 145801 33704
rect 146024 33669 146245 33741
rect 146024 33624 146141 33669
rect 146170 33624 146245 33669
rect 145881 33609 146024 33624
rect 146027 33609 146170 33624
rect 133242 33444 145684 33561
rect 145881 33519 146170 33609
rect 146325 33544 147407 36701
rect 145881 33481 146024 33519
rect 146027 33481 146170 33519
rect 145764 33459 145881 33481
rect 145910 33459 146027 33481
rect 133242 33401 145641 33444
rect 133242 33095 143065 33401
rect 145764 33399 146027 33459
rect 146250 33401 147407 33544
rect 145764 33364 145881 33399
rect 145910 33364 146027 33399
rect 145721 33321 145764 33364
rect 145806 33321 145910 33364
rect 143145 33291 145910 33321
rect 143145 33260 145777 33261
rect 145806 33260 145910 33291
rect 146107 33284 147407 33401
rect 143145 33231 145806 33260
rect 145721 33201 145806 33231
rect 143145 33175 145806 33201
rect 145990 33180 147407 33284
rect 145886 33095 147407 33180
rect 132815 30003 132948 30016
rect 132815 27080 133162 30003
rect 133242 27160 147407 33095
rect 155200 32953 158802 36017
rect 159200 32953 162802 36017
rect 163200 32953 166802 36017
rect 167200 32953 170802 36017
rect 171200 32953 174802 36017
rect 175200 32953 178802 36017
rect 132815 26760 133482 27080
rect 133562 26840 147407 27160
rect 132660 26360 133082 26680
rect 133162 26480 133762 26760
rect 133842 26560 147407 26840
rect 133162 26450 133949 26480
rect 133162 26440 133482 26450
rect 133482 26390 133739 26440
rect 133762 26390 133949 26450
rect 132660 26103 133402 26360
rect 133482 26293 133949 26390
rect 134029 26373 147407 26560
rect 133482 26270 133942 26293
rect 133482 26240 133739 26270
rect 133949 26240 134122 26293
rect 133482 26210 134122 26240
rect 133482 26183 133739 26210
rect 133739 26180 133929 26183
rect 133949 26180 134122 26210
rect 134202 26200 147407 26373
rect 133739 26120 134122 26180
rect 132660 25913 133659 26103
rect 133739 26090 134392 26120
rect 133739 26060 133929 26090
rect 134122 26060 134392 26090
rect 133739 26000 134392 26060
rect 133739 25993 133929 26000
rect 134122 25993 134392 26000
rect 132660 25720 133849 25913
rect 133929 25850 134392 25993
rect 134472 25930 147407 26200
rect 133929 25820 134628 25850
rect 133929 25800 134122 25820
rect 134122 25760 134364 25800
rect 134392 25760 134628 25820
rect 132660 25478 134042 25720
rect 134122 25584 134628 25760
rect 134122 25558 134364 25584
rect 134368 25558 134628 25584
rect 134364 25520 134628 25558
rect 132660 25440 134284 25478
rect 132660 20991 134322 25440
rect 134402 21071 134628 25520
rect 134708 20991 147407 25930
rect 132660 0 147407 20991
rect 186486 0 202338 40262
rect 248413 39946 248479 39949
rect 241286 39886 248479 39946
rect 241286 39600 241346 39886
rect 248413 39883 248479 39886
rect 210000 32953 213602 36017
rect 214000 32953 217602 36017
rect 218000 32953 221602 36017
rect 222000 32953 225602 36017
rect 226000 32953 229602 36017
rect 230000 32953 233602 36017
rect 238972 31961 241112 32654
rect 238972 30753 241079 31683
rect 241260 31680 246049 39600
rect 246349 39593 248524 39600
rect 248824 39593 251000 39600
rect 246129 31600 251220 39593
rect 251300 31680 256100 39600
rect 263800 32953 267402 36017
rect 267800 32953 271402 36017
rect 271800 32953 275402 36017
rect 275800 32953 279402 36017
rect 279800 32953 283402 36017
rect 283800 32953 287402 36017
rect 241200 879 256100 31600
rect 295086 0 310938 40262
rect 318600 32953 322202 36017
rect 322600 32953 326202 36017
rect 326600 32953 330202 36017
rect 330600 32953 334202 36017
rect 334600 32953 338202 36017
rect 338600 32953 342202 36017
rect 349886 0 365738 40262
rect 373400 32953 377002 36017
rect 377400 32953 381002 36017
rect 381400 32953 385002 36017
rect 385400 32953 389002 36017
rect 389400 32953 393002 36017
rect 393400 32953 397002 36017
rect 404686 0 420538 40262
rect 428200 32953 431802 36017
rect 432200 32953 435802 36017
rect 436200 32953 439802 36017
rect 440200 32953 443802 36017
rect 444200 32953 447802 36017
rect 448200 32953 451802 36017
rect 459486 0 475338 40262
rect 483000 32953 486602 36017
rect 487000 32953 490602 36017
rect 491000 32953 494602 36017
rect 495000 32953 498602 36017
rect 499000 32953 502602 36017
rect 503000 32953 506602 36017
rect 514286 0 530138 40262
rect 569125 40218 569191 40221
rect 569125 40155 569234 40218
rect 569174 40000 569234 40155
rect 537800 32953 541402 36017
rect 541800 32953 545402 36017
rect 545800 32953 549402 36017
rect 549800 32953 553402 36017
rect 553800 32953 557402 36017
rect 557800 32953 561402 36017
rect 569142 34830 573922 40000
rect 574222 39593 576422 40000
rect 576621 39593 578821 40000
rect 574002 34750 579041 39593
rect 579121 34830 583901 40000
rect 622942 37008 627722 40000
rect 628022 39593 630222 40000
rect 630421 39593 632621 40000
rect 627802 36928 632841 39593
rect 632921 37008 637701 40000
rect 569142 0 583952 34750
rect 591600 32953 595202 36017
rect 595600 32953 599202 36017
rect 599600 32953 603202 36017
rect 603600 32953 607202 36017
rect 607600 32953 611202 36017
rect 611600 32953 615202 36017
rect 622942 0 637752 36928
rect 645400 32953 649002 36017
rect 649400 32953 653002 36017
rect 653400 32953 657002 36017
rect 657400 32953 661002 36017
rect 661400 32953 665002 36017
rect 665400 32953 669002 36017
<< metal4 >>
rect 7 455800 4843 456094
rect 0 455546 4843 455800
rect 28653 407018 28719 525722
rect 32933 455546 33623 483254
rect 36323 455607 37013 483193
rect 37293 455546 38223 483254
rect 38503 455546 39593 483254
rect 679377 430346 680307 460054
rect 680587 430407 681277 459993
rect 688881 430346 688947 554382
<< obsm4 >>
rect 0 1032677 40466 1037600
rect 40546 1032757 76454 1037600
rect 0 1016680 40549 1032677
rect 40800 1016680 76200 1032757
rect 76534 1032677 91866 1037600
rect 91946 1032757 127854 1037600
rect 76393 1016680 91994 1032677
rect 92200 1016680 127600 1032757
rect 127934 1032677 143266 1037600
rect 143346 1032757 179254 1037600
rect 127793 1016680 143394 1032677
rect 143600 1016680 179000 1032757
rect 179334 1032677 194666 1037600
rect 194746 1032757 230654 1037600
rect 179193 1016680 194794 1032677
rect 195000 1016680 230400 1032757
rect 230734 1032677 246066 1037600
rect 246146 1032757 282254 1037600
rect 230593 1016680 246194 1032677
rect 246400 1016680 282000 1032757
rect 282334 1032677 297666 1037600
rect 297746 1032757 333654 1037600
rect 282193 1016680 297794 1032677
rect 298000 1016680 333400 1032757
rect 333734 1032677 348066 1037600
rect 348146 1032757 384054 1037600
rect 333593 1016680 348207 1032677
rect 348400 1016680 383800 1032757
rect 384134 1032677 399466 1037600
rect 399546 1032757 473054 1037600
rect 383993 1016680 399594 1032677
rect 399800 1016680 435200 1032757
rect 437200 1016680 472800 1032757
rect 473134 1032677 488466 1037600
rect 488546 1032757 524454 1037600
rect 472993 1016680 488594 1032677
rect 488800 1016680 524200 1032757
rect 524534 1032677 539866 1037600
rect 539946 1032757 575854 1037600
rect 524393 1016680 539994 1032677
rect 540200 1016680 575600 1032757
rect 575934 1032677 590266 1037600
rect 590346 1032757 626254 1037600
rect 575793 1016680 590407 1032677
rect 590600 1016680 626000 1032757
rect 626334 1032677 641666 1037600
rect 641746 1032757 677887 1037600
rect 642000 1032677 677600 1032757
rect 677967 1032677 717600 1037600
rect 626193 1016680 641794 1032677
rect 642000 1016680 717600 1032677
rect 0 1011527 40349 1016680
rect 40429 1011607 76454 1016600
rect 76534 1011527 91866 1016680
rect 91946 1011607 127854 1016600
rect 127934 1011527 143266 1016680
rect 143346 1011607 179254 1016600
rect 179334 1011527 194666 1016680
rect 194746 1011607 230654 1016600
rect 230734 1011527 246066 1016680
rect 246146 1011607 282254 1016600
rect 282334 1011527 297666 1016680
rect 297746 1011607 333654 1016600
rect 333734 1011527 348066 1016680
rect 348146 1011607 384054 1016600
rect 384134 1011527 399466 1016680
rect 399546 1011607 473054 1016600
rect 473134 1011527 488466 1016680
rect 488546 1011607 524454 1016600
rect 524534 1011527 539866 1016680
rect 539946 1011607 575854 1016600
rect 575934 1011527 590266 1016680
rect 590346 1011607 626254 1016600
rect 626334 1011527 641666 1016680
rect 641746 1011607 678129 1016600
rect 678209 1011527 717600 1016680
rect 0 1011387 40549 1011527
rect 40800 1011387 76200 1011527
rect 76393 1011387 91994 1011527
rect 92200 1011387 127600 1011527
rect 127793 1011387 143394 1011527
rect 143600 1011387 179000 1011527
rect 179193 1011387 194794 1011527
rect 195000 1011387 230400 1011527
rect 230593 1011387 246194 1011527
rect 246400 1011387 282000 1011527
rect 282193 1011387 297794 1011527
rect 298000 1011387 333400 1011527
rect 333593 1011387 348207 1011527
rect 348400 1011387 383800 1011527
rect 383993 1011387 399594 1011527
rect 399800 1011387 435200 1011527
rect 437200 1011387 472800 1011527
rect 472993 1011387 488594 1011527
rect 488800 1011387 524200 1011527
rect 524393 1011387 539994 1011527
rect 540200 1011387 575600 1011527
rect 575793 1011387 590407 1011527
rect 590600 1011387 626000 1011527
rect 626193 1011387 641794 1011527
rect 642000 1011387 717600 1011527
rect 0 1010337 40466 1011387
rect 40546 1010417 76454 1011307
rect 76534 1010337 91866 1011387
rect 91946 1010417 127854 1011307
rect 127934 1010337 143266 1011387
rect 143346 1010417 179254 1011307
rect 179334 1010337 194666 1011387
rect 194746 1010417 230654 1011307
rect 230734 1010337 246066 1011387
rect 246146 1010417 282254 1011307
rect 282334 1010337 297666 1011387
rect 297746 1010417 333654 1011307
rect 333734 1010337 348066 1011387
rect 348146 1010417 384054 1011307
rect 384134 1010337 399466 1011387
rect 399546 1010417 473054 1011307
rect 473134 1010337 488466 1011387
rect 488546 1010417 524454 1011307
rect 524534 1010337 539866 1011387
rect 539946 1010417 575854 1011307
rect 575934 1010337 590266 1011387
rect 590346 1010417 626254 1011307
rect 626334 1010337 641666 1011387
rect 641746 1010417 677896 1011307
rect 677976 1010337 717600 1011387
rect 0 1010217 40549 1010337
rect 40800 1010217 76200 1010337
rect 76393 1010217 91994 1010337
rect 92200 1010217 127600 1010337
rect 127793 1010217 143394 1010337
rect 143600 1010217 179000 1010337
rect 179193 1010217 194794 1010337
rect 195000 1010217 230400 1010337
rect 230593 1010217 246194 1010337
rect 246400 1010217 282000 1010337
rect 282193 1010217 297794 1010337
rect 298000 1010217 333400 1010337
rect 333593 1010217 348207 1010337
rect 348400 1010217 383800 1010337
rect 383993 1010217 399594 1010337
rect 399800 1010217 435200 1010337
rect 437200 1010217 472800 1010337
rect 472993 1010217 488594 1010337
rect 488800 1010217 524200 1010337
rect 524393 1010217 539994 1010337
rect 540200 1010217 575600 1010337
rect 575793 1010217 590407 1010337
rect 590600 1010217 626000 1010337
rect 626193 1010217 641794 1010337
rect 642000 1010217 717600 1010337
rect 0 1009167 40466 1010217
rect 40546 1009247 76454 1010137
rect 76534 1009167 91866 1010217
rect 91946 1009247 127854 1010137
rect 127934 1009167 143266 1010217
rect 143346 1009247 179254 1010137
rect 179334 1009167 194666 1010217
rect 194746 1009247 230654 1010137
rect 230734 1009167 246066 1010217
rect 246146 1009247 282254 1010137
rect 282334 1009167 297666 1010217
rect 297746 1009247 333654 1010137
rect 333734 1009167 348066 1010217
rect 348146 1009247 384054 1010137
rect 384134 1009167 399466 1010217
rect 399546 1009247 473054 1010137
rect 473134 1009167 488466 1010217
rect 488546 1009247 524454 1010137
rect 524534 1009167 539866 1010217
rect 539946 1009247 575854 1010137
rect 575934 1009167 590266 1010217
rect 590346 1009247 626254 1010137
rect 626334 1009167 641666 1010217
rect 641746 1009247 677925 1010137
rect 678005 1009167 717600 1010217
rect 0 1009027 40549 1009167
rect 40800 1009027 76200 1009167
rect 76393 1009027 91994 1009167
rect 92200 1009027 127600 1009167
rect 127793 1009027 143394 1009167
rect 143600 1009027 179000 1009167
rect 179193 1009027 194794 1009167
rect 195000 1009027 230400 1009167
rect 230593 1009027 246194 1009167
rect 246400 1009027 282000 1009167
rect 282193 1009027 297794 1009167
rect 298000 1009027 333400 1009167
rect 333593 1009027 348207 1009167
rect 348400 1009027 383800 1009167
rect 383993 1009027 399594 1009167
rect 399800 1009027 435200 1009167
rect 437200 1009027 472800 1009167
rect 472993 1009027 488594 1009167
rect 488800 1009027 524200 1009167
rect 524393 1009027 539994 1009167
rect 540200 1009027 575600 1009167
rect 575793 1009027 590407 1009167
rect 590600 1009027 626000 1009167
rect 626193 1009027 641794 1009167
rect 642000 1009027 717600 1009167
rect 0 1008801 35285 1009027
rect 35365 1008881 76722 1008947
rect 76802 1008901 85538 1009027
rect 0 1008145 35338 1008801
rect 35418 1008225 83488 1008821
rect 0 1007849 36409 1008145
rect 36489 1007929 76454 1008165
rect 83568 1008145 83872 1008901
rect 85618 1008881 128122 1008947
rect 128202 1008901 136938 1009027
rect 83952 1008225 134888 1008821
rect 76534 1007949 91866 1008145
rect 0 1007293 36545 1007849
rect 0 1007067 36005 1007293
rect 36625 1007273 86629 1007869
rect 86709 1007293 87013 1007949
rect 91946 1007929 127854 1008165
rect 134968 1008145 135272 1008901
rect 137018 1008881 179522 1008947
rect 179602 1008901 188338 1009027
rect 135352 1008225 186288 1008821
rect 127934 1007949 143266 1008145
rect 87093 1007273 138029 1007869
rect 138109 1007293 138413 1007949
rect 143346 1007929 179254 1008165
rect 186368 1008145 186672 1008901
rect 188418 1008881 230922 1008947
rect 231002 1008901 239738 1009027
rect 186752 1008225 237688 1008821
rect 179334 1007949 194666 1008145
rect 138493 1007273 189429 1007869
rect 189509 1007293 189813 1007949
rect 194746 1007929 230654 1008165
rect 237768 1008145 238072 1008901
rect 239818 1008881 282522 1008947
rect 282602 1008901 291338 1009027
rect 238152 1008225 289288 1008821
rect 230734 1007949 246066 1008145
rect 189893 1007273 240829 1007869
rect 240909 1007293 241213 1007949
rect 246146 1007929 282254 1008165
rect 289368 1008145 289672 1008901
rect 291418 1008881 384322 1008947
rect 384402 1008901 393138 1009027
rect 289752 1008225 391088 1008821
rect 282334 1007949 297666 1008145
rect 241293 1007273 292429 1007869
rect 292509 1007293 292813 1007949
rect 297746 1007929 333654 1008165
rect 333734 1007949 348066 1008145
rect 348146 1007929 384054 1008165
rect 391168 1008145 391472 1008901
rect 393218 1008881 435200 1008947
rect 436200 1008881 473322 1008947
rect 473402 1008901 482138 1009027
rect 391552 1008225 480088 1008821
rect 384134 1007949 399466 1008145
rect 292893 1007273 394229 1007869
rect 394309 1007293 394613 1007949
rect 399546 1007929 435200 1008165
rect 436200 1007929 473054 1008165
rect 480168 1008145 480472 1008901
rect 482218 1008881 524722 1008947
rect 524802 1008901 533538 1009027
rect 480552 1008225 531488 1008821
rect 473134 1007949 488466 1008145
rect 394693 1007273 483229 1007869
rect 483309 1007293 483613 1007949
rect 488546 1007929 524454 1008165
rect 531568 1008145 531872 1008901
rect 533618 1008881 575854 1008947
rect 575934 1008901 590266 1009027
rect 590346 1008881 626522 1008947
rect 626602 1008901 635338 1009027
rect 531952 1008225 633288 1008821
rect 524534 1007949 539866 1008145
rect 483693 1007273 534629 1007869
rect 534709 1007293 535013 1007949
rect 539946 1007929 575854 1008165
rect 575934 1007949 590266 1008145
rect 590346 1007929 626254 1008165
rect 633368 1008145 633672 1008901
rect 635418 1008881 682235 1008947
rect 633752 1008225 682182 1008821
rect 682315 1008801 717600 1009027
rect 626334 1007949 641666 1008145
rect 535093 1007273 636429 1007869
rect 636509 1007293 636813 1007949
rect 641746 1007929 681910 1008165
rect 682262 1008145 717600 1008801
rect 636893 1007273 681787 1007869
rect 681990 1007849 717600 1008145
rect 36085 1007147 76722 1007213
rect 76802 1007067 85538 1007193
rect 85618 1007147 128122 1007213
rect 128202 1007067 136938 1007193
rect 137018 1007147 179522 1007213
rect 179602 1007067 188338 1007193
rect 188418 1007147 230922 1007213
rect 231002 1007067 239738 1007193
rect 239818 1007147 282522 1007213
rect 282602 1007067 291338 1007193
rect 291418 1007147 384322 1007213
rect 384402 1007067 393138 1007193
rect 393218 1007147 435200 1007213
rect 436200 1007147 473322 1007213
rect 473402 1007067 482138 1007193
rect 482218 1007147 524722 1007213
rect 524802 1007067 533538 1007193
rect 533618 1007147 575854 1007213
rect 575934 1007067 590266 1007193
rect 590346 1007147 626522 1007213
rect 626602 1007067 635338 1007193
rect 635418 1007147 681515 1007213
rect 681867 1007193 717600 1007849
rect 681595 1007067 717600 1007193
rect 0 1006927 40549 1007067
rect 76393 1006927 91994 1007067
rect 127793 1006927 143394 1007067
rect 179193 1006927 194794 1007067
rect 230593 1006927 246194 1007067
rect 282193 1006927 297794 1007067
rect 333593 1006927 348207 1007067
rect 383993 1006927 399594 1007067
rect 472993 1006927 488594 1007067
rect 524393 1006927 539994 1007067
rect 575793 1006927 590407 1007067
rect 626193 1006927 641794 1007067
rect 677600 1006927 717600 1007067
rect 0 1005837 40466 1006927
rect 40546 1005917 76454 1006847
rect 76534 1005837 91866 1006927
rect 91946 1005917 127854 1006847
rect 127934 1005837 143266 1006927
rect 143346 1005917 179254 1006847
rect 179334 1005837 194666 1006927
rect 194746 1005917 230654 1006847
rect 230734 1005837 246066 1006927
rect 246146 1005917 282254 1006847
rect 282334 1005837 297666 1006927
rect 297746 1005917 333654 1006847
rect 333734 1005837 348066 1006927
rect 348146 1005917 384054 1006847
rect 384134 1005837 399466 1006927
rect 399546 1005917 436200 1006847
rect 437200 1005917 473054 1006847
rect 473134 1005837 488466 1006927
rect 488546 1005917 524454 1006847
rect 524534 1005837 539866 1006927
rect 539946 1005917 575854 1006847
rect 575934 1005837 590266 1006927
rect 590346 1005917 626254 1006847
rect 626334 1005837 641666 1006927
rect 641746 1005917 677895 1006847
rect 677975 1005837 717600 1006927
rect 0 1005717 40549 1005837
rect 76393 1005717 91994 1005837
rect 127793 1005717 143394 1005837
rect 179193 1005717 194794 1005837
rect 230593 1005717 246194 1005837
rect 282193 1005717 297794 1005837
rect 333593 1005717 348207 1005837
rect 383993 1005717 399594 1005837
rect 472993 1005717 488594 1005837
rect 524393 1005717 539994 1005837
rect 575793 1005717 590407 1005837
rect 626193 1005717 641794 1005837
rect 677600 1005717 717600 1005837
rect 0 1004867 40466 1005717
rect 40546 1004947 76454 1005637
rect 76534 1004867 91866 1005717
rect 91946 1004947 127854 1005637
rect 127934 1004867 143266 1005717
rect 143346 1004947 179254 1005637
rect 179334 1004867 194666 1005717
rect 194746 1004947 230654 1005637
rect 230734 1004867 246066 1005717
rect 246146 1004947 282254 1005637
rect 282334 1004867 297666 1005717
rect 297746 1004947 333654 1005637
rect 333734 1004867 348066 1005717
rect 348146 1004947 384054 1005637
rect 384134 1004867 399466 1005717
rect 399546 1004947 435200 1005637
rect 436200 1004947 473054 1005637
rect 473134 1004867 488466 1005717
rect 488546 1004947 524454 1005637
rect 524534 1004867 539866 1005717
rect 539946 1004947 575854 1005637
rect 575934 1004867 590266 1005717
rect 590346 1004947 626254 1005637
rect 626334 1004867 641666 1005717
rect 641746 1004947 677867 1005637
rect 677947 1004867 717600 1005717
rect 0 1004747 40549 1004867
rect 76393 1004747 91994 1004867
rect 127793 1004747 143394 1004867
rect 179193 1004747 194794 1004867
rect 230593 1004747 246194 1004867
rect 282193 1004747 297794 1004867
rect 333593 1004747 348207 1004867
rect 383993 1004747 399594 1004867
rect 472993 1004747 488594 1004867
rect 524393 1004747 539994 1004867
rect 575793 1004747 590407 1004867
rect 626193 1004747 641794 1004867
rect 677600 1004747 717600 1004867
rect 0 1003897 40466 1004747
rect 40546 1003977 76454 1004667
rect 76534 1003897 91866 1004747
rect 91946 1003977 127854 1004667
rect 127934 1003897 143266 1004747
rect 143346 1003977 179254 1004667
rect 179334 1003897 194666 1004747
rect 194746 1003977 230654 1004667
rect 230734 1003897 246066 1004747
rect 246146 1003977 282254 1004667
rect 282334 1003897 297666 1004747
rect 297746 1003977 333654 1004667
rect 333734 1003897 348066 1004747
rect 348146 1003977 384054 1004667
rect 384134 1003897 399466 1004747
rect 399546 1003977 473054 1004667
rect 473134 1003897 488466 1004747
rect 488546 1003977 524454 1004667
rect 524534 1003897 539866 1004747
rect 539946 1003977 575854 1004667
rect 575934 1003897 590266 1004747
rect 590346 1003977 626254 1004667
rect 626334 1003897 641666 1004747
rect 641746 1003977 677877 1004667
rect 677957 1003897 717600 1004747
rect 0 1003777 40549 1003897
rect 76393 1003777 91994 1003897
rect 127793 1003777 143394 1003897
rect 179193 1003777 194794 1003897
rect 230593 1003777 246194 1003897
rect 282193 1003777 297794 1003897
rect 333593 1003777 348207 1003897
rect 383993 1003777 399594 1003897
rect 472993 1003777 488594 1003897
rect 524393 1003777 539994 1003897
rect 575793 1003777 590407 1003897
rect 626193 1003777 641794 1003897
rect 677600 1003777 717600 1003897
rect 0 1002687 40466 1003777
rect 40546 1002767 76454 1003697
rect 76534 1002687 91866 1003777
rect 91946 1002767 127854 1003697
rect 127934 1002687 143266 1003777
rect 143346 1002767 179254 1003697
rect 179334 1002687 194666 1003777
rect 194746 1002767 230654 1003697
rect 230734 1002687 246066 1003777
rect 246146 1002767 282254 1003697
rect 282334 1002687 297666 1003777
rect 297746 1002767 333654 1003697
rect 333734 1002687 348066 1003777
rect 348146 1002767 384054 1003697
rect 384134 1002687 399466 1003777
rect 399546 1002767 473054 1003697
rect 473134 1002687 488466 1003777
rect 488546 1002767 524454 1003697
rect 524534 1002687 539866 1003777
rect 539946 1002767 575854 1003697
rect 575934 1002687 590266 1003777
rect 590346 1002767 626254 1003697
rect 626334 1002687 641666 1003777
rect 641746 1002767 677920 1003697
rect 678000 1002687 717600 1003777
rect 0 1002567 40549 1002687
rect 76393 1002567 91994 1002687
rect 127793 1002567 143394 1002687
rect 179193 1002567 194794 1002687
rect 230593 1002567 246194 1002687
rect 282193 1002567 297794 1002687
rect 333593 1002567 348207 1002687
rect 383993 1002567 399594 1002687
rect 472993 1002567 488594 1002687
rect 524393 1002567 539994 1002687
rect 575793 1002567 590407 1002687
rect 626193 1002567 641794 1002687
rect 677600 1002567 717600 1002687
rect 0 1002315 40466 1002567
rect 0 998209 28573 1002315
rect 28799 1002262 40466 1002315
rect 0 997967 20920 998209
rect 0 997600 4843 997887
rect 4923 997600 20920 997967
rect 0 970200 20920 997600
rect 0 969946 4843 970200
rect 4923 969866 20920 969994
rect 21000 969946 25993 998129
rect 26073 998005 28573 998209
rect 26073 997976 27383 998005
rect 26073 970200 26213 997976
rect 26073 969866 26213 969994
rect 26293 969946 27183 997896
rect 27263 970200 27383 997976
rect 27263 969866 27383 969994
rect 27463 969946 28353 997925
rect 28433 970200 28573 998005
rect 28433 969866 28573 969994
rect 0 963538 28573 969866
rect 28653 963618 28719 1002235
rect 0 961872 28699 963538
rect 28779 961952 29375 1002182
rect 29455 1001990 40466 1002262
rect 29435 969946 29671 1001910
rect 29751 1001867 40466 1001990
rect 29455 965013 29651 969866
rect 29731 965093 30327 1001787
rect 30407 1001595 40466 1001867
rect 29455 964709 30307 965013
rect 29455 961872 29651 964709
rect 0 961568 29651 961872
rect 0 954802 28699 961568
rect 0 954534 28573 954802
rect 0 954200 4843 954454
rect 4923 954393 20920 954534
rect 0 927000 20920 954200
rect 0 926957 4850 927000
rect 0 926746 4843 926957
rect 4923 926666 20920 927000
rect 21000 926746 25993 954454
rect 26073 954393 26213 954534
rect 26073 926666 26213 954200
rect 26293 926746 27183 954454
rect 27263 954393 27383 954534
rect 27263 926666 27383 954200
rect 27463 926746 28353 954454
rect 28433 954393 28573 954534
rect 28433 926666 28573 954200
rect 0 912334 28573 926666
rect 0 912000 4843 912254
rect 4923 912000 20920 912334
rect 0 884800 20920 912000
rect 0 884546 4843 884800
rect 4923 884466 20920 884607
rect 21000 884546 25993 912254
rect 26073 884800 26213 912334
rect 26073 884466 26213 884607
rect 26293 884546 27183 912254
rect 27263 884800 27383 912334
rect 27263 884466 27383 884607
rect 27463 884546 28353 912254
rect 28433 884800 28573 912334
rect 28433 884466 28573 884607
rect 0 870134 28573 884466
rect 0 869800 4843 870054
rect 4923 869993 20920 870134
rect 0 842600 20920 869800
rect 0 842346 4843 842600
rect 4923 842266 20920 842407
rect 21000 842346 25993 870054
rect 26073 869993 26213 870134
rect 26073 842600 26213 869800
rect 26073 842266 26213 842407
rect 26293 842346 27183 870054
rect 27263 869993 27383 870134
rect 27263 842600 27383 869800
rect 27263 842266 27383 842407
rect 27463 842346 28353 870054
rect 28433 869993 28573 870134
rect 28433 842600 28573 869800
rect 28433 842266 28573 842407
rect 28653 842346 28719 954722
rect 0 827934 28699 842266
rect 0 827600 4843 827854
rect 4923 827793 20920 827934
rect 0 800400 20920 827600
rect 0 800146 4843 800400
rect 4923 800066 20920 800194
rect 21000 800146 25993 827854
rect 26073 827793 26213 827934
rect 26073 800400 26213 827600
rect 26073 800066 26213 800194
rect 26293 800146 27183 827854
rect 27263 827793 27383 827934
rect 27263 800400 27383 827600
rect 27263 800066 27383 800194
rect 27463 800146 28353 827854
rect 28433 827793 28573 827934
rect 28433 800400 28573 827600
rect 28433 800066 28573 800194
rect 0 793738 28573 800066
rect 28653 793818 28719 827854
rect 0 792072 28699 793738
rect 28779 792152 29375 961488
rect 29455 954534 29651 961568
rect 29435 926746 29671 954454
rect 29455 912334 29651 926666
rect 29435 884546 29671 912254
rect 29455 870134 29651 884466
rect 29435 842346 29671 870054
rect 29455 827934 29651 842266
rect 29435 800146 29671 827854
rect 29455 795213 29651 800066
rect 29731 795293 30327 964629
rect 30387 963618 30453 1001515
rect 30533 1001477 40466 1001595
rect 40546 1001557 76454 1002487
rect 76534 1001477 91866 1002567
rect 91946 1001557 127854 1002487
rect 127934 1001477 143266 1002567
rect 143346 1001557 179254 1002487
rect 179334 1001477 194666 1002567
rect 194746 1001557 230654 1002487
rect 230734 1001477 246066 1002567
rect 246146 1001557 282254 1002487
rect 282334 1001477 297666 1002567
rect 297746 1001557 333654 1002487
rect 333734 1001477 348066 1002567
rect 348146 1001557 384054 1002487
rect 384134 1001477 399466 1002567
rect 399546 1001557 473054 1002487
rect 473134 1001477 488466 1002567
rect 488546 1001557 524454 1002487
rect 524534 1001477 539866 1002567
rect 539946 1001557 575854 1002487
rect 575934 1001477 590266 1002567
rect 590346 1001557 626254 1002487
rect 626334 1001477 641666 1002567
rect 641746 1001557 677905 1002487
rect 677985 1002315 717600 1002567
rect 677985 1002262 688801 1002315
rect 677985 1001595 688145 1002262
rect 677985 1001477 687067 1001595
rect 30533 1001357 40549 1001477
rect 76393 1001357 91994 1001477
rect 127793 1001357 143394 1001477
rect 179193 1001357 194794 1001477
rect 230593 1001357 246194 1001477
rect 282193 1001357 297794 1001477
rect 333593 1001357 348207 1001477
rect 383993 1001357 399594 1001477
rect 472993 1001357 488594 1001477
rect 524393 1001357 539994 1001477
rect 575793 1001357 590407 1001477
rect 626193 1001357 641794 1001477
rect 677600 1001357 687067 1001477
rect 30533 1000507 40469 1001357
rect 40549 1000587 76393 1001277
rect 76473 1000507 91914 1001357
rect 91994 1000587 127793 1001277
rect 127873 1000507 143314 1001357
rect 143394 1000587 179193 1001277
rect 179273 1000507 194714 1001357
rect 194794 1000587 230593 1001277
rect 230673 1000507 246114 1001357
rect 246194 1000587 282193 1001277
rect 282273 1000507 297714 1001357
rect 297794 1000587 333593 1001277
rect 333673 1000507 348127 1001357
rect 348207 1000587 383993 1001277
rect 384073 1000507 399514 1001357
rect 399594 1000587 435200 1001277
rect 436200 1000587 472993 1001277
rect 473073 1000507 488514 1001357
rect 488594 1000587 524393 1001277
rect 524473 1000507 539914 1001357
rect 539994 1000587 575793 1001277
rect 575873 1000507 590327 1001357
rect 590407 1000587 626193 1001277
rect 626273 1000507 641714 1001357
rect 641794 1000587 677894 1001277
rect 677974 1000507 687067 1001357
rect 30533 1000387 40549 1000507
rect 76393 1000387 91994 1000507
rect 127793 1000387 143394 1000507
rect 179193 1000387 194794 1000507
rect 230593 1000387 246194 1000507
rect 282193 1000387 297794 1000507
rect 333593 1000387 348207 1000507
rect 383993 1000387 399594 1000507
rect 472993 1000387 488594 1000507
rect 524393 1000387 539994 1000507
rect 575793 1000387 590407 1000507
rect 626193 1000387 641794 1000507
rect 677600 1000387 687067 1000507
rect 30533 999297 40466 1000387
rect 40546 999377 76454 1000307
rect 76534 999297 91866 1000387
rect 91946 999377 127854 1000307
rect 127934 999297 143266 1000387
rect 143346 999377 179254 1000307
rect 179334 999297 194666 1000387
rect 194746 999377 230654 1000307
rect 230734 999297 246066 1000387
rect 246146 999377 282254 1000307
rect 282334 999297 297666 1000387
rect 297746 999377 333654 1000307
rect 333734 999297 348066 1000387
rect 348146 999377 384054 1000307
rect 384134 999297 399466 1000387
rect 399546 999377 436200 1000307
rect 437200 999377 473054 1000307
rect 473134 999297 488466 1000387
rect 488546 999377 524454 1000307
rect 524534 999297 539866 1000387
rect 539946 999377 575854 1000307
rect 575934 999297 590266 1000387
rect 590346 999377 626254 1000307
rect 626334 999297 641666 1000387
rect 641746 999377 678357 1000307
rect 678437 999297 687067 1000387
rect 30533 999177 40549 999297
rect 76393 999177 91994 999297
rect 127793 999177 143394 999297
rect 179193 999177 194794 999297
rect 230593 999177 246194 999297
rect 282193 999177 297794 999297
rect 333593 999177 348207 999297
rect 383993 999177 399594 999297
rect 472993 999177 488594 999297
rect 524393 999177 539994 999297
rect 575793 999177 590407 999297
rect 626193 999177 641794 999297
rect 677600 999177 687067 999297
rect 30533 998437 40466 999177
rect 30533 998000 37213 998437
rect 30533 997975 33823 998000
rect 30533 997600 30673 997975
rect 31763 997957 33823 997975
rect 31763 997947 32853 997957
rect 30533 969866 30673 969994
rect 30753 969946 31683 997895
rect 31763 997600 31883 997947
rect 31763 969866 31883 969994
rect 31963 969946 32653 997867
rect 32733 997600 32853 997947
rect 32733 969866 32853 969994
rect 32933 969946 33623 997877
rect 33703 997600 33823 997957
rect 34913 997985 37213 998000
rect 33703 969866 33823 969994
rect 33903 969946 34833 997920
rect 34913 997600 35033 997985
rect 36123 997974 37213 997985
rect 34913 969866 35033 969994
rect 35113 969946 36043 997905
rect 36123 997600 36243 997974
rect 36323 969994 37013 997894
rect 37093 997600 37213 997974
rect 36123 969914 36243 969994
rect 37093 969914 37213 969994
rect 37293 969946 38223 998357
rect 38303 998150 40466 998437
rect 38303 997600 38423 998150
rect 38503 998007 39593 998070
rect 39673 998007 40466 998150
rect 40546 998007 76454 999097
rect 38503 997927 40466 998007
rect 76534 997927 91866 999177
rect 91946 998007 127854 999097
rect 127934 997927 143266 999177
rect 143346 998007 179254 999097
rect 179334 997927 194666 999177
rect 194746 998007 230654 999097
rect 230734 997927 246066 999177
rect 246146 998007 282254 999097
rect 282334 997927 297666 999177
rect 297746 998007 333654 999097
rect 333734 998007 348066 999177
rect 348146 998007 384054 999097
rect 384134 997927 399466 999177
rect 399546 998007 473054 999097
rect 473134 997927 488466 999177
rect 488546 998007 524454 999097
rect 524534 997927 539866 999177
rect 539946 998007 575854 999097
rect 575934 998007 590266 999177
rect 590346 998007 626254 999097
rect 626334 997927 641666 999177
rect 641746 998007 678070 999097
tri 677600 997927 677680 998007 ne
rect 677680 997927 678007 998007
rect 678150 997927 687067 999177
rect 38503 997680 40549 997927
rect 76393 997707 91994 997927
rect 127793 997707 143394 997927
rect 179193 997707 194794 997927
rect 230593 997707 246194 997927
rect 282193 997707 297794 997927
rect 383993 997707 399594 997927
rect 472993 997707 488594 997927
rect 524393 997707 539994 997927
rect 626193 997707 641794 997927
rect 36123 969866 37213 969914
rect 38303 969866 38423 969994
rect 38503 969946 39593 997680
tri 39593 997600 39673 997680 nw
rect 39673 997600 40549 997680
rect 677600 997134 687067 997927
rect 677600 997051 677927 997134
rect 39673 969866 39893 969994
rect 30533 963538 39893 969866
rect 30407 954802 39893 963538
rect 30387 842346 30453 954722
rect 30533 954534 39893 954802
rect 30533 954393 30673 954534
rect 30533 926666 30673 927000
rect 30753 926746 31683 954454
rect 31763 954393 31883 954534
rect 31763 926666 31883 927000
rect 31963 926746 32653 954454
rect 32733 954393 32853 954534
rect 32733 926666 32853 927000
rect 32933 926746 33623 954454
rect 33703 954393 33823 954534
rect 33903 929187 34833 954454
rect 34913 954393 35033 954534
rect 36123 954473 37213 954534
rect 33703 926666 33823 927000
rect 33903 926987 34840 929187
rect 33903 926746 34833 926987
rect 34913 926666 35033 927000
rect 35113 926746 36043 954454
rect 36123 954393 36243 954473
rect 37093 954393 37213 954473
rect 36123 926727 36243 927000
rect 36323 926807 37013 954393
rect 37093 926727 37213 927000
rect 37293 926746 38223 954454
rect 38303 954393 38423 954534
rect 36123 926666 37213 926727
rect 38303 926666 38423 927000
rect 38503 926746 39593 954454
rect 39673 954393 39893 954534
rect 677707 967266 677927 967407
rect 678007 967346 679097 997054
rect 679177 997051 679297 997134
rect 680387 997131 681477 997134
rect 679177 967266 679297 967407
rect 679377 967346 680307 997054
rect 680387 997051 680507 997131
rect 681357 997051 681477 997131
rect 680587 967407 681277 997051
rect 680387 967327 680507 967407
rect 681357 967327 681477 967407
rect 681557 967346 682487 997054
rect 682567 997051 682687 997134
rect 680387 967266 681477 967327
rect 682567 967266 682687 967407
rect 682767 967346 683697 997054
rect 683777 997051 683897 997134
rect 683777 967266 683897 967407
rect 683977 967346 684667 997054
rect 684747 997051 684867 997134
rect 684747 967266 684867 967407
rect 684947 967346 685637 997054
rect 685717 997051 685837 997134
rect 685717 967266 685837 967407
rect 685917 967346 686847 997054
rect 686927 997051 687067 997134
rect 686927 967266 687067 967407
rect 677707 966998 687067 967266
rect 687147 967078 687213 1001515
rect 687293 1001191 688145 1001595
rect 687293 1001055 687849 1001191
rect 677707 958262 687193 966998
rect 677707 951934 687067 958262
rect 677707 951806 677927 951934
rect 30533 912334 39593 926666
rect 678007 922346 679097 951854
rect 679177 951806 679297 951934
rect 680387 951886 681477 951934
rect 679177 922266 679297 922600
rect 679377 922346 680307 951854
rect 680387 951806 680507 951886
rect 681357 951806 681477 951886
rect 680387 922327 680507 922600
rect 680587 922407 681277 951806
rect 681357 922327 681477 922600
rect 681557 922346 682487 951854
rect 682567 951806 682687 951934
rect 680387 922266 681477 922327
rect 682567 922266 682687 922600
rect 682767 922346 683697 951854
rect 683777 951806 683897 951934
rect 683777 922266 683897 922600
rect 683977 922346 684667 951854
rect 684747 951806 684867 951934
rect 684747 922266 684867 922600
rect 684947 922346 685637 951854
rect 685717 951806 685837 951934
rect 685917 924795 686847 951854
rect 686927 951806 687067 951934
rect 685717 922266 685837 922600
rect 685910 922586 686847 924795
rect 685917 922346 686847 922586
rect 686927 922266 687067 922600
rect 30533 912000 30673 912334
rect 30753 912014 31683 912254
rect 30753 909805 31690 912014
rect 31763 912000 31883 912334
rect 30533 884466 30673 884607
rect 30753 884546 31683 909805
rect 31763 884466 31883 884607
rect 31963 884546 32653 912254
rect 32733 912000 32853 912334
rect 32733 884466 32853 884607
rect 32933 884546 33623 912254
rect 33703 912000 33823 912334
rect 33703 884466 33823 884607
rect 33903 884546 34833 912254
rect 34913 912000 35033 912334
rect 36123 912273 37213 912334
rect 34913 884466 35033 884607
rect 35113 884546 36043 912254
rect 36123 912000 36243 912273
rect 36323 884607 37013 912193
rect 37093 912000 37213 912273
rect 36123 884527 36243 884607
rect 37093 884527 37213 884607
rect 37293 884546 38223 912254
rect 38303 912000 38423 912334
rect 36123 884466 37213 884527
rect 38303 884466 38423 884607
rect 38503 884546 39593 912254
rect 678007 907934 687067 922266
rect 30533 870134 39593 884466
rect 677707 878066 677927 878207
rect 678007 878146 679097 907854
rect 679177 907600 679297 907934
rect 680387 907873 681477 907934
rect 679177 878066 679297 878207
rect 679377 878146 680307 907854
rect 680387 907600 680507 907873
rect 680587 878207 681277 907793
rect 681357 907600 681477 907873
rect 680387 878127 680507 878207
rect 681357 878127 681477 878207
rect 681557 878146 682487 907854
rect 682567 907600 682687 907934
rect 682767 907613 683697 907854
rect 682760 905413 683697 907613
rect 683777 907600 683897 907934
rect 680387 878066 681477 878127
rect 682567 878066 682687 878207
rect 682767 878146 683697 905413
rect 683777 878066 683897 878207
rect 683977 878146 684667 907854
rect 684747 907600 684867 907934
rect 684747 878066 684867 878207
rect 684947 878146 685637 907854
rect 685717 907600 685837 907934
rect 685717 878066 685837 878207
rect 685917 878146 686847 907854
rect 686927 907600 687067 907934
rect 686927 878066 687067 878207
rect 677707 877798 687067 878066
rect 687147 877878 687213 958182
rect 687273 957171 687869 1000975
rect 687929 967346 688165 1001111
rect 687949 960232 688145 967266
rect 688225 960312 688821 1002182
rect 688881 967078 688947 1002235
rect 689027 997251 717600 1002315
rect 689027 997134 691527 997251
rect 689027 997051 689167 997134
rect 689027 967600 689167 996800
rect 689027 967266 689167 967407
rect 689247 967346 690137 997054
rect 690217 997051 690337 997134
rect 690217 967600 690337 996800
rect 690217 967266 690337 967407
rect 690417 967346 691307 997054
rect 691387 997051 691527 997134
rect 691387 967600 691527 996800
rect 691387 967266 691527 967407
rect 691607 967346 696600 997171
rect 696680 997134 717600 997251
rect 696680 997051 712677 997134
rect 712757 996800 717600 997054
rect 696680 967600 717600 996800
rect 696680 967266 712677 967407
rect 712757 967346 717600 967600
rect 689027 966998 717600 967266
rect 688901 960232 717600 966998
rect 687949 959928 717600 960232
rect 687949 957091 688145 959928
rect 687293 956787 688145 957091
rect 30533 869993 30673 870134
rect 30533 842266 30673 842407
rect 30753 842346 31683 870054
rect 31763 869993 31883 870134
rect 31763 842266 31883 842407
rect 31963 842346 32653 870054
rect 32733 869993 32853 870134
rect 32733 842266 32853 842407
rect 32933 842346 33623 870054
rect 33703 869993 33823 870134
rect 33703 842266 33823 842407
rect 33903 842346 34833 870054
rect 34913 869993 35033 870134
rect 36123 870073 37213 870134
rect 34913 842266 35033 842407
rect 35113 842346 36043 870054
rect 36123 869993 36243 870073
rect 37093 869993 37213 870073
rect 36323 842407 37013 869993
rect 36123 842327 36243 842407
rect 37093 842327 37213 842407
rect 37293 842346 38223 870054
rect 38303 869993 38423 870134
rect 36123 842266 37213 842327
rect 38303 842266 38423 842407
rect 38503 842346 39593 870054
rect 677707 869062 687193 877798
rect 677707 862734 687067 869062
rect 677707 862606 677927 862734
rect 30407 827934 39593 842266
rect 678007 833146 679097 862654
rect 679177 862606 679297 862734
rect 680387 862686 681477 862734
rect 679177 833066 679297 833207
rect 679377 833146 680307 862654
rect 680387 862606 680507 862686
rect 681357 862606 681477 862686
rect 680587 833207 681277 862606
rect 680387 833127 680507 833207
rect 681357 833127 681477 833207
rect 681557 833146 682487 862654
rect 682567 862606 682687 862734
rect 680387 833066 681477 833127
rect 682567 833066 682687 833207
rect 682767 833146 683697 862654
rect 683777 862606 683897 862734
rect 683777 833066 683897 833207
rect 683977 833146 684667 862654
rect 684747 862606 684867 862734
rect 684747 833066 684867 833207
rect 684947 833146 685637 862654
rect 685717 862606 685837 862734
rect 685717 833066 685837 833207
rect 685917 833146 686847 862654
rect 686927 862606 687067 862734
rect 686927 833066 687067 833207
rect 29455 794909 30307 795213
rect 29455 792072 29651 794909
rect 0 791768 29651 792072
rect 0 785002 28699 791768
rect 0 784734 28573 785002
rect 0 784400 4843 784654
rect 4923 784593 20920 784734
rect 0 757200 20920 784400
rect 0 756946 4843 757200
rect 4923 756866 20920 756994
rect 21000 756946 25993 784654
rect 26073 784593 26213 784734
rect 26073 757200 26213 784400
rect 26073 756866 26213 756994
rect 26293 756946 27183 784654
rect 27263 784593 27383 784734
rect 27263 757200 27383 784400
rect 27263 756866 27383 756994
rect 27463 756946 28353 784654
rect 28433 784593 28573 784734
rect 28433 757200 28573 784400
rect 28433 756866 28573 756994
rect 0 750538 28573 756866
rect 28653 750618 28719 784922
rect 0 748872 28699 750538
rect 28779 748952 29375 791688
rect 29455 784734 29651 791768
rect 29435 756946 29671 784654
rect 29455 752013 29651 756866
rect 29731 752093 30327 794829
rect 30387 793818 30453 827854
rect 30533 827793 30673 827934
rect 30533 800066 30673 800194
rect 30753 800146 31683 827854
rect 31763 827793 31883 827934
rect 31763 800066 31883 800194
rect 31963 800146 32653 827854
rect 32733 827793 32853 827934
rect 32733 800066 32853 800194
rect 32933 800146 33623 827854
rect 33703 827793 33823 827934
rect 33703 800066 33823 800194
rect 33903 800146 34833 827854
rect 34913 827793 35033 827934
rect 36123 827873 37213 827934
rect 34913 800066 35033 800194
rect 35113 800146 36043 827854
rect 36123 827793 36243 827873
rect 37093 827793 37213 827873
rect 36323 800194 37013 827793
rect 36123 800114 36243 800194
rect 37093 800114 37213 800194
rect 37293 800146 38223 827854
rect 38303 827793 38423 827934
rect 36123 800066 37213 800114
rect 38303 800066 38423 800194
rect 38503 800146 39593 827854
rect 678007 818734 687067 833066
rect 39673 800066 39893 800194
rect 30533 793738 39893 800066
rect 30407 785002 39893 793738
rect 29455 751709 30307 752013
rect 29455 748872 29651 751709
rect 0 748568 29651 748872
rect 0 741802 28699 748568
rect 0 741534 28573 741802
rect 0 741200 4843 741454
rect 4923 741393 20920 741534
rect 0 714000 20920 741200
rect 0 713746 4843 714000
rect 4923 713666 20920 713794
rect 21000 713746 25993 741454
rect 26073 741393 26213 741534
rect 26073 714000 26213 741200
rect 26073 713666 26213 713794
rect 26293 713746 27183 741454
rect 27263 741393 27383 741534
rect 27263 714000 27383 741200
rect 27263 713666 27383 713794
rect 27463 713746 28353 741454
rect 28433 741393 28573 741534
rect 28433 714000 28573 741200
rect 28433 713666 28573 713794
rect 0 707338 28573 713666
rect 28653 707418 28719 741722
rect 0 705672 28699 707338
rect 28779 705752 29375 748488
rect 29455 741534 29651 748568
rect 29435 713746 29671 741454
rect 29455 708813 29651 713666
rect 29731 708893 30327 751629
rect 30387 750618 30453 784922
rect 30533 784734 39893 785002
rect 30533 784593 30673 784734
rect 30533 756866 30673 756994
rect 30753 756946 31683 784654
rect 31763 784593 31883 784734
rect 31763 756866 31883 756994
rect 31963 756946 32653 784654
rect 32733 784593 32853 784734
rect 32733 756866 32853 756994
rect 32933 756946 33623 784654
rect 33703 784593 33823 784734
rect 33703 756866 33823 756994
rect 33903 756946 34833 784654
rect 34913 784593 35033 784734
rect 36123 784673 37213 784734
rect 34913 756866 35033 756994
rect 35113 756946 36043 784654
rect 36123 784593 36243 784673
rect 37093 784593 37213 784673
rect 36323 756994 37013 784593
rect 36123 756914 36243 756994
rect 37093 756914 37213 756994
rect 37293 756946 38223 784654
rect 38303 784593 38423 784734
rect 36123 756866 37213 756914
rect 38303 756866 38423 756994
rect 38503 756946 39593 784654
rect 39673 784593 39893 784734
rect 677707 788866 677927 789007
rect 678007 788946 679097 818654
rect 679177 818593 679297 818734
rect 680387 818673 681477 818734
rect 679177 788866 679297 789007
rect 679377 788946 680307 818654
rect 680387 818593 680507 818673
rect 681357 818593 681477 818673
rect 680587 789007 681277 818593
rect 680387 788927 680507 789007
rect 681357 788927 681477 789007
rect 681557 788946 682487 818654
rect 682567 818593 682687 818734
rect 680387 788866 681477 788927
rect 682567 788866 682687 789007
rect 682767 788946 683697 818654
rect 683777 818593 683897 818734
rect 683777 788866 683897 789007
rect 683977 788946 684667 818654
rect 684747 818593 684867 818734
rect 684747 788866 684867 789007
rect 684947 788946 685637 818654
rect 685717 818593 685837 818734
rect 685717 788866 685837 789007
rect 685917 788946 686847 818654
rect 686927 818593 687067 818734
rect 686927 788866 687067 789007
rect 677707 788598 687067 788866
rect 687147 788678 687213 868982
rect 687273 867971 687869 956707
rect 687949 951934 688145 956787
rect 687929 922346 688165 951854
rect 687949 907934 688145 922266
rect 687929 878146 688165 907854
rect 687949 871032 688145 878066
rect 688225 871112 688821 959848
rect 688901 958262 717600 959928
rect 688881 877878 688947 958182
rect 689027 951934 717600 958262
rect 689027 951806 689167 951934
rect 689027 922266 689167 951600
rect 689247 922346 690137 951854
rect 690217 951806 690337 951934
rect 690217 922266 690337 951600
rect 690417 922346 691307 951854
rect 691387 951806 691527 951934
rect 691387 922266 691527 951600
rect 691607 922346 696600 951854
rect 696680 951806 712677 951934
rect 712757 951600 717600 951854
rect 696680 922600 717600 951600
rect 696680 922266 712677 922600
rect 712757 922346 717600 922600
rect 689027 907934 717600 922266
rect 689027 878400 689167 907934
rect 689027 878066 689167 878207
rect 689247 878146 690137 907854
rect 690217 878400 690337 907934
rect 690217 878066 690337 878207
rect 690417 878146 691307 907854
rect 691387 878400 691527 907934
rect 691387 878066 691527 878207
rect 691607 878146 696600 907854
rect 696680 907600 712677 907934
rect 712757 907643 717600 907854
rect 712750 907600 717600 907643
rect 696680 878400 717600 907600
rect 696680 878066 712677 878207
rect 712757 878146 717600 878400
rect 689027 877798 717600 878066
rect 688901 871032 717600 877798
rect 687949 870728 717600 871032
rect 687949 867891 688145 870728
rect 687293 867587 688145 867891
rect 677707 779862 687193 788598
rect 677707 773534 687067 779862
rect 677707 773406 677927 773534
rect 39673 756866 39893 756994
rect 30533 750538 39893 756866
rect 30407 741802 39893 750538
rect 29455 708509 30307 708813
rect 29455 705672 29651 708509
rect 0 705368 29651 705672
rect 0 698602 28699 705368
rect 0 698334 28573 698602
rect 0 698000 4843 698254
rect 4923 698193 20920 698334
rect 0 670800 20920 698000
rect 0 670546 4843 670800
rect 4923 670466 20920 670594
rect 21000 670546 25993 698254
rect 26073 698193 26213 698334
rect 26073 670800 26213 698000
rect 26073 670466 26213 670594
rect 26293 670546 27183 698254
rect 27263 698193 27383 698334
rect 27263 670800 27383 698000
rect 27263 670466 27383 670594
rect 27463 670546 28353 698254
rect 28433 698193 28573 698334
rect 28433 670800 28573 698000
rect 28433 670466 28573 670594
rect 0 664138 28573 670466
rect 28653 664218 28719 698522
rect 0 662472 28699 664138
rect 28779 662552 29375 705288
rect 29455 698334 29651 705368
rect 29435 670546 29671 698254
rect 29455 665613 29651 670466
rect 29731 665693 30327 708429
rect 30387 707418 30453 741722
rect 30533 741534 39893 741802
rect 30533 741393 30673 741534
rect 30533 713666 30673 713794
rect 30753 713746 31683 741454
rect 31763 741393 31883 741534
rect 31763 713666 31883 713794
rect 31963 713746 32653 741454
rect 32733 741393 32853 741534
rect 32733 713666 32853 713794
rect 32933 713746 33623 741454
rect 33703 741393 33823 741534
rect 33703 713666 33823 713794
rect 33903 713746 34833 741454
rect 34913 741393 35033 741534
rect 36123 741473 37213 741534
rect 34913 713666 35033 713794
rect 35113 713746 36043 741454
rect 36123 741393 36243 741473
rect 37093 741393 37213 741473
rect 36323 713794 37013 741393
rect 36123 713714 36243 713794
rect 37093 713714 37213 713794
rect 37293 713746 38223 741454
rect 38303 741393 38423 741534
rect 36123 713666 37213 713714
rect 38303 713666 38423 713794
rect 38503 713746 39593 741454
rect 39673 741393 39893 741534
rect 677707 743866 677927 744007
rect 678007 743946 679097 773454
rect 679177 773406 679297 773534
rect 680387 773486 681477 773534
rect 679177 743866 679297 744007
rect 679377 743946 680307 773454
rect 680387 773406 680507 773486
rect 681357 773406 681477 773486
rect 680587 744007 681277 773406
rect 680387 743927 680507 744007
rect 681357 743927 681477 744007
rect 681557 743946 682487 773454
rect 682567 773406 682687 773534
rect 680387 743866 681477 743927
rect 682567 743866 682687 744007
rect 682767 743946 683697 773454
rect 683777 773406 683897 773534
rect 683777 743866 683897 744007
rect 683977 743946 684667 773454
rect 684747 773406 684867 773534
rect 684747 743866 684867 744007
rect 684947 743946 685637 773454
rect 685717 773406 685837 773534
rect 685717 743866 685837 744007
rect 685917 743946 686847 773454
rect 686927 773406 687067 773534
rect 686927 743866 687067 744007
rect 677707 743598 687067 743866
rect 687147 743678 687213 779782
rect 687273 778771 687869 867507
rect 687949 862734 688145 867587
rect 687929 833146 688165 862654
rect 687949 818734 688145 833066
rect 687929 788946 688165 818654
rect 687949 781832 688145 788866
rect 688225 781912 688821 870648
rect 688901 869062 717600 870728
rect 688881 788678 688947 868982
rect 689027 862734 717600 869062
rect 689027 862606 689167 862734
rect 689027 833400 689167 862400
rect 689027 833066 689167 833207
rect 689247 833146 690137 862654
rect 690217 862606 690337 862734
rect 690217 833400 690337 862400
rect 690217 833066 690337 833207
rect 690417 833146 691307 862654
rect 691387 862606 691527 862734
rect 691387 833400 691527 862400
rect 691387 833066 691527 833207
rect 691607 833146 696600 862654
rect 696680 862606 712677 862734
rect 712757 862400 717600 862654
rect 696680 833400 717600 862400
rect 696680 833066 712677 833207
rect 712757 833146 717600 833400
rect 689027 818734 717600 833066
rect 689027 818593 689167 818734
rect 689027 789200 689167 818400
rect 689027 788866 689167 789007
rect 689247 788946 690137 818654
rect 690217 818593 690337 818734
rect 690217 789200 690337 818400
rect 690217 788866 690337 789007
rect 690417 788946 691307 818654
rect 691387 818593 691527 818734
rect 691387 789200 691527 818400
rect 691387 788866 691527 789007
rect 691607 788946 696600 818654
rect 696680 818593 712677 818734
rect 712757 818400 717600 818654
rect 696680 789200 717600 818400
rect 696680 788866 712677 789007
rect 712757 788946 717600 789200
rect 689027 788598 717600 788866
rect 688901 781832 717600 788598
rect 687949 781528 717600 781832
rect 687949 778691 688145 781528
rect 687293 778387 688145 778691
rect 677707 734862 687193 743598
rect 677707 728534 687067 734862
rect 677707 728406 677927 728534
rect 39673 713666 39893 713794
rect 30533 707338 39893 713666
rect 30407 698602 39893 707338
rect 29455 665309 30307 665613
rect 29455 662472 29651 665309
rect 0 662168 29651 662472
rect 0 655402 28699 662168
rect 0 655134 28573 655402
rect 0 654800 4843 655054
rect 4923 654993 20920 655134
rect 0 627600 20920 654800
rect 0 627346 4843 627600
rect 4923 627266 20920 627394
rect 21000 627346 25993 655054
rect 26073 654993 26213 655134
rect 26073 627600 26213 654800
rect 26073 627266 26213 627394
rect 26293 627346 27183 655054
rect 27263 654993 27383 655134
rect 27263 627600 27383 654800
rect 27263 627266 27383 627394
rect 27463 627346 28353 655054
rect 28433 654993 28573 655134
rect 28433 627600 28573 654800
rect 28433 627266 28573 627394
rect 0 620938 28573 627266
rect 28653 621018 28719 655322
rect 0 619272 28699 620938
rect 28779 619352 29375 662088
rect 29455 655134 29651 662168
rect 29435 627346 29671 655054
rect 29455 622413 29651 627266
rect 29731 622493 30327 665229
rect 30387 664218 30453 698522
rect 30533 698334 39893 698602
rect 30533 698193 30673 698334
rect 30533 670466 30673 670594
rect 30753 670546 31683 698254
rect 31763 698193 31883 698334
rect 31763 670466 31883 670594
rect 31963 670546 32653 698254
rect 32733 698193 32853 698334
rect 32733 670466 32853 670594
rect 32933 670546 33623 698254
rect 33703 698193 33823 698334
rect 33703 670466 33823 670594
rect 33903 670546 34833 698254
rect 34913 698193 35033 698334
rect 36123 698273 37213 698334
rect 34913 670466 35033 670594
rect 35113 670546 36043 698254
rect 36123 698193 36243 698273
rect 37093 698193 37213 698273
rect 36323 670594 37013 698193
rect 36123 670514 36243 670594
rect 37093 670514 37213 670594
rect 37293 670546 38223 698254
rect 38303 698193 38423 698334
rect 36123 670466 37213 670514
rect 38303 670466 38423 670594
rect 38503 670546 39593 698254
rect 39673 698193 39893 698334
rect 677707 698866 677927 699007
rect 678007 698946 679097 728454
rect 679177 728406 679297 728534
rect 680387 728486 681477 728534
rect 679177 698866 679297 699007
rect 679377 698946 680307 728454
rect 680387 728406 680507 728486
rect 681357 728406 681477 728486
rect 680587 699007 681277 728406
rect 680387 698927 680507 699007
rect 681357 698927 681477 699007
rect 681557 698946 682487 728454
rect 682567 728406 682687 728534
rect 680387 698866 681477 698927
rect 682567 698866 682687 699007
rect 682767 698946 683697 728454
rect 683777 728406 683897 728534
rect 683777 698866 683897 699007
rect 683977 698946 684667 728454
rect 684747 728406 684867 728534
rect 684747 698866 684867 699007
rect 684947 698946 685637 728454
rect 685717 728406 685837 728534
rect 685717 698866 685837 699007
rect 685917 698946 686847 728454
rect 686927 728406 687067 728534
rect 686927 698866 687067 699007
rect 677707 698598 687067 698866
rect 687147 698678 687213 734782
rect 687273 733771 687869 778307
rect 687949 773534 688145 778387
rect 687929 743946 688165 773454
rect 687949 736832 688145 743866
rect 688225 736912 688821 781448
rect 688901 779862 717600 781528
rect 688881 743678 688947 779782
rect 689027 773534 717600 779862
rect 689027 773406 689167 773534
rect 689027 744200 689167 773200
rect 689027 743866 689167 744007
rect 689247 743946 690137 773454
rect 690217 773406 690337 773534
rect 690217 744200 690337 773200
rect 690217 743866 690337 744007
rect 690417 743946 691307 773454
rect 691387 773406 691527 773534
rect 691387 744200 691527 773200
rect 691387 743866 691527 744007
rect 691607 743946 696600 773454
rect 696680 773406 712677 773534
rect 712757 773200 717600 773454
rect 696680 744200 717600 773200
rect 696680 743866 712677 744007
rect 712757 743946 717600 744200
rect 689027 743598 717600 743866
rect 688901 736832 717600 743598
rect 687949 736528 717600 736832
rect 687949 733691 688145 736528
rect 687293 733387 688145 733691
rect 677707 689862 687193 698598
rect 677707 683534 687067 689862
rect 677707 683406 677927 683534
rect 39673 670466 39893 670594
rect 30533 664138 39893 670466
rect 30407 655402 39893 664138
rect 29455 622109 30307 622413
rect 29455 619272 29651 622109
rect 0 618968 29651 619272
rect 0 612202 28699 618968
rect 0 611934 28573 612202
rect 0 611600 4843 611854
rect 4923 611793 20920 611934
rect 0 584400 20920 611600
rect 0 584146 4843 584400
rect 4923 584066 20920 584194
rect 21000 584146 25993 611854
rect 26073 611793 26213 611934
rect 26073 584400 26213 611600
rect 26073 584066 26213 584194
rect 26293 584146 27183 611854
rect 27263 611793 27383 611934
rect 27263 584400 27383 611600
rect 27263 584066 27383 584194
rect 27463 584146 28353 611854
rect 28433 611793 28573 611934
rect 28433 584400 28573 611600
rect 28433 584066 28573 584194
rect 0 577738 28573 584066
rect 28653 577818 28719 612122
rect 0 576072 28699 577738
rect 28779 576152 29375 618888
rect 29455 611934 29651 618968
rect 29435 584146 29671 611854
rect 29455 579213 29651 584066
rect 29731 579293 30327 622029
rect 30387 621018 30453 655322
rect 30533 655134 39893 655402
rect 30533 654993 30673 655134
rect 30533 627266 30673 627394
rect 30753 627346 31683 655054
rect 31763 654993 31883 655134
rect 31763 627266 31883 627394
rect 31963 627346 32653 655054
rect 32733 654993 32853 655134
rect 32733 627266 32853 627394
rect 32933 627346 33623 655054
rect 33703 654993 33823 655134
rect 33703 627266 33823 627394
rect 33903 627346 34833 655054
rect 34913 654993 35033 655134
rect 36123 655073 37213 655134
rect 34913 627266 35033 627394
rect 35113 627346 36043 655054
rect 36123 654993 36243 655073
rect 37093 654993 37213 655073
rect 36323 627394 37013 654993
rect 36123 627314 36243 627394
rect 37093 627314 37213 627394
rect 37293 627346 38223 655054
rect 38303 654993 38423 655134
rect 36123 627266 37213 627314
rect 38303 627266 38423 627394
rect 38503 627346 39593 655054
rect 39673 654993 39893 655134
rect 677707 653666 677927 653807
rect 678007 653746 679097 683454
rect 679177 683406 679297 683534
rect 680387 683486 681477 683534
rect 679177 653666 679297 653807
rect 679377 653746 680307 683454
rect 680387 683406 680507 683486
rect 681357 683406 681477 683486
rect 680587 653807 681277 683406
rect 680387 653727 680507 653807
rect 681357 653727 681477 653807
rect 681557 653746 682487 683454
rect 682567 683406 682687 683534
rect 680387 653666 681477 653727
rect 682567 653666 682687 653807
rect 682767 653746 683697 683454
rect 683777 683406 683897 683534
rect 683777 653666 683897 653807
rect 683977 653746 684667 683454
rect 684747 683406 684867 683534
rect 684747 653666 684867 653807
rect 684947 653746 685637 683454
rect 685717 683406 685837 683534
rect 685717 653666 685837 653807
rect 685917 653746 686847 683454
rect 686927 683406 687067 683534
rect 686927 653666 687067 653807
rect 677707 653398 687067 653666
rect 687147 653478 687213 689782
rect 687273 688771 687869 733307
rect 687949 728534 688145 733387
rect 687929 698946 688165 728454
rect 687949 691832 688145 698866
rect 688225 691912 688821 736448
rect 688901 734862 717600 736528
rect 688881 698678 688947 734782
rect 689027 728534 717600 734862
rect 689027 728406 689167 728534
rect 689027 699200 689167 728200
rect 689027 698866 689167 699007
rect 689247 698946 690137 728454
rect 690217 728406 690337 728534
rect 690217 699200 690337 728200
rect 690217 698866 690337 699007
rect 690417 698946 691307 728454
rect 691387 728406 691527 728534
rect 691387 699200 691527 728200
rect 691387 698866 691527 699007
rect 691607 698946 696600 728454
rect 696680 728406 712677 728534
rect 712757 728200 717600 728454
rect 696680 699200 717600 728200
rect 696680 698866 712677 699007
rect 712757 698946 717600 699200
rect 689027 698598 717600 698866
rect 688901 691832 717600 698598
rect 687949 691528 717600 691832
rect 687949 688691 688145 691528
rect 687293 688387 688145 688691
rect 677707 644662 687193 653398
rect 677707 638334 687067 644662
rect 677707 638206 677927 638334
rect 39673 627266 39893 627394
rect 30533 620938 39893 627266
rect 30407 612202 39893 620938
rect 29455 578909 30307 579213
rect 29455 576072 29651 578909
rect 0 575768 29651 576072
rect 0 569002 28699 575768
rect 0 568734 28573 569002
rect 0 568400 4843 568654
rect 4923 568593 20920 568734
rect 0 541200 20920 568400
rect 0 540946 4843 541200
rect 4923 540866 20920 540994
rect 21000 540946 25993 568654
rect 26073 568593 26213 568734
rect 26073 541200 26213 568400
rect 26073 540866 26213 540994
rect 26293 540946 27183 568654
rect 27263 568593 27383 568734
rect 27263 541200 27383 568400
rect 27263 540866 27383 540994
rect 27463 540946 28353 568654
rect 28433 568593 28573 568734
rect 28433 541200 28573 568400
rect 28433 540866 28573 540994
rect 0 534538 28573 540866
rect 28653 534618 28719 568922
rect 0 532872 28699 534538
rect 28779 532952 29375 575688
rect 29455 568734 29651 575768
rect 29435 540946 29671 568654
rect 29455 536013 29651 540866
rect 29731 536093 30327 578829
rect 30387 577818 30453 612122
rect 30533 611934 39893 612202
rect 30533 611793 30673 611934
rect 30533 584066 30673 584194
rect 30753 584146 31683 611854
rect 31763 611793 31883 611934
rect 31763 584066 31883 584194
rect 31963 584146 32653 611854
rect 32733 611793 32853 611934
rect 32733 584066 32853 584194
rect 32933 584146 33623 611854
rect 33703 611793 33823 611934
rect 33703 584066 33823 584194
rect 33903 584146 34833 611854
rect 34913 611793 35033 611934
rect 36123 611873 37213 611934
rect 34913 584066 35033 584194
rect 35113 584146 36043 611854
rect 36123 611793 36243 611873
rect 37093 611793 37213 611873
rect 36323 584194 37013 611793
rect 36123 584114 36243 584194
rect 37093 584114 37213 584194
rect 37293 584146 38223 611854
rect 38303 611793 38423 611934
rect 36123 584066 37213 584114
rect 38303 584066 38423 584194
rect 38503 584146 39593 611854
rect 39673 611793 39893 611934
rect 677707 608666 677927 608807
rect 678007 608746 679097 638254
rect 679177 638206 679297 638334
rect 680387 638286 681477 638334
rect 679177 608666 679297 608807
rect 679377 608746 680307 638254
rect 680387 638206 680507 638286
rect 681357 638206 681477 638286
rect 680587 608807 681277 638206
rect 680387 608727 680507 608807
rect 681357 608727 681477 608807
rect 681557 608746 682487 638254
rect 682567 638206 682687 638334
rect 680387 608666 681477 608727
rect 682567 608666 682687 608807
rect 682767 608746 683697 638254
rect 683777 638206 683897 638334
rect 683777 608666 683897 608807
rect 683977 608746 684667 638254
rect 684747 638206 684867 638334
rect 684747 608666 684867 608807
rect 684947 608746 685637 638254
rect 685717 638206 685837 638334
rect 685717 608666 685837 608807
rect 685917 608746 686847 638254
rect 686927 638206 687067 638334
rect 686927 608666 687067 608807
rect 677707 608398 687067 608666
rect 687147 608478 687213 644582
rect 687273 643571 687869 688307
rect 687949 683534 688145 688387
rect 687929 653746 688165 683454
rect 687949 646632 688145 653666
rect 688225 646712 688821 691448
rect 688901 689862 717600 691528
rect 688881 653478 688947 689782
rect 689027 683534 717600 689862
rect 689027 683406 689167 683534
rect 689027 654000 689167 683200
rect 689027 653666 689167 653807
rect 689247 653746 690137 683454
rect 690217 683406 690337 683534
rect 690217 654000 690337 683200
rect 690217 653666 690337 653807
rect 690417 653746 691307 683454
rect 691387 683406 691527 683534
rect 691387 654000 691527 683200
rect 691387 653666 691527 653807
rect 691607 653746 696600 683454
rect 696680 683406 712677 683534
rect 712757 683200 717600 683454
rect 696680 654000 717600 683200
rect 696680 653666 712677 653807
rect 712757 653746 717600 654000
rect 689027 653398 717600 653666
rect 688901 646632 717600 653398
rect 687949 646328 717600 646632
rect 687949 643491 688145 646328
rect 687293 643187 688145 643491
rect 677707 599662 687193 608398
rect 677707 593334 687067 599662
rect 677707 593206 677927 593334
rect 39673 584066 39893 584194
rect 30533 577738 39893 584066
rect 30407 569002 39893 577738
rect 29455 535709 30307 536013
rect 29455 532872 29651 535709
rect 0 532568 29651 532872
rect 0 525802 28699 532568
rect 0 525534 28573 525802
rect 0 525200 4843 525454
rect 4923 525393 20920 525534
rect 0 498000 20920 525200
rect 0 497746 4843 498000
rect 4923 497666 20920 497807
rect 21000 497746 25993 525454
rect 26073 525393 26213 525534
rect 26073 498000 26213 525200
rect 26073 497666 26213 497807
rect 26293 497746 27183 525454
rect 27263 525393 27383 525534
rect 27263 498000 27383 525200
rect 27263 497666 27383 497807
rect 27463 497746 28353 525454
rect 28433 525393 28573 525534
rect 28433 498000 28573 525200
rect 28433 497666 28573 497807
rect 0 483334 28573 497666
rect 0 483000 4843 483254
rect 4923 483193 20920 483334
rect 0 456094 20920 483000
rect 0 455800 7 456094
rect 4843 455800 20920 456094
rect 4843 455757 4850 455800
rect 4923 455466 20920 455800
rect 21000 455546 25993 483254
rect 26073 483193 26213 483334
rect 26073 455466 26213 483000
rect 26293 455546 27183 483254
rect 27263 483193 27383 483334
rect 27263 455466 27383 483000
rect 27463 455546 28353 483254
rect 28433 483193 28573 483334
rect 28433 455466 28573 483000
rect 0 441134 28573 455466
rect 0 440800 4843 441054
rect 4923 440800 20920 441134
rect 0 413600 20920 440800
rect 0 413346 4843 413600
rect 4923 413266 20920 413394
rect 21000 413346 25993 441054
rect 26073 413600 26213 441134
rect 26073 413266 26213 413394
rect 26293 413346 27183 441054
rect 27263 413600 27383 441134
rect 27263 413266 27383 413394
rect 27463 413346 28353 441054
rect 28433 413600 28573 441134
rect 28433 413266 28573 413394
rect 0 406938 28573 413266
rect 0 405272 28699 406938
rect 28779 405352 29375 532488
rect 29455 525534 29651 532568
rect 29435 497746 29671 525454
rect 29455 483334 29651 497666
rect 29435 455546 29671 483254
rect 29455 441134 29651 455466
rect 29435 413346 29671 441054
rect 29455 408413 29651 413266
rect 29731 408493 30327 535629
rect 30387 534618 30453 568922
rect 30533 568734 39893 569002
rect 30533 568593 30673 568734
rect 30533 540866 30673 540994
rect 30753 540946 31683 568654
rect 31763 568593 31883 568734
rect 31763 540866 31883 540994
rect 31963 540946 32653 568654
rect 32733 568593 32853 568734
rect 32733 540866 32853 540994
rect 32933 540946 33623 568654
rect 33703 568593 33823 568734
rect 33703 540866 33823 540994
rect 33903 540946 34833 568654
rect 34913 568593 35033 568734
rect 36123 568673 37213 568734
rect 34913 540866 35033 540994
rect 35113 540946 36043 568654
rect 36123 568593 36243 568673
rect 37093 568593 37213 568673
rect 36323 540994 37013 568593
rect 36123 540914 36243 540994
rect 37093 540914 37213 540994
rect 37293 540946 38223 568654
rect 38303 568593 38423 568734
rect 36123 540866 37213 540914
rect 38303 540866 38423 540994
rect 38503 540946 39593 568654
rect 39673 568593 39893 568734
rect 677707 563466 677927 563607
rect 678007 563546 679097 593254
rect 679177 593206 679297 593334
rect 680387 593286 681477 593334
rect 679177 563466 679297 563607
rect 679377 563546 680307 593254
rect 680387 593206 680507 593286
rect 681357 593206 681477 593286
rect 680587 563607 681277 593206
rect 680387 563527 680507 563607
rect 681357 563527 681477 563607
rect 681557 563546 682487 593254
rect 682567 593206 682687 593334
rect 680387 563466 681477 563527
rect 682567 563466 682687 563607
rect 682767 563546 683697 593254
rect 683777 593206 683897 593334
rect 683777 563466 683897 563607
rect 683977 563546 684667 593254
rect 684747 593206 684867 593334
rect 684747 563466 684867 563607
rect 684947 563546 685637 593254
rect 685717 593206 685837 593334
rect 685717 563466 685837 563607
rect 685917 563546 686847 593254
rect 686927 593206 687067 593334
rect 686927 563466 687067 563607
rect 677707 563198 687067 563466
rect 687147 563278 687213 599582
rect 687273 598571 687869 643107
rect 687949 638334 688145 643187
rect 687929 608746 688165 638254
rect 687949 601632 688145 608666
rect 688225 601712 688821 646248
rect 688901 644662 717600 646328
rect 688881 608478 688947 644582
rect 689027 638334 717600 644662
rect 689027 638206 689167 638334
rect 689027 609000 689167 638000
rect 689027 608666 689167 608807
rect 689247 608746 690137 638254
rect 690217 638206 690337 638334
rect 690217 609000 690337 638000
rect 690217 608666 690337 608807
rect 690417 608746 691307 638254
rect 691387 638206 691527 638334
rect 691387 609000 691527 638000
rect 691387 608666 691527 608807
rect 691607 608746 696600 638254
rect 696680 638206 712677 638334
rect 712757 638000 717600 638254
rect 696680 609000 717600 638000
rect 696680 608666 712677 608807
rect 712757 608746 717600 609000
rect 689027 608398 717600 608666
rect 688901 601632 717600 608398
rect 687949 601328 717600 601632
rect 687949 598491 688145 601328
rect 687293 598187 688145 598491
rect 677707 554462 687193 563198
rect 677707 548134 687067 554462
rect 677707 548006 677927 548134
rect 39673 540866 39893 540994
rect 30533 534538 39893 540866
rect 30407 525802 39893 534538
rect 29455 408109 30307 408413
rect 29455 405272 29651 408109
rect 0 404968 29651 405272
rect 0 398202 28699 404968
rect 0 397934 28573 398202
rect 0 397600 4843 397854
rect 4923 397793 20920 397934
rect 0 370400 20920 397600
rect 0 370146 4843 370400
rect 4923 370066 20920 370194
rect 21000 370146 25993 397854
rect 26073 397793 26213 397934
rect 26073 370400 26213 397600
rect 26073 370066 26213 370194
rect 26293 370146 27183 397854
rect 27263 397793 27383 397934
rect 27263 370400 27383 397600
rect 27263 370066 27383 370194
rect 27463 370146 28353 397854
rect 28433 397793 28573 397934
rect 28433 370400 28573 397600
rect 28433 370066 28573 370194
rect 0 363738 28573 370066
rect 28653 363818 28719 398122
rect 0 362072 28699 363738
rect 28779 362152 29375 404888
rect 29455 397934 29651 404968
rect 29435 370146 29671 397854
rect 29455 365213 29651 370066
rect 29731 365293 30327 408029
rect 30387 407018 30453 525722
rect 30533 525534 39893 525802
rect 30533 525393 30673 525534
rect 30533 497666 30673 497807
rect 30753 497746 31683 525454
rect 31763 525393 31883 525534
rect 31763 497666 31883 497807
rect 31963 497746 32653 525454
rect 32733 525393 32853 525534
rect 32733 497666 32853 497807
rect 32933 497746 33623 525454
rect 33703 525393 33823 525534
rect 33703 497666 33823 497807
rect 33903 497746 34833 525454
rect 34913 525393 35033 525534
rect 36123 525473 37213 525534
rect 34913 497666 35033 497807
rect 35113 497746 36043 525454
rect 36123 525393 36243 525473
rect 37093 525393 37213 525473
rect 36323 497807 37013 525393
rect 36123 497727 36243 497807
rect 37093 497727 37213 497807
rect 37293 497746 38223 525454
rect 38303 525393 38423 525534
rect 36123 497666 37213 497727
rect 38303 497666 38423 497807
rect 38503 497746 39593 525454
rect 39673 525393 39893 525534
rect 678007 518546 679097 548054
rect 679177 548006 679297 548134
rect 680387 548086 681477 548134
rect 679177 518466 679297 518607
rect 679377 518546 680307 548054
rect 680387 548006 680507 548086
rect 681357 548006 681477 548086
rect 680587 518607 681277 548006
rect 680387 518527 680507 518607
rect 681357 518527 681477 518607
rect 681557 518546 682487 548054
rect 682567 548006 682687 548134
rect 680387 518466 681477 518527
rect 682567 518466 682687 518607
rect 682767 518546 683697 548054
rect 683777 548006 683897 548134
rect 683777 518466 683897 518607
rect 683977 518546 684667 548054
rect 684747 548006 684867 548134
rect 684747 518466 684867 518607
rect 684947 518546 685637 548054
rect 685717 548006 685837 548134
rect 685717 518466 685837 518607
rect 685917 518546 686847 548054
rect 686927 548006 687067 548134
rect 686927 518466 687067 518607
rect 678007 504134 687067 518466
rect 30533 483334 39593 497666
rect 30533 483193 30673 483334
rect 30533 455466 30673 455800
rect 30753 455546 31683 483254
rect 31763 483193 31883 483334
rect 31763 455466 31883 455800
rect 31963 455546 32653 483254
rect 32733 483193 32853 483334
rect 32733 455466 32853 455800
rect 33703 483193 33823 483334
rect 33903 457987 34833 483254
rect 34913 483193 35033 483334
rect 36123 483273 37213 483334
rect 33703 455466 33823 455800
rect 33903 455787 34840 457987
rect 33903 455546 34833 455787
rect 34913 455466 35033 455800
rect 35113 455546 36043 483254
rect 36123 483193 36243 483273
rect 37093 483193 37213 483273
rect 36123 455527 36243 455800
rect 37093 455527 37213 455800
rect 38303 483193 38423 483334
rect 36123 455466 37213 455527
rect 38303 455466 38423 455800
rect 678007 474546 679097 504054
rect 679177 503993 679297 504134
rect 680387 504073 681477 504134
rect 679177 474466 679297 474800
rect 679377 474546 680307 504054
rect 680387 503993 680507 504073
rect 681357 503993 681477 504073
rect 680387 474527 680507 474800
rect 680587 474607 681277 503993
rect 681357 474527 681477 474800
rect 681557 474546 682487 504054
rect 682567 503993 682687 504134
rect 680387 474466 681477 474527
rect 682567 474466 682687 474800
rect 682767 474546 683697 504054
rect 683777 503993 683897 504134
rect 683777 474466 683897 474800
rect 683977 474546 684667 504054
rect 684747 503993 684867 504134
rect 684747 474466 684867 474800
rect 684947 474546 685637 504054
rect 685717 503993 685837 504134
rect 685917 476995 686847 504054
rect 686927 503993 687067 504134
rect 685717 474466 685837 474800
rect 685910 474786 686847 476995
rect 685917 474546 686847 474786
rect 686927 474466 687067 474800
rect 678007 460134 687067 474466
rect 30533 441134 39593 455466
rect 30533 440800 30673 441134
rect 30753 440814 31683 441054
rect 30753 438605 31690 440814
rect 31763 440800 31883 441134
rect 30533 413266 30673 413394
rect 30753 413346 31683 438605
rect 31763 413266 31883 413394
rect 31963 413346 32653 441054
rect 32733 440800 32853 441134
rect 32733 413266 32853 413394
rect 32933 413346 33623 441054
rect 33703 440800 33823 441134
rect 33703 413266 33823 413394
rect 33903 413346 34833 441054
rect 34913 440800 35033 441134
rect 36123 441073 37213 441134
rect 34913 413266 35033 413394
rect 35113 413346 36043 441054
rect 36123 440800 36243 441073
rect 36323 413394 37013 440993
rect 37093 440800 37213 441073
rect 36123 413314 36243 413394
rect 37093 413314 37213 413394
rect 37293 413346 38223 441054
rect 38303 440800 38423 441134
rect 36123 413266 37213 413314
rect 38303 413266 38423 413394
rect 38503 413346 39593 441054
rect 678007 430346 679097 460054
rect 679177 459800 679297 460134
rect 680387 460073 681477 460134
rect 679177 430266 679297 430407
rect 680387 459800 680507 460073
rect 681357 459800 681477 460073
rect 680387 430327 680507 430407
rect 681357 430327 681477 430407
rect 681557 430346 682487 460054
rect 682567 459800 682687 460134
rect 682767 459813 683697 460054
rect 682760 457613 683697 459813
rect 683777 459800 683897 460134
rect 680387 430266 681477 430327
rect 682567 430266 682687 430407
rect 682767 430346 683697 457613
rect 683777 430266 683897 430407
rect 683977 430346 684667 460054
rect 684747 459800 684867 460134
rect 684747 430266 684867 430407
rect 684947 430346 685637 460054
rect 685717 459800 685837 460134
rect 685717 430266 685837 430407
rect 685917 430346 686847 460054
rect 686927 459800 687067 460134
rect 686927 430266 687067 430407
rect 687147 430346 687213 554382
rect 687273 553371 687869 598107
rect 687949 593334 688145 598187
rect 687929 563546 688165 593254
rect 687949 556432 688145 563466
rect 688225 556512 688821 601248
rect 688901 599662 717600 601328
rect 688881 563278 688947 599582
rect 689027 593334 717600 599662
rect 689027 593206 689167 593334
rect 689027 563800 689167 593000
rect 689027 563466 689167 563607
rect 689247 563546 690137 593254
rect 690217 593206 690337 593334
rect 690217 563800 690337 593000
rect 690217 563466 690337 563607
rect 690417 563546 691307 593254
rect 691387 593206 691527 593334
rect 691387 563800 691527 593000
rect 691387 563466 691527 563607
rect 691607 563546 696600 593254
rect 696680 593206 712677 593334
rect 712757 593000 717600 593254
rect 696680 563800 717600 593000
rect 696680 563466 712677 563607
rect 712757 563546 717600 563800
rect 689027 563198 717600 563466
rect 688901 556432 717600 563198
rect 687949 556128 717600 556432
rect 687949 553291 688145 556128
rect 687293 552987 688145 553291
rect 678007 415934 687193 430266
rect 39673 413266 39893 413394
rect 30533 406938 39893 413266
rect 30407 398202 39893 406938
rect 29455 364909 30307 365213
rect 29455 362072 29651 364909
rect 0 361768 29651 362072
rect 0 355002 28699 361768
rect 0 354734 28573 355002
rect 0 354400 4843 354654
rect 4923 354593 20920 354734
rect 0 327200 20920 354400
rect 0 326946 4843 327200
rect 4923 326866 20920 326994
rect 21000 326946 25993 354654
rect 26073 354593 26213 354734
rect 26073 327200 26213 354400
rect 26073 326866 26213 326994
rect 26293 326946 27183 354654
rect 27263 354593 27383 354734
rect 27263 327200 27383 354400
rect 27263 326866 27383 326994
rect 27463 326946 28353 354654
rect 28433 354593 28573 354734
rect 28433 327200 28573 354400
rect 28433 326866 28573 326994
rect 0 320538 28573 326866
rect 28653 320618 28719 354922
rect 0 318872 28699 320538
rect 28779 318952 29375 361688
rect 29455 354734 29651 361768
rect 29435 326946 29671 354654
rect 29455 322013 29651 326866
rect 29731 322093 30327 364829
rect 30387 363818 30453 398122
rect 30533 397934 39893 398202
rect 30533 397793 30673 397934
rect 30533 370066 30673 370194
rect 30753 370146 31683 397854
rect 31763 397793 31883 397934
rect 31763 370066 31883 370194
rect 31963 370146 32653 397854
rect 32733 397793 32853 397934
rect 32733 370066 32853 370194
rect 32933 370146 33623 397854
rect 33703 397793 33823 397934
rect 33703 370066 33823 370194
rect 33903 370146 34833 397854
rect 34913 397793 35033 397934
rect 36123 397873 37213 397934
rect 34913 370066 35033 370194
rect 35113 370146 36043 397854
rect 36123 397793 36243 397873
rect 37093 397793 37213 397873
rect 36323 370194 37013 397793
rect 36123 370114 36243 370194
rect 37093 370114 37213 370194
rect 37293 370146 38223 397854
rect 38303 397793 38423 397934
rect 36123 370066 37213 370114
rect 38303 370066 38423 370194
rect 38503 370146 39593 397854
rect 39673 397793 39893 397934
rect 677707 386266 677927 386407
rect 678007 386346 679097 415854
rect 679177 415793 679297 415934
rect 680387 415873 681477 415934
rect 679177 386266 679297 386407
rect 679377 386346 680307 415854
rect 680387 415793 680507 415873
rect 681357 415793 681477 415873
rect 680587 386407 681277 415793
rect 680387 386327 680507 386407
rect 681357 386327 681477 386407
rect 681557 386346 682487 415854
rect 682567 415793 682687 415934
rect 680387 386266 681477 386327
rect 682567 386266 682687 386407
rect 682767 386346 683697 415854
rect 683777 415793 683897 415934
rect 683777 386266 683897 386407
rect 683977 386346 684667 415854
rect 684747 415793 684867 415934
rect 684747 386266 684867 386407
rect 684947 386346 685637 415854
rect 685717 415793 685837 415934
rect 685717 386266 685837 386407
rect 685917 386346 686847 415854
rect 686927 415793 687067 415934
rect 686927 386266 687067 386407
rect 677707 385998 687067 386266
rect 687147 386078 687213 415854
rect 677707 377262 687193 385998
rect 677707 370934 687067 377262
rect 677707 370806 677927 370934
rect 39673 370066 39893 370194
rect 30533 363738 39893 370066
rect 30407 355002 39893 363738
rect 29455 321709 30307 322013
rect 29455 318872 29651 321709
rect 0 318568 29651 318872
rect 0 311802 28699 318568
rect 0 311534 28573 311802
rect 0 311200 4843 311454
rect 4923 311393 20920 311534
rect 0 284000 20920 311200
rect 0 283746 4843 284000
rect 4923 283666 20920 283794
rect 21000 283746 25993 311454
rect 26073 311393 26213 311534
rect 26073 284000 26213 311200
rect 26073 283666 26213 283794
rect 26293 283746 27183 311454
rect 27263 311393 27383 311534
rect 27263 284000 27383 311200
rect 27263 283666 27383 283794
rect 27463 283746 28353 311454
rect 28433 311393 28573 311534
rect 28433 284000 28573 311200
rect 28433 283666 28573 283794
rect 0 277338 28573 283666
rect 28653 277418 28719 311722
rect 0 275672 28699 277338
rect 28779 275752 29375 318488
rect 29455 311534 29651 318568
rect 29435 283746 29671 311454
rect 29455 278813 29651 283666
rect 29731 278893 30327 321629
rect 30387 320618 30453 354922
rect 30533 354734 39893 355002
rect 30533 354593 30673 354734
rect 30533 326866 30673 326994
rect 30753 326946 31683 354654
rect 31763 354593 31883 354734
rect 31763 326866 31883 326994
rect 31963 326946 32653 354654
rect 32733 354593 32853 354734
rect 32733 326866 32853 326994
rect 32933 326946 33623 354654
rect 33703 354593 33823 354734
rect 33703 326866 33823 326994
rect 33903 326946 34833 354654
rect 34913 354593 35033 354734
rect 36123 354673 37213 354734
rect 34913 326866 35033 326994
rect 35113 326946 36043 354654
rect 36123 354593 36243 354673
rect 37093 354593 37213 354673
rect 36323 326994 37013 354593
rect 36123 326914 36243 326994
rect 37093 326914 37213 326994
rect 37293 326946 38223 354654
rect 38303 354593 38423 354734
rect 36123 326866 37213 326914
rect 38303 326866 38423 326994
rect 38503 326946 39593 354654
rect 39673 354593 39893 354734
rect 677707 341066 677927 341207
rect 678007 341146 679097 370854
rect 679177 370806 679297 370934
rect 680387 370886 681477 370934
rect 679177 341066 679297 341207
rect 679377 341146 680307 370854
rect 680387 370806 680507 370886
rect 681357 370806 681477 370886
rect 680587 341207 681277 370806
rect 680387 341127 680507 341207
rect 681357 341127 681477 341207
rect 681557 341146 682487 370854
rect 682567 370806 682687 370934
rect 680387 341066 681477 341127
rect 682567 341066 682687 341207
rect 682767 341146 683697 370854
rect 683777 370806 683897 370934
rect 683777 341066 683897 341207
rect 683977 341146 684667 370854
rect 684747 370806 684867 370934
rect 684747 341066 684867 341207
rect 684947 341146 685637 370854
rect 685717 370806 685837 370934
rect 685717 341066 685837 341207
rect 685917 341146 686847 370854
rect 686927 370806 687067 370934
rect 686927 341066 687067 341207
rect 677707 340798 687067 341066
rect 687147 340878 687213 377182
rect 687273 376171 687869 552907
rect 687949 548134 688145 552987
rect 687929 518546 688165 548054
rect 687949 504134 688145 518466
rect 687929 474546 688165 504054
rect 687949 460134 688145 474466
rect 687929 430346 688165 460054
rect 687949 415934 688145 430266
rect 687929 386346 688165 415854
rect 687949 379232 688145 386266
rect 688225 379312 688821 556048
rect 688901 554462 717600 556128
rect 689027 548134 717600 554462
rect 689027 548006 689167 548134
rect 689027 518800 689167 547800
rect 689027 518466 689167 518607
rect 689247 518546 690137 548054
rect 690217 548006 690337 548134
rect 690217 518800 690337 547800
rect 690217 518466 690337 518607
rect 690417 518546 691307 548054
rect 691387 548006 691527 548134
rect 691387 518800 691527 547800
rect 691387 518466 691527 518607
rect 691607 518546 696600 548054
rect 696680 548006 712677 548134
rect 712757 547800 717600 548054
rect 696680 518800 717600 547800
rect 696680 518466 712677 518607
rect 712757 518546 717600 518800
rect 689027 504134 717600 518466
rect 689027 503993 689167 504134
rect 689027 474466 689167 503800
rect 689247 474546 690137 504054
rect 690217 503993 690337 504134
rect 690217 474466 690337 503800
rect 690417 474546 691307 504054
rect 691387 503993 691527 504134
rect 691387 474466 691527 503800
rect 691607 474546 696600 504054
rect 696680 503993 712677 504134
rect 712757 503800 717600 504054
rect 696680 474800 717600 503800
rect 696680 474466 712677 474800
rect 712757 474546 717600 474800
rect 689027 460134 717600 474466
rect 689027 430600 689167 460134
rect 689027 430266 689167 430407
rect 689247 430346 690137 460054
rect 690217 430600 690337 460134
rect 690217 430266 690337 430407
rect 690417 430346 691307 460054
rect 691387 430600 691527 460134
rect 691387 430266 691527 430407
rect 691607 430346 696600 460054
rect 696680 459800 712677 460134
rect 712757 459843 717600 460054
rect 712750 459800 717600 459843
rect 696680 430600 717600 459800
rect 696680 430266 712677 430407
rect 712757 430346 717600 430600
rect 688901 415934 717600 430266
rect 688881 386078 688947 415854
rect 689027 415793 689167 415934
rect 689027 386600 689167 415600
rect 689027 386266 689167 386407
rect 689247 386346 690137 415854
rect 690217 415793 690337 415934
rect 690217 386600 690337 415600
rect 690217 386266 690337 386407
rect 690417 386346 691307 415854
rect 691387 415793 691527 415934
rect 691387 386600 691527 415600
rect 691387 386266 691527 386407
rect 691607 386346 696600 415854
rect 696680 415793 712677 415934
rect 712757 415600 717600 415854
rect 696680 386600 717600 415600
rect 696680 386266 712677 386407
rect 712757 386346 717600 386600
rect 689027 385998 717600 386266
rect 688901 379232 717600 385998
rect 687949 378928 717600 379232
rect 687949 376091 688145 378928
rect 687293 375787 688145 376091
rect 677707 332062 687193 340798
rect 39673 326866 39893 326994
rect 30533 320538 39893 326866
rect 677707 325734 687067 332062
rect 677707 325606 677927 325734
rect 30407 311802 39893 320538
rect 29455 278509 30307 278813
rect 29455 275672 29651 278509
rect 0 275368 29651 275672
rect 0 268602 28699 275368
rect 0 268334 28573 268602
rect 0 268000 4843 268254
rect 4923 268193 20920 268334
rect 0 240800 20920 268000
rect 0 240546 4843 240800
rect 4923 240466 20920 240594
rect 21000 240546 25993 268254
rect 26073 268193 26213 268334
rect 26073 240800 26213 268000
rect 26073 240466 26213 240594
rect 26293 240546 27183 268254
rect 27263 268193 27383 268334
rect 27263 240800 27383 268000
rect 27263 240466 27383 240594
rect 27463 240546 28353 268254
rect 28433 268193 28573 268334
rect 28433 240800 28573 268000
rect 28433 240466 28573 240594
rect 0 234138 28573 240466
rect 28653 234218 28719 268522
rect 0 232472 28699 234138
rect 28779 232552 29375 275288
rect 29455 268334 29651 275368
rect 29435 240546 29671 268254
rect 29455 235613 29651 240466
rect 29731 235693 30327 278429
rect 30387 277418 30453 311722
rect 30533 311534 39893 311802
rect 30533 311393 30673 311534
rect 30533 283666 30673 283794
rect 30753 283746 31683 311454
rect 31763 311393 31883 311534
rect 31763 283666 31883 283794
rect 31963 283746 32653 311454
rect 32733 311393 32853 311534
rect 32733 283666 32853 283794
rect 32933 283746 33623 311454
rect 33703 311393 33823 311534
rect 33703 283666 33823 283794
rect 33903 283746 34833 311454
rect 34913 311393 35033 311534
rect 36123 311473 37213 311534
rect 34913 283666 35033 283794
rect 35113 283746 36043 311454
rect 36123 311393 36243 311473
rect 37093 311393 37213 311473
rect 36323 283794 37013 311393
rect 36123 283714 36243 283794
rect 37093 283714 37213 283794
rect 37293 283746 38223 311454
rect 38303 311393 38423 311534
rect 36123 283666 37213 283714
rect 38303 283666 38423 283794
rect 38503 283746 39593 311454
rect 39673 311393 39893 311534
rect 677707 296066 677927 296207
rect 678007 296146 679097 325654
rect 679177 325606 679297 325734
rect 680387 325686 681477 325734
rect 679177 296066 679297 296207
rect 679377 296146 680307 325654
rect 680387 325606 680507 325686
rect 681357 325606 681477 325686
rect 680587 296207 681277 325606
rect 680387 296127 680507 296207
rect 681357 296127 681477 296207
rect 681557 296146 682487 325654
rect 682567 325606 682687 325734
rect 680387 296066 681477 296127
rect 682567 296066 682687 296207
rect 682767 296146 683697 325654
rect 683777 325606 683897 325734
rect 683777 296066 683897 296207
rect 683977 296146 684667 325654
rect 684747 325606 684867 325734
rect 684747 296066 684867 296207
rect 684947 296146 685637 325654
rect 685717 325606 685837 325734
rect 685717 296066 685837 296207
rect 685917 296146 686847 325654
rect 686927 325606 687067 325734
rect 686927 296066 687067 296207
rect 677707 295798 687067 296066
rect 687147 295878 687213 331982
rect 687273 330971 687869 375707
rect 687949 370934 688145 375787
rect 687929 341146 688165 370854
rect 687949 334032 688145 341066
rect 688225 334112 688821 378848
rect 688901 377262 717600 378928
rect 688881 340878 688947 377182
rect 689027 370934 717600 377262
rect 689027 370806 689167 370934
rect 689027 341400 689167 370600
rect 689027 341066 689167 341207
rect 689247 341146 690137 370854
rect 690217 370806 690337 370934
rect 690217 341400 690337 370600
rect 690217 341066 690337 341207
rect 690417 341146 691307 370854
rect 691387 370806 691527 370934
rect 691387 341400 691527 370600
rect 691387 341066 691527 341207
rect 691607 341146 696600 370854
rect 696680 370806 712677 370934
rect 712757 370600 717600 370854
rect 696680 341400 717600 370600
rect 696680 341066 712677 341207
rect 712757 341146 717600 341400
rect 689027 340798 717600 341066
rect 688901 334032 717600 340798
rect 687949 333728 717600 334032
rect 687949 330891 688145 333728
rect 687293 330587 688145 330891
rect 677707 287062 687193 295798
rect 39673 283666 39893 283794
rect 30533 277338 39893 283666
rect 677707 280734 687067 287062
rect 677707 280606 677927 280734
rect 30407 268602 39893 277338
rect 29455 235309 30307 235613
rect 29455 232472 29651 235309
rect 0 232168 29651 232472
rect 0 225402 28699 232168
rect 0 225134 28573 225402
rect 0 224800 4843 225054
rect 4923 224993 20920 225134
rect 0 197600 20920 224800
rect 0 197346 4843 197600
rect 4923 197266 20920 197394
rect 21000 197346 25993 225054
rect 26073 224993 26213 225134
rect 26073 197600 26213 224800
rect 26073 197266 26213 197394
rect 26293 197346 27183 225054
rect 27263 224993 27383 225134
rect 27263 197600 27383 224800
rect 27263 197266 27383 197394
rect 27463 197346 28353 225054
rect 28433 224993 28573 225134
rect 28433 197600 28573 224800
rect 28433 197266 28573 197394
rect 0 190938 28573 197266
rect 28653 191018 28719 225322
rect 0 189272 28699 190938
rect 28779 189352 29375 232088
rect 29455 225134 29651 232168
rect 29435 197346 29671 225054
rect 29455 192413 29651 197266
rect 29731 192493 30327 235229
rect 30387 234218 30453 268522
rect 30533 268334 39893 268602
rect 30533 268193 30673 268334
rect 30533 240466 30673 240594
rect 30753 240546 31683 268254
rect 31763 268193 31883 268334
rect 31763 240466 31883 240594
rect 31963 240546 32653 268254
rect 32733 268193 32853 268334
rect 32733 240466 32853 240594
rect 32933 240546 33623 268254
rect 33703 268193 33823 268334
rect 33703 240466 33823 240594
rect 33903 240546 34833 268254
rect 34913 268193 35033 268334
rect 36123 268273 37213 268334
rect 34913 240466 35033 240594
rect 35113 240546 36043 268254
rect 36123 268193 36243 268273
rect 37093 268193 37213 268273
rect 36323 240594 37013 268193
rect 36123 240514 36243 240594
rect 37093 240514 37213 240594
rect 37293 240546 38223 268254
rect 38303 268193 38423 268334
rect 36123 240466 37213 240514
rect 38303 240466 38423 240594
rect 38503 240546 39593 268254
rect 39673 268193 39893 268334
rect 677707 251066 677927 251207
rect 678007 251146 679097 280654
rect 679177 280606 679297 280734
rect 680387 280686 681477 280734
rect 679177 251066 679297 251207
rect 679377 251146 680307 280654
rect 680387 280606 680507 280686
rect 681357 280606 681477 280686
rect 680587 251207 681277 280606
rect 680387 251127 680507 251207
rect 681357 251127 681477 251207
rect 681557 251146 682487 280654
rect 682567 280606 682687 280734
rect 680387 251066 681477 251127
rect 682567 251066 682687 251207
rect 682767 251146 683697 280654
rect 683777 280606 683897 280734
rect 683777 251066 683897 251207
rect 683977 251146 684667 280654
rect 684747 280606 684867 280734
rect 684747 251066 684867 251207
rect 684947 251146 685637 280654
rect 685717 280606 685837 280734
rect 685717 251066 685837 251207
rect 685917 251146 686847 280654
rect 686927 280606 687067 280734
rect 686927 251066 687067 251207
rect 677707 250798 687067 251066
rect 687147 250878 687213 286982
rect 687273 285971 687869 330507
rect 687949 325734 688145 330587
rect 687929 296146 688165 325654
rect 687949 289032 688145 296066
rect 688225 289112 688821 333648
rect 688901 332062 717600 333728
rect 688881 295878 688947 331982
rect 689027 325734 717600 332062
rect 689027 325606 689167 325734
rect 689027 296400 689167 325400
rect 689027 296066 689167 296207
rect 689247 296146 690137 325654
rect 690217 325606 690337 325734
rect 690217 296400 690337 325400
rect 690217 296066 690337 296207
rect 690417 296146 691307 325654
rect 691387 325606 691527 325734
rect 691387 296400 691527 325400
rect 691387 296066 691527 296207
rect 691607 296146 696600 325654
rect 696680 325606 712677 325734
rect 712757 325400 717600 325654
rect 696680 296400 717600 325400
rect 696680 296066 712677 296207
rect 712757 296146 717600 296400
rect 689027 295798 717600 296066
rect 688901 289032 717600 295798
rect 687949 288728 717600 289032
rect 687949 285891 688145 288728
rect 687293 285587 688145 285891
rect 677707 242062 687193 250798
rect 39673 240466 39893 240594
rect 30533 234138 39893 240466
rect 677707 235734 687067 242062
rect 677707 235606 677927 235734
rect 30407 225402 39893 234138
rect 29455 192109 30307 192413
rect 29455 189272 29651 192109
rect 0 188968 29651 189272
rect 0 182202 28699 188968
rect 0 181934 28573 182202
rect 0 181600 4843 181854
rect 4923 181793 20920 181934
rect 0 154400 20920 181600
rect 0 152400 4843 154400
rect 0 125200 20920 152400
rect 0 124946 4843 125200
rect 4923 124866 20920 125007
rect 21000 124946 25993 181854
rect 26073 181793 26213 181934
rect 26073 154400 26213 181600
rect 26073 125200 26213 152400
rect 26073 124866 26213 125007
rect 26293 124946 27183 181854
rect 27263 181793 27383 181934
rect 27263 154400 27383 181600
rect 27263 125200 27383 152400
rect 27263 124866 27383 125007
rect 27463 124946 28353 181854
rect 28433 181793 28573 181934
rect 28433 154400 28573 181600
rect 28653 153400 28719 182122
rect 28433 125200 28573 152400
rect 28433 124866 28573 125007
rect 0 110534 28573 124866
rect 0 110200 4843 110454
rect 4923 110393 20920 110534
rect 0 83000 20920 110200
rect 0 82746 4843 83000
rect 4923 82666 20920 83000
rect 21000 82746 25993 110454
rect 26073 110393 26213 110534
rect 26073 82666 26213 110200
rect 26293 82746 27183 110454
rect 27263 110393 27383 110534
rect 27263 82666 27383 110200
rect 27463 82746 28353 110454
rect 28433 110393 28573 110534
rect 28433 82666 28573 110200
rect 0 68334 28573 82666
rect 0 68000 4843 68254
rect 4923 68193 20920 68334
rect 0 40800 20920 68000
rect 0 40546 4843 40800
rect 4923 40466 20920 40549
rect 0 40349 20920 40466
rect 21000 40429 25993 68254
rect 26073 68193 26213 68334
rect 26073 40800 26213 68000
rect 26073 40466 26213 40549
rect 26293 40546 27183 68254
rect 27263 68193 27383 68334
rect 27263 40800 27383 68000
rect 27263 40466 27383 40549
rect 27463 40546 28353 68254
rect 28433 68193 28573 68334
rect 28433 40800 28573 68000
rect 28433 40466 28573 40549
rect 26073 40349 28573 40466
rect 0 35285 28573 40349
rect 28653 35365 28719 152400
rect 28779 35418 29375 188888
rect 29455 181934 29651 188968
rect 29435 153400 29671 181854
rect 29435 124946 29671 152400
rect 29455 110534 29651 124866
rect 29435 82746 29671 110454
rect 29455 68334 29651 82666
rect 29435 36489 29671 68254
rect 29731 36625 30327 192029
rect 30387 191018 30453 225322
rect 30533 225134 39893 225402
rect 30533 224993 30673 225134
rect 30533 197266 30673 197394
rect 30753 197346 31683 225054
rect 31763 224993 31883 225134
rect 31763 197266 31883 197394
rect 31963 197346 32653 225054
rect 32733 224993 32853 225134
rect 32733 197266 32853 197394
rect 32933 197346 33623 225054
rect 33703 224993 33823 225134
rect 33703 197266 33823 197394
rect 33903 197346 34833 225054
rect 34913 224993 35033 225134
rect 36123 225073 37213 225134
rect 34913 197266 35033 197394
rect 35113 197346 36043 225054
rect 36123 224993 36243 225073
rect 37093 224993 37213 225073
rect 36323 197394 37013 224993
rect 36123 197314 36243 197394
rect 37093 197314 37213 197394
rect 37293 197346 38223 225054
rect 38303 224993 38423 225134
rect 36123 197266 37213 197314
rect 38303 197266 38423 197394
rect 38503 197346 39593 225054
rect 39673 224993 39893 225134
rect 677707 205866 677927 206007
rect 678007 205946 679097 235654
rect 679177 235606 679297 235734
rect 680387 235686 681477 235734
rect 679177 205866 679297 206007
rect 679377 205946 680307 235654
rect 680387 235606 680507 235686
rect 681357 235606 681477 235686
rect 680587 206007 681277 235606
rect 680387 205927 680507 206007
rect 681357 205927 681477 206007
rect 681557 205946 682487 235654
rect 682567 235606 682687 235734
rect 680387 205866 681477 205927
rect 682567 205866 682687 206007
rect 682767 205946 683697 235654
rect 683777 235606 683897 235734
rect 683777 205866 683897 206007
rect 683977 205946 684667 235654
rect 684747 235606 684867 235734
rect 684747 205866 684867 206007
rect 684947 205946 685637 235654
rect 685717 235606 685837 235734
rect 685717 205866 685837 206007
rect 685917 205946 686847 235654
rect 686927 235606 687067 235734
rect 686927 205866 687067 206007
rect 677707 205598 687067 205866
rect 687147 205678 687213 241982
rect 687273 240971 687869 285507
rect 687949 280734 688145 285587
rect 687929 251146 688165 280654
rect 687949 244032 688145 251066
rect 688225 244112 688821 288648
rect 688901 287062 717600 288728
rect 688881 250878 688947 286982
rect 689027 280734 717600 287062
rect 689027 280606 689167 280734
rect 689027 251400 689167 280400
rect 689027 251066 689167 251207
rect 689247 251146 690137 280654
rect 690217 280606 690337 280734
rect 690217 251400 690337 280400
rect 690217 251066 690337 251207
rect 690417 251146 691307 280654
rect 691387 280606 691527 280734
rect 691387 251400 691527 280400
rect 691387 251066 691527 251207
rect 691607 251146 696600 280654
rect 696680 280606 712677 280734
rect 712757 280400 717600 280654
rect 696680 251400 717600 280400
rect 696680 251066 712677 251207
rect 712757 251146 717600 251400
rect 689027 250798 717600 251066
rect 688901 244032 717600 250798
rect 687949 243728 717600 244032
rect 687949 240891 688145 243728
rect 687293 240587 688145 240891
rect 39673 197266 39893 197394
rect 30533 190938 39893 197266
rect 30407 182202 39893 190938
rect 677707 196862 687193 205598
rect 677707 190534 687067 196862
rect 677707 190406 677927 190534
rect 30387 153400 30453 182122
rect 30533 181934 39893 182202
rect 30533 181793 30673 181934
rect 30753 154400 31683 181854
rect 31763 181793 31883 181934
rect 31963 153400 32653 181854
rect 32733 181793 32853 181934
rect 29751 36409 30307 36545
rect 29455 36005 30307 36409
rect 30387 36085 30453 152400
rect 30533 124866 30673 125007
rect 30753 124946 31683 153400
rect 31763 124866 31883 125007
rect 31963 124946 32653 152400
rect 32733 124866 32853 125007
rect 32933 124946 33623 181854
rect 33703 181793 33823 181934
rect 33703 124866 33823 125007
rect 33903 124946 34833 181854
rect 34913 181793 35033 181934
rect 36123 181873 37213 181934
rect 34913 124866 35033 125007
rect 35113 124946 36043 181854
rect 36123 181793 36243 181873
rect 37093 181793 37213 181873
rect 36323 153400 37013 181793
rect 37293 154400 38223 181854
rect 38303 181793 38423 181934
rect 36323 125007 37013 152400
rect 36123 124927 36243 125007
rect 37093 124927 37213 125007
rect 37293 124946 38223 153400
rect 36123 124866 37213 124927
rect 38303 124866 38423 125007
rect 38503 124946 39593 181854
rect 39673 181793 39893 181934
rect 677707 160866 677927 161007
rect 678007 160946 679097 190454
rect 679177 190406 679297 190534
rect 680387 190486 681477 190534
rect 679177 160866 679297 161007
rect 679377 160946 680307 190454
rect 680387 190406 680507 190486
rect 681357 190406 681477 190486
rect 680587 161007 681277 190406
rect 680387 160927 680507 161007
rect 681357 160927 681477 161007
rect 681557 160946 682487 190454
rect 682567 190406 682687 190534
rect 680387 160866 681477 160927
rect 682567 160866 682687 161007
rect 682767 160946 683697 190454
rect 683777 190406 683897 190534
rect 683777 160866 683897 161007
rect 683977 160946 684667 190454
rect 684747 190406 684867 190534
rect 684747 160866 684867 161007
rect 684947 160946 685637 190454
rect 685717 190406 685837 190534
rect 685717 160866 685837 161007
rect 685917 160946 686847 190454
rect 686927 190406 687067 190534
rect 686927 160866 687067 161007
rect 677707 160598 687067 160866
rect 687147 160678 687213 196782
rect 687273 195771 687869 240507
rect 687949 235734 688145 240587
rect 687929 205946 688165 235654
rect 687949 198832 688145 205866
rect 688225 198912 688821 243648
rect 688901 242062 717600 243728
rect 688881 205678 688947 241982
rect 689027 235734 717600 242062
rect 689027 235606 689167 235734
rect 689027 206200 689167 235400
rect 689027 205866 689167 206007
rect 689247 205946 690137 235654
rect 690217 235606 690337 235734
rect 690217 206200 690337 235400
rect 690217 205866 690337 206007
rect 690417 205946 691307 235654
rect 691387 235606 691527 235734
rect 691387 206200 691527 235400
rect 691387 205866 691527 206007
rect 691607 205946 696600 235654
rect 696680 235606 712677 235734
rect 712757 235400 717600 235654
rect 696680 206200 717600 235400
rect 696680 205866 712677 206007
rect 712757 205946 717600 206200
rect 689027 205598 717600 205866
rect 688901 198832 717600 205598
rect 687949 198528 717600 198832
rect 687949 195691 688145 198528
rect 687293 195387 688145 195691
rect 677707 151862 687193 160598
rect 677707 145534 687067 151862
rect 677707 145406 677927 145534
rect 30533 110534 39593 124866
rect 677707 115666 677927 115807
rect 678007 115746 679097 145454
rect 679177 145406 679297 145534
rect 680387 145486 681477 145534
rect 679177 115666 679297 115807
rect 679377 115746 680307 145454
rect 680387 145406 680507 145486
rect 681357 145406 681477 145486
rect 680587 115807 681277 145406
rect 680387 115727 680507 115807
rect 681357 115727 681477 115807
rect 681557 115746 682487 145454
rect 682567 145406 682687 145534
rect 680387 115666 681477 115727
rect 682567 115666 682687 115807
rect 682767 115746 683697 145454
rect 683777 145406 683897 145534
rect 683777 115666 683897 115807
rect 683977 115746 684667 145454
rect 684747 145406 684867 145534
rect 684747 115666 684867 115807
rect 684947 115746 685637 145454
rect 685717 145406 685837 145534
rect 685717 115666 685837 115807
rect 685917 115746 686847 145454
rect 686927 145406 687067 145534
rect 686927 115666 687067 115807
rect 677707 115398 687067 115666
rect 687147 115478 687213 151782
rect 687273 150771 687869 195307
rect 687949 190534 688145 195387
rect 687929 160946 688165 190454
rect 687949 153832 688145 160866
rect 688225 153912 688821 198448
rect 688901 196862 717600 198528
rect 688881 160678 688947 196782
rect 689027 190534 717600 196862
rect 689027 190406 689167 190534
rect 689027 161200 689167 190200
rect 689027 160866 689167 161007
rect 689247 160946 690137 190454
rect 690217 190406 690337 190534
rect 690217 161200 690337 190200
rect 690217 160866 690337 161007
rect 690417 160946 691307 190454
rect 691387 190406 691527 190534
rect 691387 161200 691527 190200
rect 691387 160866 691527 161007
rect 691607 160946 696600 190454
rect 696680 190406 712677 190534
rect 712757 190200 717600 190454
rect 696680 161200 717600 190200
rect 696680 160866 712677 161007
rect 712757 160946 717600 161200
rect 689027 160598 717600 160866
rect 688901 153832 717600 160598
rect 687949 153528 717600 153832
rect 687949 150691 688145 153528
rect 687293 150387 688145 150691
rect 30533 110393 30673 110534
rect 30533 82666 30673 83000
rect 30753 82746 31683 110454
rect 31763 110393 31883 110534
rect 31763 82666 31883 83000
rect 31963 82746 32653 110454
rect 32733 110393 32853 110534
rect 32733 82666 32853 83000
rect 32933 82746 33623 110454
rect 33703 110393 33823 110534
rect 33703 82666 33823 83000
rect 33903 82746 34833 110454
rect 34913 110393 35033 110534
rect 36123 110473 37213 110534
rect 34913 82666 35033 83000
rect 35113 82746 36043 110454
rect 36123 110393 36243 110473
rect 37093 110393 37213 110473
rect 36123 82727 36243 83000
rect 36323 82807 37013 110393
rect 37093 82727 37213 83000
rect 37293 82746 38223 110454
rect 38303 110393 38423 110534
rect 36123 82666 37213 82727
rect 38303 82666 38423 83000
rect 38503 82746 39593 110454
rect 677707 106662 687193 115398
rect 677707 100334 687067 106662
rect 677707 100206 677927 100334
rect 30533 68334 39593 82666
rect 30533 68193 30673 68334
rect 30533 40466 30673 40549
rect 30753 40546 31683 68254
rect 31763 68193 31883 68334
rect 31763 40466 31883 40549
rect 31963 40546 32653 68254
rect 32733 68193 32853 68334
rect 32733 40466 32853 40549
rect 32933 40546 33623 68254
rect 33703 68193 33823 68334
rect 33703 40466 33823 40549
rect 33903 40546 34833 68254
rect 34913 68193 35033 68334
rect 36123 68273 37213 68334
rect 34913 40466 35033 40549
rect 35113 40546 36043 68254
rect 36123 68193 36243 68273
rect 37093 68193 37213 68273
rect 36323 40549 37013 68193
rect 36123 40469 36243 40549
rect 37093 40469 37213 40549
rect 37293 40546 38223 68254
rect 38303 68193 38423 68334
rect 36123 40466 37213 40469
rect 38303 40466 38423 40549
rect 38503 40546 39593 68254
rect 39673 40466 40000 40549
rect 30533 39673 40000 40466
rect 677051 39920 677927 40000
tri 677927 39920 678007 40000 se
rect 678007 39920 679097 100254
rect 679177 100206 679297 100334
rect 680387 100286 681477 100334
rect 679377 71000 680307 100254
rect 680387 100206 680507 100286
rect 681357 100206 681477 100286
rect 680587 70000 681277 100206
rect 186606 39673 202207 39893
rect 295206 39673 310807 39893
rect 350006 39673 365607 39893
rect 404806 39673 420407 39893
rect 459606 39673 475207 39893
rect 514406 39673 530007 39893
rect 677051 39673 679097 39920
rect 30533 38423 39450 39673
rect 39593 39593 39920 39673
tri 39920 39593 40000 39673 sw
rect 39530 38503 79054 39593
rect 79134 38423 93466 39593
rect 93546 38503 186654 39593
rect 30533 38303 40000 38423
rect 78993 38303 93607 38423
rect 30533 37213 39163 38303
rect 39243 37293 79054 38223
rect 79134 37213 93466 38303
rect 132600 38223 147600 38503
rect 186734 38423 202066 39673
rect 202146 38503 241454 39593
rect 241534 38423 255866 39593
rect 255946 38503 295254 39593
rect 295334 38423 310666 39673
rect 310746 38503 350054 39593
rect 350134 38423 365466 39673
rect 365546 38503 404854 39593
rect 404934 38423 420266 39673
rect 420346 38503 459654 39593
rect 459734 38423 475066 39673
rect 475146 38503 514454 39593
rect 514534 38423 529866 39673
rect 677134 39593 679097 39673
rect 529946 38503 569254 39593
rect 569334 38423 583666 39593
rect 583746 38503 623054 39593
rect 623134 38423 637466 39593
rect 637546 38503 677054 39593
rect 677134 39450 677927 39593
rect 678007 39530 679097 39593
rect 679177 39450 679297 40000
rect 677134 39163 679297 39450
rect 679377 39243 680307 70000
rect 680387 39626 680507 40000
rect 680587 39706 681277 69000
rect 681357 39626 681477 40000
rect 681557 39695 682487 100254
rect 682567 100206 682687 100334
rect 680387 39615 681477 39626
rect 682567 39615 682687 40000
rect 682767 39680 683697 100254
rect 683777 100206 683897 100334
rect 680387 39600 682687 39615
rect 683777 39643 683897 40000
rect 683977 39723 684667 100254
rect 684747 100206 684867 100334
rect 684947 70000 685637 100254
rect 685717 100206 685837 100334
rect 685917 71000 686847 100254
rect 686927 100206 687067 100334
rect 687147 70000 687213 106582
rect 687273 105571 687869 150307
rect 687949 145534 688145 150387
rect 687929 115746 688165 145454
rect 687949 108632 688145 115666
rect 688225 108712 688821 153448
rect 688901 151862 717600 153528
rect 688881 115478 688947 151782
rect 689027 145534 717600 151862
rect 689027 145406 689167 145534
rect 689027 116000 689167 145200
rect 689027 115666 689167 115807
rect 689247 115746 690137 145454
rect 690217 145406 690337 145534
rect 690217 116000 690337 145200
rect 690217 115666 690337 115807
rect 690417 115746 691307 145454
rect 691387 145406 691527 145534
rect 691387 116000 691527 145200
rect 691387 115666 691527 115807
rect 691607 115746 696600 145454
rect 696680 145406 712677 145534
rect 712757 145200 717600 145454
rect 696680 116000 717600 145200
rect 696680 115666 712677 115807
rect 712757 115746 717600 116000
rect 689027 115398 717600 115666
rect 688901 108632 717600 115398
rect 687949 108328 717600 108632
rect 687949 105491 688145 108328
rect 687293 105187 688145 105491
rect 684747 39653 684867 40000
rect 684947 39733 685637 69000
rect 685717 39653 685837 40000
rect 685917 39705 686847 70000
rect 684747 39643 685837 39653
rect 683777 39625 685837 39643
rect 686927 39625 687067 40000
rect 683777 39600 687067 39625
rect 680387 39163 687067 39600
rect 677134 38423 687067 39163
rect 186606 38303 202207 38423
rect 241200 38303 256007 38423
rect 295206 38303 310807 38423
rect 350006 38303 365607 38423
rect 404806 38303 420407 38423
rect 459606 38303 475207 38423
rect 514406 38303 530007 38423
rect 569193 38303 583807 38423
rect 622993 38303 637607 38423
rect 677051 38303 687067 38423
rect 93546 37293 186654 38223
rect 30533 37093 40000 37213
rect 78993 37093 93607 37213
rect 30533 36243 39626 37093
rect 39706 36323 78993 37013
rect 79073 36243 93527 37093
rect 132600 37013 147600 37293
rect 186734 37213 202066 38303
rect 202146 37293 241454 38223
rect 241534 37213 255866 38303
rect 255946 37293 295254 38223
rect 295334 37213 310666 38303
rect 310746 37293 350054 38223
rect 350134 37213 365466 38303
rect 365546 37293 404854 38223
rect 404934 37213 420266 38303
rect 420346 37293 459654 38223
rect 459734 37213 475066 38303
rect 475146 37293 514454 38223
rect 514534 37213 529866 38303
rect 529946 37293 569254 38223
rect 569334 37213 583666 38303
rect 583746 37293 623054 38223
rect 623134 37213 637466 38303
rect 637546 37293 677054 38223
rect 677134 37213 687067 38303
rect 186606 37093 202207 37213
rect 241200 37093 256007 37213
rect 295206 37093 310807 37213
rect 350006 37093 365607 37213
rect 404806 37093 420407 37213
rect 459606 37093 475207 37213
rect 514406 37093 530007 37213
rect 569193 37093 583807 37213
rect 622993 37093 637607 37213
rect 677051 37093 687067 37213
rect 93607 36323 186606 37013
rect 30533 36123 40000 36243
rect 78993 36123 93607 36243
rect 30533 36005 39615 36123
rect 29455 35338 39615 36005
rect 28799 35285 39615 35338
rect 0 35033 39615 35285
rect 39695 35113 79054 36043
rect 79134 35033 93466 36123
rect 132600 36043 147600 36323
rect 186686 36243 202127 37093
rect 202207 36323 241393 37013
rect 241473 36243 255927 37093
rect 256007 36323 295206 37013
rect 295286 36243 310727 37093
rect 310807 36323 350006 37013
rect 350086 36243 365527 37093
rect 365607 36323 404806 37013
rect 404886 36243 420327 37093
rect 420407 36323 459606 37013
rect 459686 36243 475127 37093
rect 475207 36323 514406 37013
rect 514486 36243 529927 37093
rect 530007 36323 569193 37013
rect 569273 36243 583727 37093
rect 583807 36323 622993 37013
rect 623073 36243 637527 37093
rect 637607 36323 677051 37013
rect 677131 36243 687067 37093
rect 186606 36123 202207 36243
rect 241200 36123 256007 36243
rect 295206 36123 310807 36243
rect 350006 36123 365607 36243
rect 404806 36123 420407 36243
rect 459606 36123 475207 36243
rect 514406 36123 530007 36243
rect 569193 36123 583807 36243
rect 622993 36123 637607 36243
rect 677051 36123 687067 36243
rect 93546 35113 186654 36043
rect 0 34913 40000 35033
rect 78993 34913 93607 35033
rect 0 33823 39600 34913
rect 39680 33903 79054 34833
rect 79134 33823 93466 34913
rect 132600 34833 147600 35113
rect 186734 35033 202066 36123
rect 202146 35113 241454 36043
rect 241534 35033 255866 36123
rect 255946 35113 295254 36043
rect 295334 35033 310666 36123
rect 310746 35113 350054 36043
rect 350134 35033 365466 36123
rect 365546 35113 404854 36043
rect 404934 35033 420266 36123
rect 420346 35113 459654 36043
rect 459734 35033 475066 36123
rect 475146 35113 514454 36043
rect 514534 35033 529866 36123
rect 529946 35113 569254 36043
rect 569334 35033 583666 36123
rect 583746 35113 623054 36043
rect 623134 35033 637466 36123
rect 637546 35113 677054 36043
rect 677134 36005 687067 36123
rect 687147 36085 687213 69000
rect 677134 35733 687193 36005
rect 687273 35813 687869 105107
rect 687949 100334 688145 105187
rect 687929 70000 688165 100254
rect 677134 35610 687849 35733
rect 687929 35690 688165 69000
rect 677134 35338 688145 35610
rect 688225 35418 688821 108248
rect 688901 106662 717600 108328
rect 688881 70000 688947 106582
rect 689027 100334 717600 106662
rect 689027 100206 689167 100334
rect 689027 71000 689167 100000
rect 688881 35365 688947 69000
rect 689027 39595 689167 69000
rect 689247 39675 690137 100254
rect 690217 100206 690337 100334
rect 690217 71000 690337 100000
rect 690217 39624 690337 69000
rect 690417 39704 691307 100254
rect 691387 100206 691527 100334
rect 691387 71000 691527 100000
rect 691387 39624 691527 69000
rect 690217 39595 691527 39624
rect 689027 39391 691527 39595
rect 691607 39471 696600 100254
rect 696680 100206 712677 100334
rect 712757 100000 717600 100254
rect 696680 71000 717600 100000
rect 712757 69000 717600 71000
rect 696680 40000 717600 69000
rect 696680 39633 712677 40000
rect 712757 39713 717600 40000
rect 696680 39391 717600 39633
rect 677134 35285 688801 35338
rect 689027 35285 717600 39391
rect 677134 35033 717600 35285
rect 186606 34913 202207 35033
rect 241200 34913 256007 35033
rect 295206 34913 310807 35033
rect 350006 34913 365607 35033
rect 404806 34913 420407 35033
rect 459606 34913 475207 35033
rect 514406 34913 530007 35033
rect 569193 34913 583807 35033
rect 622993 34913 637607 35033
rect 677051 34913 717600 35033
rect 93546 33903 186654 34833
rect 0 33703 40000 33823
rect 78993 33703 93607 33823
rect 0 32853 39643 33703
rect 39723 32933 79054 33623
rect 79134 32853 93466 33703
rect 132600 33623 147600 33903
rect 186734 33823 202066 34913
rect 202146 33903 241454 34833
rect 241534 33823 255866 34913
rect 255946 33903 295254 34833
rect 295334 33823 310666 34913
rect 310746 33903 350054 34833
rect 350134 33823 365466 34913
rect 365546 33903 404854 34833
rect 404934 33823 420266 34913
rect 420346 33903 459654 34833
rect 459734 33823 475066 34913
rect 475146 33903 514454 34833
rect 514534 33823 529866 34913
rect 529946 33903 569254 34833
rect 569334 33823 583666 34913
rect 583746 33903 623054 34833
rect 623134 33823 637466 34913
rect 637546 33903 677054 34833
rect 677134 33823 717600 34913
rect 186606 33703 202207 33823
rect 241200 33703 256007 33823
rect 295206 33703 310807 33823
rect 350006 33703 365607 33823
rect 404806 33703 420407 33823
rect 459606 33703 475207 33823
rect 514406 33703 530007 33823
rect 569193 33703 583807 33823
rect 622993 33703 637607 33823
rect 677051 33703 717600 33823
rect 93546 32933 186654 33623
rect 0 32733 40000 32853
rect 78993 32733 93607 32853
rect 0 31883 39653 32733
rect 39733 31963 79054 32653
rect 79134 31883 93466 32733
rect 132600 32653 147600 32933
rect 186734 32853 202066 33703
rect 202146 32933 241454 33623
rect 241534 32853 255866 33703
rect 255946 32933 295254 33623
rect 295334 32853 310666 33703
rect 310746 32933 350054 33623
rect 350134 32853 365466 33703
rect 365546 32933 404854 33623
rect 404934 32853 420266 33703
rect 420346 32933 459654 33623
rect 459734 32853 475066 33703
rect 475146 32933 514454 33623
rect 514534 32853 529866 33703
rect 529946 32933 569254 33623
rect 569334 32853 583666 33703
rect 583746 32933 623054 33623
rect 623134 32853 637466 33703
rect 637546 32933 677054 33623
rect 677134 32853 717600 33703
rect 186606 32733 202207 32853
rect 241200 32733 256007 32853
rect 295206 32733 310807 32853
rect 350006 32733 365607 32853
rect 404806 32733 420407 32853
rect 459606 32733 475207 32853
rect 514406 32733 530007 32853
rect 569193 32733 583807 32853
rect 622993 32733 637607 32853
rect 677051 32733 717600 32853
rect 93546 31963 186654 32653
rect 0 31763 40000 31883
rect 78993 31763 93607 31883
rect 0 30673 39625 31763
rect 39705 30753 79054 31683
rect 79134 30673 93466 31763
rect 132600 31683 147600 31963
rect 186734 31883 202066 32733
rect 202146 31963 241454 32653
rect 241534 31883 255866 32733
rect 255946 31963 295254 32653
rect 295334 31883 310666 32733
rect 310746 31963 350054 32653
rect 350134 31883 365466 32733
rect 365546 31963 404854 32653
rect 404934 31883 420266 32733
rect 420346 31963 459654 32653
rect 459734 31883 475066 32733
rect 475146 31963 514454 32653
rect 514534 31883 529866 32733
rect 529946 31963 569254 32653
rect 569334 31883 583666 32733
rect 583746 31963 623054 32653
rect 623134 31883 637466 32733
rect 637546 31963 677054 32653
rect 677134 31883 717600 32733
rect 186606 31763 202207 31883
rect 241200 31763 256007 31883
rect 295206 31763 310807 31883
rect 350006 31763 365607 31883
rect 404806 31763 420407 31883
rect 459606 31763 475207 31883
rect 514406 31763 530007 31883
rect 569193 31763 583807 31883
rect 622993 31763 637607 31883
rect 677051 31763 717600 31883
rect 93546 30753 186654 31683
rect 0 30533 40000 30673
rect 78993 30533 93607 30673
rect 0 30407 36005 30533
rect 0 29751 35733 30407
rect 36085 30387 79054 30453
rect 79134 30407 93466 30533
rect 132600 30453 147600 30753
rect 186734 30673 202066 31763
rect 202146 30753 241454 31683
rect 241534 30673 255866 31763
rect 255946 30753 295254 31683
rect 295334 30673 310666 31763
rect 310746 30753 350054 31683
rect 350134 30673 365466 31763
rect 365546 30753 404854 31683
rect 404934 30673 420266 31763
rect 420346 30753 459654 31683
rect 459734 30673 475066 31763
rect 475146 30753 514454 31683
rect 514534 30673 529866 31763
rect 529946 30753 569254 31683
rect 569334 30673 583666 31763
rect 583746 30753 623054 31683
rect 623134 30673 637466 31763
rect 637546 30753 677054 31683
rect 677134 30673 717600 31763
rect 186606 30533 202207 30673
rect 241200 30533 256007 30673
rect 295206 30533 310807 30673
rect 350006 30533 365607 30673
rect 404806 30533 420407 30673
rect 459606 30533 475207 30673
rect 514406 30533 530007 30673
rect 569193 30533 583807 30673
rect 622993 30533 637607 30673
rect 677051 30533 717600 30673
rect 93546 30407 192982 30453
rect 193062 30407 201798 30533
rect 93546 30387 132600 30407
rect 147600 30387 192982 30407
rect 201878 30387 301582 30453
rect 301662 30407 310398 30533
rect 310478 30387 356382 30453
rect 356462 30407 365198 30533
rect 365278 30387 411182 30453
rect 411262 30407 419998 30533
rect 420078 30387 465982 30453
rect 466062 30407 474798 30533
rect 474878 30387 520782 30453
rect 520862 30407 529598 30533
rect 529678 30387 681515 30453
rect 0 29455 35610 29751
rect 35813 29731 191507 30327
rect 0 28799 35338 29455
rect 35690 29435 79054 29671
rect 93546 29651 132600 29671
rect 147600 29651 186654 29671
rect 191587 29651 191891 30307
rect 191971 29731 300107 30327
rect 79134 29455 93466 29651
rect 93546 29455 186654 29651
rect 186734 29455 202066 29651
rect 93546 29435 132600 29455
rect 147600 29435 186654 29455
rect 0 28573 35285 28799
rect 35418 28779 194648 29375
rect 35365 28653 79054 28719
rect 93546 28699 132600 28719
rect 147600 28699 192982 28719
rect 194728 28699 195032 29455
rect 202146 29435 241454 29671
rect 241534 29455 255866 29651
rect 255946 29435 295254 29671
rect 300187 29651 300491 30307
rect 300571 29731 354907 30327
rect 295334 29455 310666 29651
rect 195112 28779 303248 29375
rect 79134 28573 93466 28699
rect 93546 28653 192982 28699
rect 132600 28573 147600 28653
rect 193062 28573 201798 28699
rect 201878 28653 301582 28719
rect 303328 28699 303632 29455
rect 310746 29435 350054 29671
rect 354987 29651 355291 30307
rect 355371 29731 409707 30327
rect 350134 29455 365466 29651
rect 303712 28779 358048 29375
rect 301662 28573 310398 28699
rect 310478 28653 356382 28719
rect 358128 28699 358432 29455
rect 365546 29435 404854 29671
rect 409787 29651 410091 30307
rect 410171 29731 464507 30327
rect 404934 29455 420266 29651
rect 358512 28779 412848 29375
rect 356462 28573 365198 28699
rect 365278 28653 411182 28719
rect 412928 28699 413232 29455
rect 420346 29435 459654 29671
rect 464587 29651 464891 30307
rect 464971 29731 519307 30327
rect 459734 29455 475066 29651
rect 413312 28779 467648 29375
rect 411262 28573 419998 28699
rect 420078 28653 465982 28719
rect 467728 28699 468032 29455
rect 475146 29435 514454 29671
rect 519387 29651 519691 30307
rect 519771 29731 680975 30327
rect 681595 30307 717600 30533
rect 681055 29751 717600 30307
rect 514534 29455 529866 29651
rect 468112 28779 522448 29375
rect 466062 28573 474798 28699
rect 474878 28653 520782 28719
rect 522528 28699 522832 29455
rect 529946 29435 569254 29671
rect 569334 29455 583666 29651
rect 583746 29435 623054 29671
rect 623134 29455 637466 29651
rect 637546 29435 681111 29671
rect 681191 29455 717600 29751
rect 522912 28779 682182 29375
rect 682262 28799 717600 29455
rect 520862 28573 529598 28699
rect 529678 28653 682235 28719
rect 682315 28573 717600 28799
rect 0 28433 47400 28573
rect 71400 28433 78800 28573
rect 78993 28433 93607 28573
rect 93800 28433 101200 28573
rect 125200 28433 155000 28573
rect 179000 28433 186400 28573
rect 186606 28433 202207 28573
rect 202400 28433 209800 28573
rect 233800 28433 256007 28573
rect 256200 28433 263600 28573
rect 287600 28433 295000 28573
rect 295206 28433 310807 28573
rect 311000 28433 318400 28573
rect 342400 28433 349800 28573
rect 350006 28433 365607 28573
rect 365800 28433 373200 28573
rect 397200 28433 404600 28573
rect 404806 28433 420407 28573
rect 420600 28433 428000 28573
rect 452000 28433 459400 28573
rect 459606 28433 475207 28573
rect 475400 28433 482800 28573
rect 506800 28433 514200 28573
rect 514406 28433 530007 28573
rect 530200 28433 537600 28573
rect 561600 28433 569000 28573
rect 569193 28433 583807 28573
rect 584000 28433 591400 28573
rect 615400 28433 622800 28573
rect 622993 28433 637607 28573
rect 637800 28433 645200 28573
rect 669200 28433 676800 28573
rect 677051 28433 717600 28573
rect 0 27383 39595 28433
rect 39675 27463 79054 28353
rect 79134 27383 93466 28433
rect 132600 28353 147600 28433
rect 93546 27463 186654 28353
rect 132600 27383 147600 27463
rect 186734 27383 202066 28433
rect 202146 27463 241454 28353
rect 241534 27383 255866 28433
rect 255946 27463 295254 28353
rect 295334 27383 310666 28433
rect 310746 27463 350054 28353
rect 350134 27383 365466 28433
rect 365546 27463 404854 28353
rect 404934 27383 420266 28433
rect 420346 27463 459654 28353
rect 459734 27383 475066 28433
rect 475146 27463 514454 28353
rect 514534 27383 529866 28433
rect 529946 27463 569254 28353
rect 569334 27383 583666 28433
rect 583746 27463 623054 28353
rect 623134 27383 637466 28433
rect 637546 27463 677054 28353
rect 677134 27383 717600 28433
rect 0 27263 47400 27383
rect 71400 27263 78800 27383
rect 78993 27263 93607 27383
rect 93800 27263 101200 27383
rect 125200 27263 155000 27383
rect 179000 27263 186400 27383
rect 186606 27263 202207 27383
rect 202400 27263 209800 27383
rect 233800 27263 256007 27383
rect 256200 27263 263600 27383
rect 287600 27263 295000 27383
rect 295206 27263 310807 27383
rect 311000 27263 318400 27383
rect 342400 27263 349800 27383
rect 350006 27263 365607 27383
rect 365800 27263 373200 27383
rect 397200 27263 404600 27383
rect 404806 27263 420407 27383
rect 420600 27263 428000 27383
rect 452000 27263 459400 27383
rect 459606 27263 475207 27383
rect 475400 27263 482800 27383
rect 506800 27263 514200 27383
rect 514406 27263 530007 27383
rect 530200 27263 537600 27383
rect 561600 27263 569000 27383
rect 569193 27263 583807 27383
rect 584000 27263 591400 27383
rect 615400 27263 622800 27383
rect 622993 27263 637607 27383
rect 637800 27263 645200 27383
rect 669200 27263 676800 27383
rect 677051 27263 717600 27383
rect 0 26213 39624 27263
rect 39704 26293 79054 27183
rect 79134 26213 93466 27263
rect 132600 27183 147600 27263
rect 93546 26293 186654 27183
rect 132600 26213 147600 26293
rect 186734 26213 202066 27263
rect 202146 26293 241454 27183
rect 241534 26213 255866 27263
rect 255946 26293 295254 27183
rect 295334 26213 310666 27263
rect 310746 26293 350054 27183
rect 350134 26213 365466 27263
rect 365546 26293 404854 27183
rect 404934 26213 420266 27263
rect 420346 26293 459654 27183
rect 459734 26213 475066 27263
rect 475146 26293 514454 27183
rect 514534 26213 529866 27263
rect 529946 26293 569254 27183
rect 569334 26213 583666 27263
rect 583746 26293 623054 27183
rect 623134 26213 637466 27263
rect 637546 26293 677054 27183
rect 677134 26213 717600 27263
rect 0 26073 47400 26213
rect 71400 26073 78800 26213
rect 78993 26073 93607 26213
rect 93800 26073 101200 26213
rect 125200 26073 155000 26213
rect 179000 26073 186400 26213
rect 186606 26073 202207 26213
rect 202400 26073 209800 26213
rect 233800 26073 256007 26213
rect 256200 26073 263600 26213
rect 287600 26073 295000 26213
rect 295206 26073 310807 26213
rect 311000 26073 318400 26213
rect 342400 26073 349800 26213
rect 350006 26073 365607 26213
rect 365800 26073 373200 26213
rect 397200 26073 404600 26213
rect 404806 26073 420407 26213
rect 420600 26073 428000 26213
rect 452000 26073 459400 26213
rect 459606 26073 475207 26213
rect 475400 26073 482800 26213
rect 506800 26073 514200 26213
rect 514406 26073 530007 26213
rect 530200 26073 537600 26213
rect 561600 26073 569000 26213
rect 569193 26073 583807 26213
rect 584000 26073 591400 26213
rect 615400 26073 622800 26213
rect 622993 26073 637607 26213
rect 637800 26073 645200 26213
rect 669200 26073 676800 26213
rect 677051 26073 717600 26213
rect 0 20920 39391 26073
rect 39471 21000 79054 25993
rect 79134 20920 93466 26073
rect 132600 25993 147600 26073
rect 93546 21000 186654 25993
rect 132600 20920 147600 21000
rect 186734 20920 202066 26073
rect 202146 21000 241454 25993
rect 241534 20920 255866 26073
rect 255946 21000 295254 25993
rect 295334 20920 310666 26073
rect 310746 21000 350054 25993
rect 350134 20920 365466 26073
rect 365546 21000 404854 25993
rect 404934 20920 420266 26073
rect 420346 21000 459654 25993
rect 459734 20920 475066 26073
rect 475146 21000 514454 25993
rect 514534 20920 529866 26073
rect 529946 21000 569254 25993
rect 569334 20920 583666 26073
rect 583746 21000 623054 25993
rect 623134 20920 637466 26073
rect 637546 21000 677171 25993
rect 677251 20920 717600 26073
rect 0 4923 47400 20920
rect 0 0 39633 4923
rect 40000 4843 47400 4923
rect 71400 4843 78800 20920
rect 78993 4923 93607 20920
rect 39713 0 79054 4843
rect 79134 0 93466 4923
rect 93800 4843 101200 20920
rect 125200 4843 155000 20920
rect 179000 4843 186400 20920
rect 186606 4923 202207 20920
rect 93546 0 186654 4843
rect 186734 0 202066 4923
rect 202400 4843 209800 20920
rect 233800 4923 256007 20920
rect 233800 4843 241200 4923
rect 202146 0 241454 4843
rect 241534 0 255866 4923
rect 256200 4843 263600 20920
rect 287600 4843 295000 20920
rect 295206 4923 310807 20920
rect 255946 0 295254 4843
rect 295334 0 310666 4923
rect 311000 4843 318400 20920
rect 342400 4843 349800 20920
rect 350006 4923 365607 20920
rect 310746 0 350054 4843
rect 350134 0 365466 4923
rect 365800 4843 373200 20920
rect 397200 4843 404600 20920
rect 404806 4923 420407 20920
rect 365546 0 404854 4843
rect 404934 0 420266 4923
rect 420600 4843 428000 20920
rect 452000 4843 459400 20920
rect 459606 4923 475207 20920
rect 420346 0 459654 4843
rect 459734 0 475066 4923
rect 475400 4843 482800 20920
rect 506800 4843 514200 20920
rect 514406 4923 530007 20920
rect 475146 0 514454 4843
rect 514534 0 529866 4923
rect 530200 4843 537600 20920
rect 561600 4843 569000 20920
rect 569193 4923 583807 20920
rect 529946 0 569254 4843
rect 569334 0 583666 4923
rect 584000 4843 591400 20920
rect 615400 4843 622800 20920
rect 622993 4923 637607 20920
rect 583746 0 623054 4843
rect 623134 0 637466 4923
rect 637800 4843 645200 20920
rect 669200 4843 676800 20920
rect 677051 4923 717600 20920
rect 637546 0 677054 4843
rect 677134 0 717600 4923
<< metal5 >>
rect 78440 1018512 90960 1031002
rect 129840 1018512 142360 1031002
rect 181240 1018512 193760 1031002
rect 232640 1018512 245160 1031002
rect 284240 1018512 296760 1031002
rect 334810 1018624 346978 1030789
rect 386040 1018512 398560 1031002
rect 475040 1018512 487560 1031002
rect 526440 1018512 538960 1031002
rect 577010 1018624 589178 1030789
rect 628240 1018512 640760 1031002
rect 6598 956440 19088 968960
rect 698512 952840 711002 965360
rect 6167 914054 19620 924934
rect 697980 909666 711433 920546
rect 6811 871210 18976 883378
rect 698512 863640 711002 876160
rect 6811 829010 18976 841178
rect 698624 819822 710789 831990
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 698624 505222 710789 517390
rect 6811 484410 18976 496578
rect 697980 461866 711433 472746
rect 6167 442854 19620 453734
rect 698624 417022 710789 429190
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 6598 313440 19088 325960
rect 698512 326640 711002 339160
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 6811 111610 18976 123778
rect 698512 101240 711002 113760
rect 6167 70054 19620 80934
rect 93607 36343 132793 36993
rect 93546 30773 132854 31663
rect 93546 28653 132854 30453
rect 80222 6811 92390 18976
rect 133840 6675 146380 19198
rect 187640 6598 200160 19088
rect 243266 6167 254146 19620
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18976
rect 624222 6811 636390 18976
<< obsm5 >>
rect 0 1032757 717600 1037600
rect 0 1016917 40800 1032757
rect 76200 1031322 92200 1032757
rect 76200 1018192 78120 1031322
rect 91280 1018192 92200 1031322
rect 76200 1016917 92200 1018192
rect 127600 1031322 143600 1032757
rect 127600 1018192 129520 1031322
rect 142680 1018192 143600 1031322
rect 127600 1016917 143600 1018192
rect 179000 1031322 195000 1032757
rect 179000 1018192 180920 1031322
rect 194080 1018192 195000 1031322
rect 179000 1016917 195000 1018192
rect 230400 1031322 246400 1032757
rect 230400 1018192 232320 1031322
rect 245480 1018192 246400 1031322
rect 230400 1016917 246400 1018192
rect 282000 1031322 298000 1032757
rect 282000 1018192 283920 1031322
rect 297080 1018192 298000 1031322
rect 282000 1016917 298000 1018192
rect 333400 1031109 348400 1032757
rect 333400 1018304 334490 1031109
rect 347298 1018304 348400 1031109
rect 333400 1016917 348400 1018304
rect 383800 1031322 399800 1032757
rect 383800 1018192 385720 1031322
rect 398880 1018192 399800 1031322
rect 383800 1016917 399800 1018192
rect 472800 1031322 488800 1032757
rect 472800 1018192 474720 1031322
rect 487880 1018192 488800 1031322
rect 472800 1016917 488800 1018192
rect 524200 1031322 540200 1032757
rect 524200 1018192 526120 1031322
rect 539280 1018192 540200 1031322
rect 524200 1016917 540200 1018192
rect 575600 1031109 590600 1032757
rect 575600 1018304 576690 1031109
rect 589498 1018304 590600 1031109
rect 575600 1016917 590600 1018304
rect 626000 1031322 642000 1032757
rect 626000 1018192 627920 1031322
rect 641080 1018192 642000 1031322
rect 626000 1016917 642000 1018192
rect 677600 1016917 717600 1032757
rect 0 1011287 40109 1016917
rect 40429 1011607 76454 1016597
rect 0 1009267 40226 1011287
rect 40546 1010437 76454 1011287
rect 40546 1009267 76454 1010117
rect 0 1006827 35049 1009267
rect 35369 1007147 76454 1008947
rect 0 1002551 40226 1006827
rect 40546 1005937 76454 1006827
rect 40546 1004968 76454 1005617
rect 40800 1004967 76200 1004968
rect 40546 1003997 76454 1004647
rect 40546 1002787 76454 1003677
rect 0 998449 28333 1002551
rect 0 997600 20683 998449
rect 26313 998245 28333 998449
rect 26313 998216 27163 998245
rect 0 970200 4843 997600
rect 0 969626 20683 970200
rect 21003 969946 25993 998129
rect 26313 969946 27163 997896
rect 27483 969946 28333 997925
rect 28653 969946 30453 1002231
rect 30773 1001257 40226 1002551
rect 40546 1001577 76454 1002467
rect 76774 1001257 91626 1016917
rect 91946 1011607 127854 1016597
rect 91946 1010437 127854 1011287
rect 91946 1009267 127854 1010117
rect 91946 1007147 127854 1008947
rect 91946 1005937 127854 1006827
rect 91946 1004968 127854 1005617
rect 92200 1004967 127600 1004968
rect 91946 1003997 127854 1004647
rect 91946 1002787 127854 1003677
rect 91946 1001577 127854 1002467
rect 128174 1001257 143026 1016917
rect 143346 1011607 179254 1016597
rect 143346 1010437 179254 1011287
rect 143346 1009267 179254 1010117
rect 143346 1007147 179254 1008947
rect 143346 1005937 179254 1006827
rect 143346 1004968 179254 1005617
rect 143600 1004967 179000 1004968
rect 143346 1003997 179254 1004647
rect 143346 1002787 179254 1003677
rect 143346 1001577 179254 1002467
rect 179574 1001257 194426 1016917
rect 194746 1011607 230654 1016597
rect 194746 1010437 230654 1011287
rect 194746 1009267 230654 1010117
rect 194746 1007147 230654 1008947
rect 194746 1005937 230654 1006827
rect 194746 1004968 230654 1005617
rect 195000 1004967 230400 1004968
rect 194746 1003997 230654 1004647
rect 194746 1002787 230654 1003677
rect 194746 1001577 230654 1002467
rect 230974 1001257 245826 1016917
rect 246146 1011607 282254 1016597
rect 246146 1010437 282254 1011287
rect 246146 1009267 282254 1010117
rect 246146 1007147 282254 1008947
rect 246146 1005937 282254 1006827
rect 246146 1004968 282254 1005617
rect 246400 1004967 282000 1004968
rect 246146 1003997 282254 1004647
rect 246146 1002787 282254 1003677
rect 246146 1001577 282254 1002467
rect 282574 1001257 297426 1016917
rect 297746 1011607 333654 1016597
rect 297746 1010437 333654 1011287
rect 297746 1009267 333654 1010117
rect 297746 1007147 333654 1008947
rect 297746 1005937 333654 1006827
rect 297746 1004968 333654 1005617
rect 333974 1004968 347826 1016917
rect 348146 1011607 384054 1016597
rect 348146 1010437 384054 1011287
rect 348146 1009267 384054 1010117
rect 348146 1007147 384054 1008947
rect 348146 1005937 384054 1006827
rect 348146 1004968 384054 1005617
rect 298000 1004967 383800 1004968
rect 297746 1003997 333654 1004647
rect 297746 1002787 333654 1003677
rect 297746 1001577 333654 1002467
rect 333974 1001257 347826 1004967
rect 348146 1003997 384054 1004647
rect 348146 1002787 384054 1003677
rect 348146 1001577 384054 1002467
rect 384374 1001257 399226 1016917
rect 399546 1011607 473054 1016597
rect 399546 1010437 473054 1011287
rect 399546 1009267 473054 1010117
rect 399546 1007147 435200 1008947
rect 436200 1007147 473054 1008947
rect 399546 1005937 436200 1006827
rect 437200 1005937 473054 1006827
rect 399546 1004968 435200 1005617
rect 399800 1004967 435200 1004968
rect 436200 1004968 473054 1005617
rect 436200 1004967 472800 1004968
rect 399546 1003997 473054 1004647
rect 399546 1002787 473054 1003677
rect 399546 1001577 473054 1002467
rect 473374 1001257 488226 1016917
rect 488546 1011607 524454 1016597
rect 488546 1010437 524454 1011287
rect 488546 1009267 524454 1010117
rect 488546 1007147 524454 1008947
rect 488546 1005937 524454 1006827
rect 488546 1004968 524454 1005617
rect 488800 1004967 524200 1004968
rect 488546 1003997 524454 1004647
rect 488546 1002787 524454 1003677
rect 488546 1001577 524454 1002467
rect 524774 1001257 539626 1016917
rect 539946 1011607 575854 1016597
rect 539946 1010437 575854 1011287
rect 539946 1009267 575854 1010117
rect 539946 1007147 575854 1008947
rect 539946 1005937 575854 1006827
rect 539946 1004968 575854 1005617
rect 576174 1004968 590026 1016917
rect 590346 1011607 626254 1016597
rect 590346 1010437 626254 1011287
rect 590346 1009267 626254 1010117
rect 590346 1007147 626254 1008947
rect 590346 1005937 626254 1006827
rect 590346 1004968 626254 1005617
rect 540200 1004967 626000 1004968
rect 539946 1003997 575854 1004647
rect 539946 1002787 575854 1003677
rect 539946 1001577 575854 1002467
rect 576174 1001257 590026 1004967
rect 590346 1003997 626254 1004647
rect 590346 1002787 626254 1003677
rect 590346 1001577 626254 1002467
rect 626574 1001257 641426 1016917
rect 641746 1011607 678129 1016597
rect 678449 1011287 717600 1016917
rect 641746 1010437 677896 1011287
rect 678216 1010437 717600 1011287
rect 641746 1009267 677925 1010117
rect 678245 1009267 717600 1010437
rect 641746 1007147 682231 1008947
rect 682551 1006827 717600 1009267
rect 641746 1005937 677895 1006827
rect 678215 1005617 717600 1006827
rect 641746 1004968 677867 1005617
rect 642000 1004967 677867 1004968
rect 678187 1004967 717600 1005617
rect 641746 1003997 677877 1004647
rect 678197 1003997 717600 1004967
rect 641746 1002787 677920 1003677
rect 678240 1002551 717600 1003997
rect 678240 1002467 686827 1002551
rect 641746 1001577 677905 1002467
rect 678225 1001257 686827 1002467
rect 30773 1000607 40229 1001257
rect 40549 1000607 76393 1001257
rect 76713 1000607 91674 1001257
rect 91994 1000607 127793 1001257
rect 128113 1000607 143074 1001257
rect 143394 1000607 179193 1001257
rect 179513 1000607 194474 1001257
rect 194794 1000607 230593 1001257
rect 230913 1000607 245874 1001257
rect 246194 1000607 282193 1001257
rect 282513 1000607 297474 1001257
rect 297794 1000607 333593 1001257
rect 333913 1000607 347887 1001257
rect 348207 1000607 383993 1001257
rect 384313 1000607 399274 1001257
rect 399594 1000607 435200 1001257
rect 436200 1000607 472993 1001257
rect 473313 1000607 488274 1001257
rect 488594 1000607 524393 1001257
rect 524713 1000607 539674 1001257
rect 539994 1000607 575793 1001257
rect 576113 1000607 590087 1001257
rect 590407 1000607 626193 1001257
rect 626513 1000607 641474 1001257
rect 641794 1000607 677894 1001257
rect 678214 1000607 686827 1001257
rect 30773 998677 40226 1000607
rect 40546 999397 76454 1000287
rect 30773 998240 36993 998677
rect 38523 998390 40226 998677
rect 30773 998215 33603 998240
rect 35133 998225 36993 998240
rect 31983 998197 33603 998215
rect 36343 998214 36993 998225
rect 31983 998187 32633 998197
rect 30773 969946 31663 997895
rect 31983 970200 32633 997867
rect 31983 969946 32632 970200
rect 32953 969946 33603 997877
rect 33923 969946 34813 997920
rect 35133 969946 36023 997905
rect 36343 969994 36993 997894
rect 37313 969946 38203 998357
rect 38523 998027 39573 998070
rect 39893 998027 40226 998390
rect 40546 998027 76454 999077
rect 76774 998027 91626 1000607
rect 91946 999397 127854 1000287
rect 91946 998027 127854 999077
rect 128174 998027 143026 1000607
rect 143346 999397 179254 1000287
rect 143346 998027 179254 999077
rect 179574 998027 194426 1000607
rect 194746 999397 230654 1000287
rect 194746 998027 230654 999077
rect 230974 998027 245826 1000607
rect 246146 999397 282254 1000287
rect 246146 998027 282254 999077
rect 282574 998027 297426 1000607
rect 297746 999397 333654 1000287
rect 297746 998027 333654 999077
rect 333974 998027 347826 1000607
rect 348146 999397 384054 1000287
rect 348146 998027 384054 999077
rect 384374 998027 399226 1000607
rect 399546 999397 436200 1000287
rect 437200 999397 473054 1000287
rect 399546 998027 473054 999077
rect 473374 998027 488226 1000607
rect 488546 999397 524454 1000287
rect 488546 998027 524454 999077
rect 524774 998027 539626 1000607
rect 539946 999397 575854 1000287
rect 539946 998027 575854 999077
rect 576174 998027 590026 1000607
rect 590346 999397 626254 1000287
rect 590346 998027 626254 999077
rect 626574 998027 641426 1000607
rect 641746 999397 678357 1000287
rect 678677 999077 686827 1000607
rect 641746 998027 678070 999077
rect 38523 997920 40226 998027
rect 38523 969946 39573 997920
tri 39573 997600 39893 997920 nw
rect 39893 997707 40226 997920
tri 677600 997707 677920 998027 ne
rect 677920 997707 678027 998027
rect 678390 997707 686827 999077
rect 39893 997600 40800 997707
rect 677600 997374 686827 997707
rect 677600 996800 677707 997374
rect 680607 997371 681257 997374
rect 36343 969626 36993 969674
rect 0 969280 39573 969626
rect 0 956120 6278 969280
rect 19408 956120 39573 969280
rect 678027 967346 679077 997054
rect 679397 967346 680287 997054
rect 680607 967407 681257 997051
rect 681577 967346 682467 997054
rect 682787 967346 683677 997054
rect 683997 967346 684647 997054
rect 684968 996800 685617 997054
rect 684967 967600 685617 996800
rect 684968 967346 685617 967600
rect 685937 967346 686827 997054
rect 687147 967346 688947 1002231
rect 689267 997491 717600 1002551
rect 689267 997374 691287 997491
rect 689267 967346 690117 997054
rect 690437 967346 691287 997054
rect 691607 967346 696597 997171
rect 696917 996800 717600 997491
rect 712757 967600 717600 996800
rect 680607 967026 681257 967087
rect 696917 967026 717600 967600
rect 0 954774 39573 956120
rect 678027 965680 717600 967026
rect 0 954200 20683 954774
rect 36343 954713 36993 954774
rect 0 927000 4843 954200
rect 0 926426 20683 927000
rect 21003 926746 25993 954454
rect 26313 926746 27163 954454
rect 27483 926746 28333 954454
rect 28653 926746 30453 954454
rect 30773 926746 31663 954454
rect 31983 954200 32632 954454
rect 31983 927000 32633 954200
rect 31983 926746 32632 927000
rect 32953 926746 33603 954454
rect 33923 926746 34813 954454
rect 35133 926746 36023 954454
rect 36343 926807 36993 954393
rect 37313 926746 38203 954454
rect 38523 926746 39573 954454
rect 678027 952520 698192 965680
rect 711322 952520 717600 965680
rect 678027 952174 717600 952520
rect 680607 952126 681257 952174
rect 36343 926426 36993 926487
rect 0 925254 39573 926426
rect 0 913734 5847 925254
rect 19940 913734 39573 925254
rect 678027 922346 679077 951854
rect 679397 922346 680287 951854
rect 680607 922407 681257 951806
rect 681577 922346 682467 951854
rect 682787 922346 683677 951854
rect 683997 922346 684647 951854
rect 684968 951600 685617 951854
rect 684967 922600 685617 951600
rect 684968 922346 685617 922600
rect 685937 922346 686827 951854
rect 687147 922346 688947 951854
rect 689267 922346 690117 951854
rect 690437 922346 691287 951854
rect 691607 922346 696597 951854
rect 696917 951600 717600 952174
rect 712757 922600 717600 951600
rect 680607 922026 681257 922087
rect 696917 922026 717600 922600
rect 0 912574 39573 913734
rect 678027 920866 717600 922026
rect 0 912000 20683 912574
rect 36343 912513 36993 912574
rect 0 884800 4843 912000
rect 0 884226 20683 884800
rect 21003 884546 25993 912254
rect 26313 884546 27163 912254
rect 27483 884546 28333 912254
rect 28653 884546 30453 912254
rect 30773 884546 31663 912254
rect 31983 912000 32632 912254
rect 31983 884546 32633 912000
rect 32953 884546 33603 912254
rect 33923 884546 34813 912254
rect 35133 884546 36023 912254
rect 36343 884607 36993 912193
rect 37313 884546 38203 912254
rect 38523 884546 39573 912254
rect 678027 909346 697660 920866
rect 711753 909346 717600 920866
rect 678027 908174 717600 909346
rect 680607 908113 681257 908174
rect 32632 884226 32633 884546
rect 36343 884226 36993 884287
rect 0 883698 39573 884226
rect 0 870890 6491 883698
rect 19296 870890 39573 883698
rect 678027 878146 679077 907854
rect 679397 878146 680287 907854
rect 680607 878207 681257 907793
rect 681577 878146 682467 907854
rect 682787 878146 683677 907854
rect 683997 878146 684647 907854
rect 684968 907600 685617 907854
rect 684967 878400 685617 907600
rect 684968 878146 685617 878400
rect 685937 878146 686827 907854
rect 687147 878146 688947 907854
rect 689267 878146 690117 907854
rect 690437 878146 691287 907854
rect 691607 878146 696597 907854
rect 696917 907600 717600 908174
rect 712757 878400 717600 907600
rect 680607 877826 681257 877887
rect 696917 877826 717600 878400
rect 0 870374 39573 870890
rect 678027 876480 717600 877826
rect 0 869800 20683 870374
rect 32632 870054 32633 870374
rect 36343 870313 36993 870374
rect 0 842600 4843 869800
rect 0 842026 20683 842600
rect 21003 842346 25993 870054
rect 26313 842346 27163 870054
rect 27483 842346 28333 870054
rect 28653 842346 30453 870054
rect 30773 842346 31663 870054
rect 31983 842346 32633 870054
rect 32953 842346 33603 870054
rect 33923 842346 34813 870054
rect 35133 842346 36023 870054
rect 36343 842407 36993 869993
rect 37313 842346 38203 870054
rect 38523 842346 39573 870054
rect 678027 863320 698192 876480
rect 711322 863320 717600 876480
rect 678027 862974 717600 863320
rect 680607 862926 681257 862974
rect 32632 842026 32633 842346
rect 36343 842026 36993 842087
rect 0 841498 39573 842026
rect 0 828690 6491 841498
rect 19296 828690 39573 841498
rect 678027 833146 679077 862654
rect 679397 833146 680287 862654
rect 680607 833207 681257 862606
rect 681577 833146 682467 862654
rect 682787 833146 683677 862654
rect 683997 833146 684647 862654
rect 684968 862400 685617 862654
rect 684967 833146 685617 862400
rect 685937 833146 686827 862654
rect 687147 833146 688947 862654
rect 689267 833146 690117 862654
rect 690437 833146 691287 862654
rect 691607 833146 696597 862654
rect 696917 862400 717600 862974
rect 712757 833400 717600 862400
rect 680607 832826 681257 832887
rect 684967 832826 684968 833146
rect 696917 832826 717600 833400
rect 0 828174 39573 828690
rect 678027 832310 717600 832826
rect 0 827600 20683 828174
rect 32632 827854 32633 828174
rect 36343 828113 36993 828174
rect 0 800400 4843 827600
rect 0 799826 20683 800400
rect 21003 800146 25993 827854
rect 26313 800146 27163 827854
rect 27483 800146 28333 827854
rect 28653 800146 30453 827854
rect 30773 800146 31663 827854
rect 31983 800400 32633 827854
rect 31983 800146 32632 800400
rect 32953 800146 33603 827854
rect 33923 800146 34813 827854
rect 35133 800146 36023 827854
rect 36343 800194 36993 827793
rect 37313 800146 38203 827854
rect 38523 800146 39573 827854
rect 678027 819502 698304 832310
rect 711109 819502 717600 832310
rect 678027 818974 717600 819502
rect 680607 818913 681257 818974
rect 684967 818654 684968 818974
rect 36343 799826 36993 799874
rect 0 799480 39573 799826
rect 0 786320 6278 799480
rect 19408 786320 39573 799480
rect 678027 788946 679077 818654
rect 679397 788946 680287 818654
rect 680607 789007 681257 818593
rect 681577 788946 682467 818654
rect 682787 788946 683677 818654
rect 683997 788946 684647 818654
rect 684967 789200 685617 818654
rect 684968 788946 685617 789200
rect 685937 788946 686827 818654
rect 687147 788946 688947 818654
rect 689267 788946 690117 818654
rect 690437 788946 691287 818654
rect 691607 788946 696597 818654
rect 696917 818400 717600 818974
rect 712757 789200 717600 818400
rect 680607 788626 681257 788687
rect 696917 788626 717600 789200
rect 0 784974 39573 786320
rect 678027 787280 717600 788626
rect 0 784400 20683 784974
rect 36343 784913 36993 784974
rect 0 757200 4843 784400
rect 0 756626 20683 757200
rect 21003 756946 25993 784654
rect 26313 756946 27163 784654
rect 27483 756946 28333 784654
rect 28653 756946 30453 784654
rect 30773 756946 31663 784654
rect 31983 784400 32632 784654
rect 31983 757200 32633 784400
rect 31983 756946 32632 757200
rect 32953 756946 33603 784654
rect 33923 756946 34813 784654
rect 35133 756946 36023 784654
rect 36343 756994 36993 784593
rect 37313 756946 38203 784654
rect 38523 756946 39573 784654
rect 678027 774120 698192 787280
rect 711322 774120 717600 787280
rect 678027 773774 717600 774120
rect 680607 773726 681257 773774
rect 36343 756626 36993 756674
rect 0 756280 39573 756626
rect 0 743120 6278 756280
rect 19408 743120 39573 756280
rect 678027 743946 679077 773454
rect 679397 743946 680287 773454
rect 680607 744007 681257 773406
rect 681577 743946 682467 773454
rect 682787 743946 683677 773454
rect 683997 743946 684647 773454
rect 684968 773200 685617 773454
rect 684967 744200 685617 773200
rect 684968 743946 685617 744200
rect 685937 743946 686827 773454
rect 687147 743946 688947 773454
rect 689267 743946 690117 773454
rect 690437 743946 691287 773454
rect 691607 743946 696597 773454
rect 696917 773200 717600 773774
rect 712757 744200 717600 773200
rect 680607 743626 681257 743687
rect 696917 743626 717600 744200
rect 0 741774 39573 743120
rect 678027 742280 717600 743626
rect 0 741200 20683 741774
rect 36343 741713 36993 741774
rect 0 714000 4843 741200
rect 0 713426 20683 714000
rect 21003 713746 25993 741454
rect 26313 713746 27163 741454
rect 27483 713746 28333 741454
rect 28653 713746 30453 741454
rect 30773 713746 31663 741454
rect 31983 741200 32632 741454
rect 31983 714000 32633 741200
rect 31983 713746 32632 714000
rect 32953 713746 33603 741454
rect 33923 713746 34813 741454
rect 35133 713746 36023 741454
rect 36343 713794 36993 741393
rect 37313 713746 38203 741454
rect 38523 713746 39573 741454
rect 678027 729120 698192 742280
rect 711322 729120 717600 742280
rect 678027 728774 717600 729120
rect 680607 728726 681257 728774
rect 36343 713426 36993 713474
rect 0 713080 39573 713426
rect 0 699920 6278 713080
rect 19408 699920 39573 713080
rect 0 698574 39573 699920
rect 678027 698946 679077 728454
rect 679397 698946 680287 728454
rect 680607 699007 681257 728406
rect 681577 698946 682467 728454
rect 682787 698946 683677 728454
rect 683997 698946 684647 728454
rect 684968 728200 685617 728454
rect 684967 699200 685617 728200
rect 684968 698946 685617 699200
rect 685937 698946 686827 728454
rect 687147 698946 688947 728454
rect 689267 698946 690117 728454
rect 690437 698946 691287 728454
rect 691607 698946 696597 728454
rect 696917 728200 717600 728774
rect 712757 699200 717600 728200
rect 680607 698626 681257 698687
rect 696917 698626 717600 699200
rect 0 698000 20683 698574
rect 36343 698513 36993 698574
rect 0 670800 4843 698000
rect 0 670226 20683 670800
rect 21003 670546 25993 698254
rect 26313 670546 27163 698254
rect 27483 670546 28333 698254
rect 28653 670546 30453 698254
rect 30773 670546 31663 698254
rect 31983 698000 32632 698254
rect 31983 670800 32633 698000
rect 31983 670546 32632 670800
rect 32953 670546 33603 698254
rect 33923 670546 34813 698254
rect 35133 670546 36023 698254
rect 36343 670594 36993 698193
rect 37313 670546 38203 698254
rect 38523 670546 39573 698254
rect 678027 697280 717600 698626
rect 678027 684120 698192 697280
rect 711322 684120 717600 697280
rect 678027 683774 717600 684120
rect 680607 683726 681257 683774
rect 36343 670226 36993 670274
rect 0 669880 39573 670226
rect 0 656720 6278 669880
rect 19408 656720 39573 669880
rect 0 655374 39573 656720
rect 0 654800 20683 655374
rect 36343 655313 36993 655374
rect 0 627600 4843 654800
rect 0 627026 20683 627600
rect 21003 627346 25993 655054
rect 26313 627346 27163 655054
rect 27483 627346 28333 655054
rect 28653 627346 30453 655054
rect 30773 627346 31663 655054
rect 31983 654800 32632 655054
rect 31983 627600 32633 654800
rect 31983 627346 32632 627600
rect 32953 627346 33603 655054
rect 33923 627346 34813 655054
rect 35133 627346 36023 655054
rect 36343 627394 36993 654993
rect 37313 627346 38203 655054
rect 38523 627346 39573 655054
rect 678027 653746 679077 683454
rect 679397 653746 680287 683454
rect 680607 653807 681257 683406
rect 681577 653746 682467 683454
rect 682787 653746 683677 683454
rect 683997 653746 684647 683454
rect 684968 683200 685617 683454
rect 684967 654000 685617 683200
rect 684968 653746 685617 654000
rect 685937 653746 686827 683454
rect 687147 653746 688947 683454
rect 689267 653746 690117 683454
rect 690437 653746 691287 683454
rect 691607 653746 696597 683454
rect 696917 683200 717600 683774
rect 712757 654000 717600 683200
rect 680607 653426 681257 653487
rect 696917 653426 717600 654000
rect 678027 652080 717600 653426
rect 678027 638920 698192 652080
rect 711322 638920 717600 652080
rect 678027 638574 717600 638920
rect 680607 638526 681257 638574
rect 36343 627026 36993 627074
rect 0 626680 39573 627026
rect 0 613520 6278 626680
rect 19408 613520 39573 626680
rect 0 612174 39573 613520
rect 0 611600 20683 612174
rect 36343 612113 36993 612174
rect 0 584400 4843 611600
rect 0 583826 20683 584400
rect 21003 584146 25993 611854
rect 26313 584146 27163 611854
rect 27483 584146 28333 611854
rect 28653 584146 30453 611854
rect 30773 584146 31663 611854
rect 31983 611600 32632 611854
rect 31983 584400 32633 611600
rect 31983 584146 32632 584400
rect 32953 584146 33603 611854
rect 33923 584146 34813 611854
rect 35133 584146 36023 611854
rect 36343 584194 36993 611793
rect 37313 584146 38203 611854
rect 38523 584146 39573 611854
rect 678027 608746 679077 638254
rect 679397 608746 680287 638254
rect 680607 608807 681257 638206
rect 681577 608746 682467 638254
rect 682787 608746 683677 638254
rect 683997 608746 684647 638254
rect 684968 638000 685617 638254
rect 684967 609000 685617 638000
rect 684968 608746 685617 609000
rect 685937 608746 686827 638254
rect 687147 608746 688947 638254
rect 689267 608746 690117 638254
rect 690437 608746 691287 638254
rect 691607 608746 696597 638254
rect 696917 638000 717600 638574
rect 712757 609000 717600 638000
rect 680607 608426 681257 608487
rect 696917 608426 717600 609000
rect 678027 607080 717600 608426
rect 678027 593920 698192 607080
rect 711322 593920 717600 607080
rect 678027 593574 717600 593920
rect 680607 593526 681257 593574
rect 36343 583826 36993 583874
rect 0 583480 39573 583826
rect 0 570320 6278 583480
rect 19408 570320 39573 583480
rect 0 568974 39573 570320
rect 0 568400 20683 568974
rect 36343 568913 36993 568974
rect 0 541200 4843 568400
rect 0 540626 20683 541200
rect 21003 540946 25993 568654
rect 26313 540946 27163 568654
rect 27483 540946 28333 568654
rect 28653 540946 30453 568654
rect 30773 540946 31663 568654
rect 31983 568400 32632 568654
rect 31983 541200 32633 568400
rect 31983 540946 32632 541200
rect 32953 540946 33603 568654
rect 33923 540946 34813 568654
rect 35133 540946 36023 568654
rect 36343 540994 36993 568593
rect 37313 540946 38203 568654
rect 38523 540946 39573 568654
rect 678027 563546 679077 593254
rect 679397 563546 680287 593254
rect 680607 563607 681257 593206
rect 681577 563546 682467 593254
rect 682787 563546 683677 593254
rect 683997 563546 684647 593254
rect 684968 593000 685617 593254
rect 684967 563800 685617 593000
rect 684968 563546 685617 563800
rect 685937 563546 686827 593254
rect 687147 563546 688947 593254
rect 689267 563546 690117 593254
rect 690437 563546 691287 593254
rect 691607 563546 696597 593254
rect 696917 593000 717600 593574
rect 712757 563800 717600 593000
rect 680607 563226 681257 563287
rect 696917 563226 717600 563800
rect 678027 561880 717600 563226
rect 678027 548720 698192 561880
rect 711322 548720 717600 561880
rect 678027 548374 717600 548720
rect 680607 548326 681257 548374
rect 36343 540626 36993 540674
rect 0 540280 39573 540626
rect 0 527120 6278 540280
rect 19408 527120 39573 540280
rect 0 525774 39573 527120
rect 0 525200 20683 525774
rect 36343 525713 36993 525774
rect 0 498000 4843 525200
rect 0 497426 20683 498000
rect 21003 497746 25993 525454
rect 26313 497746 27163 525454
rect 27483 497746 28333 525454
rect 28653 497746 30453 525454
rect 30773 497746 31663 525454
rect 31983 525200 32632 525454
rect 31983 497746 32633 525200
rect 32953 497746 33603 525454
rect 33923 497746 34813 525454
rect 35133 497746 36023 525454
rect 36343 497807 36993 525393
rect 37313 497746 38203 525454
rect 38523 497746 39573 525454
rect 678027 518546 679077 548054
rect 679397 518546 680287 548054
rect 680607 518607 681257 548006
rect 681577 518546 682467 548054
rect 682787 518546 683677 548054
rect 683997 518546 684647 548054
rect 684968 547800 685617 548054
rect 684967 518546 685617 547800
rect 685937 518546 686827 548054
rect 687147 518546 688947 548054
rect 689267 518546 690117 548054
rect 690437 518546 691287 548054
rect 691607 518546 696597 548054
rect 696917 547800 717600 548374
rect 712757 518800 717600 547800
rect 680607 518226 681257 518287
rect 684967 518226 684968 518546
rect 696917 518226 717600 518800
rect 678027 517710 717600 518226
rect 678027 504902 698304 517710
rect 711109 504902 717600 517710
rect 678027 504374 717600 504902
rect 680607 504313 681257 504374
rect 684967 504054 684968 504374
rect 32632 497426 32633 497746
rect 36343 497426 36993 497487
rect 0 496898 39573 497426
rect 0 484090 6491 496898
rect 19296 484090 39573 496898
rect 0 483574 39573 484090
rect 0 483000 20683 483574
rect 32632 483254 32633 483574
rect 36343 483513 36993 483574
rect 0 455800 4843 483000
rect 0 455226 20683 455800
rect 21003 455546 25993 483254
rect 26313 455546 27163 483254
rect 27483 455546 28333 483254
rect 28653 455546 30453 483254
rect 30773 455546 31663 483254
rect 31983 455800 32633 483254
rect 31983 455546 32632 455800
rect 32953 455546 33603 483254
rect 33923 455546 34813 483254
rect 35133 455546 36023 483254
rect 36343 455607 36993 483193
rect 37313 455546 38203 483254
rect 38523 455546 39573 483254
rect 678027 474546 679077 504054
rect 679397 474546 680287 504054
rect 680607 474607 681257 503993
rect 681577 474546 682467 504054
rect 682787 474546 683677 504054
rect 683997 474546 684647 504054
rect 684967 474800 685617 504054
rect 684968 474546 685617 474800
rect 685937 474546 686827 504054
rect 687147 474546 688947 504054
rect 689267 474546 690117 504054
rect 690437 474546 691287 504054
rect 691607 474546 696597 504054
rect 696917 503800 717600 504374
rect 712757 474800 717600 503800
rect 680607 474226 681257 474287
rect 696917 474226 717600 474800
rect 678027 473066 717600 474226
rect 678027 461546 697660 473066
rect 711753 461546 717600 473066
rect 678027 460374 717600 461546
rect 680607 460313 681257 460374
rect 36343 455226 36993 455287
rect 0 454054 39573 455226
rect 0 442534 5847 454054
rect 19940 442534 39573 454054
rect 0 441374 39573 442534
rect 0 440800 20683 441374
rect 36343 441313 36993 441374
rect 0 413600 4843 440800
rect 0 413026 20683 413600
rect 21003 413346 25993 441054
rect 26313 413346 27163 441054
rect 27483 413346 28333 441054
rect 28653 413346 30453 441054
rect 30773 413346 31663 441054
rect 31983 440800 32632 441054
rect 31983 413600 32633 440800
rect 31983 413346 32632 413600
rect 32953 413346 33603 441054
rect 33923 413346 34813 441054
rect 35133 413346 36023 441054
rect 36343 413394 36993 440993
rect 37313 413346 38203 441054
rect 38523 413346 39573 441054
rect 678027 430346 679077 460054
rect 679397 430346 680287 460054
rect 680607 430407 681257 459993
rect 681577 430346 682467 460054
rect 682787 430346 683677 460054
rect 683997 430346 684647 460054
rect 684968 459800 685617 460054
rect 684967 430346 685617 459800
rect 685937 430346 686827 460054
rect 687147 430346 688947 460054
rect 689267 430346 690117 460054
rect 690437 430346 691287 460054
rect 691607 430346 696597 460054
rect 696917 459800 717600 460374
rect 712757 430600 717600 459800
rect 680607 430026 681257 430087
rect 684967 430026 684968 430346
rect 696917 430026 717600 430600
rect 678027 429510 717600 430026
rect 678027 416702 698304 429510
rect 711109 416702 717600 429510
rect 678027 416174 717600 416702
rect 680607 416113 681257 416174
rect 684967 415854 684968 416174
rect 36343 413026 36993 413074
rect 0 412680 39573 413026
rect 0 399520 6278 412680
rect 19408 399520 39573 412680
rect 0 398174 39573 399520
rect 0 397600 20683 398174
rect 36343 398113 36993 398174
rect 0 370400 4843 397600
rect 0 369826 20683 370400
rect 21003 370146 25993 397854
rect 26313 370146 27163 397854
rect 27483 370146 28333 397854
rect 28653 370146 30453 397854
rect 30773 370146 31663 397854
rect 31983 397600 32632 397854
rect 31983 370400 32633 397600
rect 31983 370146 32632 370400
rect 32953 370146 33603 397854
rect 33923 370146 34813 397854
rect 35133 370146 36023 397854
rect 36343 370194 36993 397793
rect 37313 370146 38203 397854
rect 38523 370146 39573 397854
rect 678027 386346 679077 415854
rect 679397 386346 680287 415854
rect 680607 386407 681257 415793
rect 681577 386346 682467 415854
rect 682787 386346 683677 415854
rect 683997 386346 684647 415854
rect 684967 386600 685617 415854
rect 684968 386346 685617 386600
rect 685937 386346 686827 415854
rect 687147 386346 688947 415854
rect 689267 386346 690117 415854
rect 690437 386346 691287 415854
rect 691607 386346 696597 415854
rect 696917 415600 717600 416174
rect 712757 386600 717600 415600
rect 680607 386026 681257 386087
rect 696917 386026 717600 386600
rect 678027 384680 717600 386026
rect 678027 371520 698192 384680
rect 711322 371520 717600 384680
rect 678027 371174 717600 371520
rect 680607 371126 681257 371174
rect 36343 369826 36993 369874
rect 0 369480 39573 369826
rect 0 356320 6278 369480
rect 19408 356320 39573 369480
rect 0 354974 39573 356320
rect 0 354400 20683 354974
rect 36343 354913 36993 354974
rect 0 327200 4843 354400
rect 0 326626 20683 327200
rect 21003 326946 25993 354654
rect 26313 326946 27163 354654
rect 27483 326946 28333 354654
rect 28653 326946 30453 354654
rect 30773 326946 31663 354654
rect 31983 354400 32632 354654
rect 31983 327200 32633 354400
rect 31983 326946 32632 327200
rect 32953 326946 33603 354654
rect 33923 326946 34813 354654
rect 35133 326946 36023 354654
rect 36343 326994 36993 354593
rect 37313 326946 38203 354654
rect 38523 326946 39573 354654
rect 678027 341146 679077 370854
rect 679397 341146 680287 370854
rect 680607 341207 681257 370806
rect 681577 341146 682467 370854
rect 682787 341146 683677 370854
rect 683997 341146 684647 370854
rect 684968 370600 685617 370854
rect 684967 341400 685617 370600
rect 684968 341146 685617 341400
rect 685937 341146 686827 370854
rect 687147 341146 688947 370854
rect 689267 341146 690117 370854
rect 690437 341146 691287 370854
rect 691607 341146 696597 370854
rect 696917 370600 717600 371174
rect 712757 341400 717600 370600
rect 680607 340826 681257 340887
rect 696917 340826 717600 341400
rect 678027 339480 717600 340826
rect 36343 326626 36993 326674
rect 0 326280 39573 326626
rect 0 313120 6278 326280
rect 19408 313120 39573 326280
rect 678027 326320 698192 339480
rect 711322 326320 717600 339480
rect 678027 325974 717600 326320
rect 680607 325926 681257 325974
rect 0 311774 39573 313120
rect 0 311200 20683 311774
rect 36343 311713 36993 311774
rect 0 284000 4843 311200
rect 0 283426 20683 284000
rect 21003 283746 25993 311454
rect 26313 283746 27163 311454
rect 27483 283746 28333 311454
rect 28653 283746 30453 311454
rect 30773 283746 31663 311454
rect 31983 311200 32632 311454
rect 31983 284000 32633 311200
rect 31983 283746 32632 284000
rect 32953 283746 33603 311454
rect 33923 283746 34813 311454
rect 35133 283746 36023 311454
rect 36343 283794 36993 311393
rect 37313 283746 38203 311454
rect 38523 283746 39573 311454
rect 678027 296146 679077 325654
rect 679397 296146 680287 325654
rect 680607 296207 681257 325606
rect 681577 296146 682467 325654
rect 682787 296146 683677 325654
rect 683997 296146 684647 325654
rect 684968 325400 685617 325654
rect 684967 296400 685617 325400
rect 684968 296146 685617 296400
rect 685937 296146 686827 325654
rect 687147 296146 688947 325654
rect 689267 296146 690117 325654
rect 690437 296146 691287 325654
rect 691607 296146 696597 325654
rect 696917 325400 717600 325974
rect 712757 296400 717600 325400
rect 680607 295826 681257 295887
rect 696917 295826 717600 296400
rect 678027 294480 717600 295826
rect 36343 283426 36993 283474
rect 0 283080 39573 283426
rect 0 269920 6278 283080
rect 19408 269920 39573 283080
rect 678027 281320 698192 294480
rect 711322 281320 717600 294480
rect 678027 280974 717600 281320
rect 680607 280926 681257 280974
rect 0 268574 39573 269920
rect 0 268000 20683 268574
rect 36343 268513 36993 268574
rect 0 240800 4843 268000
rect 0 240226 20683 240800
rect 21003 240546 25993 268254
rect 26313 240546 27163 268254
rect 27483 240546 28333 268254
rect 28653 240546 30453 268254
rect 30773 240546 31663 268254
rect 31983 268000 32632 268254
rect 31983 240800 32633 268000
rect 31983 240546 32632 240800
rect 32953 240546 33603 268254
rect 33923 240546 34813 268254
rect 35133 240546 36023 268254
rect 36343 240594 36993 268193
rect 37313 240546 38203 268254
rect 38523 240546 39573 268254
rect 678027 251146 679077 280654
rect 679397 251146 680287 280654
rect 680607 251207 681257 280606
rect 681577 251146 682467 280654
rect 682787 251146 683677 280654
rect 683997 251146 684647 280654
rect 684968 280400 685617 280654
rect 684967 251400 685617 280400
rect 684968 251146 685617 251400
rect 685937 251146 686827 280654
rect 687147 251146 688947 280654
rect 689267 251146 690117 280654
rect 690437 251146 691287 280654
rect 691607 251146 696597 280654
rect 696917 280400 717600 280974
rect 712757 251400 717600 280400
rect 680607 250826 681257 250887
rect 696917 250826 717600 251400
rect 678027 249480 717600 250826
rect 36343 240226 36993 240274
rect 0 239880 39573 240226
rect 0 226720 6278 239880
rect 19408 226720 39573 239880
rect 678027 236320 698192 249480
rect 711322 236320 717600 249480
rect 678027 235974 717600 236320
rect 680607 235926 681257 235974
rect 0 225374 39573 226720
rect 0 224800 20683 225374
rect 36343 225313 36993 225374
rect 0 197600 4843 224800
rect 0 197026 20683 197600
rect 21003 197346 25993 225054
rect 26313 197346 27163 225054
rect 27483 197346 28333 225054
rect 28653 197346 30453 225054
rect 30773 197346 31663 225054
rect 31983 224800 32632 225054
rect 31983 197600 32633 224800
rect 31983 197346 32632 197600
rect 32953 197346 33603 225054
rect 33923 197346 34813 225054
rect 35133 197346 36023 225054
rect 36343 197394 36993 224993
rect 37313 197346 38203 225054
rect 38523 197346 39573 225054
rect 678027 205946 679077 235654
rect 679397 205946 680287 235654
rect 680607 206007 681257 235606
rect 681577 205946 682467 235654
rect 682787 205946 683677 235654
rect 683997 205946 684647 235654
rect 684968 235400 685617 235654
rect 684967 206200 685617 235400
rect 684968 205946 685617 206200
rect 685937 205946 686827 235654
rect 687147 205946 688947 235654
rect 689267 205946 690117 235654
rect 690437 205946 691287 235654
rect 691607 205946 696597 235654
rect 696917 235400 717600 235974
rect 712757 206200 717600 235400
rect 680607 205626 681257 205687
rect 696917 205626 717600 206200
rect 678027 204280 717600 205626
rect 36343 197026 36993 197074
rect 0 196680 39573 197026
rect 0 183520 6278 196680
rect 19408 183520 39573 196680
rect 678027 191120 698192 204280
rect 711322 191120 717600 204280
rect 678027 190774 717600 191120
rect 680607 190726 681257 190774
rect 0 182174 39573 183520
rect 0 181600 20683 182174
rect 36343 182113 36993 182174
rect 0 125200 4843 181600
rect 0 124626 20683 125200
rect 21003 124946 25993 181854
rect 26313 124946 27163 181854
rect 27483 124946 28333 181854
rect 28653 153400 30453 181854
rect 30773 154400 31663 181854
rect 31983 181600 32632 181854
rect 31983 153400 32633 181600
rect 28653 124946 30453 152400
rect 30773 124946 31663 153400
rect 31983 124946 32633 152400
rect 32953 124946 33603 181854
rect 33923 124946 34813 181854
rect 35133 124946 36023 181854
rect 36343 153400 36993 181793
rect 37313 154400 38203 181854
rect 36343 125007 36993 152400
rect 37313 124946 38203 153400
rect 38523 124946 39573 181854
rect 678027 160946 679077 190454
rect 679397 160946 680287 190454
rect 680607 161007 681257 190406
rect 681577 160946 682467 190454
rect 682787 160946 683677 190454
rect 683997 160946 684647 190454
rect 684968 190200 685617 190454
rect 684967 161200 685617 190200
rect 684968 160946 685617 161200
rect 685937 160946 686827 190454
rect 687147 160946 688947 190454
rect 689267 160946 690117 190454
rect 690437 160946 691287 190454
rect 691607 160946 696597 190454
rect 696917 190200 717600 190774
rect 712757 161200 717600 190200
rect 680607 160626 681257 160687
rect 696917 160626 717600 161200
rect 678027 159280 717600 160626
rect 678027 146120 698192 159280
rect 711322 146120 717600 159280
rect 678027 145774 717600 146120
rect 680607 145726 681257 145774
rect 32632 124626 32633 124946
rect 36343 124626 36993 124687
rect 0 124098 39573 124626
rect 0 111290 6491 124098
rect 19296 111290 39573 124098
rect 678027 115746 679077 145454
rect 679397 115746 680287 145454
rect 680607 115807 681257 145406
rect 681577 115746 682467 145454
rect 682787 115746 683677 145454
rect 683997 115746 684647 145454
rect 684968 145200 685617 145454
rect 684967 116000 685617 145200
rect 684968 115746 685617 116000
rect 685937 115746 686827 145454
rect 687147 115746 688947 145454
rect 689267 115746 690117 145454
rect 690437 115746 691287 145454
rect 691607 115746 696597 145454
rect 696917 145200 717600 145774
rect 712757 116000 717600 145200
rect 680607 115426 681257 115487
rect 696917 115426 717600 116000
rect 0 110774 39573 111290
rect 678027 114080 717600 115426
rect 0 110200 20683 110774
rect 32632 110454 32633 110774
rect 36343 110713 36993 110774
rect 0 83000 4843 110200
rect 0 82426 20683 83000
rect 21003 82746 25993 110454
rect 26313 82746 27163 110454
rect 27483 82746 28333 110454
rect 28653 82746 30453 110454
rect 30773 82746 31663 110454
rect 31983 82746 32633 110454
rect 32953 82746 33603 110454
rect 33923 82746 34813 110454
rect 35133 82746 36023 110454
rect 36343 82807 36993 110393
rect 37313 82746 38203 110454
rect 38523 82746 39573 110454
rect 678027 100920 698192 114080
rect 711322 100920 717600 114080
rect 678027 100574 717600 100920
rect 680607 100526 681257 100574
rect 32632 82426 32633 82746
rect 36343 82426 36993 82487
rect 0 81254 39573 82426
rect 0 69734 5847 81254
rect 19940 69734 39573 81254
rect 0 68574 39573 69734
rect 0 68000 20683 68574
rect 32632 68254 32633 68574
rect 36343 68513 36993 68574
rect 0 40800 4843 68000
rect 0 40109 20683 40800
rect 21003 40429 25993 68254
rect 26313 40546 27163 68254
rect 27483 40546 28333 68254
rect 26313 40109 28333 40226
rect 0 35049 28333 40109
rect 28653 35369 30453 68254
rect 30773 40546 31663 68254
rect 31983 40800 32633 68254
rect 31983 40546 32632 40800
rect 32953 40546 33603 68254
rect 33923 40546 34813 68254
rect 35133 40546 36023 68254
rect 36343 40549 36993 68193
rect 37313 40546 38203 68254
rect 38523 40546 39573 68254
rect 36343 40226 36993 40229
rect 39893 40226 40000 40800
rect 30773 39893 40000 40226
rect 676800 39893 677707 40000
rect 30773 38523 39210 39893
rect 39573 39573 39680 39893
tri 39680 39573 40000 39893 sw
rect 677374 39680 677707 39893
tri 677707 39680 678027 40000 se
rect 678027 39680 679077 100254
rect 679397 71000 680287 100254
rect 680607 70000 681257 100206
rect 677374 39573 679077 39680
rect 39530 38523 79054 39573
rect 30773 36993 38923 38523
rect 47400 38203 71400 38523
rect 39243 37313 79054 38203
rect 79374 36993 93226 39573
rect 93546 38523 132854 39573
rect 133174 38523 186654 39573
rect 101200 38203 125200 38523
rect 133174 38203 147600 38523
rect 155000 38203 179000 38523
rect 93546 37313 132854 38203
rect 133174 37313 186654 38203
rect 133174 36993 147600 37313
rect 186974 36993 201826 39573
rect 202146 38523 241454 39573
rect 209800 38203 233800 38523
rect 202146 37313 241454 38203
rect 241774 36993 255626 39573
rect 255946 38523 295254 39573
rect 263600 38203 287600 38523
rect 255946 37313 295254 38203
rect 295574 36993 310426 39573
rect 310746 38523 350054 39573
rect 318400 38203 342400 38523
rect 310746 37313 350054 38203
rect 350374 36993 365226 39573
rect 365546 38523 404854 39573
rect 373200 38203 397200 38523
rect 365546 37313 404854 38203
rect 405174 36993 420026 39573
rect 420346 38523 459654 39573
rect 428000 38203 452000 38523
rect 420346 37313 459654 38203
rect 459974 36993 474826 39573
rect 475146 38523 514454 39573
rect 482800 38203 506800 38523
rect 475146 37313 514454 38203
rect 514774 36993 529626 39573
rect 529946 38523 569254 39573
rect 537600 38203 561600 38523
rect 529946 37313 569254 38203
rect 569574 36993 583426 39573
rect 583746 38523 623054 39573
rect 591400 38203 615400 38523
rect 583746 37313 623054 38203
rect 623374 36993 637226 39573
rect 637546 38523 677054 39573
rect 677374 39210 677707 39573
rect 678027 39530 679077 39573
rect 679397 39243 680287 70000
rect 680607 39706 681257 69000
rect 681577 39695 682467 100254
rect 682787 39680 683677 100254
rect 683997 39723 684647 100254
rect 684968 100000 685617 100254
rect 684967 70000 685617 100000
rect 685937 71000 686827 100254
rect 687147 70000 688947 100254
rect 684967 39733 685617 69000
rect 685937 39705 686827 70000
rect 684967 39403 685617 39413
rect 680607 39375 681257 39386
rect 683997 39385 685617 39403
rect 680607 39360 682467 39375
rect 683997 39360 686827 39385
rect 677374 38923 679077 39210
rect 680607 38923 686827 39360
rect 645200 38203 669200 38523
rect 637546 37313 677054 38203
rect 677374 36993 686827 38923
rect 30773 36343 39386 36993
rect 39706 36343 78993 36993
rect 79313 36343 93287 36993
rect 133113 36343 186606 36993
rect 186926 36343 201887 36993
rect 202207 36343 241393 36993
rect 241713 36343 255687 36993
rect 256007 36343 295206 36993
rect 295526 36343 310487 36993
rect 310807 36343 350006 36993
rect 350326 36343 365287 36993
rect 365607 36343 404806 36993
rect 405126 36343 420087 36993
rect 420407 36343 459606 36993
rect 459926 36343 474887 36993
rect 475207 36343 514406 36993
rect 514726 36343 529687 36993
rect 530007 36343 569193 36993
rect 569513 36343 583487 36993
rect 583807 36343 622993 36993
rect 623313 36343 637287 36993
rect 637607 36343 677051 36993
rect 677371 36343 686827 36993
rect 30773 35133 39375 36343
rect 39695 35133 79054 36023
rect 30773 35049 39360 35133
rect 0 33603 39360 35049
rect 39680 33923 79054 34813
rect 0 32633 39403 33603
rect 39723 32953 79054 33603
rect 79374 32633 93226 36343
rect 133113 36023 147600 36343
rect 93546 35133 186654 36023
rect 133174 34813 147600 35133
rect 93546 33923 132854 34813
rect 133174 33923 186654 34813
rect 133174 33603 147600 33923
rect 93546 32953 132854 33603
rect 133174 32953 186654 33603
rect 133174 32633 147600 32953
rect 0 31983 39413 32633
rect 39733 32632 186400 32633
rect 39733 31983 79054 32632
rect 0 30773 39385 31983
rect 39705 30773 79054 31663
rect 0 28333 35049 30773
rect 35369 28653 79054 30453
rect 0 27163 39355 28333
rect 39675 27483 79054 28333
rect 0 26313 39384 27163
rect 39704 26313 79054 27163
rect 0 20683 39151 26313
rect 39471 21003 79054 25993
rect 79374 20683 93226 32632
rect 93546 31983 186654 32632
rect 133174 31663 147600 31983
rect 133174 30773 186654 31663
rect 133174 30453 147600 30773
rect 133174 28653 186654 30453
rect 133174 28333 147600 28653
rect 93546 27483 132854 28333
rect 133174 27483 186654 28333
rect 133174 27163 147600 27483
rect 93546 26313 132854 27163
rect 133174 26313 186654 27163
rect 133174 25993 147600 26313
rect 93546 21003 132854 25993
rect 133174 21003 186654 25993
rect 133174 20683 147600 21003
rect 186974 20683 201826 36343
rect 202146 35133 241454 36023
rect 202146 33923 241454 34813
rect 202146 32953 241454 33603
rect 241774 32633 255626 36343
rect 255946 35133 295254 36023
rect 255946 33923 295254 34813
rect 255946 32953 295254 33603
rect 202400 32632 295000 32633
rect 202146 31983 241454 32632
rect 202146 30773 241454 31663
rect 202146 28653 241454 30453
rect 202146 27483 241454 28333
rect 202146 26313 241454 27163
rect 202146 21003 241454 25993
rect 241774 20683 255626 32632
rect 255946 31983 295254 32632
rect 255946 30773 295254 31663
rect 255946 28653 295254 30453
rect 255946 27483 295254 28333
rect 255946 26313 295254 27163
rect 255946 21003 295254 25993
rect 295574 20683 310426 36343
rect 310746 35133 350054 36023
rect 310746 33923 350054 34813
rect 310746 32953 350054 33603
rect 311000 32632 349800 32633
rect 310746 31983 350054 32632
rect 310746 30773 350054 31663
rect 310746 28653 350054 30453
rect 310746 27483 350054 28333
rect 310746 26313 350054 27163
rect 310746 21003 350054 25993
rect 350374 20683 365226 36343
rect 365546 35133 404854 36023
rect 365546 33923 404854 34813
rect 365546 32953 404854 33603
rect 365800 32632 404600 32633
rect 365546 31983 404854 32632
rect 365546 30773 404854 31663
rect 365546 28653 404854 30453
rect 365546 27483 404854 28333
rect 365546 26313 404854 27163
rect 365546 21003 404854 25993
rect 405174 20683 420026 36343
rect 420346 35133 459654 36023
rect 420346 33923 459654 34813
rect 420346 32953 459654 33603
rect 420600 32632 459400 32633
rect 420346 31983 459654 32632
rect 420346 30773 459654 31663
rect 420346 28653 459654 30453
rect 420346 27483 459654 28333
rect 420346 26313 459654 27163
rect 420346 21003 459654 25993
rect 459974 20683 474826 36343
rect 475146 35133 514454 36023
rect 475146 33923 514454 34813
rect 475146 32953 514454 33603
rect 475400 32632 514200 32633
rect 475146 31983 514454 32632
rect 475146 30773 514454 31663
rect 475146 28653 514454 30453
rect 475146 27483 514454 28333
rect 475146 26313 514454 27163
rect 475146 21003 514454 25993
rect 514774 20683 529626 36343
rect 529946 35133 569254 36023
rect 529946 33923 569254 34813
rect 529946 32953 569254 33603
rect 569574 32633 583426 36343
rect 583746 35133 623054 36023
rect 583746 33923 623054 34813
rect 583746 32953 623054 33603
rect 623374 32633 637226 36343
rect 637546 35133 677054 36023
rect 677374 35049 686827 36343
rect 687147 35369 688947 69000
rect 689267 39675 690117 100254
rect 690437 39704 691287 100254
rect 691607 39471 696597 100254
rect 696917 100000 717600 100574
rect 712757 40000 717600 100000
rect 690437 39355 691287 39384
rect 689267 39151 691287 39355
rect 696917 39151 717600 40000
rect 689267 35049 717600 39151
rect 637546 33923 677054 34813
rect 637546 32953 677054 33603
rect 530200 32632 676800 32633
rect 529946 31983 569254 32632
rect 529946 30773 569254 31663
rect 529946 28653 569254 30453
rect 529946 27483 569254 28333
rect 529946 26313 569254 27163
rect 529946 21003 569254 25993
rect 569574 20683 583426 32632
rect 583746 31983 623054 32632
rect 583746 30773 623054 31663
rect 583746 28653 623054 30453
rect 583746 27483 623054 28333
rect 583746 26313 623054 27163
rect 583746 21003 623054 25993
rect 623374 20683 637226 32632
rect 637546 31983 677054 32632
rect 637546 30773 677054 31663
rect 677374 30773 717600 35049
rect 637546 28653 682231 30453
rect 682551 28333 717600 30773
rect 637546 27483 677054 28333
rect 637546 26313 677054 27163
rect 677374 26313 717600 28333
rect 637546 21003 677171 25993
rect 677491 20683 717600 26313
rect 0 4843 40000 20683
rect 78800 19296 93800 20683
rect 78800 6491 79902 19296
rect 92710 6491 93800 19296
rect 78800 4843 93800 6491
rect 132600 19518 147600 20683
rect 132600 6355 133520 19518
rect 146700 6355 147600 19518
rect 132600 4843 147600 6355
rect 186400 19408 202400 20683
rect 186400 6278 187320 19408
rect 200480 6278 202400 19408
rect 186400 4843 202400 6278
rect 241200 19940 256200 20683
rect 241200 5847 242946 19940
rect 254466 5847 256200 19940
rect 241200 4843 256200 5847
rect 295000 19408 311000 20683
rect 295000 6278 295920 19408
rect 309080 6278 311000 19408
rect 295000 4843 311000 6278
rect 349800 19408 365800 20683
rect 349800 6278 350720 19408
rect 363880 6278 365800 19408
rect 349800 4843 365800 6278
rect 404600 19408 420600 20683
rect 404600 6278 405520 19408
rect 418680 6278 420600 19408
rect 404600 4843 420600 6278
rect 459400 19408 475400 20683
rect 459400 6278 460320 19408
rect 473480 6278 475400 19408
rect 459400 4843 475400 6278
rect 514200 19408 530200 20683
rect 514200 6278 515120 19408
rect 528280 6278 530200 19408
rect 514200 4843 530200 6278
rect 569000 19296 584000 20683
rect 569000 6491 570102 19296
rect 582910 6491 584000 19296
rect 569000 4843 584000 6491
rect 622800 19296 637800 20683
rect 622800 6491 623902 19296
rect 636710 6491 637800 19296
rect 622800 4843 637800 6491
rect 676800 4843 717600 20683
rect 0 0 717600 4843
<< labels >>
rlabel metal5 s 187640 6598 200160 19088 6 clock
port 1 nsew signal input
rlabel metal2 s 187327 41713 187383 42193 6 clock_core
port 2 nsew signal output
rlabel metal2 s 194043 41713 194099 42193 6 por
port 3 nsew signal input
rlabel metal5 s 351040 6598 363560 19088 6 flash_clk
port 4 nsew signal output
rlabel metal2 s 361767 41713 361823 42193 6 flash_clk_core
port 5 nsew signal input
rlabel metal2 s 357443 41713 357499 42193 6 flash_clk_ieb_core
port 6 nsew signal input
rlabel metal2 s 364895 41713 364951 42193 6 flash_clk_oeb_core
port 7 nsew signal input
rlabel metal5 s 296240 6598 308760 19088 6 flash_csb
port 8 nsew signal output
rlabel metal2 s 306967 41713 307023 42193 6 flash_csb_core
port 9 nsew signal input
rlabel metal2 s 302643 41713 302699 42193 6 flash_csb_ieb_core
port 10 nsew signal input
rlabel metal2 s 310095 41713 310151 42193 6 flash_csb_oeb_core
port 11 nsew signal input
rlabel metal5 s 405840 6598 418360 19088 6 flash_io0
port 12 nsew signal bidirectional
rlabel metal2 s 405527 41713 405583 42193 6 flash_io0_di_core
port 13 nsew signal output
rlabel metal2 s 416567 41713 416623 42193 6 flash_io0_do_core
port 14 nsew signal input
rlabel metal2 s 415371 41713 415427 41806 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 415216 41754 415268 41806 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 415216 41806 415427 41818 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 412364 41754 412416 41806 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 412243 41713 412299 41806 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 412243 41806 412416 41818 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 409328 41754 409380 41806 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 409207 41713 409263 41806 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 409207 41806 409380 41818 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 415228 41818 415427 41834 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 412243 41818 412404 41834 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 409207 41818 409368 41834 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 415371 41834 415427 42193 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 412243 41834 412299 42193 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 409207 41834 409263 42193 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel via1 s 415216 41760 415268 41812 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel via1 s 412364 41760 412416 41812 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel via1 s 409328 41760 409380 41812 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 415210 41760 415274 41772 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 412358 41760 412422 41772 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 409322 41760 409386 41772 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 409322 41772 415274 41800 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 415210 41800 415274 41812 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 412358 41800 412422 41812 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 409322 41800 409386 41812 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal3 s 419717 44235 419783 44238 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal3 s 419490 44238 419783 44298 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal3 s 419717 44298 419783 44301 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal3 s 419490 44298 419550 44374 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal3 s 411069 44371 411135 44374 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal3 s 411069 44374 419550 44434 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal3 s 411069 44434 411135 44437 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel via2 s 419722 44240 419778 44296 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel via2 s 411074 44376 411130 44432 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 419695 41713 419751 41820 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 411047 41713 411103 41820 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 419695 41820 419764 42193 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 411047 41820 411116 42193 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 419736 42193 419764 44231 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 419722 44231 419778 44305 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 411088 42193 411116 44367 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 411074 44367 411130 44441 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal5 s 460640 6598 473160 19088 6 flash_io1
port 17 nsew signal bidirectional
rlabel metal2 s 460327 41713 460383 42193 6 flash_io1_di_core
port 18 nsew signal output
rlabel metal2 s 471367 41713 471423 42193 6 flash_io1_do_core
port 19 nsew signal input
rlabel metal2 s 470171 41713 470227 41806 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 470048 41754 470100 41806 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 470048 41806 470227 41818 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 467196 41754 467248 41806 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 467043 41713 467099 41806 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 467043 41806 467248 41818 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 464160 41754 464212 41806 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 464007 41713 464063 41806 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 464007 41806 464212 41818 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 470060 41818 470227 41834 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 467043 41818 467236 41834 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 464007 41818 464200 41834 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 470171 41834 470227 42193 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 467043 41834 467099 42193 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 464007 41834 464063 42193 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel via1 s 470048 41760 470100 41812 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel via1 s 467196 41760 467248 41812 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel via1 s 464160 41760 464212 41812 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 470042 41760 470106 41772 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 467190 41760 467254 41772 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 464154 41760 464218 41772 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 464154 41772 470106 41800 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 470042 41800 470106 41812 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 467190 41800 467254 41812 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 464154 41800 464218 41812 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal3 s 474457 44371 474523 44374 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal3 s 465809 44371 465875 44374 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal3 s 465809 44374 474523 44434 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal3 s 474457 44434 474523 44437 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal3 s 465809 44434 465875 44437 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel via2 s 474462 44376 474518 44432 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel via2 s 465814 44376 465870 44432 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 474495 41713 474551 41806 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 465847 41713 465903 41806 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 474476 41806 474551 42193 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 465828 41806 465903 42193 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 474476 42193 474504 44367 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 465828 42193 465856 44367 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 474462 44367 474518 44441 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 465814 44367 465870 44441 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal5 s 515440 6598 527960 19088 6 gpio
port 22 nsew signal bidirectional
rlabel metal2 s 515127 41713 515183 42193 6 gpio_in_core
port 23 nsew signal output
rlabel metal2 s 521843 41713 521899 42193 6 gpio_inenb_core
port 24 nsew signal input
rlabel metal2 s 520647 41713 520703 42193 6 gpio_mode0_core
port 25 nsew signal input
rlabel metal3 s 524965 44235 525031 44238 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal3 s 518801 44235 518867 44238 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal3 s 518801 44238 525031 44298 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal3 s 524965 44298 525031 44301 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal3 s 518801 44298 518867 44301 6 gpio_mode1_core
port 26 nsew signal input
rlabel via2 s 524970 44240 525026 44296 6 gpio_mode1_core
port 26 nsew signal input
rlabel via2 s 518806 44240 518862 44296 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 524971 41713 525027 42193 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 518807 41713 518863 42193 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 524984 42193 525012 44231 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 518820 42193 518848 44231 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 524970 44231 525026 44305 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 518806 44231 518862 44305 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 526167 41713 526223 42193 6 gpio_out_core
port 27 nsew signal input
rlabel metal2 s 529295 41713 529351 42193 6 gpio_outenb_core
port 28 nsew signal input
rlabel metal5 s 6167 70054 19620 80934 6 vccd_pad
port 29 nsew signal bidirectional
rlabel metal5 s 624222 6811 636390 18976 6 vdda_pad
port 30 nsew signal bidirectional
rlabel metal5 s 6811 111610 18976 123778 6 vddio_pad
port 31 nsew signal bidirectional
rlabel metal5 s 6811 871210 18976 883378 6 vddio_pad2
port 32 nsew signal bidirectional
rlabel metal5 s 80222 6811 92390 18976 6 vssa_pad
port 33 nsew signal bidirectional
rlabel metal5 s 243266 6167 254146 19620 6 vssd_pad
port 34 nsew signal bidirectional
rlabel metal5 s 334810 1018624 346978 1030789 6 vssio_pad
port 35 nsew signal bidirectional
rlabel metal5 s 570422 6811 582590 18976 6 vssio_pad2
port 36 nsew signal bidirectional
rlabel metal5 s 698512 101240 711002 113760 6 mprj_io[0]
port 37 nsew signal bidirectional
rlabel metal2 s 675407 105803 675887 105859 6 mprj_io_analog_en[0]
port 38 nsew signal input
rlabel metal2 s 675407 107091 675887 107147 6 mprj_io_analog_pol[0]
port 39 nsew signal input
rlabel metal2 s 675407 110127 675887 110183 6 mprj_io_analog_sel[0]
port 40 nsew signal input
rlabel metal2 s 675407 106447 675887 106503 6 mprj_io_dm[0]
port 41 nsew signal input
rlabel metal2 s 675407 104607 675887 104663 6 mprj_io_dm[1]
port 42 nsew signal input
rlabel metal2 s 675407 110771 675887 110827 6 mprj_io_dm[2]
port 43 nsew signal input
rlabel metal2 s 675407 111415 675887 111471 6 mprj_io_holdover[0]
port 44 nsew signal input
rlabel metal2 s 675407 114451 675887 114507 6 mprj_io_ib_mode_sel[0]
port 45 nsew signal input
rlabel metal2 s 675407 107643 675887 107699 6 mprj_io_inp_dis[0]
port 46 nsew signal input
rlabel metal2 s 675407 115095 675887 115151 6 mprj_io_oeb[0]
port 47 nsew signal input
rlabel metal2 s 675407 111967 675887 112023 6 mprj_io_out[0]
port 48 nsew signal input
rlabel metal2 s 675407 102767 675887 102823 6 mprj_io_slow_sel[0]
port 49 nsew signal input
rlabel metal2 s 675407 113807 675887 113863 6 mprj_io_vtrip_sel[0]
port 50 nsew signal input
rlabel metal2 s 675407 100927 675887 100983 6 mprj_io_in[0]
port 51 nsew signal output
rlabel metal2 s 675407 686611 675887 686667 6 mprj_analog_io[3]
port 52 nsew signal bidirectional
rlabel metal5 s 698512 684440 711002 696960 6 mprj_io[10]
port 53 nsew signal bidirectional
rlabel metal2 s 675407 689003 675887 689059 6 mprj_io_analog_en[10]
port 54 nsew signal input
rlabel metal2 s 675407 690291 675887 690347 6 mprj_io_analog_pol[10]
port 55 nsew signal input
rlabel metal2 s 675407 693327 675887 693383 6 mprj_io_analog_sel[10]
port 56 nsew signal input
rlabel metal2 s 675407 689647 675887 689703 6 mprj_io_dm[30]
port 57 nsew signal input
rlabel metal2 s 675407 687807 675887 687863 6 mprj_io_dm[31]
port 58 nsew signal input
rlabel metal2 s 675407 693971 675887 694027 6 mprj_io_dm[32]
port 59 nsew signal input
rlabel metal2 s 675407 694615 675887 694671 6 mprj_io_holdover[10]
port 60 nsew signal input
rlabel metal2 s 675407 697651 675887 697707 6 mprj_io_ib_mode_sel[10]
port 61 nsew signal input
rlabel metal2 s 675407 690843 675887 690899 6 mprj_io_inp_dis[10]
port 62 nsew signal input
rlabel metal2 s 675407 698295 675887 698351 6 mprj_io_oeb[10]
port 63 nsew signal input
rlabel metal2 s 675407 695167 675887 695223 6 mprj_io_out[10]
port 64 nsew signal input
rlabel metal2 s 675407 685967 675887 686023 6 mprj_io_slow_sel[10]
port 65 nsew signal input
rlabel metal2 s 675407 697007 675887 697063 6 mprj_io_vtrip_sel[10]
port 66 nsew signal input
rlabel metal2 s 675407 684127 675887 684183 6 mprj_io_in[10]
port 67 nsew signal output
rlabel metal2 s 675407 731611 675887 731667 6 mprj_analog_io[4]
port 68 nsew signal bidirectional
rlabel metal5 s 698512 729440 711002 741960 6 mprj_io[11]
port 69 nsew signal bidirectional
rlabel metal2 s 675407 734003 675887 734059 6 mprj_io_analog_en[11]
port 70 nsew signal input
rlabel metal2 s 675407 735291 675887 735347 6 mprj_io_analog_pol[11]
port 71 nsew signal input
rlabel metal2 s 675407 738327 675887 738383 6 mprj_io_analog_sel[11]
port 72 nsew signal input
rlabel metal2 s 675407 734647 675887 734703 6 mprj_io_dm[33]
port 73 nsew signal input
rlabel metal2 s 675407 732807 675887 732863 6 mprj_io_dm[34]
port 74 nsew signal input
rlabel metal2 s 675407 738971 675887 739027 6 mprj_io_dm[35]
port 75 nsew signal input
rlabel metal2 s 675407 739615 675887 739671 6 mprj_io_holdover[11]
port 76 nsew signal input
rlabel metal2 s 675407 742651 675887 742707 6 mprj_io_ib_mode_sel[11]
port 77 nsew signal input
rlabel metal2 s 675407 735843 675887 735899 6 mprj_io_inp_dis[11]
port 78 nsew signal input
rlabel metal2 s 675407 743295 675887 743351 6 mprj_io_oeb[11]
port 79 nsew signal input
rlabel metal2 s 675407 740167 675887 740223 6 mprj_io_out[11]
port 80 nsew signal input
rlabel metal2 s 675407 730967 675887 731023 6 mprj_io_slow_sel[11]
port 81 nsew signal input
rlabel metal2 s 675407 742007 675887 742063 6 mprj_io_vtrip_sel[11]
port 82 nsew signal input
rlabel metal2 s 675407 729127 675887 729183 6 mprj_io_in[11]
port 83 nsew signal output
rlabel metal2 s 675407 776611 675887 776667 6 mprj_analog_io[5]
port 84 nsew signal bidirectional
rlabel metal5 s 698512 774440 711002 786960 6 mprj_io[12]
port 85 nsew signal bidirectional
rlabel metal2 s 675407 779003 675887 779059 6 mprj_io_analog_en[12]
port 86 nsew signal input
rlabel metal2 s 675407 780291 675887 780347 6 mprj_io_analog_pol[12]
port 87 nsew signal input
rlabel metal2 s 675407 783327 675887 783383 6 mprj_io_analog_sel[12]
port 88 nsew signal input
rlabel metal2 s 675407 779647 675887 779703 6 mprj_io_dm[36]
port 89 nsew signal input
rlabel metal2 s 675407 777807 675887 777863 6 mprj_io_dm[37]
port 90 nsew signal input
rlabel metal2 s 675407 783971 675887 784027 6 mprj_io_dm[38]
port 91 nsew signal input
rlabel metal2 s 675407 784615 675887 784671 6 mprj_io_holdover[12]
port 92 nsew signal input
rlabel metal2 s 675407 787651 675887 787707 6 mprj_io_ib_mode_sel[12]
port 93 nsew signal input
rlabel metal2 s 675407 780843 675887 780899 6 mprj_io_inp_dis[12]
port 94 nsew signal input
rlabel metal2 s 675407 788295 675887 788351 6 mprj_io_oeb[12]
port 95 nsew signal input
rlabel metal2 s 675407 785167 675887 785223 6 mprj_io_out[12]
port 96 nsew signal input
rlabel metal2 s 675407 775967 675887 776023 6 mprj_io_slow_sel[12]
port 97 nsew signal input
rlabel metal2 s 675407 787007 675887 787063 6 mprj_io_vtrip_sel[12]
port 98 nsew signal input
rlabel metal2 s 675407 774127 675887 774183 6 mprj_io_in[12]
port 99 nsew signal output
rlabel metal2 s 675407 865811 675887 865867 6 mprj_analog_io[6]
port 100 nsew signal bidirectional
rlabel metal5 s 698512 863640 711002 876160 6 mprj_io[13]
port 101 nsew signal bidirectional
rlabel metal2 s 675407 868203 675887 868259 6 mprj_io_analog_en[13]
port 102 nsew signal input
rlabel metal2 s 675407 869491 675887 869547 6 mprj_io_analog_pol[13]
port 103 nsew signal input
rlabel metal2 s 675407 872527 675887 872583 6 mprj_io_analog_sel[13]
port 104 nsew signal input
rlabel metal2 s 675407 868847 675887 868903 6 mprj_io_dm[39]
port 105 nsew signal input
rlabel metal2 s 675407 867007 675887 867063 6 mprj_io_dm[40]
port 106 nsew signal input
rlabel metal2 s 675407 873171 675887 873227 6 mprj_io_dm[41]
port 107 nsew signal input
rlabel metal2 s 675407 873815 675887 873871 6 mprj_io_holdover[13]
port 108 nsew signal input
rlabel metal2 s 675407 876851 675887 876907 6 mprj_io_ib_mode_sel[13]
port 109 nsew signal input
rlabel metal2 s 675407 870043 675887 870099 6 mprj_io_inp_dis[13]
port 110 nsew signal input
rlabel metal2 s 675407 877495 675887 877551 6 mprj_io_oeb[13]
port 111 nsew signal input
rlabel metal2 s 675407 874367 675887 874423 6 mprj_io_out[13]
port 112 nsew signal input
rlabel metal2 s 675407 865167 675887 865223 6 mprj_io_slow_sel[13]
port 113 nsew signal input
rlabel metal2 s 675407 876207 675887 876263 6 mprj_io_vtrip_sel[13]
port 114 nsew signal input
rlabel metal2 s 675407 863327 675887 863383 6 mprj_io_in[13]
port 115 nsew signal output
rlabel metal2 s 675407 955011 675887 955067 6 mprj_analog_io[7]
port 116 nsew signal bidirectional
rlabel metal5 s 698512 952840 711002 965360 6 mprj_io[14]
port 117 nsew signal bidirectional
rlabel metal2 s 675407 957403 675887 957459 6 mprj_io_analog_en[14]
port 118 nsew signal input
rlabel metal2 s 675407 958691 675887 958747 6 mprj_io_analog_pol[14]
port 119 nsew signal input
rlabel metal2 s 675407 961727 675887 961783 6 mprj_io_analog_sel[14]
port 120 nsew signal input
rlabel metal2 s 675407 958047 675887 958103 6 mprj_io_dm[42]
port 121 nsew signal input
rlabel metal2 s 675407 956207 675887 956263 6 mprj_io_dm[43]
port 122 nsew signal input
rlabel metal2 s 675407 962371 675887 962427 6 mprj_io_dm[44]
port 123 nsew signal input
rlabel metal2 s 675407 963015 675887 963071 6 mprj_io_holdover[14]
port 124 nsew signal input
rlabel metal2 s 675407 966051 675887 966107 6 mprj_io_ib_mode_sel[14]
port 125 nsew signal input
rlabel metal2 s 675407 959243 675887 959299 6 mprj_io_inp_dis[14]
port 126 nsew signal input
rlabel metal2 s 675407 966695 675887 966751 6 mprj_io_oeb[14]
port 127 nsew signal input
rlabel metal2 s 675407 963567 675887 963623 6 mprj_io_out[14]
port 128 nsew signal input
rlabel metal2 s 675407 954367 675887 954423 6 mprj_io_slow_sel[14]
port 129 nsew signal input
rlabel metal2 s 675407 965407 675887 965463 6 mprj_io_vtrip_sel[14]
port 130 nsew signal input
rlabel metal2 s 675407 952527 675887 952583 6 mprj_io_in[14]
port 131 nsew signal output
rlabel metal2 s 638533 995407 638589 995887 6 mprj_analog_io[8]
port 132 nsew signal bidirectional
rlabel metal5 s 628240 1018512 640760 1031002 6 mprj_io[15]
port 133 nsew signal bidirectional
rlabel metal2 s 636141 995407 636197 995887 6 mprj_io_analog_en[15]
port 134 nsew signal input
rlabel metal2 s 634853 995407 634909 995887 6 mprj_io_analog_pol[15]
port 135 nsew signal input
rlabel metal2 s 631817 995407 631873 995887 6 mprj_io_analog_sel[15]
port 136 nsew signal input
rlabel metal2 s 635497 995407 635553 995887 6 mprj_io_dm[45]
port 137 nsew signal input
rlabel metal2 s 637337 995407 637393 995887 6 mprj_io_dm[46]
port 138 nsew signal input
rlabel metal2 s 631173 995407 631229 995887 6 mprj_io_dm[47]
port 139 nsew signal input
rlabel metal2 s 630529 995407 630585 995887 6 mprj_io_holdover[15]
port 140 nsew signal input
rlabel metal2 s 627493 995407 627549 995887 6 mprj_io_ib_mode_sel[15]
port 141 nsew signal input
rlabel metal2 s 634301 995407 634357 995887 6 mprj_io_inp_dis[15]
port 142 nsew signal input
rlabel metal2 s 626849 995407 626905 995887 6 mprj_io_oeb[15]
port 143 nsew signal input
rlabel metal2 s 629977 995407 630033 995887 6 mprj_io_out[15]
port 144 nsew signal input
rlabel metal2 s 639177 995407 639233 995887 6 mprj_io_slow_sel[15]
port 145 nsew signal input
rlabel metal2 s 628137 995407 628193 995887 6 mprj_io_vtrip_sel[15]
port 146 nsew signal input
rlabel metal2 s 641017 995407 641073 995887 6 mprj_io_in[15]
port 147 nsew signal output
rlabel metal2 s 536733 995407 536789 995887 6 mprj_analog_io[9]
port 148 nsew signal bidirectional
rlabel metal5 s 526440 1018512 538960 1031002 6 mprj_io[16]
port 149 nsew signal bidirectional
rlabel metal2 s 534341 995407 534397 995887 6 mprj_io_analog_en[16]
port 150 nsew signal input
rlabel metal2 s 533053 995407 533109 995887 6 mprj_io_analog_pol[16]
port 151 nsew signal input
rlabel metal2 s 530017 995407 530073 995887 6 mprj_io_analog_sel[16]
port 152 nsew signal input
rlabel metal2 s 533697 995407 533753 995887 6 mprj_io_dm[48]
port 153 nsew signal input
rlabel metal2 s 535537 995407 535593 995887 6 mprj_io_dm[49]
port 154 nsew signal input
rlabel metal2 s 529373 995407 529429 995887 6 mprj_io_dm[50]
port 155 nsew signal input
rlabel metal2 s 528729 995407 528785 995887 6 mprj_io_holdover[16]
port 156 nsew signal input
rlabel metal2 s 525693 995407 525749 995887 6 mprj_io_ib_mode_sel[16]
port 157 nsew signal input
rlabel metal2 s 532501 995407 532557 995887 6 mprj_io_inp_dis[16]
port 158 nsew signal input
rlabel metal2 s 525049 995407 525105 995887 6 mprj_io_oeb[16]
port 159 nsew signal input
rlabel metal2 s 528177 995407 528233 995887 6 mprj_io_out[16]
port 160 nsew signal input
rlabel metal2 s 537377 995407 537433 995887 6 mprj_io_slow_sel[16]
port 161 nsew signal input
rlabel metal2 s 526337 995407 526393 995887 6 mprj_io_vtrip_sel[16]
port 162 nsew signal input
rlabel metal2 s 539217 995407 539273 995887 6 mprj_io_in[16]
port 163 nsew signal output
rlabel metal2 s 485333 995407 485389 995887 6 mprj_analog_io[10]
port 164 nsew signal bidirectional
rlabel metal5 s 475040 1018512 487560 1031002 6 mprj_io[17]
port 165 nsew signal bidirectional
rlabel metal2 s 482941 995407 482997 995887 6 mprj_io_analog_en[17]
port 166 nsew signal input
rlabel metal2 s 481653 995407 481709 995887 6 mprj_io_analog_pol[17]
port 167 nsew signal input
rlabel metal2 s 478617 995407 478673 995887 6 mprj_io_analog_sel[17]
port 168 nsew signal input
rlabel metal2 s 482297 995407 482353 995887 6 mprj_io_dm[51]
port 169 nsew signal input
rlabel metal2 s 484137 995407 484193 995887 6 mprj_io_dm[52]
port 170 nsew signal input
rlabel metal2 s 477973 995407 478029 995887 6 mprj_io_dm[53]
port 171 nsew signal input
rlabel metal2 s 477329 995407 477385 995887 6 mprj_io_holdover[17]
port 172 nsew signal input
rlabel metal2 s 474293 995407 474349 995887 6 mprj_io_ib_mode_sel[17]
port 173 nsew signal input
rlabel metal2 s 481101 995407 481157 995887 6 mprj_io_inp_dis[17]
port 174 nsew signal input
rlabel metal2 s 473649 995407 473705 995887 6 mprj_io_oeb[17]
port 175 nsew signal input
rlabel metal2 s 476777 995407 476833 995887 6 mprj_io_out[17]
port 176 nsew signal input
rlabel metal2 s 485977 995407 486033 995887 6 mprj_io_slow_sel[17]
port 177 nsew signal input
rlabel metal2 s 474937 995407 474993 995887 6 mprj_io_vtrip_sel[17]
port 178 nsew signal input
rlabel metal2 s 487817 995407 487873 995887 6 mprj_io_in[17]
port 179 nsew signal output
rlabel metal2 s 396333 995407 396389 995887 6 mprj_analog_io[11]
port 180 nsew signal bidirectional
rlabel metal5 s 386040 1018512 398560 1031002 6 mprj_io[18]
port 181 nsew signal bidirectional
rlabel metal2 s 393941 995407 393997 995887 6 mprj_io_analog_en[18]
port 182 nsew signal input
rlabel metal2 s 392653 995407 392709 995887 6 mprj_io_analog_pol[18]
port 183 nsew signal input
rlabel metal2 s 389617 995407 389673 995887 6 mprj_io_analog_sel[18]
port 184 nsew signal input
rlabel metal2 s 393297 995407 393353 995887 6 mprj_io_dm[54]
port 185 nsew signal input
rlabel metal2 s 395137 995407 395193 995887 6 mprj_io_dm[55]
port 186 nsew signal input
rlabel metal2 s 388973 995407 389029 995887 6 mprj_io_dm[56]
port 187 nsew signal input
rlabel metal2 s 388329 995407 388385 995887 6 mprj_io_holdover[18]
port 188 nsew signal input
rlabel metal2 s 385293 995407 385349 995887 6 mprj_io_ib_mode_sel[18]
port 189 nsew signal input
rlabel metal2 s 392101 995407 392157 995887 6 mprj_io_inp_dis[18]
port 190 nsew signal input
rlabel metal2 s 384649 995407 384705 995887 6 mprj_io_oeb[18]
port 191 nsew signal input
rlabel metal2 s 387777 995407 387833 995887 6 mprj_io_out[18]
port 192 nsew signal input
rlabel metal2 s 396977 995407 397033 995887 6 mprj_io_slow_sel[18]
port 193 nsew signal input
rlabel metal2 s 385937 995407 385993 995887 6 mprj_io_vtrip_sel[18]
port 194 nsew signal input
rlabel metal2 s 398817 995407 398873 995887 6 mprj_io_in[18]
port 195 nsew signal output
rlabel metal5 s 698512 146440 711002 158960 6 mprj_io[1]
port 196 nsew signal bidirectional
rlabel metal2 s 675407 151003 675887 151059 6 mprj_io_analog_en[1]
port 197 nsew signal input
rlabel metal2 s 675407 152291 675887 152347 6 mprj_io_analog_pol[1]
port 198 nsew signal input
rlabel metal2 s 675407 155327 675887 155383 6 mprj_io_analog_sel[1]
port 199 nsew signal input
rlabel metal2 s 675407 151647 675887 151703 6 mprj_io_dm[3]
port 200 nsew signal input
rlabel metal2 s 675407 149807 675887 149863 6 mprj_io_dm[4]
port 201 nsew signal input
rlabel metal2 s 675407 155971 675887 156027 6 mprj_io_dm[5]
port 202 nsew signal input
rlabel metal2 s 675407 156615 675887 156671 6 mprj_io_holdover[1]
port 203 nsew signal input
rlabel metal2 s 675407 159651 675887 159707 6 mprj_io_ib_mode_sel[1]
port 204 nsew signal input
rlabel metal2 s 675407 152843 675887 152899 6 mprj_io_inp_dis[1]
port 205 nsew signal input
rlabel metal2 s 675407 160295 675887 160351 6 mprj_io_oeb[1]
port 206 nsew signal input
rlabel metal2 s 675407 157167 675887 157223 6 mprj_io_out[1]
port 207 nsew signal input
rlabel metal2 s 675407 147967 675887 148023 6 mprj_io_slow_sel[1]
port 208 nsew signal input
rlabel metal2 s 675407 159007 675887 159063 6 mprj_io_vtrip_sel[1]
port 209 nsew signal input
rlabel metal2 s 675407 146127 675887 146183 6 mprj_io_in[1]
port 210 nsew signal output
rlabel metal5 s 698512 191440 711002 203960 6 mprj_io[2]
port 211 nsew signal bidirectional
rlabel metal2 s 675407 196003 675887 196059 6 mprj_io_analog_en[2]
port 212 nsew signal input
rlabel metal2 s 675407 197291 675887 197347 6 mprj_io_analog_pol[2]
port 213 nsew signal input
rlabel metal2 s 675407 200327 675887 200383 6 mprj_io_analog_sel[2]
port 214 nsew signal input
rlabel metal2 s 675407 196647 675887 196703 6 mprj_io_dm[6]
port 215 nsew signal input
rlabel metal2 s 675407 194807 675887 194863 6 mprj_io_dm[7]
port 216 nsew signal input
rlabel metal2 s 675407 200971 675887 201027 6 mprj_io_dm[8]
port 217 nsew signal input
rlabel metal2 s 675407 201615 675887 201671 6 mprj_io_holdover[2]
port 218 nsew signal input
rlabel metal2 s 675407 204651 675887 204707 6 mprj_io_ib_mode_sel[2]
port 219 nsew signal input
rlabel metal2 s 675407 197843 675887 197899 6 mprj_io_inp_dis[2]
port 220 nsew signal input
rlabel metal2 s 675407 205295 675887 205351 6 mprj_io_oeb[2]
port 221 nsew signal input
rlabel metal2 s 675407 202167 675887 202223 6 mprj_io_out[2]
port 222 nsew signal input
rlabel metal2 s 675407 192967 675887 193023 6 mprj_io_slow_sel[2]
port 223 nsew signal input
rlabel metal2 s 675407 204007 675887 204063 6 mprj_io_vtrip_sel[2]
port 224 nsew signal input
rlabel metal2 s 675407 191127 675887 191183 6 mprj_io_in[2]
port 225 nsew signal output
rlabel metal5 s 698512 236640 711002 249160 6 mprj_io[3]
port 226 nsew signal bidirectional
rlabel metal2 s 675407 241203 675887 241259 6 mprj_io_analog_en[3]
port 227 nsew signal input
rlabel metal2 s 675407 242491 675887 242547 6 mprj_io_analog_pol[3]
port 228 nsew signal input
rlabel metal2 s 675407 245527 675887 245583 6 mprj_io_analog_sel[3]
port 229 nsew signal input
rlabel metal2 s 675407 240007 675887 240063 6 mprj_io_dm[10]
port 230 nsew signal input
rlabel metal2 s 675407 246171 675887 246227 6 mprj_io_dm[11]
port 231 nsew signal input
rlabel metal2 s 675407 241847 675887 241903 6 mprj_io_dm[9]
port 232 nsew signal input
rlabel metal2 s 675407 246815 675887 246871 6 mprj_io_holdover[3]
port 233 nsew signal input
rlabel metal2 s 675407 249851 675887 249907 6 mprj_io_ib_mode_sel[3]
port 234 nsew signal input
rlabel metal2 s 675407 243043 675887 243099 6 mprj_io_inp_dis[3]
port 235 nsew signal input
rlabel metal2 s 675407 250495 675887 250551 6 mprj_io_oeb[3]
port 236 nsew signal input
rlabel metal2 s 675407 247367 675887 247423 6 mprj_io_out[3]
port 237 nsew signal input
rlabel metal2 s 675407 238167 675887 238223 6 mprj_io_slow_sel[3]
port 238 nsew signal input
rlabel metal2 s 675407 249207 675887 249263 6 mprj_io_vtrip_sel[3]
port 239 nsew signal input
rlabel metal2 s 675407 236327 675887 236383 6 mprj_io_in[3]
port 240 nsew signal output
rlabel metal5 s 698512 281640 711002 294160 6 mprj_io[4]
port 241 nsew signal bidirectional
rlabel metal2 s 675407 286203 675887 286259 6 mprj_io_analog_en[4]
port 242 nsew signal input
rlabel metal2 s 675407 287491 675887 287547 6 mprj_io_analog_pol[4]
port 243 nsew signal input
rlabel metal2 s 675407 290527 675887 290583 6 mprj_io_analog_sel[4]
port 244 nsew signal input
rlabel metal2 s 675407 286847 675887 286903 6 mprj_io_dm[12]
port 245 nsew signal input
rlabel metal2 s 675407 285007 675887 285063 6 mprj_io_dm[13]
port 246 nsew signal input
rlabel metal2 s 675407 291171 675887 291227 6 mprj_io_dm[14]
port 247 nsew signal input
rlabel metal2 s 675407 291815 675887 291871 6 mprj_io_holdover[4]
port 248 nsew signal input
rlabel metal2 s 675407 294851 675887 294907 6 mprj_io_ib_mode_sel[4]
port 249 nsew signal input
rlabel metal2 s 675407 288043 675887 288099 6 mprj_io_inp_dis[4]
port 250 nsew signal input
rlabel metal2 s 675407 295495 675887 295551 6 mprj_io_oeb[4]
port 251 nsew signal input
rlabel metal2 s 675407 292367 675887 292423 6 mprj_io_out[4]
port 252 nsew signal input
rlabel metal2 s 675407 283167 675887 283223 6 mprj_io_slow_sel[4]
port 253 nsew signal input
rlabel metal2 s 675407 294207 675887 294263 6 mprj_io_vtrip_sel[4]
port 254 nsew signal input
rlabel metal2 s 675407 281327 675887 281383 6 mprj_io_in[4]
port 255 nsew signal output
rlabel metal5 s 698512 326640 711002 339160 6 mprj_io[5]
port 256 nsew signal bidirectional
rlabel metal2 s 675407 331203 675887 331259 6 mprj_io_analog_en[5]
port 257 nsew signal input
rlabel metal2 s 675407 332491 675887 332547 6 mprj_io_analog_pol[5]
port 258 nsew signal input
rlabel metal2 s 675407 335527 675887 335583 6 mprj_io_analog_sel[5]
port 259 nsew signal input
rlabel metal2 s 675407 331847 675887 331903 6 mprj_io_dm[15]
port 260 nsew signal input
rlabel metal2 s 675407 330007 675887 330063 6 mprj_io_dm[16]
port 261 nsew signal input
rlabel metal2 s 675407 336171 675887 336227 6 mprj_io_dm[17]
port 262 nsew signal input
rlabel metal2 s 675407 336815 675887 336871 6 mprj_io_holdover[5]
port 263 nsew signal input
rlabel metal2 s 675407 339851 675887 339907 6 mprj_io_ib_mode_sel[5]
port 264 nsew signal input
rlabel metal2 s 675407 333043 675887 333099 6 mprj_io_inp_dis[5]
port 265 nsew signal input
rlabel metal2 s 675407 340495 675887 340551 6 mprj_io_oeb[5]
port 266 nsew signal input
rlabel metal2 s 675407 337367 675887 337423 6 mprj_io_out[5]
port 267 nsew signal input
rlabel metal2 s 675407 328167 675887 328223 6 mprj_io_slow_sel[5]
port 268 nsew signal input
rlabel metal2 s 675407 339207 675887 339263 6 mprj_io_vtrip_sel[5]
port 269 nsew signal input
rlabel metal2 s 675407 326327 675887 326383 6 mprj_io_in[5]
port 270 nsew signal output
rlabel metal5 s 698512 371840 711002 384360 6 mprj_io[6]
port 271 nsew signal bidirectional
rlabel metal2 s 675407 376403 675887 376459 6 mprj_io_analog_en[6]
port 272 nsew signal input
rlabel metal2 s 675407 377691 675887 377747 6 mprj_io_analog_pol[6]
port 273 nsew signal input
rlabel metal2 s 675407 380727 675887 380783 6 mprj_io_analog_sel[6]
port 274 nsew signal input
rlabel metal2 s 675407 377047 675887 377103 6 mprj_io_dm[18]
port 275 nsew signal input
rlabel metal2 s 675407 375207 675887 375263 6 mprj_io_dm[19]
port 276 nsew signal input
rlabel metal2 s 675407 381371 675887 381427 6 mprj_io_dm[20]
port 277 nsew signal input
rlabel metal2 s 675407 382015 675887 382071 6 mprj_io_holdover[6]
port 278 nsew signal input
rlabel metal2 s 675407 385051 675887 385107 6 mprj_io_ib_mode_sel[6]
port 279 nsew signal input
rlabel metal2 s 675407 378243 675887 378299 6 mprj_io_inp_dis[6]
port 280 nsew signal input
rlabel metal2 s 675407 385695 675887 385751 6 mprj_io_oeb[6]
port 281 nsew signal input
rlabel metal2 s 675407 382567 675887 382623 6 mprj_io_out[6]
port 282 nsew signal input
rlabel metal2 s 675407 373367 675887 373423 6 mprj_io_slow_sel[6]
port 283 nsew signal input
rlabel metal2 s 675407 384407 675887 384463 6 mprj_io_vtrip_sel[6]
port 284 nsew signal input
rlabel metal2 s 675407 371527 675887 371583 6 mprj_io_in[6]
port 285 nsew signal output
rlabel metal2 s 675407 551211 675887 551267 6 mprj_analog_io[0]
port 286 nsew signal bidirectional
rlabel metal5 s 698512 549040 711002 561560 6 mprj_io[7]
port 287 nsew signal bidirectional
rlabel metal2 s 675407 553603 675887 553659 6 mprj_io_analog_en[7]
port 288 nsew signal input
rlabel metal2 s 675407 554891 675887 554947 6 mprj_io_analog_pol[7]
port 289 nsew signal input
rlabel metal2 s 675407 557927 675887 557983 6 mprj_io_analog_sel[7]
port 290 nsew signal input
rlabel metal2 s 675407 554247 675887 554303 6 mprj_io_dm[21]
port 291 nsew signal input
rlabel metal2 s 675407 552407 675887 552463 6 mprj_io_dm[22]
port 292 nsew signal input
rlabel metal2 s 675407 558571 675887 558627 6 mprj_io_dm[23]
port 293 nsew signal input
rlabel metal2 s 675407 559215 675887 559271 6 mprj_io_holdover[7]
port 294 nsew signal input
rlabel metal2 s 675407 562251 675887 562307 6 mprj_io_ib_mode_sel[7]
port 295 nsew signal input
rlabel metal2 s 675407 555443 675887 555499 6 mprj_io_inp_dis[7]
port 296 nsew signal input
rlabel metal2 s 675407 562895 675887 562951 6 mprj_io_oeb[7]
port 297 nsew signal input
rlabel metal2 s 675407 559767 675887 559823 6 mprj_io_out[7]
port 298 nsew signal input
rlabel metal2 s 675407 550567 675887 550623 6 mprj_io_slow_sel[7]
port 299 nsew signal input
rlabel metal2 s 675407 561607 675887 561663 6 mprj_io_vtrip_sel[7]
port 300 nsew signal input
rlabel metal2 s 675407 548727 675887 548783 6 mprj_io_in[7]
port 301 nsew signal output
rlabel metal2 s 675407 596411 675887 596467 6 mprj_analog_io[1]
port 302 nsew signal bidirectional
rlabel metal5 s 698512 594240 711002 606760 6 mprj_io[8]
port 303 nsew signal bidirectional
rlabel metal2 s 675407 598803 675887 598859 6 mprj_io_analog_en[8]
port 304 nsew signal input
rlabel metal2 s 675407 600091 675887 600147 6 mprj_io_analog_pol[8]
port 305 nsew signal input
rlabel metal2 s 675407 603127 675887 603183 6 mprj_io_analog_sel[8]
port 306 nsew signal input
rlabel metal2 s 675407 599447 675887 599503 6 mprj_io_dm[24]
port 307 nsew signal input
rlabel metal2 s 675407 597607 675887 597663 6 mprj_io_dm[25]
port 308 nsew signal input
rlabel metal2 s 675407 603771 675887 603827 6 mprj_io_dm[26]
port 309 nsew signal input
rlabel metal2 s 675407 604415 675887 604471 6 mprj_io_holdover[8]
port 310 nsew signal input
rlabel metal2 s 675407 607451 675887 607507 6 mprj_io_ib_mode_sel[8]
port 311 nsew signal input
rlabel metal2 s 675407 600643 675887 600699 6 mprj_io_inp_dis[8]
port 312 nsew signal input
rlabel metal2 s 675407 608095 675887 608151 6 mprj_io_oeb[8]
port 313 nsew signal input
rlabel metal2 s 675407 604967 675887 605023 6 mprj_io_out[8]
port 314 nsew signal input
rlabel metal2 s 675407 595767 675887 595823 6 mprj_io_slow_sel[8]
port 315 nsew signal input
rlabel metal2 s 675407 606807 675887 606863 6 mprj_io_vtrip_sel[8]
port 316 nsew signal input
rlabel metal2 s 675407 593927 675887 593983 6 mprj_io_in[8]
port 317 nsew signal output
rlabel metal2 s 675407 641411 675887 641467 6 mprj_analog_io[2]
port 318 nsew signal bidirectional
rlabel metal5 s 698512 639240 711002 651760 6 mprj_io[9]
port 319 nsew signal bidirectional
rlabel metal2 s 675407 643803 675887 643859 6 mprj_io_analog_en[9]
port 320 nsew signal input
rlabel metal2 s 675407 645091 675887 645147 6 mprj_io_analog_pol[9]
port 321 nsew signal input
rlabel metal2 s 675407 648127 675887 648183 6 mprj_io_analog_sel[9]
port 322 nsew signal input
rlabel metal2 s 675407 644447 675887 644503 6 mprj_io_dm[27]
port 323 nsew signal input
rlabel metal2 s 675407 642607 675887 642663 6 mprj_io_dm[28]
port 324 nsew signal input
rlabel metal2 s 675407 648771 675887 648827 6 mprj_io_dm[29]
port 325 nsew signal input
rlabel metal2 s 675407 649415 675887 649471 6 mprj_io_holdover[9]
port 326 nsew signal input
rlabel metal2 s 675407 652451 675887 652507 6 mprj_io_ib_mode_sel[9]
port 327 nsew signal input
rlabel metal2 s 675407 645643 675887 645699 6 mprj_io_inp_dis[9]
port 328 nsew signal input
rlabel metal2 s 675407 653095 675887 653151 6 mprj_io_oeb[9]
port 329 nsew signal input
rlabel metal2 s 675407 649967 675887 650023 6 mprj_io_out[9]
port 330 nsew signal input
rlabel metal2 s 675407 640767 675887 640823 6 mprj_io_slow_sel[9]
port 331 nsew signal input
rlabel metal2 s 675407 651807 675887 651863 6 mprj_io_vtrip_sel[9]
port 332 nsew signal input
rlabel metal2 s 675407 638927 675887 638983 6 mprj_io_in[9]
port 333 nsew signal output
rlabel metal2 s 294533 995407 294589 995887 6 mprj_analog_io[12]
port 334 nsew signal bidirectional
rlabel metal5 s 284240 1018512 296760 1031002 6 mprj_io[19]
port 335 nsew signal bidirectional
rlabel metal2 s 292141 995407 292197 995887 6 mprj_io_analog_en[19]
port 336 nsew signal input
rlabel metal2 s 290853 995407 290909 995887 6 mprj_io_analog_pol[19]
port 337 nsew signal input
rlabel metal2 s 287817 995407 287873 995887 6 mprj_io_analog_sel[19]
port 338 nsew signal input
rlabel metal2 s 291497 995407 291553 995887 6 mprj_io_dm[57]
port 339 nsew signal input
rlabel metal2 s 293337 995407 293393 995887 6 mprj_io_dm[58]
port 340 nsew signal input
rlabel metal2 s 287173 995407 287229 995887 6 mprj_io_dm[59]
port 341 nsew signal input
rlabel metal2 s 286529 995407 286585 995887 6 mprj_io_holdover[19]
port 342 nsew signal input
rlabel metal2 s 283493 995407 283549 995887 6 mprj_io_ib_mode_sel[19]
port 343 nsew signal input
rlabel metal2 s 290301 995407 290357 995887 6 mprj_io_inp_dis[19]
port 344 nsew signal input
rlabel metal2 s 282849 995407 282905 995887 6 mprj_io_oeb[19]
port 345 nsew signal input
rlabel metal2 s 285977 995407 286033 995887 6 mprj_io_out[19]
port 346 nsew signal input
rlabel metal2 s 295177 995407 295233 995887 6 mprj_io_slow_sel[19]
port 347 nsew signal input
rlabel metal2 s 284137 995407 284193 995887 6 mprj_io_vtrip_sel[19]
port 348 nsew signal input
rlabel metal2 s 297017 995407 297073 995887 6 mprj_io_in[19]
port 349 nsew signal output
rlabel metal2 s 41713 624133 42193 624189 6 mprj_analog_io[22]
port 350 nsew signal bidirectional
rlabel metal5 s 6598 613840 19088 626360 6 mprj_io[29]
port 351 nsew signal bidirectional
rlabel metal2 s 41713 621741 42193 621797 6 mprj_io_analog_en[29]
port 352 nsew signal input
rlabel metal2 s 41713 620453 42193 620509 6 mprj_io_analog_pol[29]
port 353 nsew signal input
rlabel metal2 s 41713 617417 42193 617473 6 mprj_io_analog_sel[29]
port 354 nsew signal input
rlabel metal2 s 41713 621097 42193 621153 6 mprj_io_dm[87]
port 355 nsew signal input
rlabel metal2 s 41713 622937 42193 622993 6 mprj_io_dm[88]
port 356 nsew signal input
rlabel metal2 s 41713 616773 42193 616829 6 mprj_io_dm[89]
port 357 nsew signal input
rlabel metal2 s 41713 616129 42193 616185 6 mprj_io_holdover[29]
port 358 nsew signal input
rlabel metal2 s 41713 613093 42193 613149 6 mprj_io_ib_mode_sel[29]
port 359 nsew signal input
rlabel metal2 s 41713 619901 42193 619957 6 mprj_io_inp_dis[29]
port 360 nsew signal input
rlabel metal2 s 41713 612449 42193 612505 6 mprj_io_oeb[29]
port 361 nsew signal input
rlabel metal2 s 41713 615577 42193 615633 6 mprj_io_out[29]
port 362 nsew signal input
rlabel metal2 s 41713 624777 42193 624833 6 mprj_io_slow_sel[29]
port 363 nsew signal input
rlabel metal2 s 41713 613737 42193 613793 6 mprj_io_vtrip_sel[29]
port 364 nsew signal input
rlabel metal2 s 41713 626617 42193 626673 6 mprj_io_in[29]
port 365 nsew signal output
rlabel metal2 s 41713 580933 42193 580989 6 mprj_analog_io[23]
port 366 nsew signal bidirectional
rlabel metal5 s 6598 570640 19088 583160 6 mprj_io[30]
port 367 nsew signal bidirectional
rlabel metal2 s 41713 578541 42193 578597 6 mprj_io_analog_en[30]
port 368 nsew signal input
rlabel metal2 s 41713 577253 42193 577309 6 mprj_io_analog_pol[30]
port 369 nsew signal input
rlabel metal2 s 41713 574217 42193 574273 6 mprj_io_analog_sel[30]
port 370 nsew signal input
rlabel metal2 s 41713 577897 42193 577953 6 mprj_io_dm[90]
port 371 nsew signal input
rlabel metal2 s 41713 579737 42193 579793 6 mprj_io_dm[91]
port 372 nsew signal input
rlabel metal2 s 41713 573573 42193 573629 6 mprj_io_dm[92]
port 373 nsew signal input
rlabel metal2 s 41713 572929 42193 572985 6 mprj_io_holdover[30]
port 374 nsew signal input
rlabel metal2 s 41713 569893 42193 569949 6 mprj_io_ib_mode_sel[30]
port 375 nsew signal input
rlabel metal2 s 41713 576701 42193 576757 6 mprj_io_inp_dis[30]
port 376 nsew signal input
rlabel metal2 s 41713 569249 42193 569305 6 mprj_io_oeb[30]
port 377 nsew signal input
rlabel metal2 s 41713 572377 42193 572433 6 mprj_io_out[30]
port 378 nsew signal input
rlabel metal2 s 41713 581577 42193 581633 6 mprj_io_slow_sel[30]
port 379 nsew signal input
rlabel metal2 s 41713 570537 42193 570593 6 mprj_io_vtrip_sel[30]
port 380 nsew signal input
rlabel metal2 s 41713 583417 42193 583473 6 mprj_io_in[30]
port 381 nsew signal output
rlabel metal2 s 41713 537733 42193 537789 6 mprj_analog_io[24]
port 382 nsew signal bidirectional
rlabel metal5 s 6598 527440 19088 539960 6 mprj_io[31]
port 383 nsew signal bidirectional
rlabel metal2 s 41713 535341 42193 535397 6 mprj_io_analog_en[31]
port 384 nsew signal input
rlabel metal2 s 41713 534053 42193 534109 6 mprj_io_analog_pol[31]
port 385 nsew signal input
rlabel metal2 s 41713 531017 42193 531073 6 mprj_io_analog_sel[31]
port 386 nsew signal input
rlabel metal2 s 41713 534697 42193 534753 6 mprj_io_dm[93]
port 387 nsew signal input
rlabel metal2 s 41713 536537 42193 536593 6 mprj_io_dm[94]
port 388 nsew signal input
rlabel metal2 s 41713 530373 42193 530429 6 mprj_io_dm[95]
port 389 nsew signal input
rlabel metal2 s 41713 529729 42193 529785 6 mprj_io_holdover[31]
port 390 nsew signal input
rlabel metal2 s 41713 526693 42193 526749 6 mprj_io_ib_mode_sel[31]
port 391 nsew signal input
rlabel metal2 s 41713 533501 42193 533557 6 mprj_io_inp_dis[31]
port 392 nsew signal input
rlabel metal2 s 41713 526049 42193 526105 6 mprj_io_oeb[31]
port 393 nsew signal input
rlabel metal2 s 41713 529177 42193 529233 6 mprj_io_out[31]
port 394 nsew signal input
rlabel metal2 s 41713 538377 42193 538433 6 mprj_io_slow_sel[31]
port 395 nsew signal input
rlabel metal2 s 41713 527337 42193 527393 6 mprj_io_vtrip_sel[31]
port 396 nsew signal input
rlabel metal2 s 41713 540217 42193 540273 6 mprj_io_in[31]
port 397 nsew signal output
rlabel metal2 s 41713 410133 42193 410189 6 mprj_analog_io[25]
port 398 nsew signal bidirectional
rlabel metal5 s 6598 399840 19088 412360 6 mprj_io[32]
port 399 nsew signal bidirectional
rlabel metal2 s 41713 407741 42193 407797 6 mprj_io_analog_en[32]
port 400 nsew signal input
rlabel metal2 s 41713 406453 42193 406509 6 mprj_io_analog_pol[32]
port 401 nsew signal input
rlabel metal2 s 41713 403417 42193 403473 6 mprj_io_analog_sel[32]
port 402 nsew signal input
rlabel metal2 s 41713 407097 42193 407153 6 mprj_io_dm[96]
port 403 nsew signal input
rlabel metal2 s 41713 408937 42193 408993 6 mprj_io_dm[97]
port 404 nsew signal input
rlabel metal2 s 41713 402773 42193 402829 6 mprj_io_dm[98]
port 405 nsew signal input
rlabel metal2 s 41713 402129 42193 402185 6 mprj_io_holdover[32]
port 406 nsew signal input
rlabel metal2 s 41713 399093 42193 399149 6 mprj_io_ib_mode_sel[32]
port 407 nsew signal input
rlabel metal2 s 41713 405901 42193 405957 6 mprj_io_inp_dis[32]
port 408 nsew signal input
rlabel metal2 s 41713 398449 42193 398505 6 mprj_io_oeb[32]
port 409 nsew signal input
rlabel metal2 s 41713 401577 42193 401633 6 mprj_io_out[32]
port 410 nsew signal input
rlabel metal2 s 41713 410777 42193 410833 6 mprj_io_slow_sel[32]
port 411 nsew signal input
rlabel metal2 s 41713 399737 42193 399793 6 mprj_io_vtrip_sel[32]
port 412 nsew signal input
rlabel metal2 s 41713 412617 42193 412673 6 mprj_io_in[32]
port 413 nsew signal output
rlabel metal2 s 41713 366933 42193 366989 6 mprj_analog_io[26]
port 414 nsew signal bidirectional
rlabel metal5 s 6598 356640 19088 369160 6 mprj_io[33]
port 415 nsew signal bidirectional
rlabel metal2 s 41713 364541 42193 364597 6 mprj_io_analog_en[33]
port 416 nsew signal input
rlabel metal2 s 41713 363253 42193 363309 6 mprj_io_analog_pol[33]
port 417 nsew signal input
rlabel metal2 s 41713 360217 42193 360273 6 mprj_io_analog_sel[33]
port 418 nsew signal input
rlabel metal2 s 41713 365737 42193 365793 6 mprj_io_dm[100]
port 419 nsew signal input
rlabel metal2 s 41713 359573 42193 359629 6 mprj_io_dm[101]
port 420 nsew signal input
rlabel metal2 s 41713 363897 42193 363953 6 mprj_io_dm[99]
port 421 nsew signal input
rlabel metal2 s 41713 358929 42193 358985 6 mprj_io_holdover[33]
port 422 nsew signal input
rlabel metal2 s 41713 355893 42193 355949 6 mprj_io_ib_mode_sel[33]
port 423 nsew signal input
rlabel metal2 s 41713 362701 42193 362757 6 mprj_io_inp_dis[33]
port 424 nsew signal input
rlabel metal2 s 41713 355249 42193 355305 6 mprj_io_oeb[33]
port 425 nsew signal input
rlabel metal2 s 41713 358377 42193 358433 6 mprj_io_out[33]
port 426 nsew signal input
rlabel metal2 s 41713 367577 42193 367633 6 mprj_io_slow_sel[33]
port 427 nsew signal input
rlabel metal2 s 41713 356537 42193 356593 6 mprj_io_vtrip_sel[33]
port 428 nsew signal input
rlabel metal2 s 41713 369417 42193 369473 6 mprj_io_in[33]
port 429 nsew signal output
rlabel metal2 s 41713 323733 42193 323789 6 mprj_analog_io[27]
port 430 nsew signal bidirectional
rlabel metal5 s 6598 313440 19088 325960 6 mprj_io[34]
port 431 nsew signal bidirectional
rlabel metal2 s 41713 321341 42193 321397 6 mprj_io_analog_en[34]
port 432 nsew signal input
rlabel metal2 s 41713 320053 42193 320109 6 mprj_io_analog_pol[34]
port 433 nsew signal input
rlabel metal2 s 41713 317017 42193 317073 6 mprj_io_analog_sel[34]
port 434 nsew signal input
rlabel metal2 s 41713 320697 42193 320753 6 mprj_io_dm[102]
port 435 nsew signal input
rlabel metal2 s 41713 322537 42193 322593 6 mprj_io_dm[103]
port 436 nsew signal input
rlabel metal2 s 41713 316373 42193 316429 6 mprj_io_dm[104]
port 437 nsew signal input
rlabel metal2 s 41713 315729 42193 315785 6 mprj_io_holdover[34]
port 438 nsew signal input
rlabel metal2 s 41713 312693 42193 312749 6 mprj_io_ib_mode_sel[34]
port 439 nsew signal input
rlabel metal2 s 41713 319501 42193 319557 6 mprj_io_inp_dis[34]
port 440 nsew signal input
rlabel metal2 s 41713 312049 42193 312105 6 mprj_io_oeb[34]
port 441 nsew signal input
rlabel metal2 s 41713 315177 42193 315233 6 mprj_io_out[34]
port 442 nsew signal input
rlabel metal2 s 41713 324377 42193 324433 6 mprj_io_slow_sel[34]
port 443 nsew signal input
rlabel metal2 s 41713 313337 42193 313393 6 mprj_io_vtrip_sel[34]
port 444 nsew signal input
rlabel metal2 s 41713 326217 42193 326273 6 mprj_io_in[34]
port 445 nsew signal output
rlabel metal2 s 41713 280533 42193 280589 6 mprj_analog_io[28]
port 446 nsew signal bidirectional
rlabel metal5 s 6598 270240 19088 282760 6 mprj_io[35]
port 447 nsew signal bidirectional
rlabel metal2 s 41713 278141 42193 278197 6 mprj_io_analog_en[35]
port 448 nsew signal input
rlabel metal2 s 41713 276853 42193 276909 6 mprj_io_analog_pol[35]
port 449 nsew signal input
rlabel metal2 s 41713 273817 42193 273873 6 mprj_io_analog_sel[35]
port 450 nsew signal input
rlabel metal2 s 41713 277497 42193 277553 6 mprj_io_dm[105]
port 451 nsew signal input
rlabel metal2 s 41713 279337 42193 279393 6 mprj_io_dm[106]
port 452 nsew signal input
rlabel metal2 s 41713 273173 42193 273229 6 mprj_io_dm[107]
port 453 nsew signal input
rlabel metal2 s 41713 272529 42193 272585 6 mprj_io_holdover[35]
port 454 nsew signal input
rlabel metal2 s 41713 269493 42193 269549 6 mprj_io_ib_mode_sel[35]
port 455 nsew signal input
rlabel metal2 s 41713 276301 42193 276357 6 mprj_io_inp_dis[35]
port 456 nsew signal input
rlabel metal2 s 41713 268849 42193 268905 6 mprj_io_oeb[35]
port 457 nsew signal input
rlabel metal2 s 41713 271977 42193 272033 6 mprj_io_out[35]
port 458 nsew signal input
rlabel metal2 s 41713 281177 42193 281233 6 mprj_io_slow_sel[35]
port 459 nsew signal input
rlabel metal2 s 41713 270137 42193 270193 6 mprj_io_vtrip_sel[35]
port 460 nsew signal input
rlabel metal2 s 41713 283017 42193 283073 6 mprj_io_in[35]
port 461 nsew signal output
rlabel metal5 s 6598 227040 19088 239560 6 mprj_io[36]
port 462 nsew signal bidirectional
rlabel metal2 s 41713 234941 42193 234997 6 mprj_io_analog_en[36]
port 463 nsew signal input
rlabel metal2 s 41713 233653 42193 233709 6 mprj_io_analog_pol[36]
port 464 nsew signal input
rlabel metal2 s 41713 230617 42193 230673 6 mprj_io_analog_sel[36]
port 465 nsew signal input
rlabel metal2 s 41713 234297 42193 234353 6 mprj_io_dm[108]
port 466 nsew signal input
rlabel metal2 s 41713 236137 42193 236193 6 mprj_io_dm[109]
port 467 nsew signal input
rlabel metal2 s 41713 229973 42193 230029 6 mprj_io_dm[110]
port 468 nsew signal input
rlabel metal2 s 41713 229329 42193 229385 6 mprj_io_holdover[36]
port 469 nsew signal input
rlabel metal2 s 41713 226293 42193 226349 6 mprj_io_ib_mode_sel[36]
port 470 nsew signal input
rlabel metal2 s 41713 233101 42193 233157 6 mprj_io_inp_dis[36]
port 471 nsew signal input
rlabel metal2 s 41713 225649 42193 225705 6 mprj_io_oeb[36]
port 472 nsew signal input
rlabel metal2 s 41713 228777 42193 228833 6 mprj_io_out[36]
port 473 nsew signal input
rlabel metal2 s 41713 237977 42193 238033 6 mprj_io_slow_sel[36]
port 474 nsew signal input
rlabel metal2 s 41713 226937 42193 226993 6 mprj_io_vtrip_sel[36]
port 475 nsew signal input
rlabel metal2 s 41713 239817 42193 239873 6 mprj_io_in[36]
port 476 nsew signal output
rlabel metal5 s 6598 183840 19088 196360 6 mprj_io[37]
port 477 nsew signal bidirectional
rlabel metal2 s 41713 191741 42193 191797 6 mprj_io_analog_en[37]
port 478 nsew signal input
rlabel metal2 s 41713 190453 42193 190509 6 mprj_io_analog_pol[37]
port 479 nsew signal input
rlabel metal2 s 41713 187417 42193 187473 6 mprj_io_analog_sel[37]
port 480 nsew signal input
rlabel metal2 s 41713 191097 42193 191153 6 mprj_io_dm[111]
port 481 nsew signal input
rlabel metal2 s 41713 192937 42193 192993 6 mprj_io_dm[112]
port 482 nsew signal input
rlabel metal2 s 41713 186773 42193 186829 6 mprj_io_dm[113]
port 483 nsew signal input
rlabel metal2 s 41713 186129 42193 186185 6 mprj_io_holdover[37]
port 484 nsew signal input
rlabel metal2 s 41713 183093 42193 183149 6 mprj_io_ib_mode_sel[37]
port 485 nsew signal input
rlabel metal2 s 41713 189901 42193 189957 6 mprj_io_inp_dis[37]
port 486 nsew signal input
rlabel metal2 s 41713 182449 42193 182505 6 mprj_io_oeb[37]
port 487 nsew signal input
rlabel metal2 s 41713 185577 42193 185633 6 mprj_io_out[37]
port 488 nsew signal input
rlabel metal2 s 41713 194777 42193 194833 6 mprj_io_slow_sel[37]
port 489 nsew signal input
rlabel metal2 s 41713 183737 42193 183793 6 mprj_io_vtrip_sel[37]
port 490 nsew signal input
rlabel metal2 s 41713 196617 42193 196673 6 mprj_io_in[37]
port 491 nsew signal output
rlabel metal2 s 242933 995407 242989 995887 6 mprj_analog_io[13]
port 492 nsew signal bidirectional
rlabel metal5 s 232640 1018512 245160 1031002 6 mprj_io[20]
port 493 nsew signal bidirectional
rlabel metal2 s 240541 995407 240597 995887 6 mprj_io_analog_en[20]
port 494 nsew signal input
rlabel metal2 s 239253 995407 239309 995887 6 mprj_io_analog_pol[20]
port 495 nsew signal input
rlabel metal2 s 236217 995407 236273 995887 6 mprj_io_analog_sel[20]
port 496 nsew signal input
rlabel metal2 s 239897 995407 239953 995887 6 mprj_io_dm[60]
port 497 nsew signal input
rlabel metal2 s 241737 995407 241793 995887 6 mprj_io_dm[61]
port 498 nsew signal input
rlabel metal2 s 235573 995407 235629 995887 6 mprj_io_dm[62]
port 499 nsew signal input
rlabel metal2 s 234929 995407 234985 995887 6 mprj_io_holdover[20]
port 500 nsew signal input
rlabel metal2 s 231893 995407 231949 995887 6 mprj_io_ib_mode_sel[20]
port 501 nsew signal input
rlabel metal2 s 238701 995407 238757 995887 6 mprj_io_inp_dis[20]
port 502 nsew signal input
rlabel metal2 s 231249 995407 231305 995887 6 mprj_io_oeb[20]
port 503 nsew signal input
rlabel metal2 s 234377 995407 234433 995887 6 mprj_io_out[20]
port 504 nsew signal input
rlabel metal2 s 243577 995407 243633 995887 6 mprj_io_slow_sel[20]
port 505 nsew signal input
rlabel metal2 s 232537 995407 232593 995887 6 mprj_io_vtrip_sel[20]
port 506 nsew signal input
rlabel metal2 s 245417 995407 245473 995887 6 mprj_io_in[20]
port 507 nsew signal output
rlabel metal2 s 191533 995407 191589 995887 6 mprj_analog_io[14]
port 508 nsew signal bidirectional
rlabel metal5 s 181240 1018512 193760 1031002 6 mprj_io[21]
port 509 nsew signal bidirectional
rlabel metal2 s 189141 995407 189197 995887 6 mprj_io_analog_en[21]
port 510 nsew signal input
rlabel metal2 s 187853 995407 187909 995887 6 mprj_io_analog_pol[21]
port 511 nsew signal input
rlabel metal2 s 184817 995407 184873 995887 6 mprj_io_analog_sel[21]
port 512 nsew signal input
rlabel metal2 s 188497 995407 188553 995887 6 mprj_io_dm[63]
port 513 nsew signal input
rlabel metal2 s 190337 995407 190393 995887 6 mprj_io_dm[64]
port 514 nsew signal input
rlabel metal2 s 184173 995407 184229 995887 6 mprj_io_dm[65]
port 515 nsew signal input
rlabel metal2 s 183529 995407 183585 995887 6 mprj_io_holdover[21]
port 516 nsew signal input
rlabel metal2 s 180493 995407 180549 995887 6 mprj_io_ib_mode_sel[21]
port 517 nsew signal input
rlabel metal2 s 187301 995407 187357 995887 6 mprj_io_inp_dis[21]
port 518 nsew signal input
rlabel metal2 s 179849 995407 179905 995887 6 mprj_io_oeb[21]
port 519 nsew signal input
rlabel metal2 s 182977 995407 183033 995887 6 mprj_io_out[21]
port 520 nsew signal input
rlabel metal2 s 192177 995407 192233 995887 6 mprj_io_slow_sel[21]
port 521 nsew signal input
rlabel metal2 s 181137 995407 181193 995887 6 mprj_io_vtrip_sel[21]
port 522 nsew signal input
rlabel metal2 s 194017 995407 194073 995887 6 mprj_io_in[21]
port 523 nsew signal output
rlabel metal2 s 140133 995407 140189 995887 6 mprj_analog_io[15]
port 524 nsew signal bidirectional
rlabel metal5 s 129840 1018512 142360 1031002 6 mprj_io[22]
port 525 nsew signal bidirectional
rlabel metal2 s 137741 995407 137797 995887 6 mprj_io_analog_en[22]
port 526 nsew signal input
rlabel metal2 s 136453 995407 136509 995887 6 mprj_io_analog_pol[22]
port 527 nsew signal input
rlabel metal2 s 133417 995407 133473 995887 6 mprj_io_analog_sel[22]
port 528 nsew signal input
rlabel metal2 s 137097 995407 137153 995887 6 mprj_io_dm[66]
port 529 nsew signal input
rlabel metal2 s 138937 995407 138993 995887 6 mprj_io_dm[67]
port 530 nsew signal input
rlabel metal2 s 132773 995407 132829 995887 6 mprj_io_dm[68]
port 531 nsew signal input
rlabel metal2 s 132129 995407 132185 995887 6 mprj_io_holdover[22]
port 532 nsew signal input
rlabel metal2 s 129093 995407 129149 995887 6 mprj_io_ib_mode_sel[22]
port 533 nsew signal input
rlabel metal2 s 135901 995407 135957 995887 6 mprj_io_inp_dis[22]
port 534 nsew signal input
rlabel metal2 s 128449 995407 128505 995887 6 mprj_io_oeb[22]
port 535 nsew signal input
rlabel metal2 s 131577 995407 131633 995887 6 mprj_io_out[22]
port 536 nsew signal input
rlabel metal2 s 140777 995407 140833 995887 6 mprj_io_slow_sel[22]
port 537 nsew signal input
rlabel metal2 s 129737 995407 129793 995887 6 mprj_io_vtrip_sel[22]
port 538 nsew signal input
rlabel metal2 s 142617 995407 142673 995887 6 mprj_io_in[22]
port 539 nsew signal output
rlabel metal2 s 88733 995407 88789 995887 6 mprj_analog_io[16]
port 540 nsew signal bidirectional
rlabel metal5 s 78440 1018512 90960 1031002 6 mprj_io[23]
port 541 nsew signal bidirectional
rlabel metal2 s 86341 995407 86397 995887 6 mprj_io_analog_en[23]
port 542 nsew signal input
rlabel metal2 s 85053 995407 85109 995887 6 mprj_io_analog_pol[23]
port 543 nsew signal input
rlabel metal2 s 82017 995407 82073 995887 6 mprj_io_analog_sel[23]
port 544 nsew signal input
rlabel metal2 s 85697 995407 85753 995887 6 mprj_io_dm[69]
port 545 nsew signal input
rlabel metal2 s 87537 995407 87593 995887 6 mprj_io_dm[70]
port 546 nsew signal input
rlabel metal2 s 81373 995407 81429 995887 6 mprj_io_dm[71]
port 547 nsew signal input
rlabel metal2 s 80729 995407 80785 995887 6 mprj_io_holdover[23]
port 548 nsew signal input
rlabel metal2 s 77693 995407 77749 995887 6 mprj_io_ib_mode_sel[23]
port 549 nsew signal input
rlabel metal2 s 84501 995407 84557 995887 6 mprj_io_inp_dis[23]
port 550 nsew signal input
rlabel metal2 s 77049 995407 77105 995887 6 mprj_io_oeb[23]
port 551 nsew signal input
rlabel metal2 s 80177 995407 80233 995887 6 mprj_io_out[23]
port 552 nsew signal input
rlabel metal2 s 89377 995407 89433 995887 6 mprj_io_slow_sel[23]
port 553 nsew signal input
rlabel metal2 s 78337 995407 78393 995887 6 mprj_io_vtrip_sel[23]
port 554 nsew signal input
rlabel metal2 s 91217 995407 91273 995887 6 mprj_io_in[23]
port 555 nsew signal output
rlabel metal2 s 41713 966733 42193 966789 6 mprj_analog_io[17]
port 556 nsew signal bidirectional
rlabel metal5 s 6598 956440 19088 968960 6 mprj_io[24]
port 557 nsew signal bidirectional
rlabel metal2 s 41713 964341 42193 964397 6 mprj_io_analog_en[24]
port 558 nsew signal input
rlabel metal2 s 41713 963053 42193 963109 6 mprj_io_analog_pol[24]
port 559 nsew signal input
rlabel metal2 s 41713 960017 42193 960073 6 mprj_io_analog_sel[24]
port 560 nsew signal input
rlabel metal2 s 41713 963697 42193 963753 6 mprj_io_dm[72]
port 561 nsew signal input
rlabel metal2 s 41713 965537 42193 965593 6 mprj_io_dm[73]
port 562 nsew signal input
rlabel metal2 s 41713 959373 42193 959429 6 mprj_io_dm[74]
port 563 nsew signal input
rlabel metal2 s 41713 958729 42193 958785 6 mprj_io_holdover[24]
port 564 nsew signal input
rlabel metal2 s 41713 955693 42193 955749 6 mprj_io_ib_mode_sel[24]
port 565 nsew signal input
rlabel metal2 s 41713 962501 42193 962557 6 mprj_io_inp_dis[24]
port 566 nsew signal input
rlabel metal2 s 41713 955049 42193 955105 6 mprj_io_oeb[24]
port 567 nsew signal input
rlabel metal2 s 41713 958177 42193 958233 6 mprj_io_out[24]
port 568 nsew signal input
rlabel metal2 s 41713 967377 42193 967433 6 mprj_io_slow_sel[24]
port 569 nsew signal input
rlabel metal2 s 41713 956337 42193 956393 6 mprj_io_vtrip_sel[24]
port 570 nsew signal input
rlabel metal2 s 41713 969217 42193 969273 6 mprj_io_in[24]
port 571 nsew signal output
rlabel metal2 s 41713 796933 42193 796989 6 mprj_analog_io[18]
port 572 nsew signal bidirectional
rlabel metal5 s 6598 786640 19088 799160 6 mprj_io[25]
port 573 nsew signal bidirectional
rlabel metal2 s 41713 794541 42193 794597 6 mprj_io_analog_en[25]
port 574 nsew signal input
rlabel metal2 s 41713 793253 42193 793309 6 mprj_io_analog_pol[25]
port 575 nsew signal input
rlabel metal2 s 41713 790217 42193 790273 6 mprj_io_analog_sel[25]
port 576 nsew signal input
rlabel metal2 s 41713 793897 42193 793953 6 mprj_io_dm[75]
port 577 nsew signal input
rlabel metal2 s 41713 795737 42193 795793 6 mprj_io_dm[76]
port 578 nsew signal input
rlabel metal2 s 41713 789573 42193 789629 6 mprj_io_dm[77]
port 579 nsew signal input
rlabel metal2 s 41713 788929 42193 788985 6 mprj_io_holdover[25]
port 580 nsew signal input
rlabel metal2 s 41713 785893 42193 785949 6 mprj_io_ib_mode_sel[25]
port 581 nsew signal input
rlabel metal2 s 41713 792701 42193 792757 6 mprj_io_inp_dis[25]
port 582 nsew signal input
rlabel metal2 s 41713 785249 42193 785305 6 mprj_io_oeb[25]
port 583 nsew signal input
rlabel metal2 s 41713 788377 42193 788433 6 mprj_io_out[25]
port 584 nsew signal input
rlabel metal2 s 41713 797577 42193 797633 6 mprj_io_slow_sel[25]
port 585 nsew signal input
rlabel metal2 s 41713 786537 42193 786593 6 mprj_io_vtrip_sel[25]
port 586 nsew signal input
rlabel metal2 s 41713 799417 42193 799473 6 mprj_io_in[25]
port 587 nsew signal output
rlabel metal2 s 41713 753733 42193 753789 6 mprj_analog_io[19]
port 588 nsew signal bidirectional
rlabel metal5 s 6598 743440 19088 755960 6 mprj_io[26]
port 589 nsew signal bidirectional
rlabel metal2 s 41713 751341 42193 751397 6 mprj_io_analog_en[26]
port 590 nsew signal input
rlabel metal2 s 41713 750053 42193 750109 6 mprj_io_analog_pol[26]
port 591 nsew signal input
rlabel metal2 s 41713 747017 42193 747073 6 mprj_io_analog_sel[26]
port 592 nsew signal input
rlabel metal2 s 41713 750697 42193 750753 6 mprj_io_dm[78]
port 593 nsew signal input
rlabel metal2 s 41713 752537 42193 752593 6 mprj_io_dm[79]
port 594 nsew signal input
rlabel metal2 s 41713 746373 42193 746429 6 mprj_io_dm[80]
port 595 nsew signal input
rlabel metal2 s 41713 745729 42193 745785 6 mprj_io_holdover[26]
port 596 nsew signal input
rlabel metal2 s 41713 742693 42193 742749 6 mprj_io_ib_mode_sel[26]
port 597 nsew signal input
rlabel metal2 s 41713 749501 42193 749557 6 mprj_io_inp_dis[26]
port 598 nsew signal input
rlabel metal2 s 41713 742049 42193 742105 6 mprj_io_oeb[26]
port 599 nsew signal input
rlabel metal2 s 41713 745177 42193 745233 6 mprj_io_out[26]
port 600 nsew signal input
rlabel metal2 s 41713 754377 42193 754433 6 mprj_io_slow_sel[26]
port 601 nsew signal input
rlabel metal2 s 41713 743337 42193 743393 6 mprj_io_vtrip_sel[26]
port 602 nsew signal input
rlabel metal2 s 41713 756217 42193 756273 6 mprj_io_in[26]
port 603 nsew signal output
rlabel metal2 s 41713 710533 42193 710589 6 mprj_analog_io[20]
port 604 nsew signal bidirectional
rlabel metal5 s 6598 700240 19088 712760 6 mprj_io[27]
port 605 nsew signal bidirectional
rlabel metal2 s 41713 708141 42193 708197 6 mprj_io_analog_en[27]
port 606 nsew signal input
rlabel metal2 s 41713 706853 42193 706909 6 mprj_io_analog_pol[27]
port 607 nsew signal input
rlabel metal2 s 41713 703817 42193 703873 6 mprj_io_analog_sel[27]
port 608 nsew signal input
rlabel metal2 s 41713 707497 42193 707553 6 mprj_io_dm[81]
port 609 nsew signal input
rlabel metal2 s 41713 709337 42193 709393 6 mprj_io_dm[82]
port 610 nsew signal input
rlabel metal2 s 41713 703173 42193 703229 6 mprj_io_dm[83]
port 611 nsew signal input
rlabel metal2 s 41713 702529 42193 702585 6 mprj_io_holdover[27]
port 612 nsew signal input
rlabel metal2 s 41713 699493 42193 699549 6 mprj_io_ib_mode_sel[27]
port 613 nsew signal input
rlabel metal2 s 41713 706301 42193 706357 6 mprj_io_inp_dis[27]
port 614 nsew signal input
rlabel metal2 s 41713 698849 42193 698905 6 mprj_io_oeb[27]
port 615 nsew signal input
rlabel metal2 s 41713 701977 42193 702033 6 mprj_io_out[27]
port 616 nsew signal input
rlabel metal2 s 41713 711177 42193 711233 6 mprj_io_slow_sel[27]
port 617 nsew signal input
rlabel metal2 s 41713 700137 42193 700193 6 mprj_io_vtrip_sel[27]
port 618 nsew signal input
rlabel metal2 s 41713 713017 42193 713073 6 mprj_io_in[27]
port 619 nsew signal output
rlabel metal2 s 41713 667333 42193 667389 6 mprj_analog_io[21]
port 620 nsew signal bidirectional
rlabel metal5 s 6598 657040 19088 669560 6 mprj_io[28]
port 621 nsew signal bidirectional
rlabel metal2 s 41713 664941 42193 664997 6 mprj_io_analog_en[28]
port 622 nsew signal input
rlabel metal2 s 41713 663653 42193 663709 6 mprj_io_analog_pol[28]
port 623 nsew signal input
rlabel metal2 s 41713 660617 42193 660673 6 mprj_io_analog_sel[28]
port 624 nsew signal input
rlabel metal2 s 41713 664297 42193 664353 6 mprj_io_dm[84]
port 625 nsew signal input
rlabel metal2 s 41713 666137 42193 666193 6 mprj_io_dm[85]
port 626 nsew signal input
rlabel metal2 s 41713 659973 42193 660029 6 mprj_io_dm[86]
port 627 nsew signal input
rlabel metal2 s 41713 659329 42193 659385 6 mprj_io_holdover[28]
port 628 nsew signal input
rlabel metal2 s 41713 656293 42193 656349 6 mprj_io_ib_mode_sel[28]
port 629 nsew signal input
rlabel metal2 s 41713 663101 42193 663157 6 mprj_io_inp_dis[28]
port 630 nsew signal input
rlabel metal2 s 41713 655649 42193 655705 6 mprj_io_oeb[28]
port 631 nsew signal input
rlabel metal2 s 41713 658777 42193 658833 6 mprj_io_out[28]
port 632 nsew signal input
rlabel metal2 s 41713 667977 42193 668033 6 mprj_io_slow_sel[28]
port 633 nsew signal input
rlabel metal2 s 41713 656937 42193 656993 6 mprj_io_vtrip_sel[28]
port 634 nsew signal input
rlabel metal2 s 41713 669817 42193 669873 6 mprj_io_in[28]
port 635 nsew signal output
rlabel metal2 s 145091 39706 145143 40000 6 porb_h
port 636 nsew signal input
rlabel metal2 s 145103 40000 145131 40174 6 porb_h
port 636 nsew signal input
rlabel metal2 s 145103 40174 145144 40202 6 porb_h
port 636 nsew signal input
rlabel metal2 s 527455 41713 527511 42193 6 porb_h
port 636 nsew signal input
rlabel metal2 s 523131 41713 523187 42193 6 porb_h
port 636 nsew signal input
rlabel metal2 s 472655 41713 472711 41806 6 porb_h
port 636 nsew signal input
rlabel metal2 s 468331 41713 468387 41806 6 porb_h
port 636 nsew signal input
rlabel metal2 s 472636 41806 472711 42193 6 porb_h
port 636 nsew signal input
rlabel metal2 s 468312 41806 468387 42193 6 porb_h
port 636 nsew signal input
rlabel metal2 s 417855 41713 417911 41820 6 porb_h
port 636 nsew signal input
rlabel metal2 s 413531 41713 413587 41820 6 porb_h
port 636 nsew signal input
rlabel metal2 s 527468 42193 527496 44134 6 porb_h
port 636 nsew signal input
rlabel metal2 s 523144 42193 523172 44134 6 porb_h
port 636 nsew signal input
rlabel metal2 s 527456 44134 527508 44198 6 porb_h
port 636 nsew signal input
rlabel metal2 s 523132 44134 523184 44198 6 porb_h
port 636 nsew signal input
rlabel metal2 s 527468 44198 527496 46854 6 porb_h
port 636 nsew signal input
rlabel metal2 s 472636 42193 472664 44270 6 porb_h
port 636 nsew signal input
rlabel metal2 s 468312 42193 468340 44270 6 porb_h
port 636 nsew signal input
rlabel metal2 s 417855 41820 417924 42193 6 porb_h
port 636 nsew signal input
rlabel metal2 s 413531 41820 413600 42193 6 porb_h
port 636 nsew signal input
rlabel metal2 s 363055 41713 363111 42193 6 porb_h
port 636 nsew signal input
rlabel metal2 s 358731 41713 358787 42193 6 porb_h
port 636 nsew signal input
rlabel metal2 s 308255 41713 308311 41806 6 porb_h
port 636 nsew signal input
rlabel metal2 s 303931 41713 303987 41806 6 porb_h
port 636 nsew signal input
rlabel metal2 s 308232 41806 308311 42193 6 porb_h
port 636 nsew signal input
rlabel metal2 s 303908 41806 303987 42193 6 porb_h
port 636 nsew signal input
rlabel metal2 s 199655 41713 199711 42193 6 porb_h
port 636 nsew signal input
rlabel metal2 s 195331 41713 195387 42193 6 porb_h
port 636 nsew signal input
rlabel metal2 s 417896 42193 417924 44270 6 porb_h
port 636 nsew signal input
rlabel metal2 s 413572 42193 413600 44270 6 porb_h
port 636 nsew signal input
rlabel metal2 s 363064 42193 363092 44270 6 porb_h
port 636 nsew signal input
rlabel metal2 s 358740 42193 358768 44202 6 porb_h
port 636 nsew signal input
rlabel metal2 s 308232 42193 308260 44202 6 porb_h
port 636 nsew signal input
rlabel metal2 s 303908 42193 303936 44202 6 porb_h
port 636 nsew signal input
rlabel metal2 s 199672 42193 199700 44134 6 porb_h
port 636 nsew signal input
rlabel metal2 s 195348 42193 195376 44134 6 porb_h
port 636 nsew signal input
rlabel metal2 s 145116 40202 145144 44134 6 porb_h
port 636 nsew signal input
rlabel metal2 s 199660 44134 199712 44198 6 porb_h
port 636 nsew signal input
rlabel metal2 s 195336 44134 195388 44198 6 porb_h
port 636 nsew signal input
rlabel metal2 s 145104 44134 145156 44198 6 porb_h
port 636 nsew signal input
rlabel metal2 s 143632 44134 143684 44198 6 porb_h
port 636 nsew signal input
rlabel metal2 s 358728 44202 358780 44266 6 porb_h
port 636 nsew signal input
rlabel metal2 s 308220 44202 308272 44266 6 porb_h
port 636 nsew signal input
rlabel metal2 s 303896 44202 303948 44266 6 porb_h
port 636 nsew signal input
rlabel metal2 s 472624 44270 472676 44334 6 porb_h
port 636 nsew signal input
rlabel metal2 s 468300 44270 468352 44334 6 porb_h
port 636 nsew signal input
rlabel metal2 s 417884 44270 417936 44334 6 porb_h
port 636 nsew signal input
rlabel metal2 s 413560 44270 413612 44334 6 porb_h
port 636 nsew signal input
rlabel metal2 s 363052 44270 363104 44334 6 porb_h
port 636 nsew signal input
rlabel metal2 s 199672 44198 199700 44406 6 porb_h
port 636 nsew signal input
rlabel metal2 s 199660 44406 199712 44470 6 porb_h
port 636 nsew signal input
rlabel metal2 s 143644 44198 143672 45562 6 porb_h
port 636 nsew signal input
rlabel metal2 s 143632 45562 143684 45626 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42340 45562 42392 45626 6 porb_h
port 636 nsew signal input
rlabel metal2 s 527456 46854 527508 46918 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673644 46922 673696 46986 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673656 46986 673684 108394 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675392 108394 675444 108458 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673644 108394 673696 108458 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 108458 675432 108931 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 108931 675887 108945 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 108945 675887 108973 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 108973 675887 108987 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 113255 675887 113269 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 108973 675340 113269 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 113269 675887 113297 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 113297 675887 113311 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 113311 675432 113698 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675392 113698 675444 113762 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673644 113698 673696 113762 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673656 113762 673684 139318 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673656 139318 673776 139346 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 154059 675340 154090 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673748 139346 673776 154090 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 154131 675887 154142 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675300 154090 675352 154142 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675300 154142 675887 154154 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673736 154090 673788 154154 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 154154 675887 154170 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 154170 675887 154187 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 158455 675887 158494 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 154170 675340 158494 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 158494 675887 158511 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 158511 675432 158522 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 158522 675432 158578 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675392 158578 675444 158642 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673736 158578 673788 158642 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673748 158642 673776 199038 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42352 45626 42380 184303 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 184289 42193 184303 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 184303 42380 184331 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 184331 42288 188822 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 184331 42193 184345 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 188613 42193 188669 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41800 188669 41828 188822 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41800 188822 42380 188850 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42352 188850 42380 197270 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42340 197270 42392 197334 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42340 197474 42392 197538 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675392 199038 675444 199102 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673736 199038 673788 199102 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 199102 675432 199131 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 199131 675887 199158 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 199158 675887 199186 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 199186 675887 199187 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 203455 675887 203469 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 199186 675340 203458 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675300 203458 675352 203469 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675300 203469 675887 203497 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 203497 675887 203511 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675300 203497 675352 203522 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673736 203458 673788 203522 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 203522 675340 203580 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673748 203522 673776 243782 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42352 197538 42380 227582 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 227489 42193 227545 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41800 227545 41828 227582 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41800 227582 42380 227610 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 227610 42288 231827 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 231813 42193 231827 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 231827 42380 231855 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675392 243782 675444 243846 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673736 243782 673788 243846 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 243846 675432 244331 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 244331 675887 244345 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 244345 675887 244373 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 244373 675887 244387 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 248655 675887 248662 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 244373 675340 248662 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 248662 675887 248690 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 248690 675887 248711 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 248711 675432 249086 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675392 249086 675444 249150 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673736 249086 673788 249150 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673748 249150 673776 288798 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42352 231855 42380 264946 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 231855 42193 231869 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 264946 42380 264974 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 264974 42288 270830 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 270689 42193 270745 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41892 270745 41920 270830 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41892 270830 42288 270858 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 270858 42288 275182 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 275013 42193 275069 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41722 275069 41828 275074 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41800 275074 41828 275182 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41800 275182 42380 275210 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675392 288798 675444 288862 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673736 288798 673788 288862 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 288862 675432 289326 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 289326 675432 289331 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 289331 675887 289354 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 289354 675887 289387 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 293655 675887 293678 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 289354 675340 293678 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 293678 675887 293694 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675300 293694 675887 293706 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 293706 675887 293711 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675300 293706 675352 293758 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673828 293694 673880 293758 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 293758 675340 293789 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673840 293758 673868 334222 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42352 275210 42380 303586 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 303586 42380 303614 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 303614 42288 313806 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41800 313806 42288 313834 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 313834 42288 318227 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41800 313834 41828 313889 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 313889 42193 313945 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 318213 42193 318227 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 318227 42380 318255 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42352 318255 42380 332574 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 318255 42193 318269 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 332574 42380 332602 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675392 334222 675444 334286 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673828 334222 673880 334286 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 334286 675432 334331 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 334331 675887 334342 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 334342 675887 334370 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 334370 675887 334387 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 334370 675340 338150 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 338150 675432 338178 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 338178 675432 338655 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 338655 675887 338711 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 338711 675432 338778 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675392 338778 675444 338842 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673644 338778 673696 338842 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673656 338842 673684 379034 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 332602 42288 356646 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41984 356646 42288 356674 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 356674 42288 361406 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41984 356674 42012 357089 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 357089 42193 357145 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41722 361406 42288 361413 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 361413 42288 361434 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675392 379034 675444 379098 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673644 379034 673696 379098 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 379098 675432 379531 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 379531 675887 379545 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 379545 675887 379573 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 379573 675887 379587 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 383855 675887 383860 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 383860 675887 383911 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 383911 675432 383982 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 379573 675340 383982 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 383982 675432 384010 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 361434 42288 400302 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 361434 42193 361469 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 400289 42193 400302 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 400302 42288 400330 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 400330 42288 405198 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 400330 42193 400345 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 404613 42193 404669 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41722 404669 41828 404682 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41800 404682 41828 405198 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41800 405198 42380 405226 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42352 405226 42380 419506 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 419506 42380 419534 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 419534 42288 527870 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41708 527870 42288 527898 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 527898 42288 532086 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41708 527898 42193 527917 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 527917 42193 527945 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41892 532086 42380 532114 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 556731 675887 556759 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 556759 675887 556787 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 556787 675432 557262 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675392 557262 675444 557326 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675208 557262 675260 557326 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 561055 675887 561068 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 561068 675887 561111 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 561111 675432 561206 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675220 557326 675248 561206 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675392 561206 675444 561270 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675208 561206 675260 561270 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673736 561206 673788 561270 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673748 561270 673776 601802 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42352 532114 42380 571254 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41892 532114 41920 532213 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 532213 42193 532269 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 571089 42193 571145 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41722 571145 41828 571146 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41800 571146 41828 571254 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41800 571254 42380 571282 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 571282 42288 575427 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 575413 42193 575427 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 575427 42380 575455 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675392 601802 675444 601866 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675208 601802 675260 601866 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673736 601802 673788 601866 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 601866 675432 601931 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 601931 675887 601959 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 601959 675887 601987 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675220 601866 675248 605746 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675392 605746 675444 605810 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675208 605746 675260 605810 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673736 605746 673788 605810 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 605810 675432 606255 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 606255 675887 606283 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 606283 675887 606311 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673748 605810 673776 646410 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42352 575455 42380 612706 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 575455 42193 575469 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 612706 42380 612734 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 612734 42288 614303 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 614289 42193 614303 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 614303 42288 614331 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 614331 42288 618718 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 614331 42193 614345 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 618613 42193 618669 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41800 618669 41828 618718 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41800 618718 42380 618746 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675392 646410 675444 646474 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673736 646410 673788 646474 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 646474 675432 646931 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 646931 675887 646959 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 646959 675887 646987 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673748 646474 673776 651102 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675392 651102 675444 651166 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673736 651102 673788 651166 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 651166 675432 651255 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 651255 675887 651283 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 651283 675887 651311 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673748 651166 673776 692038 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42352 618746 42380 651346 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 651346 42380 651374 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 651374 42288 657614 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41722 657478 41920 657489 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 657489 42193 657545 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41892 657545 41920 657614 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41892 657614 42288 657642 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 657642 42288 661966 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 661813 42193 661869 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41800 661869 41828 661966 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41800 661966 42380 661994 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42352 661994 42380 689986 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 689986 42380 690014 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675392 692038 675444 692102 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675208 692038 675260 692102 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673736 692038 673788 692102 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 692102 675432 692131 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 692131 675887 692172 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 692172 675887 692187 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675220 692102 675248 695914 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675392 695914 675444 695978 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675208 695914 675260 695978 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673736 695914 673788 695978 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 695978 675432 696455 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 696455 675887 696483 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 696483 675887 696511 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673748 695978 673776 736986 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 690014 42288 700590 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41892 700590 42288 700618 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 700618 42288 704942 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41892 700618 41920 700689 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 700689 42193 700745 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41722 700745 41920 700754 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41892 704942 42380 704970 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42352 704970 42380 718830 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41892 704970 41920 705013 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 705013 42193 705069 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42340 718830 42392 718894 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42340 719034 42392 719098 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675392 736986 675444 737050 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675208 736986 675260 737050 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673736 736986 673788 737050 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 737050 675432 737131 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 737131 675887 737159 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 737159 675887 737187 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675220 737050 675248 740930 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675392 740930 675444 740994 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675208 740930 675260 740994 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673736 740930 673788 740994 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 740994 675432 741455 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 741455 675887 741483 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 741483 675887 741511 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673748 740994 673776 781594 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42352 719098 42380 743446 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42340 743446 42392 743510 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41788 743446 41840 743510 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42352 743510 42380 747866 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41800 743510 41828 743889 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 743889 42193 743945 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42340 747866 42392 747930 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41972 747866 42024 747930 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42352 747930 42380 749278 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41984 747930 42012 748213 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 748213 42193 748269 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42352 749278 42472 749306 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42444 749306 42472 756366 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42432 756366 42484 756430 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42432 756570 42484 756634 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675392 781594 675444 781658 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675208 781594 675260 781658 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673736 781594 673788 781658 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 781658 675432 782131 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 782131 675887 782159 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 782159 675887 782187 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675220 781658 675248 785946 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675392 785946 675444 786010 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675208 785946 675260 786010 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673828 785946 673880 786010 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 786010 675432 786455 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 786455 675887 786483 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 786483 675887 786511 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673840 786010 673868 871286 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42444 756634 42472 786966 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42432 786966 42484 787030 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41788 786966 41840 787030 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42444 787030 42472 787630 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41800 787030 41828 787086 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41722 787086 41828 787089 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 787089 42193 787145 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42444 787630 42564 787658 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42536 787658 42564 791930 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 791413 42193 791469 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41800 791469 41828 791930 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42524 791930 42576 791994 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41788 791930 41840 791994 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 871331 675887 871345 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675300 871286 675352 871345 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675300 871345 675887 871350 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673828 871286 673880 871350 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 871350 675887 871373 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 871373 675887 871387 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 875655 675887 875669 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 871373 675340 875669 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 875669 675887 875697 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 875697 675887 875711 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 875711 675432 875774 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675392 875774 675444 875838 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673644 875774 673696 875838 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673656 875838 673684 960026 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42536 791994 42564 941146 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 941146 42564 941174 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42260 941174 42288 956814 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41800 956814 42564 956842 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675392 960026 675444 960090 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673644 960026 673696 960090 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 960090 675432 960531 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 960531 675887 960545 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 960545 675887 960573 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 960573 675887 960587 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675407 964855 675887 964869 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 960573 675340 964869 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42536 956842 42564 961114 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41800 956842 41828 956889 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 956889 42193 956945 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42524 961114 42576 961178 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41788 961114 41840 961178 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675312 964869 675887 964897 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 964897 675887 964911 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675404 964911 675432 965262 6 porb_h
port 636 nsew signal input
rlabel metal2 s 675392 965262 675444 965326 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673828 965262 673880 965326 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673840 965326 673868 990082 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42536 961178 42564 969598 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41800 961178 41828 961213 6 porb_h
port 636 nsew signal input
rlabel metal2 s 41713 961213 42193 961269 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42352 969598 42564 969626 6 porb_h
port 636 nsew signal input
rlabel metal2 s 673828 990082 673880 990146 6 porb_h
port 636 nsew signal input
rlabel metal2 s 634728 990082 634780 990146 6 porb_h
port 636 nsew signal input
rlabel metal2 s 634740 990146 634768 990558 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42352 969626 42380 990218 6 porb_h
port 636 nsew signal input
rlabel metal2 s 78864 990218 78916 990282 6 porb_h
port 636 nsew signal input
rlabel metal2 s 42340 990218 42392 990282 6 porb_h
port 636 nsew signal input
rlabel metal2 s 274468 990542 274680 990558 6 porb_h
port 636 nsew signal input
rlabel metal2 s 78876 990282 78904 990558 6 porb_h
port 636 nsew signal input
rlabel metal2 s 634728 990558 634780 990622 6 porb_h
port 636 nsew signal input
rlabel metal2 s 632980 990558 633032 990622 6 porb_h
port 636 nsew signal input
rlabel metal2 s 628656 990558 628708 990622 6 porb_h
port 636 nsew signal input
rlabel metal2 s 531228 990558 531280 990622 6 porb_h
port 636 nsew signal input
rlabel metal2 s 526904 990558 526956 990622 6 porb_h
port 636 nsew signal input
rlabel metal2 s 479800 990558 479852 990622 6 porb_h
port 636 nsew signal input
rlabel metal2 s 475476 990558 475528 990622 6 porb_h
port 636 nsew signal input
rlabel metal2 s 390836 990558 390888 990622 6 porb_h
port 636 nsew signal input
rlabel metal2 s 386512 990558 386564 990622 6 porb_h
port 636 nsew signal input
rlabel metal2 s 274456 990558 274680 990570 6 porb_h
port 636 nsew signal input
rlabel metal2 s 632992 990622 633020 995407 6 porb_h
port 636 nsew signal input
rlabel metal2 s 628668 990622 628696 995407 6 porb_h
port 636 nsew signal input
rlabel metal2 s 531240 990622 531268 995407 6 porb_h
port 636 nsew signal input
rlabel metal2 s 526916 990622 526944 995407 6 porb_h
port 636 nsew signal input
rlabel metal2 s 479812 990622 479840 995407 6 porb_h
port 636 nsew signal input
rlabel metal2 s 475488 990622 475516 995407 6 porb_h
port 636 nsew signal input
rlabel metal2 s 632992 995407 633069 995466 6 porb_h
port 636 nsew signal input
rlabel metal2 s 628668 995407 628745 995466 6 porb_h
port 636 nsew signal input
rlabel metal2 s 633013 995466 633069 995887 6 porb_h
port 636 nsew signal input
rlabel metal2 s 628689 995466 628745 995887 6 porb_h
port 636 nsew signal input
rlabel metal2 s 531213 995407 531269 995887 6 porb_h
port 636 nsew signal input
rlabel metal2 s 526889 995407 526945 995887 6 porb_h
port 636 nsew signal input
rlabel metal2 s 479812 995407 479869 995452 6 porb_h
port 636 nsew signal input
rlabel metal2 s 475488 995407 475545 995452 6 porb_h
port 636 nsew signal input
rlabel metal2 s 390848 990622 390876 995407 6 porb_h
port 636 nsew signal input
rlabel metal2 s 386524 990622 386552 995407 6 porb_h
port 636 nsew signal input
rlabel metal2 s 288992 990626 289044 990690 6 porb_h
port 636 nsew signal input
rlabel metal2 s 284668 990626 284720 990690 6 porb_h
port 636 nsew signal input
rlabel metal2 s 274732 990626 274784 990644 6 porb_h
port 636 nsew signal input
rlabel metal2 s 274652 990570 274680 990644 6 porb_h
port 636 nsew signal input
rlabel metal2 s 274456 990570 274508 990622 6 porb_h
port 636 nsew signal input
rlabel metal2 s 237380 990558 237432 990622 6 porb_h
port 636 nsew signal input
rlabel metal2 s 233056 990558 233108 990622 6 porb_h
port 636 nsew signal input
rlabel metal2 s 186044 990558 186096 990622 6 porb_h
port 636 nsew signal input
rlabel metal2 s 181720 990558 181772 990622 6 porb_h
port 636 nsew signal input
rlabel metal2 s 134616 990558 134668 990622 6 porb_h
port 636 nsew signal input
rlabel metal2 s 130292 990558 130344 990622 6 porb_h
port 636 nsew signal input
rlabel metal2 s 83188 990558 83240 990622 6 porb_h
port 636 nsew signal input
rlabel metal2 s 78864 990558 78916 990622 6 porb_h
port 636 nsew signal input
rlabel metal2 s 274652 990644 274784 990672 6 porb_h
port 636 nsew signal input
rlabel metal2 s 274732 990672 274784 990690 6 porb_h
port 636 nsew signal input
rlabel metal2 s 289004 990690 289032 995407 6 porb_h
port 636 nsew signal input
rlabel metal2 s 284680 990690 284708 995407 6 porb_h
port 636 nsew signal input
rlabel metal2 s 237392 990622 237420 995407 6 porb_h
port 636 nsew signal input
rlabel metal2 s 233068 990622 233096 995407 6 porb_h
port 636 nsew signal input
rlabel metal2 s 390813 995407 390876 995452 6 porb_h
port 636 nsew signal input
rlabel metal2 s 386489 995407 386552 995452 6 porb_h
port 636 nsew signal input
rlabel metal2 s 479813 995452 479869 995887 6 porb_h
port 636 nsew signal input
rlabel metal2 s 475489 995452 475545 995887 6 porb_h
port 636 nsew signal input
rlabel metal2 s 390813 995452 390869 995887 6 porb_h
port 636 nsew signal input
rlabel metal2 s 386489 995452 386545 995887 6 porb_h
port 636 nsew signal input
rlabel metal2 s 289004 995407 289069 995452 6 porb_h
port 636 nsew signal input
rlabel metal2 s 284680 995407 284745 995452 6 porb_h
port 636 nsew signal input
rlabel metal2 s 289013 995452 289069 995887 6 porb_h
port 636 nsew signal input
rlabel metal2 s 284689 995452 284745 995887 6 porb_h
port 636 nsew signal input
rlabel metal2 s 237392 995407 237469 995466 6 porb_h
port 636 nsew signal input
rlabel metal2 s 233068 995407 233145 995466 6 porb_h
port 636 nsew signal input
rlabel metal2 s 186056 990622 186084 995407 6 porb_h
port 636 nsew signal input
rlabel metal2 s 181732 990622 181760 995407 6 porb_h
port 636 nsew signal input
rlabel metal2 s 134628 990622 134656 995407 6 porb_h
port 636 nsew signal input
rlabel metal2 s 130304 990622 130332 995407 6 porb_h
port 636 nsew signal input
rlabel metal2 s 83200 990622 83228 995407 6 porb_h
port 636 nsew signal input
rlabel metal2 s 78876 990622 78904 995407 6 porb_h
port 636 nsew signal input
rlabel metal2 s 186013 995407 186084 995466 6 porb_h
port 636 nsew signal input
rlabel metal2 s 181689 995407 181760 995466 6 porb_h
port 636 nsew signal input
rlabel metal2 s 237413 995466 237469 995887 6 porb_h
port 636 nsew signal input
rlabel metal2 s 233089 995466 233145 995887 6 porb_h
port 636 nsew signal input
rlabel metal2 s 186013 995466 186069 995887 6 porb_h
port 636 nsew signal input
rlabel metal2 s 181689 995466 181745 995887 6 porb_h
port 636 nsew signal input
rlabel metal2 s 134613 995407 134669 995887 6 porb_h
port 636 nsew signal input
rlabel metal2 s 130289 995407 130345 995887 6 porb_h
port 636 nsew signal input
rlabel metal2 s 83200 995407 83269 995452 6 porb_h
port 636 nsew signal input
rlabel metal2 s 78876 995407 78945 995452 6 porb_h
port 636 nsew signal input
rlabel metal2 s 83213 995452 83269 995887 6 porb_h
port 636 nsew signal input
rlabel metal2 s 78889 995452 78945 995887 6 porb_h
port 636 nsew signal input
rlabel via1 s 527456 44140 527508 44192 6 porb_h
port 636 nsew signal input
rlabel via1 s 523132 44140 523184 44192 6 porb_h
port 636 nsew signal input
rlabel via1 s 199660 44140 199712 44192 6 porb_h
port 636 nsew signal input
rlabel via1 s 195336 44140 195388 44192 6 porb_h
port 636 nsew signal input
rlabel via1 s 145104 44140 145156 44192 6 porb_h
port 636 nsew signal input
rlabel via1 s 143632 44140 143684 44192 6 porb_h
port 636 nsew signal input
rlabel via1 s 472624 44276 472676 44328 6 porb_h
port 636 nsew signal input
rlabel via1 s 468300 44276 468352 44328 6 porb_h
port 636 nsew signal input
rlabel via1 s 417884 44276 417936 44328 6 porb_h
port 636 nsew signal input
rlabel via1 s 413560 44276 413612 44328 6 porb_h
port 636 nsew signal input
rlabel via1 s 363052 44276 363104 44328 6 porb_h
port 636 nsew signal input
rlabel via1 s 358728 44208 358780 44260 6 porb_h
port 636 nsew signal input
rlabel via1 s 308220 44208 308272 44260 6 porb_h
port 636 nsew signal input
rlabel via1 s 303896 44208 303948 44260 6 porb_h
port 636 nsew signal input
rlabel via1 s 199660 44412 199712 44464 6 porb_h
port 636 nsew signal input
rlabel via1 s 143632 45568 143684 45620 6 porb_h
port 636 nsew signal input
rlabel via1 s 42340 45568 42392 45620 6 porb_h
port 636 nsew signal input
rlabel via1 s 527456 46860 527508 46912 6 porb_h
port 636 nsew signal input
rlabel via1 s 673644 46928 673696 46980 6 porb_h
port 636 nsew signal input
rlabel via1 s 675392 108400 675444 108452 6 porb_h
port 636 nsew signal input
rlabel via1 s 673644 108400 673696 108452 6 porb_h
port 636 nsew signal input
rlabel via1 s 675392 113704 675444 113756 6 porb_h
port 636 nsew signal input
rlabel via1 s 673644 113704 673696 113756 6 porb_h
port 636 nsew signal input
rlabel via1 s 675300 154096 675352 154148 6 porb_h
port 636 nsew signal input
rlabel via1 s 673736 154096 673788 154148 6 porb_h
port 636 nsew signal input
rlabel via1 s 675392 158584 675444 158636 6 porb_h
port 636 nsew signal input
rlabel via1 s 673736 158584 673788 158636 6 porb_h
port 636 nsew signal input
rlabel via1 s 42340 197276 42392 197328 6 porb_h
port 636 nsew signal input
rlabel via1 s 42340 197480 42392 197532 6 porb_h
port 636 nsew signal input
rlabel via1 s 675392 199044 675444 199096 6 porb_h
port 636 nsew signal input
rlabel via1 s 673736 199044 673788 199096 6 porb_h
port 636 nsew signal input
rlabel via1 s 675300 203464 675352 203516 6 porb_h
port 636 nsew signal input
rlabel via1 s 673736 203464 673788 203516 6 porb_h
port 636 nsew signal input
rlabel via1 s 675392 243788 675444 243840 6 porb_h
port 636 nsew signal input
rlabel via1 s 673736 243788 673788 243840 6 porb_h
port 636 nsew signal input
rlabel via1 s 675392 249092 675444 249144 6 porb_h
port 636 nsew signal input
rlabel via1 s 673736 249092 673788 249144 6 porb_h
port 636 nsew signal input
rlabel via1 s 675392 288804 675444 288856 6 porb_h
port 636 nsew signal input
rlabel via1 s 673736 288804 673788 288856 6 porb_h
port 636 nsew signal input
rlabel via1 s 675300 293700 675352 293752 6 porb_h
port 636 nsew signal input
rlabel via1 s 673828 293700 673880 293752 6 porb_h
port 636 nsew signal input
rlabel via1 s 675392 334228 675444 334280 6 porb_h
port 636 nsew signal input
rlabel via1 s 673828 334228 673880 334280 6 porb_h
port 636 nsew signal input
rlabel via1 s 675392 338784 675444 338836 6 porb_h
port 636 nsew signal input
rlabel via1 s 673644 338784 673696 338836 6 porb_h
port 636 nsew signal input
rlabel via1 s 675392 379040 675444 379092 6 porb_h
port 636 nsew signal input
rlabel via1 s 673644 379040 673696 379092 6 porb_h
port 636 nsew signal input
rlabel via1 s 675392 557268 675444 557320 6 porb_h
port 636 nsew signal input
rlabel via1 s 675208 557268 675260 557320 6 porb_h
port 636 nsew signal input
rlabel via1 s 675392 561212 675444 561264 6 porb_h
port 636 nsew signal input
rlabel via1 s 675208 561212 675260 561264 6 porb_h
port 636 nsew signal input
rlabel via1 s 673736 561212 673788 561264 6 porb_h
port 636 nsew signal input
rlabel via1 s 675392 601808 675444 601860 6 porb_h
port 636 nsew signal input
rlabel via1 s 675208 601808 675260 601860 6 porb_h
port 636 nsew signal input
rlabel via1 s 673736 601808 673788 601860 6 porb_h
port 636 nsew signal input
rlabel via1 s 675392 605752 675444 605804 6 porb_h
port 636 nsew signal input
rlabel via1 s 675208 605752 675260 605804 6 porb_h
port 636 nsew signal input
rlabel via1 s 673736 605752 673788 605804 6 porb_h
port 636 nsew signal input
rlabel via1 s 675392 646416 675444 646468 6 porb_h
port 636 nsew signal input
rlabel via1 s 673736 646416 673788 646468 6 porb_h
port 636 nsew signal input
rlabel via1 s 675392 651108 675444 651160 6 porb_h
port 636 nsew signal input
rlabel via1 s 673736 651108 673788 651160 6 porb_h
port 636 nsew signal input
rlabel via1 s 675392 692044 675444 692096 6 porb_h
port 636 nsew signal input
rlabel via1 s 675208 692044 675260 692096 6 porb_h
port 636 nsew signal input
rlabel via1 s 673736 692044 673788 692096 6 porb_h
port 636 nsew signal input
rlabel via1 s 675392 695920 675444 695972 6 porb_h
port 636 nsew signal input
rlabel via1 s 675208 695920 675260 695972 6 porb_h
port 636 nsew signal input
rlabel via1 s 673736 695920 673788 695972 6 porb_h
port 636 nsew signal input
rlabel via1 s 42340 718836 42392 718888 6 porb_h
port 636 nsew signal input
rlabel via1 s 42340 719040 42392 719092 6 porb_h
port 636 nsew signal input
rlabel via1 s 675392 736992 675444 737044 6 porb_h
port 636 nsew signal input
rlabel via1 s 675208 736992 675260 737044 6 porb_h
port 636 nsew signal input
rlabel via1 s 673736 736992 673788 737044 6 porb_h
port 636 nsew signal input
rlabel via1 s 675392 740936 675444 740988 6 porb_h
port 636 nsew signal input
rlabel via1 s 675208 740936 675260 740988 6 porb_h
port 636 nsew signal input
rlabel via1 s 673736 740936 673788 740988 6 porb_h
port 636 nsew signal input
rlabel via1 s 42340 743452 42392 743504 6 porb_h
port 636 nsew signal input
rlabel via1 s 41788 743452 41840 743504 6 porb_h
port 636 nsew signal input
rlabel via1 s 42340 747872 42392 747924 6 porb_h
port 636 nsew signal input
rlabel via1 s 41972 747872 42024 747924 6 porb_h
port 636 nsew signal input
rlabel via1 s 42432 756372 42484 756424 6 porb_h
port 636 nsew signal input
rlabel via1 s 42432 756576 42484 756628 6 porb_h
port 636 nsew signal input
rlabel via1 s 675392 781600 675444 781652 6 porb_h
port 636 nsew signal input
rlabel via1 s 675208 781600 675260 781652 6 porb_h
port 636 nsew signal input
rlabel via1 s 673736 781600 673788 781652 6 porb_h
port 636 nsew signal input
rlabel via1 s 675392 785952 675444 786004 6 porb_h
port 636 nsew signal input
rlabel via1 s 675208 785952 675260 786004 6 porb_h
port 636 nsew signal input
rlabel via1 s 673828 785952 673880 786004 6 porb_h
port 636 nsew signal input
rlabel via1 s 42432 786972 42484 787024 6 porb_h
port 636 nsew signal input
rlabel via1 s 41788 786972 41840 787024 6 porb_h
port 636 nsew signal input
rlabel via1 s 42524 791936 42576 791988 6 porb_h
port 636 nsew signal input
rlabel via1 s 41788 791936 41840 791988 6 porb_h
port 636 nsew signal input
rlabel via1 s 675300 871292 675352 871344 6 porb_h
port 636 nsew signal input
rlabel via1 s 673828 871292 673880 871344 6 porb_h
port 636 nsew signal input
rlabel via1 s 675392 875780 675444 875832 6 porb_h
port 636 nsew signal input
rlabel via1 s 673644 875780 673696 875832 6 porb_h
port 636 nsew signal input
rlabel via1 s 675392 960032 675444 960084 6 porb_h
port 636 nsew signal input
rlabel via1 s 673644 960032 673696 960084 6 porb_h
port 636 nsew signal input
rlabel via1 s 42524 961120 42576 961172 6 porb_h
port 636 nsew signal input
rlabel via1 s 41788 961120 41840 961172 6 porb_h
port 636 nsew signal input
rlabel via1 s 675392 965268 675444 965320 6 porb_h
port 636 nsew signal input
rlabel via1 s 673828 965268 673880 965320 6 porb_h
port 636 nsew signal input
rlabel via1 s 673828 990088 673880 990140 6 porb_h
port 636 nsew signal input
rlabel via1 s 634728 990088 634780 990140 6 porb_h
port 636 nsew signal input
rlabel via1 s 78864 990224 78916 990276 6 porb_h
port 636 nsew signal input
rlabel via1 s 42340 990224 42392 990276 6 porb_h
port 636 nsew signal input
rlabel via1 s 634728 990564 634780 990616 6 porb_h
port 636 nsew signal input
rlabel via1 s 632980 990564 633032 990616 6 porb_h
port 636 nsew signal input
rlabel via1 s 628656 990564 628708 990616 6 porb_h
port 636 nsew signal input
rlabel via1 s 531228 990564 531280 990616 6 porb_h
port 636 nsew signal input
rlabel via1 s 526904 990564 526956 990616 6 porb_h
port 636 nsew signal input
rlabel via1 s 479800 990564 479852 990616 6 porb_h
port 636 nsew signal input
rlabel via1 s 475476 990564 475528 990616 6 porb_h
port 636 nsew signal input
rlabel via1 s 390836 990564 390888 990616 6 porb_h
port 636 nsew signal input
rlabel via1 s 386512 990564 386564 990616 6 porb_h
port 636 nsew signal input
rlabel via1 s 274456 990564 274508 990616 6 porb_h
port 636 nsew signal input
rlabel via1 s 237380 990564 237432 990616 6 porb_h
port 636 nsew signal input
rlabel via1 s 233056 990564 233108 990616 6 porb_h
port 636 nsew signal input
rlabel via1 s 186044 990564 186096 990616 6 porb_h
port 636 nsew signal input
rlabel via1 s 181720 990564 181772 990616 6 porb_h
port 636 nsew signal input
rlabel via1 s 134616 990564 134668 990616 6 porb_h
port 636 nsew signal input
rlabel via1 s 130292 990564 130344 990616 6 porb_h
port 636 nsew signal input
rlabel via1 s 83188 990564 83240 990616 6 porb_h
port 636 nsew signal input
rlabel via1 s 78864 990564 78916 990616 6 porb_h
port 636 nsew signal input
rlabel via1 s 288992 990632 289044 990684 6 porb_h
port 636 nsew signal input
rlabel via1 s 284668 990632 284720 990684 6 porb_h
port 636 nsew signal input
rlabel via1 s 274732 990632 274784 990684 6 porb_h
port 636 nsew signal input
rlabel metal1 s 527450 44140 527514 44152 6 porb_h
port 636 nsew signal input
rlabel metal1 s 523126 44140 523190 44152 6 porb_h
port 636 nsew signal input
rlabel metal1 s 523126 44152 527514 44180 6 porb_h
port 636 nsew signal input
rlabel metal1 s 527450 44180 527514 44192 6 porb_h
port 636 nsew signal input
rlabel metal1 s 523126 44180 523190 44192 6 porb_h
port 636 nsew signal input
rlabel metal1 s 199654 44140 199718 44152 6 porb_h
port 636 nsew signal input
rlabel metal1 s 195330 44140 195394 44152 6 porb_h
port 636 nsew signal input
rlabel metal1 s 145098 44140 145162 44152 6 porb_h
port 636 nsew signal input
rlabel metal1 s 143626 44140 143690 44152 6 porb_h
port 636 nsew signal input
rlabel metal1 s 143626 44152 199718 44180 6 porb_h
port 636 nsew signal input
rlabel metal1 s 199654 44180 199718 44192 6 porb_h
port 636 nsew signal input
rlabel metal1 s 195330 44180 195394 44192 6 porb_h
port 636 nsew signal input
rlabel metal1 s 145098 44180 145162 44192 6 porb_h
port 636 nsew signal input
rlabel metal1 s 143626 44180 143690 44192 6 porb_h
port 636 nsew signal input
rlabel metal1 s 523144 44192 523172 44288 6 porb_h
port 636 nsew signal input
rlabel metal1 s 358722 44208 358786 44220 6 porb_h
port 636 nsew signal input
rlabel metal1 s 308214 44208 308278 44220 6 porb_h
port 636 nsew signal input
rlabel metal1 s 303890 44208 303954 44220 6 porb_h
port 636 nsew signal input
rlabel metal1 s 303890 44220 361574 44248 6 porb_h
port 636 nsew signal input
rlabel metal1 s 472618 44276 472682 44288 6 porb_h
port 636 nsew signal input
rlabel metal1 s 468294 44276 468358 44288 6 porb_h
port 636 nsew signal input
rlabel metal1 s 417878 44276 417942 44288 6 porb_h
port 636 nsew signal input
rlabel metal1 s 413554 44276 413618 44288 6 porb_h
port 636 nsew signal input
rlabel metal1 s 363046 44276 363110 44288 6 porb_h
port 636 nsew signal input
rlabel metal1 s 361546 44248 361574 44288 6 porb_h
port 636 nsew signal input
rlabel metal1 s 358722 44248 358786 44260 6 porb_h
port 636 nsew signal input
rlabel metal1 s 308214 44248 308278 44260 6 porb_h
port 636 nsew signal input
rlabel metal1 s 303890 44248 303954 44260 6 porb_h
port 636 nsew signal input
rlabel metal1 s 206986 44220 284294 44248 6 porb_h
port 636 nsew signal input
rlabel metal1 s 361546 44288 523172 44316 6 porb_h
port 636 nsew signal input
rlabel metal1 s 303908 44260 303936 44288 6 porb_h
port 636 nsew signal input
rlabel metal1 s 284266 44248 284294 44288 6 porb_h
port 636 nsew signal input
rlabel metal1 s 284266 44288 303936 44316 6 porb_h
port 636 nsew signal input
rlabel metal1 s 472618 44316 472682 44328 6 porb_h
port 636 nsew signal input
rlabel metal1 s 468294 44316 468358 44328 6 porb_h
port 636 nsew signal input
rlabel metal1 s 417878 44316 417942 44328 6 porb_h
port 636 nsew signal input
rlabel metal1 s 413554 44316 413618 44328 6 porb_h
port 636 nsew signal input
rlabel metal1 s 363046 44316 363110 44328 6 porb_h
port 636 nsew signal input
rlabel metal1 s 206986 44248 207014 44424 6 porb_h
port 636 nsew signal input
rlabel metal1 s 199654 44412 199718 44424 6 porb_h
port 636 nsew signal input
rlabel metal1 s 199654 44424 207014 44452 6 porb_h
port 636 nsew signal input
rlabel metal1 s 199654 44452 199718 44464 6 porb_h
port 636 nsew signal input
rlabel metal1 s 143626 45568 143690 45580 6 porb_h
port 636 nsew signal input
rlabel metal1 s 42334 45568 42398 45580 6 porb_h
port 636 nsew signal input
rlabel metal1 s 42334 45580 143690 45608 6 porb_h
port 636 nsew signal input
rlabel metal1 s 143626 45608 143690 45620 6 porb_h
port 636 nsew signal input
rlabel metal1 s 42334 45608 42398 45620 6 porb_h
port 636 nsew signal input
rlabel metal1 s 527450 46860 527514 46912 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673638 46928 673702 46940 6 porb_h
port 636 nsew signal input
rlabel metal1 s 527468 46912 527496 46940 6 porb_h
port 636 nsew signal input
rlabel metal1 s 527468 46940 673702 46968 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673638 46968 673702 46980 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 108400 675450 108412 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673638 108400 673702 108412 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673638 108412 675450 108440 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 108440 675450 108452 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673638 108440 673702 108452 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 113704 675450 113716 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673638 113704 673702 113716 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673638 113716 675450 113744 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 113744 675450 113756 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673638 113744 673702 113756 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675294 154096 675358 154108 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 154096 673794 154108 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 154108 675358 154136 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675294 154136 675358 154148 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 154136 673794 154148 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 158584 675450 158596 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 158584 673794 158596 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 158596 675450 158624 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 158624 675450 158636 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 158624 673794 158636 6 porb_h
port 636 nsew signal input
rlabel metal1 s 42334 197276 42398 197328 6 porb_h
port 636 nsew signal input
rlabel metal1 s 42352 197328 42380 197480 6 porb_h
port 636 nsew signal input
rlabel metal1 s 42334 197480 42398 197532 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 199044 675450 199056 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 199044 673794 199056 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 199056 675450 199084 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 199084 675450 199096 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 199084 673794 199096 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675294 203464 675358 203476 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 203464 673794 203476 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 203476 675358 203504 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675294 203504 675358 203516 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 203504 673794 203516 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 243788 675450 243800 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 243788 673794 243800 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 243800 675450 243828 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 243828 675450 243840 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 243828 673794 243840 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 249092 675450 249104 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 249092 673794 249104 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 249104 675450 249132 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 249132 675450 249144 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 249132 673794 249144 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 288804 675450 288816 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 288804 673794 288816 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 288816 675450 288844 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 288844 675450 288856 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 288844 673794 288856 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675294 293700 675358 293712 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673822 293700 673886 293712 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673822 293712 675358 293740 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675294 293740 675358 293752 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673822 293740 673886 293752 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 334228 675450 334240 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673822 334228 673886 334240 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673822 334240 675450 334268 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 334268 675450 334280 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673822 334268 673886 334280 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 338784 675450 338796 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673638 338784 673702 338796 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673638 338796 675450 338824 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 338824 675450 338836 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673638 338824 673702 338836 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 379040 675450 379052 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673638 379040 673702 379052 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673638 379052 675450 379080 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 379080 675450 379092 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673638 379080 673702 379092 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 557268 675450 557280 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675202 557268 675266 557280 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675202 557280 675450 557308 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 557308 675450 557320 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675202 557308 675266 557320 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 561212 675450 561224 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675202 561212 675266 561224 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 561212 673794 561224 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 561224 675450 561252 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 561252 675450 561264 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675202 561252 675266 561264 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 561252 673794 561264 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 601808 675450 601820 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675202 601808 675266 601820 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 601808 673794 601820 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 601820 675450 601848 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 601848 675450 601860 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675202 601848 675266 601860 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 601848 673794 601860 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 605752 675450 605764 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675202 605752 675266 605764 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 605752 673794 605764 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 605764 675450 605792 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 605792 675450 605804 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675202 605792 675266 605804 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 605792 673794 605804 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 646416 675450 646428 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 646416 673794 646428 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 646428 675450 646456 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 646456 675450 646468 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 646456 673794 646468 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 651108 675450 651120 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 651108 673794 651120 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 651120 675450 651148 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 651148 675450 651160 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 651148 673794 651160 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 692044 675450 692056 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675202 692044 675266 692056 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 692044 673794 692056 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 692056 675450 692084 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 692084 675450 692096 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675202 692084 675266 692096 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 692084 673794 692096 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 695920 675450 695932 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675202 695920 675266 695932 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 695920 673794 695932 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 695932 675450 695960 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 695960 675450 695972 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675202 695960 675266 695972 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 695960 673794 695972 6 porb_h
port 636 nsew signal input
rlabel metal1 s 42334 718836 42398 718888 6 porb_h
port 636 nsew signal input
rlabel metal1 s 42352 718888 42380 719040 6 porb_h
port 636 nsew signal input
rlabel metal1 s 42334 719040 42398 719092 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 736992 675450 737004 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675202 736992 675266 737004 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 736992 673794 737004 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 737004 675450 737032 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 737032 675450 737044 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675202 737032 675266 737044 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 737032 673794 737044 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 740936 675450 740948 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675202 740936 675266 740948 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 740936 673794 740948 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 740948 675450 740976 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 740976 675450 740988 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675202 740976 675266 740988 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 740976 673794 740988 6 porb_h
port 636 nsew signal input
rlabel metal1 s 42334 743452 42398 743464 6 porb_h
port 636 nsew signal input
rlabel metal1 s 41782 743452 41846 743464 6 porb_h
port 636 nsew signal input
rlabel metal1 s 41782 743464 42398 743492 6 porb_h
port 636 nsew signal input
rlabel metal1 s 42334 743492 42398 743504 6 porb_h
port 636 nsew signal input
rlabel metal1 s 41782 743492 41846 743504 6 porb_h
port 636 nsew signal input
rlabel metal1 s 42334 747872 42398 747884 6 porb_h
port 636 nsew signal input
rlabel metal1 s 41966 747872 42030 747884 6 porb_h
port 636 nsew signal input
rlabel metal1 s 41966 747884 42398 747912 6 porb_h
port 636 nsew signal input
rlabel metal1 s 42334 747912 42398 747924 6 porb_h
port 636 nsew signal input
rlabel metal1 s 41966 747912 42030 747924 6 porb_h
port 636 nsew signal input
rlabel metal1 s 42426 756372 42490 756424 6 porb_h
port 636 nsew signal input
rlabel metal1 s 42444 756424 42472 756576 6 porb_h
port 636 nsew signal input
rlabel metal1 s 42426 756576 42490 756628 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 781600 675450 781612 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675202 781600 675266 781612 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 781600 673794 781612 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 781612 675450 781640 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 781640 675450 781652 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675202 781640 675266 781652 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673730 781640 673794 781652 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 785952 675450 785964 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675202 785952 675266 785964 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673822 785952 673886 785964 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673822 785964 675450 785992 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 785992 675450 786004 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675202 785992 675266 786004 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673822 785992 673886 786004 6 porb_h
port 636 nsew signal input
rlabel metal1 s 42426 786972 42490 786984 6 porb_h
port 636 nsew signal input
rlabel metal1 s 41782 786972 41846 786984 6 porb_h
port 636 nsew signal input
rlabel metal1 s 41782 786984 42490 787012 6 porb_h
port 636 nsew signal input
rlabel metal1 s 42426 787012 42490 787024 6 porb_h
port 636 nsew signal input
rlabel metal1 s 41782 787012 41846 787024 6 porb_h
port 636 nsew signal input
rlabel metal1 s 42518 791936 42582 791948 6 porb_h
port 636 nsew signal input
rlabel metal1 s 41782 791936 41846 791948 6 porb_h
port 636 nsew signal input
rlabel metal1 s 41782 791948 42582 791976 6 porb_h
port 636 nsew signal input
rlabel metal1 s 42518 791976 42582 791988 6 porb_h
port 636 nsew signal input
rlabel metal1 s 41782 791976 41846 791988 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675294 871292 675358 871304 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673822 871292 673886 871304 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673822 871304 675358 871332 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675294 871332 675358 871344 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673822 871332 673886 871344 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 875780 675450 875792 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673638 875780 673702 875792 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673638 875792 675450 875820 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 875820 675450 875832 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673638 875820 673702 875832 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 960032 675450 960044 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673638 960032 673702 960044 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673638 960044 675450 960072 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 960072 675450 960084 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673638 960072 673702 960084 6 porb_h
port 636 nsew signal input
rlabel metal1 s 42518 961120 42582 961132 6 porb_h
port 636 nsew signal input
rlabel metal1 s 41782 961120 41846 961132 6 porb_h
port 636 nsew signal input
rlabel metal1 s 41782 961132 42582 961160 6 porb_h
port 636 nsew signal input
rlabel metal1 s 42518 961160 42582 961172 6 porb_h
port 636 nsew signal input
rlabel metal1 s 41782 961160 41846 961172 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 965268 675450 965280 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673822 965268 673886 965280 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673822 965280 675450 965308 6 porb_h
port 636 nsew signal input
rlabel metal1 s 675386 965308 675450 965320 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673822 965308 673886 965320 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673822 990088 673886 990100 6 porb_h
port 636 nsew signal input
rlabel metal1 s 634722 990088 634786 990100 6 porb_h
port 636 nsew signal input
rlabel metal1 s 634722 990100 673886 990128 6 porb_h
port 636 nsew signal input
rlabel metal1 s 673822 990128 673886 990140 6 porb_h
port 636 nsew signal input
rlabel metal1 s 634722 990128 634786 990140 6 porb_h
port 636 nsew signal input
rlabel metal1 s 78858 990224 78922 990236 6 porb_h
port 636 nsew signal input
rlabel metal1 s 42334 990224 42398 990236 6 porb_h
port 636 nsew signal input
rlabel metal1 s 42334 990236 78922 990264 6 porb_h
port 636 nsew signal input
rlabel metal1 s 78858 990264 78922 990276 6 porb_h
port 636 nsew signal input
rlabel metal1 s 42334 990264 42398 990276 6 porb_h
port 636 nsew signal input
rlabel metal1 s 634722 990564 634786 990576 6 porb_h
port 636 nsew signal input
rlabel metal1 s 632974 990564 633038 990576 6 porb_h
port 636 nsew signal input
rlabel metal1 s 628650 990564 628714 990576 6 porb_h
port 636 nsew signal input
rlabel metal1 s 531222 990564 531286 990576 6 porb_h
port 636 nsew signal input
rlabel metal1 s 526898 990564 526962 990576 6 porb_h
port 636 nsew signal input
rlabel metal1 s 479794 990564 479858 990576 6 porb_h
port 636 nsew signal input
rlabel metal1 s 475470 990564 475534 990576 6 porb_h
port 636 nsew signal input
rlabel metal1 s 390830 990564 390894 990576 6 porb_h
port 636 nsew signal input
rlabel metal1 s 386506 990564 386570 990576 6 porb_h
port 636 nsew signal input
rlabel metal1 s 386506 990576 634786 990604 6 porb_h
port 636 nsew signal input
rlabel metal1 s 634722 990604 634786 990616 6 porb_h
port 636 nsew signal input
rlabel metal1 s 632974 990604 633038 990616 6 porb_h
port 636 nsew signal input
rlabel metal1 s 628650 990604 628714 990616 6 porb_h
port 636 nsew signal input
rlabel metal1 s 531222 990604 531286 990616 6 porb_h
port 636 nsew signal input
rlabel metal1 s 526898 990604 526962 990616 6 porb_h
port 636 nsew signal input
rlabel metal1 s 479794 990604 479858 990616 6 porb_h
port 636 nsew signal input
rlabel metal1 s 475470 990604 475534 990616 6 porb_h
port 636 nsew signal input
rlabel metal1 s 390830 990604 390894 990616 6 porb_h
port 636 nsew signal input
rlabel metal1 s 386506 990604 386570 990616 6 porb_h
port 636 nsew signal input
rlabel metal1 s 274450 990564 274514 990576 6 porb_h
port 636 nsew signal input
rlabel metal1 s 237374 990564 237438 990576 6 porb_h
port 636 nsew signal input
rlabel metal1 s 233050 990564 233114 990576 6 porb_h
port 636 nsew signal input
rlabel metal1 s 186038 990564 186102 990576 6 porb_h
port 636 nsew signal input
rlabel metal1 s 181714 990564 181778 990576 6 porb_h
port 636 nsew signal input
rlabel metal1 s 134610 990564 134674 990576 6 porb_h
port 636 nsew signal input
rlabel metal1 s 130286 990564 130350 990576 6 porb_h
port 636 nsew signal input
rlabel metal1 s 83182 990564 83246 990576 6 porb_h
port 636 nsew signal input
rlabel metal1 s 78858 990564 78922 990576 6 porb_h
port 636 nsew signal input
rlabel metal1 s 78858 990576 274514 990604 6 porb_h
port 636 nsew signal input
rlabel metal1 s 274450 990604 274514 990616 6 porb_h
port 636 nsew signal input
rlabel metal1 s 237374 990604 237438 990616 6 porb_h
port 636 nsew signal input
rlabel metal1 s 233050 990604 233114 990616 6 porb_h
port 636 nsew signal input
rlabel metal1 s 186038 990604 186102 990616 6 porb_h
port 636 nsew signal input
rlabel metal1 s 181714 990604 181778 990616 6 porb_h
port 636 nsew signal input
rlabel metal1 s 134610 990604 134674 990616 6 porb_h
port 636 nsew signal input
rlabel metal1 s 130286 990604 130350 990616 6 porb_h
port 636 nsew signal input
rlabel metal1 s 83182 990604 83246 990616 6 porb_h
port 636 nsew signal input
rlabel metal1 s 78858 990604 78922 990616 6 porb_h
port 636 nsew signal input
rlabel metal1 s 386524 990616 386552 990644 6 porb_h
port 636 nsew signal input
rlabel metal1 s 288986 990632 289050 990644 6 porb_h
port 636 nsew signal input
rlabel metal1 s 284662 990632 284726 990644 6 porb_h
port 636 nsew signal input
rlabel metal1 s 274726 990632 274790 990644 6 porb_h
port 636 nsew signal input
rlabel metal1 s 274726 990644 386552 990672 6 porb_h
port 636 nsew signal input
rlabel metal1 s 288986 990672 289050 990684 6 porb_h
port 636 nsew signal input
rlabel metal1 s 284662 990672 284726 990684 6 porb_h
port 636 nsew signal input
rlabel metal1 s 274726 990672 274790 990684 6 porb_h
port 636 nsew signal input
rlabel metal5 s 133840 6675 146380 19198 6 resetb
port 637 nsew signal input
rlabel metal3 s 141820 37046 141966 37818 6 resetb_core_h
port 638 nsew signal output
rlabel metal3 s 141667 37818 141966 37911 6 resetb_core_h
port 638 nsew signal output
rlabel metal3 s 141873 37911 141966 37971 6 resetb_core_h
port 638 nsew signal output
rlabel metal3 s 141667 37911 141820 37971 6 resetb_core_h
port 638 nsew signal output
rlabel metal3 s 141667 37971 141873 38031 6 resetb_core_h
port 638 nsew signal output
rlabel metal3 s 141667 38031 141813 40000 6 resetb_core_h
port 638 nsew signal output
rlabel metal5 s 93607 36343 132793 36993 6 vdda
port 639 nsew signal bidirectional
rlabel metal5 s 93546 28653 132854 30453 6 vssa
port 640 nsew signal bidirectional
rlabel metal5 s 93546 30773 132854 31663 6 vssd
port 641 nsew signal bidirectional
rlabel metal5 s 697980 909666 711433 920546 6 vccd1_pad
port 642 nsew signal bidirectional
rlabel metal5 s 698624 819822 710789 831990 6 vdda1_pad
port 643 nsew signal bidirectional
rlabel metal5 s 698624 505222 710789 517390 6 vdda1_pad2
port 644 nsew signal bidirectional
rlabel metal5 s 577010 1018624 589178 1030789 6 vssa1_pad
port 645 nsew signal bidirectional
rlabel metal5 s 698624 417022 710789 429190 6 vssa1_pad2
port 646 nsew signal bidirectional
rlabel metal4 s 679377 430346 680307 460054 6 vccd1
port 647 nsew signal bidirectional
rlabel metal4 s 680587 430407 681277 459993 6 vdda1
port 648 nsew signal bidirectional
rlabel metal4 s 688881 430346 688947 554382 6 vssa1
port 649 nsew signal bidirectional
rlabel metal3 s 678000 469900 685920 474700 6 vssd1
port 650 nsew signal bidirectional
rlabel metal5 s 697980 461866 711433 472746 6 vssd1_pad
port 651 nsew signal bidirectional
rlabel metal5 s 6167 914054 19620 924934 6 vccd2_pad
port 652 nsew signal bidirectional
rlabel metal5 s 6811 484410 18976 496578 6 vdda2_pad
port 653 nsew signal bidirectional
rlabel metal5 s 6811 829010 18976 841178 6 vssa2_pad
port 654 nsew signal bidirectional
rlabel metal4 s 38503 455546 39593 483254 6 vccd
port 655 nsew signal bidirectional
rlabel metal4 s 37293 455546 38223 483254 6 vccd2
port 656 nsew signal bidirectional
rlabel metal4 s 36323 455607 37013 483193 6 vdda2
port 657 nsew signal bidirectional
rlabel metal4 s 32933 455546 33623 483254 6 vddio
port 658 nsew signal bidirectional
rlabel metal4 s 28653 407018 28719 525722 6 vssa2
port 659 nsew signal bidirectional
rlabel metal3 s 31680 440900 39600 445700 6 vssd2
port 660 nsew signal bidirectional
rlabel metal5 s 6167 442854 19620 453734 6 vssd2_pad
port 661 nsew signal bidirectional
rlabel metal4 s 0 455546 4843 455800 6 vssio
port 662 nsew signal bidirectional
rlabel metal4 s 7 455800 4843 456094 6 vssio
port 662 nsew signal bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 717600 1037600
string LEFview TRUE
string GDS_FILE /project/openlane/chip_io/runs/chip_io/results/magic/chip_io.gds
string GDS_END 36507134
string GDS_START 36076962
<< end >>

