VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravel
  CLASS BLOCK ;
  FOREIGN caravel ;
  ORIGIN 0.000 0.000 ;
  SIZE 3200.000 BY 5300.000 ;
  OBS
      LAYER li1 ;
        RECT 0.220 0.220 3199.780 5299.705 ;
      LAYER met1 ;
        RECT 0.000 0.000 3200.000 5300.000 ;
      LAYER met2 ;
        RECT 0.000 0.000 3200.000 5300.000 ;
      LAYER met3 ;
        RECT 0.000 0.000 3200.000 5300.000 ;
      LAYER met4 ;
        RECT 0.000 0.000 3200.000 5300.000 ;
      LAYER met5 ;
        RECT 0.000 0.000 3200.000 5300.000 ;
  END
END caravel
END LIBRARY

