magic
tech sky130A
magscale 1 2
timestamp 1607580681
<< metal1 >>
rect 439216 1005745 439222 1005797
rect 439274 1005785 439280 1005797
rect 466576 1005785 466582 1005797
rect 439274 1005757 466582 1005785
rect 439274 1005745 439280 1005757
rect 466576 1005745 466582 1005757
rect 466634 1005745 466640 1005797
rect 371824 1005711 371830 1005723
rect 370786 1005683 371830 1005711
rect 92368 1005523 92374 1005575
rect 92426 1005563 92432 1005575
rect 370786 1005563 370814 1005683
rect 371824 1005671 371830 1005683
rect 371882 1005671 371888 1005723
rect 440656 1005671 440662 1005723
rect 440714 1005711 440720 1005723
rect 446416 1005711 446422 1005723
rect 440714 1005683 446422 1005711
rect 440714 1005671 440720 1005683
rect 446416 1005671 446422 1005683
rect 446474 1005671 446480 1005723
rect 383632 1005637 383638 1005649
rect 92426 1005535 108638 1005563
rect 92426 1005523 92432 1005535
rect 108610 1005501 108638 1005535
rect 357922 1005535 370814 1005563
rect 370882 1005609 383638 1005637
rect 357922 1005501 357950 1005535
rect 108592 1005449 108598 1005501
rect 108650 1005449 108656 1005501
rect 357904 1005449 357910 1005501
rect 357962 1005449 357968 1005501
rect 365008 1005449 365014 1005501
rect 365066 1005489 365072 1005501
rect 370882 1005489 370910 1005609
rect 383632 1005597 383638 1005609
rect 383690 1005597 383696 1005649
rect 466480 1005563 466486 1005575
rect 430786 1005535 466486 1005563
rect 430786 1005501 430814 1005535
rect 466480 1005523 466486 1005535
rect 466538 1005523 466544 1005575
rect 380560 1005489 380566 1005501
rect 365066 1005461 370910 1005489
rect 370978 1005461 380566 1005489
rect 365066 1005449 365072 1005461
rect 93616 1005375 93622 1005427
rect 93674 1005415 93680 1005427
rect 114160 1005415 114166 1005427
rect 93674 1005387 114166 1005415
rect 93674 1005375 93680 1005387
rect 114160 1005375 114166 1005387
rect 114218 1005375 114224 1005427
rect 298096 1005375 298102 1005427
rect 298154 1005415 298160 1005427
rect 308752 1005415 308758 1005427
rect 298154 1005387 308758 1005415
rect 298154 1005375 298160 1005387
rect 308752 1005375 308758 1005387
rect 308810 1005375 308816 1005427
rect 364144 1005375 364150 1005427
rect 364202 1005415 364208 1005427
rect 370978 1005415 371006 1005461
rect 380560 1005449 380566 1005461
rect 380618 1005449 380624 1005501
rect 430768 1005449 430774 1005501
rect 430826 1005449 430832 1005501
rect 430864 1005449 430870 1005501
rect 430922 1005489 430928 1005501
rect 446320 1005489 446326 1005501
rect 430922 1005461 446326 1005489
rect 430922 1005449 430928 1005461
rect 446320 1005449 446326 1005461
rect 446378 1005449 446384 1005501
rect 446416 1005449 446422 1005501
rect 446474 1005489 446480 1005501
rect 471856 1005489 471862 1005501
rect 446474 1005461 471862 1005489
rect 446474 1005449 446480 1005461
rect 471856 1005449 471862 1005461
rect 471914 1005449 471920 1005501
rect 364202 1005387 371006 1005415
rect 364202 1005375 364208 1005387
rect 371056 1005375 371062 1005427
rect 371114 1005415 371120 1005427
rect 380464 1005415 380470 1005427
rect 371114 1005387 380470 1005415
rect 371114 1005375 371120 1005387
rect 380464 1005375 380470 1005387
rect 380522 1005375 380528 1005427
rect 439216 1005415 439222 1005427
rect 429154 1005387 439222 1005415
rect 298384 1005301 298390 1005353
rect 298442 1005341 298448 1005353
rect 309616 1005341 309622 1005353
rect 298442 1005313 309622 1005341
rect 298442 1005301 298448 1005313
rect 309616 1005301 309622 1005313
rect 309674 1005301 309680 1005353
rect 366736 1005301 366742 1005353
rect 366794 1005341 366800 1005353
rect 380368 1005341 380374 1005353
rect 366794 1005313 380374 1005341
rect 366794 1005301 366800 1005313
rect 380368 1005301 380374 1005313
rect 380426 1005301 380432 1005353
rect 424528 1005301 424534 1005353
rect 424586 1005341 424592 1005353
rect 429154 1005341 429182 1005387
rect 439216 1005375 439222 1005387
rect 439274 1005375 439280 1005427
rect 439408 1005375 439414 1005427
rect 439466 1005415 439472 1005427
rect 470896 1005415 470902 1005427
rect 439466 1005387 470902 1005415
rect 439466 1005375 439472 1005387
rect 470896 1005375 470902 1005387
rect 470954 1005375 470960 1005427
rect 501136 1005375 501142 1005427
rect 501194 1005415 501200 1005427
rect 518320 1005415 518326 1005427
rect 501194 1005387 518326 1005415
rect 501194 1005375 501200 1005387
rect 518320 1005375 518326 1005387
rect 518378 1005375 518384 1005427
rect 460816 1005341 460822 1005353
rect 424586 1005313 429182 1005341
rect 437314 1005313 460822 1005341
rect 424586 1005301 424592 1005313
rect 217264 1005227 217270 1005279
rect 217322 1005267 217328 1005279
rect 218896 1005267 218902 1005279
rect 217322 1005239 218902 1005267
rect 217322 1005227 217328 1005239
rect 218896 1005227 218902 1005239
rect 218954 1005227 218960 1005279
rect 298288 1005227 298294 1005279
rect 298346 1005267 298352 1005279
rect 307984 1005267 307990 1005279
rect 298346 1005239 307990 1005267
rect 298346 1005227 298352 1005239
rect 307984 1005227 307990 1005239
rect 308042 1005227 308048 1005279
rect 318640 1005227 318646 1005279
rect 318698 1005267 318704 1005279
rect 331120 1005267 331126 1005279
rect 318698 1005239 331126 1005267
rect 318698 1005227 318704 1005239
rect 331120 1005227 331126 1005239
rect 331178 1005227 331184 1005279
rect 365776 1005227 365782 1005279
rect 365834 1005267 365840 1005279
rect 380272 1005267 380278 1005279
rect 365834 1005239 380278 1005267
rect 365834 1005227 365840 1005239
rect 380272 1005227 380278 1005239
rect 380330 1005227 380336 1005279
rect 425296 1005227 425302 1005279
rect 425354 1005267 425360 1005279
rect 437314 1005267 437342 1005313
rect 460816 1005301 460822 1005313
rect 460874 1005301 460880 1005353
rect 554512 1005301 554518 1005353
rect 554570 1005341 554576 1005353
rect 572848 1005341 572854 1005353
rect 554570 1005313 572854 1005341
rect 554570 1005301 554576 1005313
rect 572848 1005301 572854 1005313
rect 572906 1005301 572912 1005353
rect 439024 1005267 439030 1005279
rect 425354 1005239 437342 1005267
rect 437794 1005239 439030 1005267
rect 425354 1005227 425360 1005239
rect 93712 1005153 93718 1005205
rect 93770 1005193 93776 1005205
rect 115216 1005193 115222 1005205
rect 93770 1005165 115222 1005193
rect 93770 1005153 93776 1005165
rect 115216 1005153 115222 1005165
rect 115274 1005153 115280 1005205
rect 299920 1005153 299926 1005205
rect 299978 1005193 299984 1005205
rect 315184 1005193 315190 1005205
rect 299978 1005165 315190 1005193
rect 299978 1005153 299984 1005165
rect 315184 1005153 315190 1005165
rect 315242 1005153 315248 1005205
rect 325456 1005153 325462 1005205
rect 325514 1005193 325520 1005205
rect 331216 1005193 331222 1005205
rect 325514 1005165 331222 1005193
rect 325514 1005153 325520 1005165
rect 331216 1005153 331222 1005165
rect 331274 1005153 331280 1005205
rect 363472 1005153 363478 1005205
rect 363530 1005193 363536 1005205
rect 371056 1005193 371062 1005205
rect 363530 1005165 371062 1005193
rect 363530 1005153 363536 1005165
rect 371056 1005153 371062 1005165
rect 371114 1005153 371120 1005205
rect 371824 1005153 371830 1005205
rect 371882 1005193 371888 1005205
rect 380176 1005193 380182 1005205
rect 371882 1005165 380182 1005193
rect 371882 1005153 371888 1005165
rect 380176 1005153 380182 1005165
rect 380234 1005153 380240 1005205
rect 426064 1005153 426070 1005205
rect 426122 1005193 426128 1005205
rect 437584 1005193 437590 1005205
rect 426122 1005165 437590 1005193
rect 426122 1005153 426128 1005165
rect 437584 1005153 437590 1005165
rect 437642 1005153 437648 1005205
rect 433168 1005079 433174 1005131
rect 433226 1005119 433232 1005131
rect 437794 1005119 437822 1005239
rect 439024 1005227 439030 1005239
rect 439082 1005227 439088 1005279
rect 471472 1005267 471478 1005279
rect 439138 1005239 471478 1005267
rect 437872 1005153 437878 1005205
rect 437930 1005193 437936 1005205
rect 439138 1005193 439166 1005239
rect 471472 1005227 471478 1005239
rect 471530 1005227 471536 1005279
rect 504592 1005227 504598 1005279
rect 504650 1005267 504656 1005279
rect 521392 1005267 521398 1005279
rect 504650 1005239 521398 1005267
rect 504650 1005227 504656 1005239
rect 521392 1005227 521398 1005239
rect 521450 1005227 521456 1005279
rect 555760 1005227 555766 1005279
rect 555818 1005267 555824 1005279
rect 573040 1005267 573046 1005279
rect 555818 1005239 573046 1005267
rect 555818 1005227 555824 1005239
rect 573040 1005227 573046 1005239
rect 573098 1005227 573104 1005279
rect 437930 1005165 439166 1005193
rect 437930 1005153 437936 1005165
rect 439216 1005153 439222 1005205
rect 439274 1005193 439280 1005205
rect 471664 1005193 471670 1005205
rect 439274 1005165 471670 1005193
rect 439274 1005153 439280 1005165
rect 471664 1005153 471670 1005165
rect 471722 1005153 471728 1005205
rect 500752 1005153 500758 1005205
rect 500810 1005193 500816 1005205
rect 512560 1005193 512566 1005205
rect 500810 1005165 512566 1005193
rect 500810 1005153 500816 1005165
rect 512560 1005153 512566 1005165
rect 512618 1005153 512624 1005205
rect 518320 1005153 518326 1005205
rect 518378 1005193 518384 1005205
rect 521584 1005193 521590 1005205
rect 518378 1005165 521590 1005193
rect 518378 1005153 518384 1005165
rect 521584 1005153 521590 1005165
rect 521642 1005153 521648 1005205
rect 553744 1005153 553750 1005205
rect 553802 1005193 553808 1005205
rect 572944 1005193 572950 1005205
rect 553802 1005165 572950 1005193
rect 553802 1005153 553808 1005165
rect 572944 1005153 572950 1005165
rect 573002 1005153 573008 1005205
rect 433226 1005091 437822 1005119
rect 433226 1005079 433232 1005091
rect 435568 1005005 435574 1005057
rect 435626 1005045 435632 1005057
rect 440656 1005045 440662 1005057
rect 435626 1005017 440662 1005045
rect 435626 1005005 435632 1005017
rect 440656 1005005 440662 1005017
rect 440714 1005005 440720 1005057
rect 359920 1003969 359926 1004021
rect 359978 1004009 359984 1004021
rect 380080 1004009 380086 1004021
rect 359978 1003981 380086 1004009
rect 359978 1003969 359984 1003981
rect 380080 1003969 380086 1003981
rect 380138 1003969 380144 1004021
rect 423376 1003895 423382 1003947
rect 423434 1003935 423440 1003947
rect 453328 1003935 453334 1003947
rect 423434 1003907 453334 1003935
rect 423434 1003895 423440 1003907
rect 453328 1003895 453334 1003907
rect 453386 1003895 453392 1003947
rect 359056 1003821 359062 1003873
rect 359114 1003861 359120 1003873
rect 377488 1003861 377494 1003873
rect 359114 1003833 377494 1003861
rect 359114 1003821 359120 1003833
rect 377488 1003821 377494 1003833
rect 377546 1003821 377552 1003873
rect 426448 1003821 426454 1003873
rect 426506 1003861 426512 1003873
rect 463696 1003861 463702 1003873
rect 426506 1003833 463702 1003861
rect 426506 1003821 426512 1003833
rect 463696 1003821 463702 1003833
rect 463754 1003821 463760 1003873
rect 552592 1003821 552598 1003873
rect 552650 1003861 552656 1003873
rect 572656 1003861 572662 1003873
rect 552650 1003833 572662 1003861
rect 552650 1003821 552656 1003833
rect 572656 1003821 572662 1003833
rect 572714 1003821 572720 1003873
rect 358384 1003747 358390 1003799
rect 358442 1003787 358448 1003799
rect 377392 1003787 377398 1003799
rect 358442 1003759 377398 1003787
rect 358442 1003747 358448 1003759
rect 377392 1003747 377398 1003759
rect 377450 1003747 377456 1003799
rect 422512 1003747 422518 1003799
rect 422570 1003787 422576 1003799
rect 461008 1003787 461014 1003799
rect 422570 1003759 461014 1003787
rect 422570 1003747 422576 1003759
rect 461008 1003747 461014 1003759
rect 461066 1003747 461072 1003799
rect 499984 1003747 499990 1003799
rect 500042 1003787 500048 1003799
rect 515536 1003787 515542 1003799
rect 500042 1003759 515542 1003787
rect 500042 1003747 500048 1003759
rect 515536 1003747 515542 1003759
rect 515594 1003747 515600 1003799
rect 556528 1003747 556534 1003799
rect 556586 1003787 556592 1003799
rect 574000 1003787 574006 1003799
rect 556586 1003759 574006 1003787
rect 556586 1003747 556592 1003759
rect 574000 1003747 574006 1003759
rect 574058 1003747 574064 1003799
rect 360688 1003673 360694 1003725
rect 360746 1003713 360752 1003725
rect 377296 1003713 377302 1003725
rect 360746 1003685 377302 1003713
rect 360746 1003673 360752 1003685
rect 377296 1003673 377302 1003685
rect 377354 1003673 377360 1003725
rect 428080 1003673 428086 1003725
rect 428138 1003713 428144 1003725
rect 472048 1003713 472054 1003725
rect 428138 1003685 472054 1003713
rect 428138 1003673 428144 1003685
rect 472048 1003673 472054 1003685
rect 472106 1003673 472112 1003725
rect 551728 1003673 551734 1003725
rect 551786 1003713 551792 1003725
rect 572752 1003713 572758 1003725
rect 551786 1003685 572758 1003713
rect 551786 1003673 551792 1003685
rect 572752 1003673 572758 1003685
rect 572810 1003673 572816 1003725
rect 559216 1002637 559222 1002689
rect 559274 1002677 559280 1002689
rect 566320 1002677 566326 1002689
rect 559274 1002649 566326 1002677
rect 559274 1002637 559280 1002649
rect 566320 1002637 566326 1002649
rect 566378 1002637 566384 1002689
rect 559984 1002563 559990 1002615
rect 560042 1002603 560048 1002615
rect 566128 1002603 566134 1002615
rect 560042 1002575 566134 1002603
rect 560042 1002563 560048 1002575
rect 566128 1002563 566134 1002575
rect 566186 1002563 566192 1002615
rect 144016 1002489 144022 1002541
rect 144074 1002529 144080 1002541
rect 150352 1002529 150358 1002541
rect 144074 1002501 150358 1002529
rect 144074 1002489 144080 1002501
rect 150352 1002489 150358 1002501
rect 150410 1002489 150416 1002541
rect 299632 1002489 299638 1002541
rect 299690 1002529 299696 1002541
rect 307600 1002529 307606 1002541
rect 299690 1002501 307606 1002529
rect 299690 1002489 299696 1002501
rect 307600 1002489 307606 1002501
rect 307658 1002489 307664 1002541
rect 503440 1002489 503446 1002541
rect 503498 1002529 503504 1002541
rect 515440 1002529 515446 1002541
rect 503498 1002501 515446 1002529
rect 503498 1002489 503504 1002501
rect 515440 1002489 515446 1002501
rect 515498 1002489 515504 1002541
rect 562192 1002489 562198 1002541
rect 562250 1002529 562256 1002541
rect 567568 1002529 567574 1002541
rect 562250 1002501 567574 1002529
rect 562250 1002489 562256 1002501
rect 567568 1002489 567574 1002501
rect 567626 1002489 567632 1002541
rect 246544 1002415 246550 1002467
rect 246602 1002455 246608 1002467
rect 254032 1002455 254038 1002467
rect 246602 1002427 254038 1002455
rect 246602 1002415 246608 1002427
rect 254032 1002415 254038 1002427
rect 254090 1002415 254096 1002467
rect 299536 1002415 299542 1002467
rect 299594 1002455 299600 1002467
rect 305584 1002455 305590 1002467
rect 299594 1002427 305590 1002455
rect 299594 1002415 299600 1002427
rect 305584 1002415 305590 1002427
rect 305642 1002415 305648 1002467
rect 502768 1002415 502774 1002467
rect 502826 1002455 502832 1002467
rect 513520 1002455 513526 1002467
rect 502826 1002427 513526 1002455
rect 502826 1002415 502832 1002427
rect 513520 1002415 513526 1002427
rect 513578 1002415 513584 1002467
rect 564592 1002415 564598 1002467
rect 564650 1002455 564656 1002467
rect 568720 1002455 568726 1002467
rect 564650 1002427 568726 1002455
rect 564650 1002415 564656 1002427
rect 568720 1002415 568726 1002427
rect 568778 1002415 568784 1002467
rect 143920 1002341 143926 1002393
rect 143978 1002381 143984 1002393
rect 153616 1002381 153622 1002393
rect 143978 1002353 153622 1002381
rect 143978 1002341 143984 1002353
rect 153616 1002341 153622 1002353
rect 153674 1002341 153680 1002393
rect 299824 1002341 299830 1002393
rect 299882 1002381 299888 1002393
rect 306544 1002381 306550 1002393
rect 299882 1002353 306550 1002381
rect 299882 1002341 299888 1002353
rect 306544 1002341 306550 1002353
rect 306602 1002341 306608 1002393
rect 505072 1002341 505078 1002393
rect 505130 1002381 505136 1002393
rect 521488 1002381 521494 1002393
rect 505130 1002353 521494 1002381
rect 505130 1002341 505136 1002353
rect 521488 1002341 521494 1002353
rect 521546 1002341 521552 1002393
rect 560464 1002341 560470 1002393
rect 560522 1002381 560528 1002393
rect 564784 1002381 564790 1002393
rect 560522 1002353 564790 1002381
rect 560522 1002341 560528 1002353
rect 564784 1002341 564790 1002353
rect 564842 1002341 564848 1002393
rect 143728 1002267 143734 1002319
rect 143786 1002307 143792 1002319
rect 178480 1002307 178486 1002319
rect 143786 1002279 178486 1002307
rect 143786 1002267 143792 1002279
rect 178480 1002267 178486 1002279
rect 178538 1002267 178544 1002319
rect 246736 1002267 246742 1002319
rect 246794 1002307 246800 1002319
rect 253168 1002307 253174 1002319
rect 246794 1002279 253174 1002307
rect 246794 1002267 246800 1002279
rect 253168 1002267 253174 1002279
rect 253226 1002267 253232 1002319
rect 299728 1002267 299734 1002319
rect 299786 1002307 299792 1002319
rect 304720 1002307 304726 1002319
rect 299786 1002279 304726 1002307
rect 299786 1002267 299792 1002279
rect 304720 1002267 304726 1002279
rect 304778 1002267 304784 1002319
rect 446320 1002267 446326 1002319
rect 446378 1002307 446384 1002319
rect 446378 1002279 446462 1002307
rect 446378 1002267 446384 1002279
rect 446434 1002233 446462 1002279
rect 489520 1002267 489526 1002319
rect 489578 1002307 489584 1002319
rect 519184 1002307 519190 1002319
rect 489578 1002279 519190 1002307
rect 489578 1002267 489584 1002279
rect 519184 1002267 519190 1002279
rect 519242 1002267 519248 1002319
rect 561520 1002267 561526 1002319
rect 561578 1002307 561584 1002319
rect 564688 1002307 564694 1002319
rect 561578 1002279 564694 1002307
rect 561578 1002267 561584 1002279
rect 564688 1002267 564694 1002279
rect 564746 1002267 564752 1002319
rect 460912 1002233 460918 1002245
rect 446434 1002205 460918 1002233
rect 460912 1002193 460918 1002205
rect 460970 1002193 460976 1002245
rect 466576 1002193 466582 1002245
rect 466634 1002233 466640 1002245
rect 471952 1002233 471958 1002245
rect 466634 1002205 471958 1002233
rect 466634 1002193 466640 1002205
rect 471952 1002193 471958 1002205
rect 472010 1002193 472016 1002245
rect 573040 1002193 573046 1002245
rect 573098 1002233 573104 1002245
rect 573904 1002233 573910 1002245
rect 573098 1002205 573910 1002233
rect 573098 1002193 573104 1002205
rect 573904 1002193 573910 1002205
rect 573962 1002193 573968 1002245
rect 572944 1001823 572950 1001875
rect 573002 1001863 573008 1001875
rect 573232 1001863 573238 1001875
rect 573002 1001835 573238 1001863
rect 573002 1001823 573008 1001835
rect 573232 1001823 573238 1001835
rect 573290 1001823 573296 1001875
rect 513520 1001601 513526 1001653
rect 513578 1001641 513584 1001653
rect 518320 1001641 518326 1001653
rect 513578 1001613 518326 1001641
rect 513578 1001601 513584 1001613
rect 518320 1001601 518326 1001613
rect 518378 1001601 518384 1001653
rect 515440 1001527 515446 1001579
rect 515498 1001567 515504 1001579
rect 516880 1001567 516886 1001579
rect 515498 1001539 516886 1001567
rect 515498 1001527 515504 1001539
rect 516880 1001527 516886 1001539
rect 516938 1001527 516944 1001579
rect 566128 1001453 566134 1001505
rect 566186 1001493 566192 1001505
rect 567760 1001493 567766 1001505
rect 566186 1001465 567766 1001493
rect 566186 1001453 566192 1001465
rect 567760 1001453 567766 1001465
rect 567818 1001453 567824 1001505
rect 572848 1001305 572854 1001357
rect 572906 1001345 572912 1001357
rect 574480 1001345 574486 1001357
rect 572906 1001317 574486 1001345
rect 572906 1001305 572912 1001317
rect 574480 1001305 574486 1001317
rect 574538 1001305 574544 1001357
rect 511024 1001231 511030 1001283
rect 511082 1001271 511088 1001283
rect 516688 1001271 516694 1001283
rect 511082 1001243 516694 1001271
rect 511082 1001231 511088 1001243
rect 516688 1001231 516694 1001243
rect 516746 1001231 516752 1001283
rect 434128 1001083 434134 1001135
rect 434186 1001123 434192 1001135
rect 472624 1001123 472630 1001135
rect 434186 1001095 472630 1001123
rect 434186 1001083 434192 1001095
rect 472624 1001083 472630 1001095
rect 472682 1001083 472688 1001135
rect 463696 1001009 463702 1001061
rect 463754 1001049 463760 1001061
rect 471760 1001049 471766 1001061
rect 463754 1001021 471766 1001049
rect 463754 1001009 463760 1001021
rect 471760 1001009 471766 1001021
rect 471818 1001009 471824 1001061
rect 509392 1001009 509398 1001061
rect 509450 1001049 509456 1001061
rect 516688 1001049 516694 1001061
rect 509450 1001021 516694 1001049
rect 509450 1001009 509456 1001021
rect 516688 1001009 516694 1001021
rect 516746 1001009 516752 1001061
rect 432496 1000935 432502 1000987
rect 432554 1000975 432560 1000987
rect 472624 1000975 472630 1000987
rect 432554 1000947 472630 1000975
rect 432554 1000935 432560 1000947
rect 472624 1000935 472630 1000947
rect 472682 1000935 472688 1000987
rect 428944 1000861 428950 1000913
rect 429002 1000901 429008 1000913
rect 472528 1000901 472534 1000913
rect 429002 1000873 472534 1000901
rect 429002 1000861 429008 1000873
rect 472528 1000861 472534 1000873
rect 472586 1000861 472592 1000913
rect 143824 1000787 143830 1000839
rect 143882 1000827 143888 1000839
rect 160240 1000827 160246 1000839
rect 143882 1000799 160246 1000827
rect 143882 1000787 143888 1000799
rect 160240 1000787 160246 1000799
rect 160298 1000787 160304 1000839
rect 195088 1000787 195094 1000839
rect 195146 1000827 195152 1000839
rect 208432 1000827 208438 1000839
rect 195146 1000799 208438 1000827
rect 195146 1000787 195152 1000799
rect 208432 1000787 208438 1000799
rect 208490 1000787 208496 1000839
rect 361552 1000787 361558 1000839
rect 361610 1000827 361616 1000839
rect 383440 1000827 383446 1000839
rect 361610 1000799 383446 1000827
rect 361610 1000787 361616 1000799
rect 383440 1000787 383446 1000799
rect 383498 1000787 383504 1000839
rect 427312 1000787 427318 1000839
rect 427370 1000827 427376 1000839
rect 472336 1000827 472342 1000839
rect 427370 1000799 472342 1000827
rect 427370 1000787 427376 1000799
rect 472336 1000787 472342 1000799
rect 472394 1000787 472400 1000839
rect 507760 1000713 507766 1000765
rect 507818 1000753 507824 1000765
rect 516688 1000753 516694 1000765
rect 507818 1000725 516694 1000753
rect 507818 1000713 507824 1000725
rect 516688 1000713 516694 1000725
rect 516746 1000713 516752 1000765
rect 453328 1000417 453334 1000469
rect 453386 1000457 453392 1000469
rect 463696 1000457 463702 1000469
rect 453386 1000429 463702 1000457
rect 453386 1000417 453392 1000429
rect 463696 1000417 463702 1000429
rect 463754 1000417 463760 1000469
rect 460816 1000343 460822 1000395
rect 460874 1000383 460880 1000395
rect 472144 1000383 472150 1000395
rect 460874 1000355 472150 1000383
rect 460874 1000343 460880 1000355
rect 472144 1000343 472150 1000355
rect 472202 1000343 472208 1000395
rect 380464 999899 380470 999951
rect 380522 999939 380528 999951
rect 383248 999939 383254 999951
rect 380522 999911 383254 999939
rect 380522 999899 380528 999911
rect 383248 999899 383254 999911
rect 383306 999899 383312 999951
rect 610576 999677 610582 999729
rect 610634 999717 610640 999729
rect 625744 999717 625750 999729
rect 610634 999689 625750 999717
rect 610634 999677 610640 999689
rect 625744 999677 625750 999689
rect 625802 999677 625808 999729
rect 93040 999603 93046 999655
rect 93098 999643 93104 999655
rect 127408 999643 127414 999655
rect 93098 999615 127414 999643
rect 93098 999603 93104 999615
rect 127408 999603 127414 999615
rect 127466 999603 127472 999655
rect 298096 999603 298102 999655
rect 298154 999643 298160 999655
rect 298480 999643 298486 999655
rect 298154 999615 298486 999643
rect 298154 999603 298160 999615
rect 298480 999603 298486 999615
rect 298538 999603 298544 999655
rect 377296 999603 377302 999655
rect 377354 999643 377360 999655
rect 383152 999643 383158 999655
rect 377354 999615 383158 999643
rect 377354 999603 377360 999615
rect 383152 999603 383158 999615
rect 383210 999603 383216 999655
rect 613456 999603 613462 999655
rect 613514 999643 613520 999655
rect 625456 999643 625462 999655
rect 613514 999615 625462 999643
rect 613514 999603 613520 999615
rect 625456 999603 625462 999615
rect 625514 999603 625520 999655
rect 144208 999529 144214 999581
rect 144266 999569 144272 999581
rect 158608 999569 158614 999581
rect 144266 999541 158614 999569
rect 144266 999529 144272 999541
rect 158608 999529 158614 999541
rect 158666 999529 158672 999581
rect 246640 999529 246646 999581
rect 246698 999569 246704 999581
rect 262096 999569 262102 999581
rect 246698 999541 262102 999569
rect 246698 999529 246704 999541
rect 262096 999529 262102 999541
rect 262154 999529 262160 999581
rect 380176 999529 380182 999581
rect 380234 999569 380240 999581
rect 383344 999569 383350 999581
rect 380234 999541 383350 999569
rect 380234 999529 380240 999541
rect 383344 999529 383350 999541
rect 383402 999529 383408 999581
rect 497584 999529 497590 999581
rect 497642 999569 497648 999581
rect 516688 999569 516694 999581
rect 497642 999541 516694 999569
rect 497642 999529 497648 999541
rect 516688 999529 516694 999541
rect 516746 999529 516752 999581
rect 604720 999529 604726 999581
rect 604778 999569 604784 999581
rect 625552 999569 625558 999581
rect 604778 999541 625558 999569
rect 604778 999529 604784 999541
rect 625552 999529 625558 999541
rect 625610 999529 625616 999581
rect 144112 999455 144118 999507
rect 144170 999495 144176 999507
rect 155152 999495 155158 999507
rect 144170 999467 155158 999495
rect 144170 999455 144176 999467
rect 155152 999455 155158 999467
rect 155210 999455 155216 999507
rect 250480 999455 250486 999507
rect 250538 999495 250544 999507
rect 263056 999495 263062 999507
rect 250538 999467 263062 999495
rect 250538 999455 250544 999467
rect 263056 999455 263062 999467
rect 263114 999455 263120 999507
rect 298096 999455 298102 999507
rect 298154 999495 298160 999507
rect 311152 999495 311158 999507
rect 298154 999467 311158 999495
rect 298154 999455 298160 999467
rect 311152 999455 311158 999467
rect 311210 999455 311216 999507
rect 380368 999455 380374 999507
rect 380426 999495 380432 999507
rect 382960 999495 382966 999507
rect 380426 999467 382966 999495
rect 380426 999455 380432 999467
rect 382960 999455 382966 999467
rect 383018 999455 383024 999507
rect 506320 999455 506326 999507
rect 506378 999495 506384 999507
rect 516784 999495 516790 999507
rect 506378 999467 516790 999495
rect 506378 999455 506384 999467
rect 516784 999455 516790 999467
rect 516842 999455 516848 999507
rect 564688 999455 564694 999507
rect 564746 999495 564752 999507
rect 564746 999467 567518 999495
rect 564746 999455 564752 999467
rect 143728 999381 143734 999433
rect 143786 999421 143792 999433
rect 156880 999421 156886 999433
rect 143786 999393 156886 999421
rect 143786 999381 143792 999393
rect 156880 999381 156886 999393
rect 156938 999381 156944 999433
rect 246544 999381 246550 999433
rect 246602 999421 246608 999433
rect 259600 999421 259606 999433
rect 246602 999393 259606 999421
rect 246602 999381 246608 999393
rect 259600 999381 259606 999393
rect 259658 999381 259664 999433
rect 299440 999381 299446 999433
rect 299498 999421 299504 999433
rect 310288 999421 310294 999433
rect 299498 999393 310294 999421
rect 299498 999381 299504 999393
rect 310288 999381 310294 999393
rect 310346 999381 310352 999433
rect 380560 999381 380566 999433
rect 380618 999421 380624 999433
rect 383536 999421 383542 999433
rect 380618 999393 383542 999421
rect 380618 999381 380624 999393
rect 383536 999381 383542 999393
rect 383594 999381 383600 999433
rect 399952 999381 399958 999433
rect 400010 999421 400016 999433
rect 400010 999393 459326 999421
rect 400010 999381 400016 999393
rect 459298 999347 459326 999393
rect 540304 999381 540310 999433
rect 540362 999421 540368 999433
rect 561520 999421 561526 999433
rect 540362 999393 561526 999421
rect 540362 999381 540368 999393
rect 561520 999381 561526 999393
rect 561578 999381 561584 999433
rect 566320 999381 566326 999433
rect 566378 999421 566384 999433
rect 567490 999421 567518 999467
rect 593296 999455 593302 999507
rect 593354 999495 593360 999507
rect 625840 999495 625846 999507
rect 593354 999467 625846 999495
rect 593354 999455 593360 999467
rect 625840 999455 625846 999467
rect 625898 999455 625904 999507
rect 566378 999393 567422 999421
rect 567490 999393 570590 999421
rect 566378 999381 566384 999393
rect 460816 999347 460822 999359
rect 459298 999319 460822 999347
rect 460816 999307 460822 999319
rect 460874 999307 460880 999359
rect 502384 999307 502390 999359
rect 502442 999347 502448 999359
rect 516688 999347 516694 999359
rect 502442 999319 516694 999347
rect 502442 999307 502448 999319
rect 516688 999307 516694 999319
rect 516746 999307 516752 999359
rect 516880 999307 516886 999359
rect 516938 999347 516944 999359
rect 520912 999347 520918 999359
rect 516938 999319 520918 999347
rect 516938 999307 516944 999319
rect 520912 999307 520918 999319
rect 520970 999307 520976 999359
rect 567394 999347 567422 999393
rect 570448 999347 570454 999359
rect 567394 999319 570454 999347
rect 570448 999307 570454 999319
rect 570506 999307 570512 999359
rect 570562 999347 570590 999393
rect 590512 999381 590518 999433
rect 590570 999421 590576 999433
rect 625648 999421 625654 999433
rect 590570 999393 625654 999421
rect 590570 999381 590576 999393
rect 625648 999381 625654 999393
rect 625706 999381 625712 999433
rect 570640 999347 570646 999359
rect 570562 999319 570646 999347
rect 570640 999307 570646 999319
rect 570698 999307 570704 999359
rect 461008 999233 461014 999285
rect 461066 999273 461072 999285
rect 471568 999273 471574 999285
rect 461066 999245 471574 999273
rect 461066 999233 461072 999245
rect 471568 999233 471574 999245
rect 471626 999233 471632 999285
rect 515536 999233 515542 999285
rect 515594 999273 515600 999285
rect 523408 999273 523414 999285
rect 515594 999245 523414 999273
rect 515594 999233 515600 999245
rect 523408 999233 523414 999245
rect 523466 999233 523472 999285
rect 356272 998049 356278 998101
rect 356330 998089 356336 998101
rect 368752 998089 368758 998101
rect 356330 998061 368758 998089
rect 356330 998049 356336 998061
rect 368752 998049 368758 998061
rect 368810 998049 368816 998101
rect 357040 997975 357046 998027
rect 357098 998015 357104 998027
rect 368656 998015 368662 998027
rect 357098 997987 368662 998015
rect 357098 997975 357104 997987
rect 368656 997975 368662 997987
rect 368714 997975 368720 998027
rect 555280 997975 555286 998027
rect 555338 998015 555344 998027
rect 570736 998015 570742 998027
rect 555338 997987 570742 998015
rect 555338 997975 555344 997987
rect 570736 997975 570742 997987
rect 570794 997975 570800 998027
rect 320944 997901 320950 997953
rect 321002 997941 321008 997953
rect 367888 997941 367894 997953
rect 321002 997913 367894 997941
rect 321002 997901 321008 997913
rect 367888 997901 367894 997913
rect 367946 997941 367952 997953
rect 381712 997941 381718 997953
rect 367946 997913 381718 997941
rect 367946 997901 367952 997913
rect 381712 997901 381718 997913
rect 381770 997901 381776 997953
rect 561520 997901 561526 997953
rect 561578 997941 561584 997953
rect 616336 997941 616342 997953
rect 561578 997913 616342 997941
rect 561578 997901 561584 997913
rect 616336 997901 616342 997913
rect 616394 997901 616400 997953
rect 331120 997827 331126 997879
rect 331178 997867 331184 997879
rect 369040 997867 369046 997879
rect 331178 997839 369046 997867
rect 331178 997827 331184 997839
rect 369040 997827 369046 997839
rect 369098 997827 369104 997879
rect 557296 997827 557302 997879
rect 557354 997867 557360 997879
rect 593296 997867 593302 997879
rect 557354 997839 593302 997867
rect 557354 997827 557360 997839
rect 593296 997827 593302 997839
rect 593354 997827 593360 997879
rect 574000 997753 574006 997805
rect 574058 997793 574064 997805
rect 590512 997793 590518 997805
rect 574058 997765 590518 997793
rect 574058 997753 574064 997765
rect 590512 997753 590518 997765
rect 590570 997753 590576 997805
rect 567760 997679 567766 997731
rect 567818 997719 567824 997731
rect 604720 997719 604726 997731
rect 567818 997691 604726 997719
rect 567818 997679 567824 997691
rect 604720 997679 604726 997691
rect 604778 997679 604784 997731
rect 573904 997605 573910 997657
rect 573962 997645 573968 997657
rect 613456 997645 613462 997657
rect 573962 997617 613462 997645
rect 573962 997605 573968 997617
rect 613456 997605 613462 997617
rect 613514 997605 613520 997657
rect 564784 997531 564790 997583
rect 564842 997571 564848 997583
rect 610576 997571 610582 997583
rect 564842 997543 610582 997571
rect 564842 997531 564848 997543
rect 610576 997531 610582 997543
rect 610634 997531 610640 997583
rect 460912 996939 460918 996991
rect 460970 996979 460976 996991
rect 472240 996979 472246 996991
rect 460970 996951 472246 996979
rect 460970 996939 460976 996951
rect 472240 996939 472246 996951
rect 472298 996939 472304 996991
rect 377392 996865 377398 996917
rect 377450 996905 377456 996917
rect 382864 996905 382870 996917
rect 377450 996877 382870 996905
rect 377450 996865 377456 996877
rect 382864 996865 382870 996877
rect 382922 996865 382928 996917
rect 201616 996643 201622 996695
rect 201674 996683 201680 996695
rect 201674 996655 205790 996683
rect 201674 996643 201680 996655
rect 195760 996495 195766 996547
rect 195818 996535 195824 996547
rect 205648 996535 205654 996547
rect 195818 996507 205654 996535
rect 195818 996495 195824 996507
rect 205648 996495 205654 996507
rect 205706 996495 205712 996547
rect 205762 996535 205790 996655
rect 377488 996569 377494 996621
rect 377546 996609 377552 996621
rect 382768 996609 382774 996621
rect 377546 996581 382774 996609
rect 377546 996569 377552 996581
rect 382768 996569 382774 996581
rect 382826 996569 382832 996621
rect 510256 996569 510262 996621
rect 510314 996609 510320 996621
rect 521008 996609 521014 996621
rect 510314 996581 521014 996609
rect 510314 996569 510320 996581
rect 521008 996569 521014 996581
rect 521066 996569 521072 996621
rect 211696 996535 211702 996547
rect 205762 996507 211702 996535
rect 211696 996495 211702 996507
rect 211754 996495 211760 996547
rect 298192 996495 298198 996547
rect 298250 996535 298256 996547
rect 374512 996535 374518 996547
rect 298250 996507 374518 996535
rect 298250 996495 298256 996507
rect 374512 996495 374518 996507
rect 374570 996495 374576 996547
rect 508624 996495 508630 996547
rect 508682 996535 508688 996547
rect 521200 996535 521206 996547
rect 508682 996507 521206 996535
rect 508682 996495 508688 996507
rect 521200 996495 521206 996507
rect 521258 996495 521264 996547
rect 320176 996421 320182 996473
rect 320234 996461 320240 996473
rect 367120 996461 367126 996473
rect 320234 996433 367126 996461
rect 320234 996421 320240 996433
rect 367120 996421 367126 996433
rect 367178 996421 367184 996473
rect 144304 996273 144310 996325
rect 144362 996313 144368 996325
rect 162256 996313 162262 996325
rect 144362 996285 162262 996313
rect 144362 996273 144368 996285
rect 162256 996273 162262 996285
rect 162314 996313 162320 996325
rect 162314 996285 177182 996313
rect 162314 996273 162320 996285
rect 115312 996125 115318 996177
rect 115370 996165 115376 996177
rect 126736 996165 126742 996177
rect 115370 996137 126742 996165
rect 115370 996125 115376 996137
rect 126736 996125 126742 996137
rect 126794 996125 126800 996177
rect 115216 996051 115222 996103
rect 115274 996091 115280 996103
rect 163120 996091 163126 996103
rect 115274 996063 163126 996091
rect 115274 996051 115280 996063
rect 163120 996051 163126 996063
rect 163178 996091 163184 996103
rect 177040 996091 177046 996103
rect 163178 996063 177046 996091
rect 163178 996051 163184 996063
rect 177040 996051 177046 996063
rect 177098 996051 177104 996103
rect 177154 996091 177182 996285
rect 511120 996199 511126 996251
rect 511178 996239 511184 996251
rect 511178 996211 513566 996239
rect 511178 996199 511184 996211
rect 198544 996125 198550 996177
rect 198602 996165 198608 996177
rect 203632 996165 203638 996177
rect 198602 996137 203638 996165
rect 198602 996125 198608 996137
rect 203632 996125 203638 996137
rect 203690 996125 203696 996177
rect 214096 996125 214102 996177
rect 214154 996165 214160 996177
rect 214154 996137 258302 996165
rect 214154 996125 214160 996137
rect 213328 996091 213334 996103
rect 177154 996063 213334 996091
rect 213328 996051 213334 996063
rect 213386 996091 213392 996103
rect 258274 996091 258302 996137
rect 266800 996125 266806 996177
rect 266858 996165 266864 996177
rect 318640 996165 318646 996177
rect 266858 996137 318646 996165
rect 266858 996125 266864 996137
rect 318640 996125 318646 996137
rect 318698 996125 318704 996177
rect 371536 996125 371542 996177
rect 371594 996165 371600 996177
rect 436336 996165 436342 996177
rect 371594 996137 436342 996165
rect 371594 996125 371600 996137
rect 436336 996125 436342 996137
rect 436394 996125 436400 996177
rect 436432 996125 436438 996177
rect 436490 996165 436496 996177
rect 513424 996165 513430 996177
rect 436490 996137 513430 996165
rect 436490 996125 436496 996137
rect 513424 996125 513430 996137
rect 513482 996125 513488 996177
rect 513538 996165 513566 996211
rect 562768 996165 562774 996177
rect 513538 996137 562774 996165
rect 562768 996125 562774 996137
rect 562826 996125 562832 996177
rect 265936 996091 265942 996103
rect 213386 996063 226046 996091
rect 258274 996063 265942 996091
rect 213386 996051 213392 996063
rect 120976 995977 120982 996029
rect 121034 996017 121040 996029
rect 164560 996017 164566 996029
rect 121034 995989 164566 996017
rect 121034 995977 121040 995989
rect 164560 995977 164566 995989
rect 164618 995977 164624 996029
rect 198640 995977 198646 996029
rect 198698 996017 198704 996029
rect 202960 996017 202966 996029
rect 198698 995989 202966 996017
rect 198698 995977 198704 995989
rect 202960 995977 202966 995989
rect 203018 995977 203024 996029
rect 213040 995977 213046 996029
rect 213098 996017 213104 996029
rect 216880 996017 216886 996029
rect 213098 995989 216886 996017
rect 213098 995977 213104 995989
rect 216880 995977 216886 995989
rect 216938 995977 216944 996029
rect 226018 996017 226046 996063
rect 265936 996051 265942 996063
rect 265994 996091 266000 996103
rect 317104 996091 317110 996103
rect 265994 996063 317110 996091
rect 265994 996051 266000 996063
rect 317104 996051 317110 996063
rect 317162 996091 317168 996103
rect 320944 996091 320950 996103
rect 317162 996063 320950 996091
rect 317162 996051 317168 996063
rect 320944 996051 320950 996063
rect 321002 996051 321008 996103
rect 381712 996051 381718 996103
rect 381770 996091 381776 996103
rect 440656 996091 440662 996103
rect 381770 996063 440662 996091
rect 381770 996051 381776 996063
rect 440656 996051 440662 996063
rect 440714 996051 440720 996103
rect 563536 996091 563542 996103
rect 511906 996063 563542 996091
rect 265072 996017 265078 996029
rect 226018 995989 265078 996017
rect 265072 995977 265078 995989
rect 265130 996017 265136 996029
rect 316336 996017 316342 996029
rect 265130 995989 316342 996017
rect 265130 995977 265136 995989
rect 316336 995977 316342 995989
rect 316394 996017 316400 996029
rect 320176 996017 320182 996029
rect 316394 995989 320182 996017
rect 316394 995977 316400 995989
rect 320176 995977 320182 995989
rect 320234 995977 320240 996029
rect 367120 995977 367126 996029
rect 367178 996017 367184 996029
rect 434128 996017 434134 996029
rect 367178 995989 434134 996017
rect 367178 995977 367184 995989
rect 434128 995977 434134 995989
rect 434186 996017 434192 996029
rect 439408 996017 439414 996029
rect 434186 995989 439414 996017
rect 434186 995977 434192 995989
rect 439408 995977 439414 995989
rect 439466 995977 439472 996029
rect 470896 995977 470902 996029
rect 470954 996017 470960 996029
rect 470954 995989 476606 996017
rect 470954 995977 470960 995989
rect 100624 995943 100630 995955
rect 82306 995915 100630 995943
rect 82306 995807 82334 995915
rect 100624 995903 100630 995915
rect 100682 995903 100688 995955
rect 144112 995943 144118 995955
rect 132418 995915 144118 995943
rect 94672 995829 94678 995881
rect 94730 995869 94736 995881
rect 99952 995869 99958 995881
rect 94730 995841 99958 995869
rect 94730 995829 94736 995841
rect 99952 995829 99958 995841
rect 100010 995829 100016 995881
rect 113488 995869 113494 995881
rect 106690 995841 113494 995869
rect 82288 995755 82294 995807
rect 82346 995755 82352 995807
rect 87856 995755 87862 995807
rect 87914 995795 87920 995807
rect 102160 995795 102166 995807
rect 87914 995767 102166 995795
rect 87914 995755 87920 995767
rect 102160 995755 102166 995767
rect 102218 995755 102224 995807
rect 106480 995755 106486 995807
rect 106538 995795 106544 995807
rect 106690 995795 106718 995841
rect 113488 995829 113494 995841
rect 113546 995829 113552 995881
rect 132418 995807 132446 995915
rect 144112 995903 144118 995915
rect 144170 995903 144176 995955
rect 152080 995943 152086 995955
rect 144226 995915 152086 995943
rect 144226 995869 144254 995915
rect 152080 995903 152086 995915
rect 152138 995903 152144 995955
rect 164176 995903 164182 995955
rect 164234 995943 164240 995955
rect 215632 995943 215638 995955
rect 164234 995915 215638 995943
rect 164234 995903 164240 995915
rect 215632 995903 215638 995915
rect 215690 995903 215696 995955
rect 218896 995903 218902 995955
rect 218954 995943 218960 995955
rect 266992 995943 266998 995955
rect 218954 995915 266998 995943
rect 218954 995903 218960 995915
rect 266992 995903 266998 995915
rect 267050 995903 267056 995955
rect 370576 995903 370582 995955
rect 370634 995943 370640 995955
rect 374608 995943 374614 995955
rect 370634 995915 374614 995943
rect 370634 995903 370640 995915
rect 374608 995903 374614 995915
rect 374666 995903 374672 995955
rect 383344 995903 383350 995955
rect 383402 995943 383408 995955
rect 383402 995915 389246 995943
rect 383402 995903 383408 995915
rect 133666 995841 144254 995869
rect 133666 995807 133694 995841
rect 177040 995829 177046 995881
rect 177098 995869 177104 995881
rect 214096 995869 214102 995881
rect 177098 995841 214102 995869
rect 177098 995829 177104 995841
rect 214096 995829 214102 995841
rect 214154 995829 214160 995881
rect 246736 995869 246742 995881
rect 240898 995841 246742 995869
rect 240898 995807 240926 995841
rect 246736 995829 246742 995841
rect 246794 995829 246800 995881
rect 253360 995829 253366 995881
rect 253418 995869 253424 995881
rect 259120 995869 259126 995881
rect 253418 995841 259126 995869
rect 253418 995829 253424 995841
rect 259120 995829 259126 995841
rect 259178 995829 259184 995881
rect 299440 995869 299446 995881
rect 283714 995841 299446 995869
rect 283714 995807 283742 995841
rect 299440 995829 299446 995841
rect 299498 995829 299504 995881
rect 382960 995829 382966 995881
rect 383018 995869 383024 995881
rect 383018 995841 386078 995869
rect 383018 995829 383024 995841
rect 386050 995807 386078 995841
rect 106538 995767 106718 995795
rect 106538 995755 106544 995767
rect 113296 995755 113302 995807
rect 113354 995795 113360 995807
rect 118096 995795 118102 995807
rect 113354 995767 118102 995795
rect 113354 995755 113360 995767
rect 118096 995755 118102 995767
rect 118154 995755 118160 995807
rect 132400 995755 132406 995807
rect 132458 995755 132464 995807
rect 133648 995755 133654 995807
rect 133706 995755 133712 995807
rect 142960 995755 142966 995807
rect 143018 995795 143024 995807
rect 143728 995795 143734 995807
rect 143018 995767 143734 995795
rect 143018 995755 143024 995767
rect 143728 995755 143734 995767
rect 143786 995755 143792 995807
rect 164080 995755 164086 995807
rect 164138 995795 164144 995807
rect 165616 995795 165622 995807
rect 164138 995767 165622 995795
rect 164138 995755 164144 995767
rect 165616 995755 165622 995767
rect 165674 995755 165680 995807
rect 178480 995755 178486 995807
rect 178538 995795 178544 995807
rect 185200 995795 185206 995807
rect 178538 995767 185206 995795
rect 178538 995755 178544 995767
rect 185200 995755 185206 995767
rect 185258 995755 185264 995807
rect 190576 995755 190582 995807
rect 190634 995795 190640 995807
rect 204976 995795 204982 995807
rect 190634 995767 204982 995795
rect 190634 995755 190640 995767
rect 204976 995755 204982 995767
rect 205034 995755 205040 995807
rect 240880 995755 240886 995807
rect 240938 995755 240944 995807
rect 245680 995755 245686 995807
rect 245738 995795 245744 995807
rect 246544 995795 246550 995807
rect 245738 995767 246550 995795
rect 245738 995755 245744 995767
rect 246544 995755 246550 995767
rect 246602 995755 246608 995807
rect 283696 995755 283702 995807
rect 283754 995755 283760 995807
rect 297328 995755 297334 995807
rect 297386 995795 297392 995807
rect 298096 995795 298102 995807
rect 297386 995767 298102 995795
rect 297386 995755 297392 995767
rect 298096 995755 298102 995767
rect 298154 995755 298160 995807
rect 371344 995755 371350 995807
rect 371402 995795 371408 995807
rect 374416 995795 374422 995807
rect 371402 995767 374422 995795
rect 371402 995755 371408 995767
rect 374416 995755 374422 995767
rect 374474 995755 374480 995807
rect 383632 995755 383638 995807
rect 383690 995795 383696 995807
rect 384400 995795 384406 995807
rect 383690 995767 384406 995795
rect 383690 995755 383696 995767
rect 384400 995755 384406 995767
rect 384458 995755 384464 995807
rect 386032 995755 386038 995807
rect 386090 995755 386096 995807
rect 389218 995795 389246 995915
rect 471856 995903 471862 995955
rect 471914 995943 471920 995955
rect 471914 995915 474398 995943
rect 471914 995903 471920 995915
rect 389392 995795 389398 995807
rect 389218 995767 389398 995795
rect 389392 995755 389398 995767
rect 389450 995755 389456 995807
rect 396592 995755 396598 995807
rect 396650 995795 396656 995807
rect 399952 995795 399958 995807
rect 396650 995767 399958 995795
rect 396650 995755 396656 995767
rect 399952 995755 399958 995767
rect 400010 995755 400016 995807
rect 438736 995755 438742 995807
rect 438794 995795 438800 995807
rect 444880 995795 444886 995807
rect 438794 995767 444886 995795
rect 438794 995755 438800 995767
rect 444880 995755 444886 995767
rect 444938 995755 444944 995807
rect 472624 995755 472630 995807
rect 472682 995795 472688 995807
rect 473296 995795 473302 995807
rect 472682 995767 473302 995795
rect 472682 995755 472688 995767
rect 473296 995755 473302 995767
rect 473354 995755 473360 995807
rect 91504 995681 91510 995733
rect 91562 995721 91568 995733
rect 105328 995721 105334 995733
rect 91562 995693 105334 995721
rect 91562 995681 91568 995693
rect 105328 995681 105334 995693
rect 105386 995681 105392 995733
rect 127408 995681 127414 995733
rect 127466 995721 127472 995733
rect 134320 995721 134326 995733
rect 127466 995693 134326 995721
rect 127466 995681 127472 995693
rect 134320 995681 134326 995693
rect 134378 995681 134384 995733
rect 141040 995681 141046 995733
rect 141098 995721 141104 995733
rect 143824 995721 143830 995733
rect 141098 995693 143830 995721
rect 141098 995681 141104 995693
rect 143824 995681 143830 995693
rect 143882 995681 143888 995733
rect 163984 995681 163990 995733
rect 164042 995721 164048 995733
rect 166288 995721 166294 995733
rect 164042 995693 166294 995721
rect 164042 995681 164048 995693
rect 166288 995681 166294 995693
rect 166346 995681 166352 995733
rect 194416 995681 194422 995733
rect 194474 995721 194480 995733
rect 195088 995721 195094 995733
rect 194474 995693 195094 995721
rect 194474 995681 194480 995693
rect 195088 995681 195094 995693
rect 195146 995681 195152 995733
rect 198640 995681 198646 995733
rect 198698 995721 198704 995733
rect 206608 995721 206614 995733
rect 198698 995693 206614 995721
rect 198698 995681 198704 995693
rect 206608 995681 206614 995693
rect 206666 995681 206672 995733
rect 243184 995681 243190 995733
rect 243242 995721 243248 995733
rect 246640 995721 246646 995733
rect 243242 995693 246646 995721
rect 243242 995681 243248 995693
rect 246640 995681 246646 995693
rect 246698 995681 246704 995733
rect 294832 995681 294838 995733
rect 294890 995721 294896 995733
rect 298192 995721 298198 995733
rect 294890 995693 298198 995721
rect 294890 995681 294896 995693
rect 298192 995681 298198 995693
rect 298250 995681 298256 995733
rect 383536 995681 383542 995733
rect 383594 995721 383600 995733
rect 387472 995721 387478 995733
rect 383594 995693 387478 995721
rect 383594 995681 383600 995693
rect 387472 995681 387478 995693
rect 387530 995681 387536 995733
rect 472528 995681 472534 995733
rect 472586 995721 472592 995733
rect 474064 995721 474070 995733
rect 472586 995693 474070 995721
rect 472586 995681 472592 995693
rect 474064 995681 474070 995693
rect 474122 995681 474128 995733
rect 474370 995721 474398 995915
rect 476578 995795 476606 995989
rect 511120 995943 511126 995955
rect 478594 995915 511126 995943
rect 478594 995795 478622 995915
rect 511120 995903 511126 995915
rect 511178 995903 511184 995955
rect 511906 995881 511934 996063
rect 563536 996051 563542 996063
rect 563594 996051 563600 996103
rect 513424 995977 513430 996029
rect 513482 996017 513488 996029
rect 564784 996017 564790 996029
rect 513482 995989 564790 996017
rect 513482 995977 513488 995989
rect 564784 995977 564790 995989
rect 564842 995977 564848 996029
rect 521104 995903 521110 995955
rect 521162 995943 521168 995955
rect 521162 995915 529886 995943
rect 521162 995903 521168 995915
rect 511888 995869 511894 995881
rect 476578 995767 478622 995795
rect 478690 995841 511894 995869
rect 478690 995721 478718 995841
rect 511888 995829 511894 995841
rect 511946 995829 511952 995881
rect 523888 995829 523894 995881
rect 523946 995869 523952 995881
rect 523946 995841 529694 995869
rect 523946 995829 523952 995841
rect 524080 995755 524086 995807
rect 524138 995795 524144 995807
rect 528400 995795 528406 995807
rect 524138 995767 528406 995795
rect 524138 995755 524144 995767
rect 528400 995755 528406 995767
rect 528458 995755 528464 995807
rect 474370 995693 478718 995721
rect 523984 995681 523990 995733
rect 524042 995721 524048 995733
rect 528976 995721 528982 995733
rect 524042 995693 528982 995721
rect 524042 995681 524048 995693
rect 528976 995681 528982 995693
rect 529034 995681 529040 995733
rect 529666 995721 529694 995841
rect 529858 995807 529886 995915
rect 625456 995903 625462 995955
rect 625514 995943 625520 995955
rect 625514 995915 630686 995943
rect 625514 995903 625520 995915
rect 625648 995829 625654 995881
rect 625706 995869 625712 995881
rect 625706 995841 630206 995869
rect 625706 995829 625712 995841
rect 630178 995807 630206 995841
rect 529840 995755 529846 995807
rect 529898 995755 529904 995807
rect 537136 995755 537142 995807
rect 537194 995795 537200 995807
rect 540304 995795 540310 995807
rect 537194 995767 540310 995795
rect 537194 995755 537200 995767
rect 540304 995755 540310 995767
rect 540362 995755 540368 995807
rect 625840 995755 625846 995807
rect 625898 995795 625904 995807
rect 627088 995795 627094 995807
rect 625898 995767 627094 995795
rect 625898 995755 625904 995767
rect 627088 995755 627094 995767
rect 627146 995755 627152 995807
rect 630160 995755 630166 995807
rect 630218 995755 630224 995807
rect 630658 995795 630686 995915
rect 630928 995795 630934 995807
rect 630658 995767 630934 995795
rect 630928 995755 630934 995767
rect 630986 995755 630992 995807
rect 532816 995721 532822 995733
rect 529666 995693 532822 995721
rect 532816 995681 532822 995693
rect 532874 995681 532880 995733
rect 625744 995681 625750 995733
rect 625802 995721 625808 995733
rect 626512 995721 626518 995733
rect 625802 995693 626518 995721
rect 625802 995681 625808 995693
rect 626512 995681 626518 995693
rect 626570 995681 626576 995733
rect 139312 995607 139318 995659
rect 139370 995647 139376 995659
rect 143920 995647 143926 995659
rect 139370 995619 143926 995647
rect 139370 995607 139376 995619
rect 143920 995607 143926 995619
rect 143978 995607 143984 995659
rect 184336 995607 184342 995659
rect 184394 995647 184400 995659
rect 195760 995647 195766 995659
rect 184394 995619 195766 995647
rect 184394 995607 184400 995619
rect 195760 995607 195766 995619
rect 195818 995607 195824 995659
rect 201712 995607 201718 995659
rect 201770 995647 201776 995659
rect 206992 995647 206998 995659
rect 201770 995619 206998 995647
rect 201770 995607 201776 995619
rect 206992 995607 206998 995619
rect 207050 995607 207056 995659
rect 286768 995607 286774 995659
rect 286826 995647 286832 995659
rect 298384 995647 298390 995659
rect 286826 995619 298390 995647
rect 286826 995607 286832 995619
rect 298384 995607 298390 995619
rect 298442 995607 298448 995659
rect 383440 995607 383446 995659
rect 383498 995647 383504 995659
rect 384976 995647 384982 995659
rect 383498 995619 384982 995647
rect 383498 995607 383504 995619
rect 384976 995607 384982 995619
rect 385034 995607 385040 995659
rect 472336 995607 472342 995659
rect 472394 995647 472400 995659
rect 477712 995647 477718 995659
rect 472394 995619 477718 995647
rect 472394 995607 472400 995619
rect 477712 995607 477718 995619
rect 477770 995607 477776 995659
rect 479440 995607 479446 995659
rect 479498 995647 479504 995659
rect 479498 995619 483998 995647
rect 479498 995607 479504 995619
rect 137968 995533 137974 995585
rect 138026 995573 138032 995585
rect 144016 995573 144022 995585
rect 138026 995545 144022 995573
rect 138026 995533 138032 995545
rect 144016 995533 144022 995545
rect 144074 995533 144080 995585
rect 287536 995533 287542 995585
rect 287594 995573 287600 995585
rect 298480 995573 298486 995585
rect 287594 995545 298486 995573
rect 287594 995533 287600 995545
rect 298480 995533 298486 995545
rect 298538 995533 298544 995585
rect 383248 995533 383254 995585
rect 383306 995573 383312 995585
rect 391696 995573 391702 995585
rect 383306 995545 391702 995573
rect 383306 995533 383312 995545
rect 391696 995533 391702 995545
rect 391754 995533 391760 995585
rect 472720 995533 472726 995585
rect 472778 995573 472784 995585
rect 474640 995573 474646 995585
rect 472778 995545 474646 995573
rect 472778 995533 472784 995545
rect 474640 995533 474646 995545
rect 474698 995533 474704 995585
rect 81616 995459 81622 995511
rect 81674 995499 81680 995511
rect 102160 995499 102166 995511
rect 81674 995471 102166 995499
rect 81674 995459 81680 995471
rect 102160 995459 102166 995471
rect 102218 995459 102224 995511
rect 236464 995459 236470 995511
rect 236522 995499 236528 995511
rect 254800 995499 254806 995511
rect 236522 995471 254806 995499
rect 236522 995459 236528 995471
rect 254800 995459 254806 995471
rect 254858 995459 254864 995511
rect 287920 995459 287926 995511
rect 287978 995499 287984 995511
rect 299824 995499 299830 995511
rect 287978 995471 299830 995499
rect 287978 995459 287984 995471
rect 299824 995459 299830 995471
rect 299882 995459 299888 995511
rect 383152 995459 383158 995511
rect 383210 995499 383216 995511
rect 388048 995499 388054 995511
rect 383210 995471 388054 995499
rect 383210 995459 383216 995471
rect 388048 995459 388054 995471
rect 388106 995459 388112 995511
rect 471760 995459 471766 995511
rect 471818 995499 471824 995511
rect 483856 995499 483862 995511
rect 471818 995471 483862 995499
rect 471818 995459 471824 995471
rect 483856 995459 483862 995471
rect 483914 995459 483920 995511
rect 483970 995499 483998 995619
rect 523792 995607 523798 995659
rect 523850 995647 523856 995659
rect 525424 995647 525430 995659
rect 523850 995619 525430 995647
rect 523850 995607 523856 995619
rect 525424 995607 525430 995619
rect 525482 995607 525488 995659
rect 563536 995607 563542 995659
rect 563594 995647 563600 995659
rect 567376 995647 567382 995659
rect 563594 995619 567382 995647
rect 563594 995607 563600 995619
rect 567376 995607 567382 995619
rect 567434 995607 567440 995659
rect 625552 995607 625558 995659
rect 625610 995647 625616 995659
rect 629584 995647 629590 995659
rect 625610 995619 629590 995647
rect 625610 995607 625616 995619
rect 629584 995607 629590 995619
rect 629642 995607 629648 995659
rect 523696 995533 523702 995585
rect 523754 995573 523760 995585
rect 524752 995573 524758 995585
rect 523754 995545 524758 995573
rect 523754 995533 523760 995545
rect 524752 995533 524758 995545
rect 524810 995533 524816 995585
rect 562768 995533 562774 995585
rect 562826 995573 562832 995585
rect 567472 995573 567478 995585
rect 562826 995545 567478 995573
rect 562826 995533 562832 995545
rect 567472 995533 567478 995545
rect 567530 995533 567536 995585
rect 629200 995499 629206 995511
rect 483970 995471 629206 995499
rect 629200 995459 629206 995471
rect 629258 995459 629264 995511
rect 89776 995385 89782 995437
rect 89834 995425 89840 995437
rect 92080 995425 92086 995437
rect 89834 995397 92086 995425
rect 89834 995385 89840 995397
rect 92080 995385 92086 995397
rect 92138 995385 92144 995437
rect 126736 995385 126742 995437
rect 126794 995425 126800 995437
rect 144304 995425 144310 995437
rect 126794 995397 144310 995425
rect 126794 995385 126800 995397
rect 144304 995385 144310 995397
rect 144362 995385 144368 995437
rect 235792 995385 235798 995437
rect 235850 995425 235856 995437
rect 247600 995425 247606 995437
rect 235850 995397 247606 995425
rect 235850 995385 235856 995397
rect 247600 995385 247606 995397
rect 247658 995385 247664 995437
rect 284368 995385 284374 995437
rect 284426 995425 284432 995437
rect 299920 995425 299926 995437
rect 284426 995397 299926 995425
rect 284426 995385 284432 995397
rect 299920 995385 299926 995397
rect 299978 995385 299984 995437
rect 382864 995385 382870 995437
rect 382922 995425 382928 995437
rect 393040 995425 393046 995437
rect 382922 995397 393046 995425
rect 382922 995385 382928 995397
rect 393040 995385 393046 995397
rect 393098 995385 393104 995437
rect 460816 995385 460822 995437
rect 460874 995425 460880 995437
rect 630736 995425 630742 995437
rect 460874 995397 630742 995425
rect 460874 995385 460880 995397
rect 630736 995385 630742 995397
rect 630794 995385 630800 995437
rect 471568 995311 471574 995363
rect 471626 995351 471632 995363
rect 479440 995351 479446 995363
rect 471626 995323 479446 995351
rect 471626 995311 471632 995323
rect 479440 995311 479446 995323
rect 479498 995311 479504 995363
rect 518512 995311 518518 995363
rect 518570 995351 518576 995363
rect 533680 995351 533686 995363
rect 518570 995323 533686 995351
rect 518570 995311 518576 995323
rect 533680 995311 533686 995323
rect 533738 995311 533744 995363
rect 472144 995237 472150 995289
rect 472202 995277 472208 995289
rect 478624 995277 478630 995289
rect 472202 995249 478630 995277
rect 472202 995237 472208 995249
rect 478624 995237 478630 995249
rect 478682 995237 478688 995289
rect 521008 995237 521014 995289
rect 521066 995277 521072 995289
rect 537376 995277 537382 995289
rect 521066 995249 537382 995277
rect 521066 995237 521072 995249
rect 537376 995237 537382 995249
rect 537434 995237 537440 995289
rect 537520 995237 537526 995289
rect 537578 995277 537584 995289
rect 645136 995277 645142 995289
rect 537578 995249 645142 995277
rect 537578 995237 537584 995249
rect 645136 995237 645142 995249
rect 645194 995237 645200 995289
rect 69136 995163 69142 995215
rect 69194 995203 69200 995215
rect 343888 995203 343894 995215
rect 69194 995175 343894 995203
rect 69194 995163 69200 995175
rect 343888 995163 343894 995175
rect 343946 995163 343952 995215
rect 374512 995163 374518 995215
rect 374570 995203 374576 995215
rect 649936 995203 649942 995215
rect 374570 995175 649942 995203
rect 374570 995163 374576 995175
rect 649936 995163 649942 995175
rect 649994 995163 650000 995215
rect 262192 995089 262198 995141
rect 262250 995129 262256 995141
rect 645232 995129 645238 995141
rect 262250 995101 645238 995129
rect 262250 995089 262256 995101
rect 645232 995089 645238 995101
rect 645290 995089 645296 995141
rect 89008 995015 89014 995067
rect 89066 995055 89072 995067
rect 570256 995055 570262 995067
rect 89066 995027 570262 995055
rect 89066 995015 89072 995027
rect 570256 995015 570262 995027
rect 570314 995015 570320 995067
rect 616336 995015 616342 995067
rect 616394 995055 616400 995067
rect 640336 995055 640342 995067
rect 616394 995027 640342 995055
rect 616394 995015 616400 995027
rect 640336 995015 640342 995027
rect 640394 995015 640400 995067
rect 382768 994941 382774 994993
rect 382826 994981 382832 994993
rect 395152 994981 395158 994993
rect 382826 994953 395158 994981
rect 382826 994941 382832 994953
rect 395152 994941 395158 994953
rect 395210 994941 395216 994993
rect 463696 994941 463702 994993
rect 463754 994981 463760 994993
rect 482704 994981 482710 994993
rect 463754 994953 482710 994981
rect 463754 994941 463760 994953
rect 482704 994941 482710 994953
rect 482762 994941 482768 994993
rect 523408 994941 523414 994993
rect 523466 994981 523472 994993
rect 537520 994981 537526 994993
rect 523466 994953 537526 994981
rect 523466 994941 523472 994953
rect 537520 994941 537526 994953
rect 537578 994941 537584 994993
rect 471664 994867 471670 994919
rect 471722 994907 471728 994919
rect 481648 994907 481654 994919
rect 471722 994879 481654 994907
rect 471722 994867 471728 994879
rect 481648 994867 481654 994879
rect 481706 994867 481712 994919
rect 519184 994867 519190 994919
rect 519242 994907 519248 994919
rect 530320 994907 530326 994919
rect 519242 994879 530326 994907
rect 519242 994867 519248 994879
rect 530320 994867 530326 994879
rect 530378 994867 530384 994919
rect 158416 994571 158422 994623
rect 158474 994611 158480 994623
rect 178480 994611 178486 994623
rect 158474 994583 178486 994611
rect 158474 994571 158480 994583
rect 178480 994571 178486 994583
rect 178538 994571 178544 994623
rect 141232 994497 141238 994549
rect 141290 994537 141296 994549
rect 146992 994537 146998 994549
rect 141290 994509 146998 994537
rect 141290 994497 141296 994509
rect 146992 994497 146998 994509
rect 147050 994497 147056 994549
rect 574480 994127 574486 994179
rect 574538 994167 574544 994179
rect 635248 994167 635254 994179
rect 574538 994139 635254 994167
rect 574538 994127 574544 994139
rect 635248 994127 635254 994139
rect 635306 994127 635312 994179
rect 572752 993979 572758 994031
rect 572810 994019 572816 994031
rect 636112 994019 636118 994031
rect 572810 993991 636118 994019
rect 572810 993979 572816 993991
rect 636112 993979 636118 993991
rect 636170 993979 636176 994031
rect 180496 993905 180502 993957
rect 180554 993945 180560 993957
rect 201712 993945 201718 993957
rect 180554 993917 201718 993945
rect 180554 993905 180560 993917
rect 201712 993905 201718 993917
rect 201770 993905 201776 993957
rect 234928 993905 234934 993957
rect 234986 993945 234992 993957
rect 250480 993945 250486 993957
rect 234986 993917 250486 993945
rect 234986 993905 234992 993917
rect 250480 993905 250486 993917
rect 250538 993905 250544 993957
rect 570640 993905 570646 993957
rect 570698 993945 570704 993957
rect 639184 993945 639190 993957
rect 570698 993917 639190 993945
rect 570698 993905 570704 993917
rect 639184 993905 639190 993917
rect 639242 993905 639248 993957
rect 182992 993831 182998 993883
rect 183050 993871 183056 993883
rect 207280 993871 207286 993883
rect 183050 993843 207286 993871
rect 183050 993831 183056 993843
rect 207280 993831 207286 993843
rect 207338 993831 207344 993883
rect 232144 993831 232150 993883
rect 232202 993871 232208 993883
rect 253360 993871 253366 993883
rect 232202 993843 253366 993871
rect 232202 993831 232208 993843
rect 253360 993831 253366 993843
rect 253418 993831 253424 993883
rect 368656 993831 368662 993883
rect 368714 993871 368720 993883
rect 392656 993871 392662 993883
rect 368714 993843 392662 993871
rect 368714 993831 368720 993843
rect 392656 993831 392662 993843
rect 392714 993831 392720 993883
rect 572656 993831 572662 993883
rect 572714 993871 572720 993883
rect 634864 993871 634870 993883
rect 572714 993843 634870 993871
rect 572714 993831 572720 993843
rect 634864 993831 634870 993843
rect 634922 993831 634928 993883
rect 77680 993757 77686 993809
rect 77738 993797 77744 993809
rect 100720 993797 100726 993809
rect 77738 993769 100726 993797
rect 77738 993757 77744 993769
rect 100720 993757 100726 993769
rect 100778 993757 100784 993809
rect 129328 993757 129334 993809
rect 129386 993797 129392 993809
rect 152560 993797 152566 993809
rect 129386 993769 152566 993797
rect 129386 993757 129392 993769
rect 152560 993757 152566 993769
rect 152618 993757 152624 993809
rect 181360 993757 181366 993809
rect 181418 993797 181424 993809
rect 212656 993797 212662 993809
rect 181418 993769 212662 993797
rect 181418 993757 181424 993769
rect 212656 993757 212662 993769
rect 212714 993757 212720 993809
rect 234352 993757 234358 993809
rect 234410 993797 234416 993809
rect 261424 993797 261430 993809
rect 234410 993769 261430 993797
rect 234410 993757 234416 993769
rect 261424 993757 261430 993769
rect 261482 993757 261488 993809
rect 512752 993757 512758 993809
rect 512810 993797 512816 993809
rect 534352 993797 534358 993809
rect 512810 993769 534358 993797
rect 512810 993757 512816 993769
rect 534352 993757 534358 993769
rect 534410 993757 534416 993809
rect 570736 993757 570742 993809
rect 570794 993797 570800 993809
rect 637360 993797 637366 993809
rect 570794 993769 637366 993797
rect 570794 993757 570800 993769
rect 637360 993757 637366 993769
rect 637418 993757 637424 993809
rect 80176 993683 80182 993735
rect 80234 993723 80240 993735
rect 107248 993723 107254 993735
rect 80234 993695 107254 993723
rect 80234 993683 80240 993695
rect 107248 993683 107254 993695
rect 107306 993683 107312 993735
rect 128464 993683 128470 993735
rect 128522 993723 128528 993735
rect 159568 993723 159574 993735
rect 128522 993695 159574 993723
rect 128522 993683 128528 993695
rect 159568 993683 159574 993695
rect 159626 993683 159632 993735
rect 179824 993683 179830 993735
rect 179882 993723 179888 993735
rect 211024 993723 211030 993735
rect 179882 993695 211030 993723
rect 179882 993683 179888 993695
rect 211024 993683 211030 993695
rect 211082 993683 211088 993735
rect 232528 993683 232534 993735
rect 232586 993723 232592 993735
rect 264016 993723 264022 993735
rect 232586 993695 264022 993723
rect 232586 993683 232592 993695
rect 264016 993683 264022 993695
rect 264074 993683 264080 993735
rect 368752 993683 368758 993735
rect 368810 993723 368816 993735
rect 393712 993723 393718 993735
rect 368810 993695 393718 993723
rect 368810 993683 368816 993695
rect 393712 993683 393718 993695
rect 393770 993683 393776 993735
rect 506608 993683 506614 993735
rect 506666 993723 506672 993735
rect 538960 993723 538966 993735
rect 506666 993695 538966 993723
rect 506666 993683 506672 993695
rect 538960 993683 538966 993695
rect 539018 993683 539024 993735
rect 557968 993683 557974 993735
rect 558026 993723 558032 993735
rect 641008 993723 641014 993735
rect 558026 993695 641014 993723
rect 558026 993683 558032 993695
rect 641008 993683 641014 993695
rect 641066 993683 641072 993735
rect 77296 993609 77302 993661
rect 77354 993649 77360 993661
rect 108208 993649 108214 993661
rect 77354 993621 108214 993649
rect 77354 993609 77360 993621
rect 108208 993609 108214 993621
rect 108266 993609 108272 993661
rect 129712 993609 129718 993661
rect 129770 993649 129776 993661
rect 161200 993649 161206 993661
rect 129770 993621 161206 993649
rect 129770 993609 129776 993621
rect 161200 993609 161206 993621
rect 161258 993609 161264 993661
rect 185392 993609 185398 993661
rect 185450 993649 185456 993661
rect 236752 993649 236758 993661
rect 185450 993621 236758 993649
rect 185450 993609 185456 993621
rect 236752 993609 236758 993621
rect 236810 993649 236816 993661
rect 279280 993649 279286 993661
rect 236810 993621 279286 993649
rect 236810 993609 236816 993621
rect 279280 993609 279286 993621
rect 279338 993609 279344 993661
rect 282832 993609 282838 993661
rect 282890 993649 282896 993661
rect 313840 993649 313846 993661
rect 282890 993621 313846 993649
rect 282890 993609 282896 993621
rect 313840 993609 313846 993621
rect 313898 993609 313904 993661
rect 362320 993609 362326 993661
rect 362378 993649 362384 993661
rect 398800 993649 398806 993661
rect 362378 993621 398806 993649
rect 362378 993609 362384 993621
rect 398800 993609 398806 993621
rect 398858 993609 398864 993661
rect 429712 993609 429718 993661
rect 429770 993649 429776 993661
rect 487792 993649 487798 993661
rect 429770 993621 487798 993649
rect 429770 993609 429776 993621
rect 487792 993609 487798 993621
rect 487850 993609 487856 993661
rect 530320 993609 530326 993661
rect 530378 993649 530384 993661
rect 630832 993649 630838 993661
rect 530378 993621 630838 993649
rect 530378 993609 530384 993621
rect 630832 993609 630838 993621
rect 630890 993649 630896 993661
rect 632368 993649 632374 993661
rect 630890 993621 632374 993649
rect 630890 993609 630896 993621
rect 632368 993609 632374 993621
rect 632426 993609 632432 993661
rect 638896 993609 638902 993661
rect 638954 993649 638960 993661
rect 643600 993649 643606 993661
rect 638954 993621 643606 993649
rect 638954 993609 638960 993621
rect 643600 993609 643606 993621
rect 643658 993609 643664 993661
rect 469456 993535 469462 993587
rect 469514 993575 469520 993587
rect 479152 993575 479158 993587
rect 469514 993547 479158 993575
rect 469514 993535 469520 993547
rect 479152 993535 479158 993547
rect 479210 993575 479216 993587
rect 489520 993575 489526 993587
rect 479210 993547 489526 993575
rect 479210 993535 479216 993547
rect 489520 993535 489526 993547
rect 489578 993535 489584 993587
rect 331216 992129 331222 992181
rect 331274 992169 331280 992181
rect 332560 992169 332566 992181
rect 331274 992141 332566 992169
rect 331274 992129 331280 992141
rect 332560 992129 332566 992141
rect 332618 992129 332624 992181
rect 285136 991611 285142 991663
rect 285194 991651 285200 991663
rect 298576 991651 298582 991663
rect 285194 991623 298582 991651
rect 285194 991611 285200 991623
rect 298576 991611 298582 991623
rect 298634 991611 298640 991663
rect 241936 990871 241942 990923
rect 241994 990911 242000 990923
rect 246448 990911 246454 990923
rect 241994 990883 246454 990911
rect 241994 990871 242000 990883
rect 246448 990871 246454 990883
rect 246506 990871 246512 990923
rect 629200 990871 629206 990923
rect 629258 990911 629264 990923
rect 642160 990911 642166 990923
rect 629258 990883 642166 990911
rect 629258 990871 629264 990883
rect 642160 990871 642166 990883
rect 642218 990871 642224 990923
rect 640336 989465 640342 989517
rect 640394 989505 640400 989517
rect 650224 989505 650230 989517
rect 640394 989477 650230 989505
rect 640394 989465 640400 989477
rect 650224 989465 650230 989477
rect 650282 989465 650288 989517
rect 645232 988503 645238 988555
rect 645290 988543 645296 988555
rect 650032 988543 650038 988555
rect 645290 988515 650038 988543
rect 645290 988503 645296 988515
rect 650032 988503 650038 988515
rect 650090 988503 650096 988555
rect 604720 988207 604726 988259
rect 604778 988247 604784 988259
rect 618544 988247 618550 988259
rect 604778 988219 618550 988247
rect 604778 988207 604784 988219
rect 618544 988207 618550 988219
rect 618602 988207 618608 988259
rect 69136 987877 69142 987889
rect 67714 987849 69142 987877
rect 64912 987763 64918 987815
rect 64970 987803 64976 987815
rect 67714 987803 67742 987849
rect 69136 987837 69142 987849
rect 69194 987837 69200 987889
rect 241936 987877 241942 987889
rect 239074 987849 241942 987877
rect 64970 987775 67742 987803
rect 64970 987763 64976 987775
rect 223120 987763 223126 987815
rect 223178 987803 223184 987815
rect 235600 987803 235606 987815
rect 223178 987775 235606 987803
rect 223178 987763 223184 987775
rect 235600 987763 235606 987775
rect 235658 987763 235664 987815
rect 236272 987763 236278 987815
rect 236330 987803 236336 987815
rect 239074 987803 239102 987849
rect 241936 987837 241942 987849
rect 241994 987837 242000 987889
rect 236330 987775 239102 987803
rect 236330 987763 236336 987775
rect 518416 987763 518422 987815
rect 518474 987803 518480 987815
rect 527632 987803 527638 987815
rect 518474 987775 527638 987803
rect 518474 987763 518480 987775
rect 527632 987763 527638 987775
rect 527690 987763 527696 987815
rect 570256 987763 570262 987815
rect 570314 987803 570320 987815
rect 576304 987803 576310 987815
rect 570314 987775 576310 987803
rect 570314 987763 570320 987775
rect 576304 987763 576310 987775
rect 576362 987763 576368 987815
rect 645136 987763 645142 987815
rect 645194 987803 645200 987815
rect 649360 987803 649366 987815
rect 645194 987775 649366 987803
rect 645194 987763 645200 987775
rect 649360 987763 649366 987775
rect 649418 987763 649424 987815
rect 219472 987171 219478 987223
rect 219530 987211 219536 987223
rect 221872 987211 221878 987223
rect 219530 987183 221878 987211
rect 219530 987171 219536 987183
rect 221872 987171 221878 987183
rect 221930 987171 221936 987223
rect 374416 986505 374422 986557
rect 374474 986545 374480 986557
rect 397840 986545 397846 986557
rect 374474 986517 397846 986545
rect 374474 986505 374480 986517
rect 397840 986505 397846 986517
rect 397898 986505 397904 986557
rect 570352 986505 570358 986557
rect 570410 986545 570416 986557
rect 592432 986545 592438 986557
rect 570410 986517 592438 986545
rect 570410 986505 570416 986517
rect 592432 986505 592438 986517
rect 592490 986505 592496 986557
rect 630736 986505 630742 986557
rect 630794 986545 630800 986557
rect 639376 986545 639382 986557
rect 630794 986517 639382 986545
rect 630794 986505 630800 986517
rect 639376 986505 639382 986517
rect 639434 986505 639440 986557
rect 326800 986431 326806 986483
rect 326858 986471 326864 986483
rect 349168 986471 349174 986483
rect 326858 986443 349174 986471
rect 326858 986431 326864 986443
rect 349168 986431 349174 986443
rect 349226 986431 349232 986483
rect 377296 986431 377302 986483
rect 377354 986471 377360 986483
rect 414064 986471 414070 986483
rect 377354 986443 414070 986471
rect 377354 986431 377360 986443
rect 414064 986431 414070 986443
rect 414122 986431 414128 986483
rect 445072 986431 445078 986483
rect 445130 986471 445136 986483
rect 478960 986471 478966 986483
rect 445130 986443 478966 986471
rect 445130 986431 445136 986443
rect 478960 986431 478966 986443
rect 479018 986431 479024 986483
rect 521296 986431 521302 986483
rect 521354 986471 521360 986483
rect 543760 986471 543766 986483
rect 521354 986443 543766 986471
rect 521354 986431 521360 986443
rect 543760 986431 543766 986443
rect 543818 986431 543824 986483
rect 573136 986431 573142 986483
rect 573194 986471 573200 986483
rect 608752 986471 608758 986483
rect 573194 986443 608758 986471
rect 573194 986431 573200 986443
rect 608752 986431 608758 986443
rect 608810 986431 608816 986483
rect 622000 986431 622006 986483
rect 622058 986471 622064 986483
rect 641104 986471 641110 986483
rect 622058 986443 641110 986471
rect 622058 986431 622064 986443
rect 641104 986431 641110 986443
rect 641162 986431 641168 986483
rect 73456 986357 73462 986409
rect 73514 986397 73520 986409
rect 93616 986397 93622 986409
rect 73514 986369 93622 986397
rect 73514 986357 73520 986369
rect 93616 986357 93622 986369
rect 93674 986357 93680 986409
rect 138256 986357 138262 986409
rect 138314 986397 138320 986409
rect 164080 986397 164086 986409
rect 138314 986369 164086 986397
rect 138314 986357 138320 986369
rect 164080 986357 164086 986369
rect 164138 986357 164144 986409
rect 273712 986357 273718 986409
rect 273770 986397 273776 986409
rect 300496 986397 300502 986409
rect 273770 986369 300502 986397
rect 273770 986357 273776 986369
rect 300496 986357 300502 986369
rect 300554 986357 300560 986409
rect 323920 986357 323926 986409
rect 323978 986397 323984 986409
rect 365392 986397 365398 986409
rect 323978 986369 365398 986397
rect 323978 986357 323984 986369
rect 365392 986357 365398 986369
rect 365450 986357 365456 986409
rect 374608 986357 374614 986409
rect 374666 986397 374672 986409
rect 430288 986397 430294 986409
rect 374666 986369 430294 986397
rect 374666 986357 374672 986369
rect 430288 986357 430294 986369
rect 430346 986357 430352 986409
rect 440656 986357 440662 986409
rect 440714 986397 440720 986409
rect 495184 986397 495190 986409
rect 440714 986369 495190 986397
rect 440714 986357 440720 986369
rect 495184 986357 495190 986369
rect 495242 986357 495248 986409
rect 518608 986357 518614 986409
rect 518666 986397 518672 986409
rect 560080 986397 560086 986409
rect 518666 986369 560086 986397
rect 518666 986357 518672 986369
rect 560080 986357 560086 986369
rect 560138 986357 560144 986409
rect 570544 986357 570550 986409
rect 570602 986397 570608 986409
rect 624976 986397 624982 986409
rect 570602 986369 624982 986397
rect 570602 986357 570608 986369
rect 624976 986357 624982 986369
rect 625034 986357 625040 986409
rect 630736 986357 630742 986409
rect 630794 986397 630800 986409
rect 631024 986397 631030 986409
rect 630794 986369 631030 986397
rect 630794 986357 630800 986369
rect 631024 986357 631030 986369
rect 631082 986357 631088 986409
rect 203152 986283 203158 986335
rect 203210 986323 203216 986335
rect 213040 986323 213046 986335
rect 203210 986295 213046 986323
rect 203210 986283 203216 986295
rect 213040 986283 213046 986295
rect 213098 986283 213104 986335
rect 273616 986135 273622 986187
rect 273674 986175 273680 986187
rect 284272 986175 284278 986187
rect 273674 986147 284278 986175
rect 273674 986135 273680 986147
rect 284272 986135 284278 986147
rect 284330 986135 284336 986187
rect 154480 985987 154486 986039
rect 154538 986027 154544 986039
rect 163984 986027 163990 986039
rect 154538 985999 163990 986027
rect 154538 985987 154544 985999
rect 163984 985987 163990 985999
rect 164042 985987 164048 986039
rect 89584 985839 89590 985891
rect 89642 985879 89648 985891
rect 93712 985879 93718 985891
rect 89642 985851 93718 985879
rect 89642 985839 89648 985851
rect 93712 985839 93718 985851
rect 93770 985839 93776 985891
rect 45040 985469 45046 985521
rect 45098 985509 45104 985521
rect 45098 985481 47774 985509
rect 45098 985469 45104 985481
rect 47746 985287 47774 985481
rect 80752 985469 80758 985521
rect 80810 985509 80816 985521
rect 100816 985509 100822 985521
rect 80810 985481 100822 985509
rect 80810 985469 80816 985481
rect 100816 985469 100822 985481
rect 100874 985469 100880 985521
rect 120880 985469 120886 985521
rect 120938 985509 120944 985521
rect 146800 985509 146806 985521
rect 120938 985481 146806 985509
rect 120938 985469 120944 985481
rect 146800 985469 146806 985481
rect 146858 985469 146864 985521
rect 201520 985509 201526 985521
rect 191362 985481 201526 985509
rect 50512 985395 50518 985447
rect 50570 985435 50576 985447
rect 122032 985435 122038 985447
rect 50570 985407 122038 985435
rect 50570 985395 50576 985407
rect 122032 985395 122038 985407
rect 122090 985395 122096 985447
rect 146992 985395 146998 985447
rect 147050 985435 147056 985447
rect 191362 985435 191390 985481
rect 201520 985469 201526 985481
rect 201578 985469 201584 985521
rect 201616 985469 201622 985521
rect 201674 985509 201680 985521
rect 218896 985509 218902 985521
rect 201674 985481 218902 985509
rect 201674 985469 201680 985481
rect 218896 985469 218902 985481
rect 218954 985469 218960 985521
rect 147050 985407 191390 985435
rect 147050 985395 147056 985407
rect 239152 985395 239158 985447
rect 239210 985435 239216 985447
rect 251824 985435 251830 985447
rect 239210 985407 251830 985435
rect 239210 985395 239216 985407
rect 251824 985395 251830 985407
rect 251882 985395 251888 985447
rect 47824 985321 47830 985373
rect 47882 985361 47888 985373
rect 186928 985361 186934 985373
rect 47882 985333 186934 985361
rect 47882 985321 47888 985333
rect 186928 985321 186934 985333
rect 186986 985321 186992 985373
rect 218992 985321 218998 985373
rect 219050 985361 219056 985373
rect 219050 985333 239006 985361
rect 219050 985321 219056 985333
rect 80560 985287 80566 985299
rect 47746 985259 80566 985287
rect 80560 985247 80566 985259
rect 80618 985247 80624 985299
rect 238978 985287 239006 985333
rect 279376 985321 279382 985373
rect 279434 985361 279440 985373
rect 285136 985361 285142 985373
rect 279434 985333 285142 985361
rect 279434 985321 279440 985333
rect 285136 985321 285142 985333
rect 285194 985321 285200 985373
rect 239152 985287 239158 985299
rect 238978 985259 239158 985287
rect 239152 985247 239158 985259
rect 239210 985247 239216 985299
rect 45136 985173 45142 985225
rect 45194 985213 45200 985225
rect 239056 985213 239062 985225
rect 45194 985185 239062 985213
rect 45194 985173 45200 985185
rect 239056 985173 239062 985185
rect 239114 985173 239120 985225
rect 239536 985173 239542 985225
rect 239594 985213 239600 985225
rect 316720 985213 316726 985225
rect 239594 985185 316726 985213
rect 239594 985173 239600 985185
rect 316720 985173 316726 985185
rect 316778 985173 316784 985225
rect 44944 985099 44950 985151
rect 45002 985139 45008 985151
rect 239152 985139 239158 985151
rect 45002 985111 239158 985139
rect 45002 985099 45008 985111
rect 239152 985099 239158 985111
rect 239210 985099 239216 985151
rect 239728 985099 239734 985151
rect 239786 985139 239792 985151
rect 381616 985139 381622 985151
rect 239786 985111 381622 985139
rect 239786 985099 239792 985111
rect 381616 985099 381622 985111
rect 381674 985099 381680 985151
rect 444880 985099 444886 985151
rect 444938 985139 444944 985151
rect 462736 985139 462742 985151
rect 444938 985111 462742 985139
rect 444938 985099 444944 985111
rect 462736 985099 462742 985111
rect 462794 985099 462800 985151
rect 44848 985025 44854 985077
rect 44906 985065 44912 985077
rect 239056 985065 239062 985077
rect 44906 985037 239062 985065
rect 44906 985025 44912 985037
rect 239056 985025 239062 985037
rect 239114 985025 239120 985077
rect 239440 985025 239446 985077
rect 239498 985065 239504 985077
rect 446512 985065 446518 985077
rect 239498 985037 446518 985065
rect 239498 985025 239504 985037
rect 446512 985025 446518 985037
rect 446570 985025 446576 985077
rect 42928 984951 42934 985003
rect 42986 984991 42992 985003
rect 511408 984991 511414 985003
rect 42986 984963 511414 984991
rect 42986 984951 42992 984963
rect 511408 984951 511414 984963
rect 511466 984951 511472 985003
rect 642256 984951 642262 985003
rect 642314 984991 642320 985003
rect 642314 984963 645182 984991
rect 642314 984951 642320 984963
rect 645154 984917 645182 984963
rect 649456 984917 649462 984929
rect 645154 984889 649462 984917
rect 649456 984877 649462 984889
rect 649514 984877 649520 984929
rect 65008 983841 65014 983893
rect 65066 983881 65072 983893
rect 94960 983881 94966 983893
rect 65066 983853 94966 983881
rect 65066 983841 65072 983853
rect 94960 983841 94966 983853
rect 95018 983841 95024 983893
rect 47440 983767 47446 983819
rect 47498 983807 47504 983819
rect 118096 983807 118102 983819
rect 47498 983779 118102 983807
rect 47498 983767 47504 983779
rect 118096 983767 118102 983779
rect 118154 983767 118160 983819
rect 618544 983767 618550 983819
rect 618602 983807 618608 983819
rect 649648 983807 649654 983819
rect 618602 983779 649654 983807
rect 618602 983767 618608 983779
rect 649648 983767 649654 983779
rect 649706 983767 649712 983819
rect 44752 983693 44758 983745
rect 44810 983733 44816 983745
rect 115216 983733 115222 983745
rect 44810 983705 115222 983733
rect 44810 983693 44816 983705
rect 115216 983693 115222 983705
rect 115274 983693 115280 983745
rect 568720 983693 568726 983745
rect 568778 983733 568784 983745
rect 652240 983733 652246 983745
rect 568778 983705 652246 983733
rect 568778 983693 568784 983705
rect 652240 983693 652246 983705
rect 652298 983693 652304 983745
rect 44560 983619 44566 983671
rect 44618 983659 44624 983671
rect 115312 983659 115318 983671
rect 44618 983631 115318 983659
rect 44618 983619 44624 983631
rect 115312 983619 115318 983631
rect 115370 983619 115376 983671
rect 567472 983619 567478 983671
rect 567530 983659 567536 983671
rect 658000 983659 658006 983671
rect 567530 983631 658006 983659
rect 567530 983619 567536 983631
rect 658000 983619 658006 983631
rect 658058 983619 658064 983671
rect 65104 983545 65110 983597
rect 65162 983585 65168 983597
rect 145264 983585 145270 983597
rect 65162 983557 145270 983585
rect 65162 983545 65168 983557
rect 145264 983545 145270 983557
rect 145322 983545 145328 983597
rect 567376 983545 567382 983597
rect 567434 983585 567440 983597
rect 658096 983585 658102 983597
rect 567434 983557 658102 983585
rect 567434 983545 567440 983557
rect 658096 983545 658102 983557
rect 658154 983545 658160 983597
rect 65200 983471 65206 983523
rect 65258 983511 65264 983523
rect 195376 983511 195382 983523
rect 65258 983483 195382 983511
rect 65258 983471 65264 983483
rect 195376 983471 195382 983483
rect 195434 983471 195440 983523
rect 217360 983471 217366 983523
rect 217418 983511 217424 983523
rect 236272 983511 236278 983523
rect 217418 983483 236278 983511
rect 217418 983471 217424 983483
rect 236272 983471 236278 983483
rect 236330 983471 236336 983523
rect 544240 983471 544246 983523
rect 544298 983511 544304 983523
rect 650896 983511 650902 983523
rect 544298 983483 650902 983511
rect 544298 983471 544304 983483
rect 650896 983471 650902 983483
rect 650954 983471 650960 983523
rect 273616 982287 273622 982339
rect 273674 982327 273680 982339
rect 279376 982327 279382 982339
rect 273674 982299 279382 982327
rect 273674 982287 273680 982299
rect 279376 982287 279382 982299
rect 279434 982287 279440 982339
rect 643600 981769 643606 981821
rect 643658 981809 643664 981821
rect 649840 981809 649846 981821
rect 643658 981781 649846 981809
rect 643658 981769 643664 981781
rect 649840 981769 649846 981781
rect 649898 981769 649904 981821
rect 639376 981325 639382 981377
rect 639434 981365 639440 981377
rect 650128 981365 650134 981377
rect 639434 981337 650134 981365
rect 639434 981325 639440 981337
rect 650128 981325 650134 981337
rect 650186 981325 650192 981377
rect 130384 981029 130390 981081
rect 130442 981069 130448 981081
rect 130442 981041 151166 981069
rect 130442 981029 130448 981041
rect 106480 980995 106486 981007
rect 80674 980967 106486 980995
rect 64720 980807 64726 980859
rect 64778 980847 64784 980859
rect 80674 980847 80702 980967
rect 106480 980955 106486 980967
rect 106538 980955 106544 981007
rect 106576 980955 106582 981007
rect 106634 980995 106640 981007
rect 106634 980967 110846 980995
rect 106634 980955 106640 980967
rect 110818 980921 110846 980967
rect 130384 980921 130390 980933
rect 110818 980893 130390 980921
rect 130384 980881 130390 980893
rect 130442 980881 130448 980933
rect 151138 980921 151166 981041
rect 161296 980955 161302 981007
rect 161354 980955 161360 981007
rect 161314 980921 161342 980955
rect 178480 980921 178486 980933
rect 151138 980893 161342 980921
rect 168418 980893 178486 980921
rect 64778 980819 80702 980847
rect 110818 980819 126494 980847
rect 64778 980807 64784 980819
rect 106480 980773 106486 980785
rect 80674 980745 106486 980773
rect 64816 980659 64822 980711
rect 64874 980699 64880 980711
rect 80674 980699 80702 980745
rect 106480 980733 106486 980745
rect 106538 980733 106544 980785
rect 106576 980733 106582 980785
rect 106634 980773 106640 980785
rect 110818 980773 110846 980819
rect 106634 980745 110846 980773
rect 106634 980733 106640 980745
rect 64874 980671 80702 980699
rect 126466 980699 126494 980819
rect 146896 980807 146902 980859
rect 146954 980847 146960 980859
rect 168418 980847 168446 980893
rect 178480 980881 178486 980893
rect 178538 980881 178544 980933
rect 146954 980819 168446 980847
rect 146954 980807 146960 980819
rect 171280 980807 171286 980859
rect 171338 980847 171344 980859
rect 171338 980819 207326 980847
rect 171338 980807 171344 980819
rect 146800 980773 146806 980785
rect 131074 980745 146806 980773
rect 131074 980699 131102 980745
rect 146800 980733 146806 980745
rect 146858 980733 146864 980785
rect 178480 980733 178486 980785
rect 178538 980733 178544 980785
rect 207298 980773 207326 980819
rect 238960 980807 238966 980859
rect 239018 980847 239024 980859
rect 247600 980847 247606 980859
rect 239018 980819 247606 980847
rect 239018 980807 239024 980819
rect 247600 980807 247606 980819
rect 247658 980807 247664 980859
rect 247696 980807 247702 980859
rect 247754 980847 247760 980859
rect 247754 980819 259166 980847
rect 247754 980807 247760 980819
rect 217360 980773 217366 980785
rect 207298 980745 217366 980773
rect 217360 980733 217366 980745
rect 217418 980733 217424 980785
rect 217552 980773 217558 980785
rect 217474 980745 217558 980773
rect 126466 980671 131102 980699
rect 178498 980699 178526 980733
rect 217474 980699 217502 980745
rect 217552 980733 217558 980745
rect 217610 980733 217616 980785
rect 217648 980733 217654 980785
rect 217706 980773 217712 980785
rect 218896 980773 218902 980785
rect 217706 980745 218902 980773
rect 217706 980733 217712 980745
rect 218896 980733 218902 980745
rect 218954 980733 218960 980785
rect 178498 980671 217502 980699
rect 259138 980699 259166 980819
rect 630832 980807 630838 980859
rect 630890 980807 630896 980859
rect 273616 980733 273622 980785
rect 273674 980733 273680 980785
rect 273634 980699 273662 980733
rect 259138 980671 273662 980699
rect 630850 980699 630878 980807
rect 630928 980733 630934 980785
rect 630986 980773 630992 980785
rect 675088 980773 675094 980785
rect 630986 980745 675094 980773
rect 630986 980733 630992 980745
rect 675088 980733 675094 980745
rect 675146 980733 675152 980785
rect 675280 980699 675286 980711
rect 630850 980671 675286 980699
rect 64874 980659 64880 980671
rect 675280 980659 675286 980671
rect 675338 980659 675344 980711
rect 53296 970595 53302 970647
rect 53354 970635 53360 970647
rect 59536 970635 59542 970647
rect 53354 970607 59542 970635
rect 53354 970595 53360 970607
rect 59536 970595 59542 970607
rect 59594 970595 59600 970647
rect 42160 967265 42166 967317
rect 42218 967305 42224 967317
rect 42928 967305 42934 967317
rect 42218 967277 42934 967305
rect 42218 967265 42224 967277
rect 42928 967265 42934 967277
rect 42986 967265 42992 967317
rect 42064 961345 42070 961397
rect 42122 961385 42128 961397
rect 42544 961385 42550 961397
rect 42122 961357 42550 961385
rect 42122 961345 42128 961357
rect 42544 961345 42550 961357
rect 42602 961345 42608 961397
rect 42160 960679 42166 960731
rect 42218 960719 42224 960731
rect 42352 960719 42358 960731
rect 42218 960691 42358 960719
rect 42218 960679 42224 960691
rect 42352 960679 42358 960691
rect 42410 960679 42416 960731
rect 673936 958977 673942 959029
rect 673994 959017 674000 959029
rect 675472 959017 675478 959029
rect 673994 958989 675478 959017
rect 673994 958977 674000 958989
rect 675472 958977 675478 958989
rect 675530 958977 675536 959029
rect 675088 958385 675094 958437
rect 675146 958425 675152 958437
rect 675376 958425 675382 958437
rect 675146 958397 675382 958425
rect 675146 958385 675152 958397
rect 675376 958385 675382 958397
rect 675434 958385 675440 958437
rect 675184 956979 675190 957031
rect 675242 957019 675248 957031
rect 675472 957019 675478 957031
rect 675242 956991 675478 957019
rect 675242 956979 675248 956991
rect 675472 956979 675478 956991
rect 675530 956979 675536 957031
rect 43120 956165 43126 956217
rect 43178 956205 43184 956217
rect 59536 956205 59542 956217
rect 43178 956177 59542 956205
rect 43178 956165 43184 956177
rect 59536 956165 59542 956177
rect 59594 956165 59600 956217
rect 42064 955277 42070 955329
rect 42122 955317 42128 955329
rect 42928 955317 42934 955329
rect 42122 955289 42934 955317
rect 42122 955277 42128 955289
rect 42928 955277 42934 955289
rect 42986 955277 42992 955329
rect 669520 954685 669526 954737
rect 669578 954725 669584 954737
rect 675376 954725 675382 954737
rect 669578 954697 675382 954725
rect 669578 954685 669584 954697
rect 675376 954685 675382 954697
rect 675434 954685 675440 954737
rect 42160 954611 42166 954663
rect 42218 954651 42224 954663
rect 42832 954651 42838 954663
rect 42218 954623 42838 954651
rect 42218 954611 42224 954623
rect 42832 954611 42838 954623
rect 42890 954611 42896 954663
rect 674128 953871 674134 953923
rect 674186 953911 674192 953923
rect 675472 953911 675478 953923
rect 674186 953883 675478 953911
rect 674186 953871 674192 953883
rect 675472 953871 675478 953883
rect 675530 953871 675536 953923
rect 674032 952021 674038 952073
rect 674090 952061 674096 952073
rect 675472 952061 675478 952073
rect 674090 952033 675478 952061
rect 674090 952021 674096 952033
rect 675472 952021 675478 952033
rect 675530 952021 675536 952073
rect 649552 951799 649558 951851
rect 649610 951839 649616 951851
rect 653776 951839 653782 951851
rect 649610 951811 653782 951839
rect 649610 951799 649616 951811
rect 653776 951799 653782 951811
rect 653834 951799 653840 951851
rect 42352 948543 42358 948595
rect 42410 948583 42416 948595
rect 42640 948583 42646 948595
rect 42410 948555 42646 948583
rect 42410 948543 42416 948555
rect 42640 948543 42646 948555
rect 42698 948543 42704 948595
rect 42352 947729 42358 947781
rect 42410 947769 42416 947781
rect 47536 947769 47542 947781
rect 42410 947741 47542 947769
rect 42410 947729 42416 947741
rect 47536 947729 47542 947741
rect 47594 947729 47600 947781
rect 42160 947655 42166 947707
rect 42218 947695 42224 947707
rect 50320 947695 50326 947707
rect 42218 947667 50326 947695
rect 42218 947655 42224 947667
rect 50320 947655 50326 947667
rect 50378 947655 50384 947707
rect 655216 944843 655222 944895
rect 655274 944883 655280 944895
rect 674704 944883 674710 944895
rect 655274 944855 674710 944883
rect 655274 944843 655280 944855
rect 674704 944843 674710 944855
rect 674762 944843 674768 944895
rect 655120 944621 655126 944673
rect 655178 944661 655184 944673
rect 674704 944661 674710 944673
rect 655178 944633 674710 944661
rect 655178 944621 655184 944633
rect 674704 944621 674710 944633
rect 674762 944621 674768 944673
rect 50320 944547 50326 944599
rect 50378 944587 50384 944599
rect 59536 944587 59542 944599
rect 50378 944559 59542 944587
rect 50378 944547 50384 944559
rect 59536 944547 59542 944559
rect 59594 944547 59600 944599
rect 672304 942327 672310 942379
rect 672362 942367 672368 942379
rect 674704 942367 674710 942379
rect 672362 942339 674710 942367
rect 672362 942327 672368 942339
rect 674704 942327 674710 942339
rect 674762 942327 674768 942379
rect 658096 942179 658102 942231
rect 658154 942219 658160 942231
rect 674704 942219 674710 942231
rect 658154 942191 674710 942219
rect 658154 942179 658160 942191
rect 674704 942179 674710 942191
rect 674762 942179 674768 942231
rect 654352 942031 654358 942083
rect 654410 942071 654416 942083
rect 674608 942071 674614 942083
rect 654410 942043 674614 942071
rect 654410 942031 654416 942043
rect 674608 942031 674614 942043
rect 674666 942031 674672 942083
rect 652240 941883 652246 941935
rect 652298 941923 652304 941935
rect 674800 941923 674806 941935
rect 652298 941895 674806 941923
rect 652298 941883 652304 941895
rect 674800 941883 674806 941895
rect 674858 941883 674864 941935
rect 658000 939071 658006 939123
rect 658058 939111 658064 939123
rect 674704 939111 674710 939123
rect 658058 939083 674710 939111
rect 658058 939071 658064 939083
rect 674704 939071 674710 939083
rect 674762 939071 674768 939123
rect 42352 930931 42358 930983
rect 42410 930971 42416 930983
rect 44560 930971 44566 930983
rect 42410 930943 44566 930971
rect 42410 930931 42416 930943
rect 44560 930931 44566 930943
rect 44618 930931 44624 930983
rect 47536 930191 47542 930243
rect 47594 930231 47600 930243
rect 59536 930231 59542 930243
rect 47594 930203 59542 930231
rect 47594 930191 47600 930203
rect 59536 930191 59542 930203
rect 59594 930191 59600 930243
rect 654448 927453 654454 927505
rect 654506 927493 654512 927505
rect 666736 927493 666742 927505
rect 654506 927465 666742 927493
rect 654506 927453 654512 927465
rect 666736 927453 666742 927465
rect 666794 927453 666800 927505
rect 649552 927379 649558 927431
rect 649610 927419 649616 927431
rect 679792 927419 679798 927431
rect 649610 927391 679798 927419
rect 649610 927379 649616 927391
rect 679792 927379 679798 927391
rect 679850 927379 679856 927431
rect 654448 915835 654454 915887
rect 654506 915875 654512 915887
rect 660976 915875 660982 915887
rect 654506 915847 660982 915875
rect 654506 915835 654512 915847
rect 660976 915835 660982 915847
rect 661034 915835 661040 915887
rect 47440 912949 47446 913001
rect 47498 912989 47504 913001
rect 59536 912989 59542 913001
rect 47498 912961 59542 912989
rect 47498 912949 47504 912961
rect 59536 912949 59542 912961
rect 59594 912949 59600 913001
rect 53200 901479 53206 901531
rect 53258 901519 53264 901531
rect 58192 901519 58198 901531
rect 53258 901491 58198 901519
rect 53258 901479 53264 901491
rect 58192 901479 58198 901491
rect 58250 901479 58256 901531
rect 654448 901479 654454 901531
rect 654506 901519 654512 901531
rect 663952 901519 663958 901531
rect 654506 901491 663958 901519
rect 654506 901479 654512 901491
rect 663952 901479 663958 901491
rect 664010 901479 664016 901531
rect 50416 884163 50422 884215
rect 50474 884203 50480 884215
rect 59536 884203 59542 884215
rect 50474 884175 59542 884203
rect 50474 884163 50480 884175
rect 59536 884163 59542 884175
rect 59594 884163 59600 884215
rect 654448 878391 654454 878443
rect 654506 878431 654512 878443
rect 660880 878431 660886 878443
rect 654506 878403 660886 878431
rect 654506 878391 654512 878403
rect 660880 878391 660886 878403
rect 660938 878391 660944 878443
rect 674992 872101 674998 872153
rect 675050 872141 675056 872153
rect 675472 872141 675478 872153
rect 675050 872113 675478 872141
rect 675050 872101 675056 872113
rect 675472 872101 675478 872113
rect 675530 872101 675536 872153
rect 674512 871657 674518 871709
rect 674570 871697 674576 871709
rect 675184 871697 675190 871709
rect 674570 871669 675190 871697
rect 674570 871657 674576 871669
rect 675184 871657 675190 871669
rect 675242 871697 675248 871709
rect 675376 871697 675382 871709
rect 675242 871669 675382 871697
rect 675242 871657 675248 871669
rect 675376 871657 675382 871669
rect 675434 871657 675440 871709
rect 674320 868993 674326 869045
rect 674378 869033 674384 869045
rect 675472 869033 675478 869045
rect 674378 869005 675478 869033
rect 674378 868993 674384 869005
rect 675472 868993 675478 869005
rect 675530 868993 675536 869045
rect 674224 868327 674230 868379
rect 674282 868367 674288 868379
rect 675376 868367 675382 868379
rect 674282 868339 675382 868367
rect 674282 868327 674288 868339
rect 675376 868327 675382 868339
rect 675434 868327 675440 868379
rect 673648 867809 673654 867861
rect 673706 867849 673712 867861
rect 675376 867849 675382 867861
rect 673706 867821 675382 867849
rect 673706 867809 673712 867821
rect 675376 867809 675382 867821
rect 675434 867809 675440 867861
rect 654448 866921 654454 866973
rect 654506 866961 654512 866973
rect 669616 866961 669622 866973
rect 654506 866933 669622 866961
rect 654506 866921 654512 866933
rect 669616 866921 669622 866933
rect 669674 866921 669680 866973
rect 666640 865293 666646 865345
rect 666698 865333 666704 865345
rect 675376 865333 675382 865345
rect 666698 865305 675382 865333
rect 666698 865293 666704 865305
rect 675376 865293 675382 865305
rect 675434 865293 675440 865345
rect 674896 863961 674902 864013
rect 674954 864001 674960 864013
rect 674992 864001 674998 864013
rect 674954 863973 674998 864001
rect 674954 863961 674960 863973
rect 674992 863961 674998 863973
rect 675050 863961 675056 864013
rect 50320 858263 50326 858315
rect 50378 858303 50384 858315
rect 59536 858303 59542 858315
rect 50378 858275 59542 858303
rect 50378 858263 50384 858275
rect 59536 858263 59542 858275
rect 59594 858263 59600 858315
rect 654448 855377 654454 855429
rect 654506 855417 654512 855429
rect 661168 855417 661174 855429
rect 654506 855389 661174 855417
rect 654506 855377 654512 855389
rect 661168 855377 661174 855389
rect 661226 855377 661232 855429
rect 675184 846645 675190 846697
rect 675242 846685 675248 846697
rect 675376 846685 675382 846697
rect 675242 846657 675382 846685
rect 675242 846645 675248 846657
rect 675376 846645 675382 846657
rect 675434 846645 675440 846697
rect 53392 843833 53398 843885
rect 53450 843873 53456 843885
rect 59536 843873 59542 843885
rect 53450 843845 59542 843873
rect 53450 843833 53456 843845
rect 59536 843833 59542 843845
rect 59594 843833 59600 843885
rect 674800 843833 674806 843885
rect 674858 843873 674864 843885
rect 674896 843873 674902 843885
rect 674858 843845 674902 843873
rect 674858 843833 674864 843845
rect 674896 843833 674902 843845
rect 674954 843833 674960 843885
rect 654448 832363 654454 832415
rect 654506 832403 654512 832415
rect 666832 832403 666838 832415
rect 654506 832375 666838 832403
rect 654506 832363 654512 832375
rect 666832 832363 666838 832375
rect 666890 832363 666896 832415
rect 50608 829477 50614 829529
rect 50666 829517 50672 829529
rect 59536 829517 59542 829529
rect 50666 829489 59542 829517
rect 50666 829477 50672 829489
rect 59536 829477 59542 829489
rect 59594 829477 59600 829529
rect 675376 826591 675382 826643
rect 675434 826631 675440 826643
rect 675568 826631 675574 826643
rect 675434 826603 675574 826631
rect 675434 826591 675440 826603
rect 675568 826591 675574 826603
rect 675626 826591 675632 826643
rect 42352 823853 42358 823905
rect 42410 823893 42416 823905
rect 50416 823893 50422 823905
rect 42410 823865 50422 823893
rect 42410 823853 42416 823865
rect 50416 823853 50422 823865
rect 50474 823853 50480 823905
rect 42352 822225 42358 822277
rect 42410 822265 42416 822277
rect 53200 822265 53206 822277
rect 42410 822237 53206 822265
rect 42410 822225 42416 822237
rect 53200 822225 53206 822237
rect 53258 822225 53264 822277
rect 42448 821855 42454 821907
rect 42506 821895 42512 821907
rect 58960 821895 58966 821907
rect 42506 821867 58966 821895
rect 42506 821855 42512 821867
rect 58960 821855 58966 821867
rect 59018 821855 59024 821907
rect 654448 820819 654454 820871
rect 654506 820859 654512 820871
rect 663760 820859 663766 820871
rect 654506 820831 663766 820859
rect 654506 820819 654512 820831
rect 663760 820819 663766 820831
rect 663818 820819 663824 820871
rect 47536 815047 47542 815099
rect 47594 815087 47600 815099
rect 59536 815087 59542 815099
rect 47594 815059 59542 815087
rect 47594 815047 47600 815059
rect 59536 815047 59542 815059
rect 59594 815047 59600 815099
rect 654448 809275 654454 809327
rect 654506 809315 654512 809327
rect 664048 809315 664054 809327
rect 654506 809287 664054 809315
rect 654506 809275 654512 809287
rect 664048 809275 664054 809287
rect 664106 809275 664112 809327
rect 650128 809201 650134 809253
rect 650186 809241 650192 809253
rect 653776 809241 653782 809253
rect 650186 809213 653782 809241
rect 650186 809201 650192 809213
rect 653776 809201 653782 809213
rect 653834 809201 653840 809253
rect 42256 805131 42262 805183
rect 42314 805171 42320 805183
rect 44752 805171 44758 805183
rect 42314 805143 44758 805171
rect 42314 805131 42320 805143
rect 44752 805131 44758 805143
rect 44810 805131 44816 805183
rect 42352 804391 42358 804443
rect 42410 804431 42416 804443
rect 42928 804431 42934 804443
rect 42410 804403 42934 804431
rect 42410 804391 42416 804403
rect 42928 804391 42934 804403
rect 42986 804391 42992 804443
rect 42448 804095 42454 804147
rect 42506 804135 42512 804147
rect 42736 804135 42742 804147
rect 42506 804107 42742 804135
rect 42506 804095 42512 804107
rect 42736 804095 42742 804107
rect 42794 804095 42800 804147
rect 40144 803429 40150 803481
rect 40202 803469 40208 803481
rect 42448 803469 42454 803481
rect 40202 803441 42454 803469
rect 40202 803429 40208 803441
rect 42448 803429 42454 803441
rect 42506 803429 42512 803481
rect 41968 802393 41974 802445
rect 42026 802433 42032 802445
rect 42832 802433 42838 802445
rect 42026 802405 42838 802433
rect 42026 802393 42032 802405
rect 42832 802393 42838 802405
rect 42890 802393 42896 802445
rect 43024 801579 43030 801631
rect 43082 801619 43088 801631
rect 43408 801619 43414 801631
rect 43082 801591 43414 801619
rect 43082 801579 43088 801591
rect 43408 801579 43414 801591
rect 43466 801579 43472 801631
rect 43024 801431 43030 801483
rect 43082 801471 43088 801483
rect 44848 801471 44854 801483
rect 43082 801443 44854 801471
rect 43082 801431 43088 801443
rect 44848 801431 44854 801443
rect 44906 801431 44912 801483
rect 53200 800617 53206 800669
rect 53258 800657 53264 800669
rect 59536 800657 59542 800669
rect 53258 800629 59542 800657
rect 53258 800617 53264 800629
rect 59536 800617 59542 800629
rect 59594 800617 59600 800669
rect 41680 800543 41686 800595
rect 41738 800583 41744 800595
rect 43504 800583 43510 800595
rect 41738 800555 43510 800583
rect 41738 800543 41744 800555
rect 43504 800543 43510 800555
rect 43562 800543 43568 800595
rect 41584 800469 41590 800521
rect 41642 800509 41648 800521
rect 43312 800509 43318 800521
rect 41642 800481 43318 800509
rect 41642 800469 41648 800481
rect 43312 800469 43318 800481
rect 43370 800469 43376 800521
rect 41872 800173 41878 800225
rect 41930 800173 41936 800225
rect 41890 799781 41918 800173
rect 41872 799729 41878 799781
rect 41930 799729 41936 799781
rect 42160 798027 42166 798079
rect 42218 798067 42224 798079
rect 42448 798067 42454 798079
rect 42218 798039 42454 798067
rect 42218 798027 42224 798039
rect 42448 798027 42454 798039
rect 42506 798027 42512 798079
rect 42064 797287 42070 797339
rect 42122 797327 42128 797339
rect 43024 797327 43030 797339
rect 42122 797299 43030 797327
rect 42122 797287 42128 797299
rect 43024 797287 43030 797299
rect 43082 797287 43088 797339
rect 43024 797139 43030 797191
rect 43082 797179 43088 797191
rect 43312 797179 43318 797191
rect 43082 797151 43318 797179
rect 43082 797139 43088 797151
rect 43312 797139 43318 797151
rect 43370 797139 43376 797191
rect 42160 796251 42166 796303
rect 42218 796291 42224 796303
rect 43120 796291 43126 796303
rect 42218 796263 43126 796291
rect 42218 796251 42224 796263
rect 43120 796251 43126 796263
rect 43178 796251 43184 796303
rect 43120 796103 43126 796155
rect 43178 796143 43184 796155
rect 43408 796143 43414 796155
rect 43178 796115 43414 796143
rect 43178 796103 43184 796115
rect 43408 796103 43414 796115
rect 43466 796103 43472 796155
rect 42160 794993 42166 795045
rect 42218 795033 42224 795045
rect 42736 795033 42742 795045
rect 42218 795005 42742 795033
rect 42218 794993 42224 795005
rect 42736 794993 42742 795005
rect 42794 794993 42800 795045
rect 42160 793809 42166 793861
rect 42218 793849 42224 793861
rect 42448 793849 42454 793861
rect 42218 793821 42454 793849
rect 42218 793809 42224 793821
rect 42448 793809 42454 793821
rect 42506 793809 42512 793861
rect 42160 793143 42166 793195
rect 42218 793183 42224 793195
rect 42832 793183 42838 793195
rect 42218 793155 42838 793183
rect 42218 793143 42224 793155
rect 42832 793143 42838 793155
rect 42890 793143 42896 793195
rect 43024 793069 43030 793121
rect 43082 793069 43088 793121
rect 42832 792995 42838 793047
rect 42890 793035 42896 793047
rect 43042 793035 43070 793069
rect 42890 793007 43070 793035
rect 42890 792995 42896 793007
rect 42736 792921 42742 792973
rect 42794 792961 42800 792973
rect 43024 792961 43030 792973
rect 42794 792933 43030 792961
rect 42794 792921 42800 792933
rect 43024 792921 43030 792933
rect 43082 792921 43088 792973
rect 42256 792107 42262 792159
rect 42314 792147 42320 792159
rect 43120 792147 43126 792159
rect 42314 792119 43126 792147
rect 42314 792107 42320 792119
rect 43120 792107 43126 792119
rect 43178 792107 43184 792159
rect 42160 791959 42166 792011
rect 42218 791999 42224 792011
rect 42448 791999 42454 792011
rect 42218 791971 42454 791999
rect 42218 791959 42224 791971
rect 42448 791959 42454 791971
rect 42506 791959 42512 792011
rect 43120 791959 43126 792011
rect 43178 791999 43184 792011
rect 43504 791999 43510 792011
rect 43178 791971 43510 791999
rect 43178 791959 43184 791971
rect 43504 791959 43510 791971
rect 43562 791959 43568 792011
rect 674704 791959 674710 792011
rect 674762 791999 674768 792011
rect 674896 791999 674902 792011
rect 674762 791971 674902 791999
rect 674762 791959 674768 791971
rect 674896 791959 674902 791971
rect 674954 791959 674960 792011
rect 42256 790109 42262 790161
rect 42314 790149 42320 790161
rect 42832 790149 42838 790161
rect 42314 790121 42838 790149
rect 42314 790109 42320 790121
rect 42832 790109 42838 790121
rect 42890 790109 42896 790161
rect 42160 789887 42166 789939
rect 42218 789927 42224 789939
rect 43024 789927 43030 789939
rect 42218 789899 43030 789927
rect 42218 789887 42224 789899
rect 43024 789887 43030 789899
rect 43082 789887 43088 789939
rect 42160 789443 42166 789495
rect 42218 789483 42224 789495
rect 42928 789483 42934 789495
rect 42218 789455 42934 789483
rect 42218 789443 42224 789455
rect 42928 789443 42934 789455
rect 42986 789443 42992 789495
rect 42160 787001 42166 787053
rect 42218 787041 42224 787053
rect 43120 787041 43126 787053
rect 42218 787013 43126 787041
rect 42218 787001 42224 787013
rect 43120 787001 43126 787013
rect 43178 787001 43184 787053
rect 42160 786409 42166 786461
rect 42218 786449 42224 786461
rect 42736 786449 42742 786461
rect 42218 786421 42742 786449
rect 42218 786409 42224 786421
rect 42736 786409 42742 786421
rect 42794 786409 42800 786461
rect 654448 786261 654454 786313
rect 654506 786301 654512 786313
rect 669712 786301 669718 786313
rect 654506 786273 669718 786301
rect 654506 786261 654512 786273
rect 669712 786261 669718 786273
rect 669770 786261 669776 786313
rect 42064 785743 42070 785795
rect 42122 785783 42128 785795
rect 42448 785783 42454 785795
rect 42122 785755 42454 785783
rect 42122 785743 42128 785755
rect 42448 785743 42454 785755
rect 42506 785743 42512 785795
rect 674512 784929 674518 784981
rect 674570 784969 674576 784981
rect 675376 784969 675382 784981
rect 674570 784941 675382 784969
rect 674570 784929 674576 784941
rect 675376 784929 675382 784941
rect 675434 784929 675440 784981
rect 672880 783449 672886 783501
rect 672938 783489 672944 783501
rect 675280 783489 675286 783501
rect 672938 783461 675286 783489
rect 672938 783449 672944 783461
rect 675280 783449 675286 783461
rect 675338 783449 675344 783501
rect 674992 782857 674998 782909
rect 675050 782897 675056 782909
rect 675280 782897 675286 782909
rect 675050 782869 675286 782897
rect 675050 782857 675056 782869
rect 675280 782857 675286 782869
rect 675338 782857 675344 782909
rect 672784 782191 672790 782243
rect 672842 782231 672848 782243
rect 674608 782231 674614 782243
rect 672842 782203 674614 782231
rect 672842 782191 672848 782203
rect 674608 782191 674614 782203
rect 674666 782231 674672 782243
rect 675280 782231 675286 782243
rect 674666 782203 675286 782231
rect 674666 782191 674672 782203
rect 675280 782191 675286 782203
rect 675338 782191 675344 782243
rect 663856 780563 663862 780615
rect 663914 780603 663920 780615
rect 675088 780603 675094 780615
rect 663914 780575 675094 780603
rect 663914 780563 663920 780575
rect 675088 780563 675094 780575
rect 675146 780563 675152 780615
rect 42736 780415 42742 780467
rect 42794 780455 42800 780467
rect 50608 780455 50614 780467
rect 42794 780427 50614 780455
rect 42794 780415 42800 780427
rect 50608 780415 50614 780427
rect 50666 780415 50672 780467
rect 674896 780415 674902 780467
rect 674954 780455 674960 780467
rect 675472 780455 675478 780467
rect 674954 780427 675478 780455
rect 674954 780415 674960 780427
rect 675472 780415 675478 780427
rect 675530 780415 675536 780467
rect 42448 779897 42454 779949
rect 42506 779937 42512 779949
rect 47536 779937 47542 779949
rect 42506 779909 47542 779937
rect 42506 779897 42512 779909
rect 47536 779897 47542 779909
rect 47594 779897 47600 779949
rect 672496 779749 672502 779801
rect 672554 779789 672560 779801
rect 675376 779789 675382 779801
rect 672554 779761 675382 779789
rect 672554 779749 672560 779761
rect 675376 779749 675382 779761
rect 675434 779749 675440 779801
rect 672208 779305 672214 779357
rect 672266 779345 672272 779357
rect 675472 779345 675478 779357
rect 672266 779317 675478 779345
rect 672266 779305 672272 779317
rect 675472 779305 675478 779317
rect 675530 779305 675536 779357
rect 42736 778861 42742 778913
rect 42794 778901 42800 778913
rect 53392 778901 53398 778913
rect 42794 778873 53398 778901
rect 42794 778861 42800 778873
rect 53392 778861 53398 778873
rect 53450 778861 53456 778913
rect 672592 778565 672598 778617
rect 672650 778605 672656 778617
rect 675376 778605 675382 778617
rect 672650 778577 675382 778605
rect 672650 778565 672656 778577
rect 675376 778565 675382 778577
rect 675434 778565 675440 778617
rect 672016 777603 672022 777655
rect 672074 777643 672080 777655
rect 675472 777643 675478 777655
rect 672074 777615 675478 777643
rect 672074 777603 672080 777615
rect 675472 777603 675478 777615
rect 675530 777603 675536 777655
rect 675088 777011 675094 777063
rect 675146 777051 675152 777063
rect 675376 777051 675382 777063
rect 675146 777023 675382 777051
rect 675146 777011 675152 777023
rect 675376 777011 675382 777023
rect 675434 777011 675440 777063
rect 674224 775457 674230 775509
rect 674282 775497 674288 775509
rect 675376 775497 675382 775509
rect 674282 775469 675382 775497
rect 674282 775457 674288 775469
rect 675376 775457 675382 775469
rect 675434 775457 675440 775509
rect 654448 774717 654454 774769
rect 654506 774757 654512 774769
rect 669808 774757 669814 774769
rect 654506 774729 669814 774757
rect 654506 774717 654512 774729
rect 669808 774717 669814 774729
rect 669866 774717 669872 774769
rect 674320 773607 674326 773659
rect 674378 773647 674384 773659
rect 675376 773647 675382 773659
rect 674378 773619 675382 773647
rect 674378 773607 674384 773619
rect 675376 773607 675382 773619
rect 675434 773607 675440 773659
rect 53392 771831 53398 771883
rect 53450 771871 53456 771883
rect 59536 771871 59542 771883
rect 53450 771843 59542 771871
rect 53450 771831 53456 771843
rect 59536 771831 59542 771843
rect 59594 771831 59600 771883
rect 660976 767465 660982 767517
rect 661034 767505 661040 767517
rect 674416 767505 674422 767517
rect 661034 767477 674422 767505
rect 661034 767465 661040 767477
rect 674416 767465 674422 767477
rect 674474 767465 674480 767517
rect 666736 766873 666742 766925
rect 666794 766913 666800 766925
rect 674704 766913 674710 766925
rect 666794 766885 674710 766913
rect 666794 766873 666800 766885
rect 674704 766873 674710 766885
rect 674762 766873 674768 766925
rect 663952 765837 663958 765889
rect 664010 765877 664016 765889
rect 674416 765877 674422 765889
rect 664010 765849 674422 765877
rect 664010 765837 664016 765849
rect 674416 765837 674422 765849
rect 674474 765837 674480 765889
rect 672304 765245 672310 765297
rect 672362 765285 672368 765297
rect 674704 765285 674710 765297
rect 672362 765257 674710 765285
rect 672362 765245 672368 765257
rect 674704 765245 674710 765257
rect 674762 765245 674768 765297
rect 654448 763247 654454 763299
rect 654506 763287 654512 763299
rect 661072 763287 661078 763299
rect 654506 763259 661078 763287
rect 654506 763247 654512 763259
rect 661072 763247 661078 763259
rect 661130 763247 661136 763299
rect 672688 763247 672694 763299
rect 672746 763287 672752 763299
rect 674704 763287 674710 763299
rect 672746 763259 674710 763287
rect 672746 763247 672752 763259
rect 674704 763247 674710 763259
rect 674762 763247 674768 763299
rect 672400 762507 672406 762559
rect 672458 762547 672464 762559
rect 674704 762547 674710 762559
rect 672458 762519 674710 762547
rect 672458 762507 672464 762519
rect 674704 762507 674710 762519
rect 674762 762507 674768 762559
rect 42736 762211 42742 762263
rect 42794 762251 42800 762263
rect 44848 762251 44854 762263
rect 42794 762223 44854 762251
rect 42794 762211 42800 762223
rect 44848 762211 44854 762223
rect 44906 762211 44912 762263
rect 38992 760287 38998 760339
rect 39050 760327 39056 760339
rect 42736 760327 42742 760339
rect 39050 760299 42742 760327
rect 39050 760287 39056 760299
rect 42736 760287 42742 760299
rect 42794 760287 42800 760339
rect 43120 759325 43126 759377
rect 43178 759365 43184 759377
rect 43408 759365 43414 759377
rect 43178 759337 43414 759365
rect 43178 759325 43184 759337
rect 43408 759325 43414 759337
rect 43466 759325 43472 759377
rect 43024 757771 43030 757823
rect 43082 757811 43088 757823
rect 44944 757811 44950 757823
rect 43082 757783 44950 757811
rect 43082 757771 43088 757783
rect 44944 757771 44950 757783
rect 45002 757771 45008 757823
rect 50416 757475 50422 757527
rect 50474 757515 50480 757527
rect 59536 757515 59542 757527
rect 50474 757487 59542 757515
rect 50474 757475 50480 757487
rect 59536 757475 59542 757487
rect 59594 757475 59600 757527
rect 42448 757253 42454 757305
rect 42506 757293 42512 757305
rect 43600 757293 43606 757305
rect 42506 757265 43606 757293
rect 42506 757253 42512 757265
rect 43600 757253 43606 757265
rect 43658 757253 43664 757305
rect 41968 757105 41974 757157
rect 42026 757145 42032 757157
rect 43792 757145 43798 757157
rect 42026 757117 43798 757145
rect 42026 757105 42032 757117
rect 43792 757105 43798 757117
rect 43850 757105 43856 757157
rect 42064 757031 42070 757083
rect 42122 757071 42128 757083
rect 43504 757071 43510 757083
rect 42122 757043 43510 757071
rect 42122 757031 42128 757043
rect 43504 757031 43510 757043
rect 43562 757031 43568 757083
rect 41776 756957 41782 757009
rect 41834 756957 41840 757009
rect 41872 756957 41878 757009
rect 41930 756957 41936 757009
rect 41794 756787 41822 756957
rect 41890 756923 41918 756957
rect 43696 756923 43702 756935
rect 41890 756895 43702 756923
rect 43696 756883 43702 756895
rect 43754 756883 43760 756935
rect 41776 756735 41782 756787
rect 41834 756735 41840 756787
rect 42064 754885 42070 754937
rect 42122 754925 42128 754937
rect 42736 754925 42742 754937
rect 42122 754897 42742 754925
rect 42122 754885 42128 754897
rect 42736 754885 42742 754897
rect 42794 754885 42800 754937
rect 42448 754293 42454 754345
rect 42506 754333 42512 754345
rect 42928 754333 42934 754345
rect 42506 754305 42934 754333
rect 42506 754293 42512 754305
rect 42928 754293 42934 754305
rect 42986 754293 42992 754345
rect 42160 754071 42166 754123
rect 42218 754111 42224 754123
rect 43024 754111 43030 754123
rect 42218 754083 43030 754111
rect 42218 754071 42224 754083
rect 43024 754071 43030 754083
rect 43082 754071 43088 754123
rect 42064 753035 42070 753087
rect 42122 753075 42128 753087
rect 43408 753075 43414 753087
rect 42122 753047 43414 753075
rect 42122 753035 42128 753047
rect 43408 753035 43414 753047
rect 43466 753035 43472 753087
rect 43216 752221 43222 752273
rect 43274 752261 43280 752273
rect 43600 752261 43606 752273
rect 43274 752233 43606 752261
rect 43274 752221 43280 752233
rect 43600 752221 43606 752233
rect 43658 752221 43664 752273
rect 43120 751851 43126 751903
rect 43178 751851 43184 751903
rect 42928 751777 42934 751829
rect 42986 751817 42992 751829
rect 43138 751817 43166 751851
rect 42986 751789 43166 751817
rect 42986 751777 42992 751789
rect 43120 751629 43126 751681
rect 43178 751669 43184 751681
rect 43408 751669 43414 751681
rect 43178 751641 43414 751669
rect 43178 751629 43184 751641
rect 43408 751629 43414 751641
rect 43466 751629 43472 751681
rect 42064 751185 42070 751237
rect 42122 751225 42128 751237
rect 42928 751225 42934 751237
rect 42122 751197 42934 751225
rect 42122 751185 42128 751197
rect 42928 751185 42934 751197
rect 42986 751185 42992 751237
rect 42736 750963 42742 751015
rect 42794 751003 42800 751015
rect 43600 751003 43606 751015
rect 42794 750975 43606 751003
rect 42794 750963 42800 750975
rect 43600 750963 43606 750975
rect 43658 750963 43664 751015
rect 42160 750371 42166 750423
rect 42218 750411 42224 750423
rect 43120 750411 43126 750423
rect 42218 750383 43126 750411
rect 42218 750371 42224 750383
rect 43120 750371 43126 750383
rect 43178 750371 43184 750423
rect 43120 750223 43126 750275
rect 43178 750263 43184 750275
rect 43504 750263 43510 750275
rect 43178 750235 43510 750263
rect 43178 750223 43184 750235
rect 43504 750223 43510 750235
rect 43562 750223 43568 750275
rect 42064 749927 42070 749979
rect 42122 749967 42128 749979
rect 43024 749967 43030 749979
rect 42122 749939 43030 749967
rect 42122 749927 42128 749939
rect 43024 749927 43030 749939
rect 43082 749927 43088 749979
rect 42256 748891 42262 748943
rect 42314 748931 42320 748943
rect 42736 748931 42742 748943
rect 42314 748903 42742 748931
rect 42314 748891 42320 748903
rect 42736 748891 42742 748903
rect 42794 748891 42800 748943
rect 649648 748817 649654 748869
rect 649706 748857 649712 748869
rect 679696 748857 679702 748869
rect 649706 748829 679702 748857
rect 649706 748817 649712 748829
rect 679696 748817 679702 748829
rect 679754 748817 679760 748869
rect 42064 746079 42070 746131
rect 42122 746119 42128 746131
rect 43120 746119 43126 746131
rect 42122 746091 43126 746119
rect 42122 746079 42128 746091
rect 43120 746079 43126 746091
rect 43178 746079 43184 746131
rect 672784 745931 672790 745983
rect 672842 745971 672848 745983
rect 674992 745971 674998 745983
rect 672842 745943 674998 745971
rect 672842 745931 672848 745943
rect 674992 745931 674998 745943
rect 675050 745931 675056 745983
rect 674704 745857 674710 745909
rect 674762 745897 674768 745909
rect 674896 745897 674902 745909
rect 674762 745869 674902 745897
rect 674762 745857 674768 745869
rect 674896 745857 674902 745869
rect 674954 745857 674960 745909
rect 42160 745635 42166 745687
rect 42218 745675 42224 745687
rect 42448 745675 42454 745687
rect 42218 745647 42454 745675
rect 42218 745635 42224 745647
rect 42448 745635 42454 745647
rect 42506 745635 42512 745687
rect 42160 743785 42166 743837
rect 42218 743825 42224 743837
rect 42832 743825 42838 743837
rect 42218 743797 42838 743825
rect 42218 743785 42224 743797
rect 42832 743785 42838 743797
rect 42890 743785 42896 743837
rect 42064 743045 42070 743097
rect 42122 743085 42128 743097
rect 42928 743085 42934 743097
rect 42122 743057 42934 743085
rect 42122 743045 42128 743057
rect 42928 743045 42934 743057
rect 42986 743045 42992 743097
rect 47536 743045 47542 743097
rect 47594 743085 47600 743097
rect 59536 743085 59542 743097
rect 47594 743057 59542 743085
rect 47594 743045 47600 743057
rect 59536 743045 59542 743057
rect 59594 743045 59600 743097
rect 42160 742601 42166 742653
rect 42218 742641 42224 742653
rect 42736 742641 42742 742653
rect 42218 742613 42742 742641
rect 42218 742601 42224 742613
rect 42736 742601 42742 742613
rect 42794 742601 42800 742653
rect 674032 741565 674038 741617
rect 674090 741605 674096 741617
rect 674416 741605 674422 741617
rect 674090 741577 674422 741605
rect 674090 741565 674096 741577
rect 674416 741565 674422 741577
rect 674474 741565 674480 741617
rect 672304 738087 672310 738139
rect 672362 738127 672368 738139
rect 674992 738127 674998 738139
rect 672362 738099 674998 738127
rect 672362 738087 672368 738099
rect 674992 738087 674998 738099
rect 675050 738127 675056 738139
rect 675472 738127 675478 738139
rect 675050 738099 675478 738127
rect 675050 738087 675056 738099
rect 675472 738087 675478 738099
rect 675530 738087 675536 738139
rect 674896 738013 674902 738065
rect 674954 738053 674960 738065
rect 674954 738025 675038 738053
rect 674954 738013 674960 738025
rect 675010 737991 675038 738025
rect 674992 737939 674998 737991
rect 675050 737939 675056 737991
rect 674896 737865 674902 737917
rect 674954 737905 674960 737917
rect 675376 737905 675382 737917
rect 674954 737877 675382 737905
rect 674954 737865 674960 737877
rect 675376 737865 675382 737877
rect 675434 737865 675440 737917
rect 660976 737347 660982 737399
rect 661034 737387 661040 737399
rect 675184 737387 675190 737399
rect 661034 737359 675190 737387
rect 661034 737347 661040 737359
rect 675184 737347 675190 737359
rect 675242 737347 675248 737399
rect 654448 737273 654454 737325
rect 654506 737313 654512 737325
rect 663952 737313 663958 737325
rect 654506 737285 663958 737313
rect 654506 737273 654512 737285
rect 663952 737273 663958 737285
rect 664010 737273 664016 737325
rect 42640 737199 42646 737251
rect 42698 737239 42704 737251
rect 53392 737239 53398 737251
rect 42698 737211 53398 737239
rect 42698 737199 42704 737211
rect 53392 737199 53398 737211
rect 53450 737199 53456 737251
rect 42352 736681 42358 736733
rect 42410 736721 42416 736733
rect 50416 736721 50422 736733
rect 42410 736693 50422 736721
rect 42410 736681 42416 736693
rect 50416 736681 50422 736693
rect 50474 736681 50480 736733
rect 674512 735645 674518 735697
rect 674570 735685 674576 735697
rect 675472 735685 675478 735697
rect 674570 735657 675478 735685
rect 674570 735645 674576 735657
rect 675472 735645 675478 735657
rect 675530 735645 675536 735697
rect 42352 735423 42358 735475
rect 42410 735463 42416 735475
rect 58960 735463 58966 735475
rect 42410 735435 58966 735463
rect 42410 735423 42416 735435
rect 58960 735423 58966 735435
rect 59018 735423 59024 735475
rect 672112 733573 672118 733625
rect 672170 733613 672176 733625
rect 675472 733613 675478 733625
rect 672170 733585 675478 733613
rect 672170 733573 672176 733585
rect 675472 733573 675478 733585
rect 675530 733573 675536 733625
rect 674128 732315 674134 732367
rect 674186 732355 674192 732367
rect 675472 732355 675478 732367
rect 674186 732327 675478 732355
rect 674186 732315 674192 732327
rect 675472 732315 675478 732327
rect 675530 732315 675536 732367
rect 675184 732019 675190 732071
rect 675242 732059 675248 732071
rect 675376 732059 675382 732071
rect 675242 732031 675382 732059
rect 675242 732019 675248 732031
rect 675376 732019 675382 732031
rect 675434 732019 675440 732071
rect 674704 730465 674710 730517
rect 674762 730505 674768 730517
rect 675472 730505 675478 730517
rect 674762 730477 675478 730505
rect 674762 730465 674768 730477
rect 675472 730465 675478 730477
rect 675530 730465 675536 730517
rect 50416 728615 50422 728667
rect 50474 728655 50480 728667
rect 58384 728655 58390 728667
rect 50474 728627 58390 728655
rect 50474 728615 50480 728627
rect 58384 728615 58390 728627
rect 58442 728615 58448 728667
rect 674608 728615 674614 728667
rect 674666 728655 674672 728667
rect 675472 728655 675478 728667
rect 674666 728627 675478 728655
rect 674666 728615 674672 728627
rect 675472 728615 675478 728627
rect 675530 728615 675536 728667
rect 669616 722473 669622 722525
rect 669674 722513 669680 722525
rect 674416 722513 674422 722525
rect 669674 722485 674422 722513
rect 669674 722473 669680 722485
rect 674416 722473 674422 722485
rect 674474 722473 674480 722525
rect 660880 721733 660886 721785
rect 660938 721773 660944 721785
rect 674416 721773 674422 721785
rect 660938 721745 674422 721773
rect 660938 721733 660944 721745
rect 674416 721733 674422 721745
rect 674474 721733 674480 721785
rect 661168 720845 661174 720897
rect 661226 720885 661232 720897
rect 674416 720885 674422 720897
rect 661226 720857 674422 720885
rect 661226 720845 661232 720857
rect 674416 720845 674422 720857
rect 674474 720845 674480 720897
rect 671920 719143 671926 719195
rect 671978 719183 671984 719195
rect 674416 719183 674422 719195
rect 671978 719155 674422 719183
rect 671978 719143 671984 719155
rect 674416 719143 674422 719155
rect 674474 719143 674480 719195
rect 672400 717663 672406 717715
rect 672458 717703 672464 717715
rect 674416 717703 674422 717715
rect 672458 717675 674422 717703
rect 672458 717663 672464 717675
rect 674416 717663 674422 717675
rect 674474 717663 674480 717715
rect 43312 717219 43318 717271
rect 43370 717259 43376 717271
rect 44944 717259 44950 717271
rect 43370 717231 44950 717259
rect 43370 717219 43376 717231
rect 44944 717219 44950 717231
rect 45002 717219 45008 717271
rect 40144 715887 40150 715939
rect 40202 715927 40208 715939
rect 41872 715927 41878 715939
rect 40202 715899 41878 715927
rect 40202 715887 40208 715899
rect 41872 715887 41878 715899
rect 41930 715887 41936 715939
rect 672688 715295 672694 715347
rect 672746 715335 672752 715347
rect 673648 715335 673654 715347
rect 672746 715307 673654 715335
rect 672746 715295 672752 715307
rect 673648 715295 673654 715307
rect 673706 715295 673712 715347
rect 53392 714259 53398 714311
rect 53450 714299 53456 714311
rect 58384 714299 58390 714311
rect 53450 714271 58390 714299
rect 53450 714259 53456 714271
rect 58384 714259 58390 714271
rect 58442 714259 58448 714311
rect 654448 714259 654454 714311
rect 654506 714299 654512 714311
rect 666928 714299 666934 714311
rect 654506 714271 666934 714299
rect 654506 714259 654512 714271
rect 666928 714259 666934 714271
rect 666986 714259 666992 714311
rect 41584 714037 41590 714089
rect 41642 714037 41648 714089
rect 41680 714037 41686 714089
rect 41738 714077 41744 714089
rect 43504 714077 43510 714089
rect 41738 714049 43510 714077
rect 41738 714037 41744 714049
rect 43504 714037 43510 714049
rect 43562 714037 43568 714089
rect 41602 713559 41630 714037
rect 41776 713963 41782 714015
rect 41834 714003 41840 714015
rect 43600 714003 43606 714015
rect 41834 713975 43606 714003
rect 41834 713963 41840 713975
rect 43600 713963 43606 713975
rect 43658 713963 43664 714015
rect 41776 713559 41782 713571
rect 41602 713531 41782 713559
rect 41776 713519 41782 713531
rect 41834 713519 41840 713571
rect 42928 711743 42934 711795
rect 42986 711783 42992 711795
rect 42986 711755 43550 711783
rect 42986 711743 42992 711755
rect 43522 711425 43550 711755
rect 43504 711373 43510 711425
rect 43562 711373 43568 711425
rect 43216 711225 43222 711277
rect 43274 711265 43280 711277
rect 43696 711265 43702 711277
rect 43274 711237 43702 711265
rect 43274 711225 43280 711237
rect 43696 711225 43702 711237
rect 43754 711225 43760 711277
rect 42160 710781 42166 710833
rect 42218 710821 42224 710833
rect 45136 710821 45142 710833
rect 42218 710793 45142 710821
rect 42218 710781 42224 710793
rect 45136 710781 45142 710793
rect 45194 710781 45200 710833
rect 672880 710485 672886 710537
rect 672938 710525 672944 710537
rect 674416 710525 674422 710537
rect 672938 710497 674422 710525
rect 672938 710485 672944 710497
rect 674416 710485 674422 710497
rect 674474 710485 674480 710537
rect 42160 709893 42166 709945
rect 42218 709933 42224 709945
rect 42352 709933 42358 709945
rect 42218 709905 42358 709933
rect 42218 709893 42224 709905
rect 42352 709893 42358 709905
rect 42410 709893 42416 709945
rect 672016 709893 672022 709945
rect 672074 709933 672080 709945
rect 674800 709933 674806 709945
rect 672074 709905 674806 709933
rect 672074 709893 672080 709905
rect 674800 709893 674806 709905
rect 674858 709893 674864 709945
rect 672208 709005 672214 709057
rect 672266 709045 672272 709057
rect 674416 709045 674422 709057
rect 672266 709017 674422 709045
rect 672266 709005 672272 709017
rect 674416 709005 674422 709017
rect 674474 709005 674480 709057
rect 42544 707895 42550 707947
rect 42602 707935 42608 707947
rect 43408 707935 43414 707947
rect 42602 707907 43414 707935
rect 42602 707895 42608 707907
rect 43408 707895 43414 707907
rect 43466 707895 43472 707947
rect 42160 707377 42166 707429
rect 42218 707417 42224 707429
rect 43024 707417 43030 707429
rect 42218 707389 43030 707417
rect 42218 707377 42224 707389
rect 43024 707377 43030 707389
rect 43082 707377 43088 707429
rect 672496 707377 672502 707429
rect 672554 707417 672560 707429
rect 674416 707417 674422 707429
rect 672554 707389 674422 707417
rect 672554 707377 672560 707389
rect 674416 707377 674422 707389
rect 674474 707377 674480 707429
rect 43024 707229 43030 707281
rect 43082 707269 43088 707281
rect 43600 707269 43606 707281
rect 43082 707241 43606 707269
rect 43082 707229 43088 707241
rect 43600 707229 43606 707241
rect 43658 707229 43664 707281
rect 672592 706785 672598 706837
rect 672650 706825 672656 706837
rect 674800 706825 674806 706837
rect 672650 706797 674806 706825
rect 672650 706785 672656 706797
rect 674800 706785 674806 706797
rect 674858 706785 674864 706837
rect 42928 706415 42934 706467
rect 42986 706455 42992 706467
rect 43504 706455 43510 706467
rect 42986 706427 43510 706455
rect 42986 706415 42992 706427
rect 43504 706415 43510 706427
rect 43562 706415 43568 706467
rect 42160 705823 42166 705875
rect 42218 705823 42224 705875
rect 42178 705641 42206 705823
rect 42256 705641 42262 705653
rect 42178 705613 42262 705641
rect 42256 705601 42262 705613
rect 42314 705601 42320 705653
rect 42832 703643 42838 703655
rect 42082 703615 42838 703643
rect 42082 703581 42110 703615
rect 42832 703603 42838 703615
rect 42890 703603 42896 703655
rect 42064 703529 42070 703581
rect 42122 703529 42128 703581
rect 42160 702863 42166 702915
rect 42218 702903 42224 702915
rect 43024 702903 43030 702915
rect 42218 702875 43030 702903
rect 42218 702863 42224 702875
rect 43024 702863 43030 702875
rect 43082 702863 43088 702915
rect 649744 702715 649750 702767
rect 649802 702755 649808 702767
rect 679696 702755 679702 702767
rect 649802 702727 679702 702755
rect 649802 702715 649808 702727
rect 679696 702715 679702 702727
rect 679754 702715 679760 702767
rect 42160 702271 42166 702323
rect 42218 702311 42224 702323
rect 42544 702311 42550 702323
rect 42218 702283 42550 702311
rect 42218 702271 42224 702283
rect 42544 702271 42550 702283
rect 42602 702271 42608 702323
rect 42064 700569 42070 700621
rect 42122 700609 42128 700621
rect 42928 700609 42934 700621
rect 42122 700581 42934 700609
rect 42122 700569 42128 700581
rect 42928 700569 42934 700581
rect 42986 700569 42992 700621
rect 42160 700051 42166 700103
rect 42218 700091 42224 700103
rect 42832 700091 42838 700103
rect 42218 700063 42838 700091
rect 42218 700051 42224 700063
rect 42832 700051 42838 700063
rect 42890 700051 42896 700103
rect 42352 699829 42358 699881
rect 42410 699869 42416 699881
rect 57808 699869 57814 699881
rect 42410 699841 57814 699869
rect 42410 699829 42416 699841
rect 57808 699829 57814 699841
rect 57866 699829 57872 699881
rect 672304 699829 672310 699881
rect 672362 699869 672368 699881
rect 672592 699869 672598 699881
rect 672362 699841 672598 699869
rect 672362 699829 672368 699841
rect 672592 699829 672598 699841
rect 672650 699829 672656 699881
rect 42640 693983 42646 694035
rect 42698 694023 42704 694035
rect 53392 694023 53398 694035
rect 42698 693995 53398 694023
rect 42698 693983 42704 693995
rect 53392 693983 53398 693995
rect 53450 693983 53456 694035
rect 672208 692873 672214 692925
rect 672266 692913 672272 692925
rect 675376 692913 675382 692925
rect 672266 692885 675382 692913
rect 672266 692873 672272 692885
rect 675376 692873 675382 692885
rect 675434 692873 675440 692925
rect 672592 692651 672598 692703
rect 672650 692691 672656 692703
rect 675472 692691 675478 692703
rect 672650 692663 675478 692691
rect 672650 692651 672656 692663
rect 675472 692651 675478 692663
rect 675530 692651 675536 692703
rect 42640 692429 42646 692481
rect 42698 692469 42704 692481
rect 50416 692469 50422 692481
rect 42698 692441 50422 692469
rect 42698 692429 42704 692441
rect 50416 692429 50422 692441
rect 50474 692429 50480 692481
rect 654448 691245 654454 691297
rect 654506 691285 654512 691297
rect 661264 691285 661270 691297
rect 654506 691257 661270 691285
rect 654506 691245 654512 691257
rect 661264 691245 661270 691257
rect 661322 691245 661328 691297
rect 674320 690653 674326 690705
rect 674378 690693 674384 690705
rect 675472 690693 675478 690705
rect 674378 690665 675478 690693
rect 674378 690653 674384 690665
rect 675472 690653 675478 690665
rect 675530 690653 675536 690705
rect 675088 689765 675094 689817
rect 675146 689805 675152 689817
rect 675376 689805 675382 689817
rect 675146 689777 675382 689805
rect 675146 689765 675152 689777
rect 675376 689765 675382 689777
rect 675434 689765 675440 689817
rect 674416 689321 674422 689373
rect 674474 689361 674480 689373
rect 675376 689361 675382 689373
rect 674474 689333 675382 689361
rect 674474 689321 674480 689333
rect 675376 689321 675382 689333
rect 675434 689321 675440 689373
rect 672016 688581 672022 688633
rect 672074 688621 672080 688633
rect 675472 688621 675478 688633
rect 672074 688593 675478 688621
rect 672074 688581 672080 688593
rect 675472 688581 675478 688593
rect 675530 688581 675536 688633
rect 674224 687323 674230 687375
rect 674282 687363 674288 687375
rect 675472 687363 675478 687375
rect 674282 687335 675478 687363
rect 674282 687323 674288 687335
rect 675472 687323 675478 687335
rect 675530 687323 675536 687375
rect 669616 686213 669622 686265
rect 669674 686253 669680 686265
rect 675376 686253 675382 686265
rect 669674 686225 675382 686253
rect 669674 686213 669680 686225
rect 675376 686213 675382 686225
rect 675434 686213 675440 686265
rect 50416 685473 50422 685525
rect 50474 685513 50480 685525
rect 59536 685513 59542 685525
rect 50474 685485 59542 685513
rect 50474 685473 50480 685485
rect 59536 685473 59542 685485
rect 59594 685473 59600 685525
rect 674800 685473 674806 685525
rect 674858 685513 674864 685525
rect 675472 685513 675478 685525
rect 674858 685485 675478 685513
rect 674858 685473 674864 685485
rect 675472 685473 675478 685485
rect 675530 685473 675536 685525
rect 674896 683623 674902 683675
rect 674954 683663 674960 683675
rect 675472 683663 675478 683675
rect 674954 683635 675478 683663
rect 674954 683623 674960 683635
rect 675472 683623 675478 683635
rect 675530 683623 675536 683675
rect 663760 677333 663766 677385
rect 663818 677373 663824 677385
rect 674416 677373 674422 677385
rect 663818 677345 674422 677373
rect 663818 677333 663824 677345
rect 674416 677333 674422 677345
rect 674474 677333 674480 677385
rect 666832 676445 666838 676497
rect 666890 676485 666896 676497
rect 674416 676485 674422 676497
rect 666890 676457 674422 676485
rect 666890 676445 666896 676457
rect 674416 676445 674422 676457
rect 674474 676445 674480 676497
rect 42736 676337 42742 676349
rect 42658 676309 42742 676337
rect 42658 676053 42686 676309
rect 42736 676297 42742 676309
rect 42794 676297 42800 676349
rect 42640 676001 42646 676053
rect 42698 676001 42704 676053
rect 664048 675705 664054 675757
rect 664106 675745 664112 675757
rect 674416 675745 674422 675757
rect 664106 675717 674422 675745
rect 664106 675705 664112 675717
rect 674416 675705 674422 675717
rect 674474 675705 674480 675757
rect 42352 675631 42358 675683
rect 42410 675671 42416 675683
rect 47728 675671 47734 675683
rect 42410 675643 47734 675671
rect 42410 675631 42416 675643
rect 47728 675631 47734 675643
rect 47786 675631 47792 675683
rect 671920 674817 671926 674869
rect 671978 674857 671984 674869
rect 674416 674857 674422 674869
rect 671978 674829 674422 674857
rect 671978 674817 671984 674829
rect 674416 674817 674422 674829
rect 674474 674817 674480 674869
rect 41872 674521 41878 674573
rect 41930 674561 41936 674573
rect 43120 674561 43126 674573
rect 41930 674533 43126 674561
rect 41930 674521 41936 674533
rect 43120 674521 43126 674533
rect 43178 674521 43184 674573
rect 672496 674003 672502 674055
rect 672554 674043 672560 674055
rect 674416 674043 674422 674055
rect 672554 674015 674422 674043
rect 672554 674003 672560 674015
rect 674416 674003 674422 674015
rect 674474 674003 674480 674055
rect 43312 673781 43318 673833
rect 43370 673821 43376 673833
rect 45040 673821 45046 673833
rect 43370 673793 45046 673821
rect 43370 673781 43376 673793
rect 45040 673781 45046 673793
rect 45098 673781 45104 673833
rect 40240 672375 40246 672427
rect 40298 672415 40304 672427
rect 41872 672415 41878 672427
rect 40298 672387 41878 672415
rect 40298 672375 40304 672387
rect 41872 672375 41878 672387
rect 41930 672375 41936 672427
rect 42064 671931 42070 671983
rect 42122 671971 42128 671983
rect 42448 671971 42454 671983
rect 42122 671943 42454 671971
rect 42122 671931 42128 671943
rect 42448 671931 42454 671943
rect 42506 671931 42512 671983
rect 53392 671043 53398 671095
rect 53450 671083 53456 671095
rect 59440 671083 59446 671095
rect 53450 671055 59446 671083
rect 53450 671043 53456 671055
rect 59440 671043 59446 671055
rect 59498 671043 59504 671095
rect 672400 670969 672406 671021
rect 672458 671009 672464 671021
rect 675184 671009 675190 671021
rect 672458 670981 675190 671009
rect 672458 670969 672464 670981
rect 675184 670969 675190 670981
rect 675242 670969 675248 671021
rect 41296 670895 41302 670947
rect 41354 670935 41360 670947
rect 42928 670935 42934 670947
rect 41354 670907 42934 670935
rect 41354 670895 41360 670907
rect 42928 670895 42934 670907
rect 42986 670895 42992 670947
rect 43216 670895 43222 670947
rect 43274 670935 43280 670947
rect 43600 670935 43606 670947
rect 43274 670907 43606 670935
rect 43274 670895 43280 670907
rect 43600 670895 43606 670907
rect 43658 670895 43664 670947
rect 42256 670747 42262 670799
rect 42314 670787 42320 670799
rect 43408 670787 43414 670799
rect 42314 670759 43414 670787
rect 42314 670747 42320 670759
rect 43408 670747 43414 670759
rect 43466 670747 43472 670799
rect 41968 670673 41974 670725
rect 42026 670713 42032 670725
rect 43120 670713 43126 670725
rect 42026 670685 43126 670713
rect 42026 670673 42032 670685
rect 43120 670673 43126 670685
rect 43178 670673 43184 670725
rect 41776 670599 41782 670651
rect 41834 670599 41840 670651
rect 41872 670599 41878 670651
rect 41930 670599 41936 670651
rect 41794 670355 41822 670599
rect 41890 670565 41918 670599
rect 42928 670565 42934 670577
rect 41890 670537 42934 670565
rect 42928 670525 42934 670537
rect 42986 670525 42992 670577
rect 41776 670303 41782 670355
rect 41834 670303 41840 670355
rect 42160 668527 42166 668579
rect 42218 668567 42224 668579
rect 42928 668567 42934 668579
rect 42218 668539 42934 668567
rect 42218 668527 42224 668539
rect 42928 668527 42934 668539
rect 42986 668527 42992 668579
rect 42928 668379 42934 668431
rect 42986 668419 42992 668431
rect 43216 668419 43222 668431
rect 42986 668391 43222 668419
rect 42986 668379 42992 668391
rect 43216 668379 43222 668391
rect 43274 668379 43280 668431
rect 654448 668157 654454 668209
rect 654506 668197 654512 668209
rect 664048 668197 664054 668209
rect 654506 668169 664054 668197
rect 654506 668157 654512 668169
rect 664048 668157 664054 668169
rect 664106 668157 664112 668209
rect 649840 668083 649846 668135
rect 649898 668123 649904 668135
rect 652240 668123 652246 668135
rect 649898 668095 652246 668123
rect 649898 668083 649904 668095
rect 652240 668083 652246 668095
rect 652298 668083 652304 668135
rect 42160 667861 42166 667913
rect 42218 667901 42224 667913
rect 43312 667901 43318 667913
rect 42218 667873 43318 667901
rect 42218 667861 42224 667873
rect 43312 667861 43318 667873
rect 43370 667861 43376 667913
rect 42160 665345 42166 665397
rect 42218 665385 42224 665397
rect 42928 665385 42934 665397
rect 42218 665357 42934 665385
rect 42218 665345 42224 665357
rect 42928 665345 42934 665357
rect 42986 665345 42992 665397
rect 42928 665197 42934 665249
rect 42986 665237 42992 665249
rect 43408 665237 43414 665249
rect 42986 665209 43414 665237
rect 42986 665197 42992 665209
rect 43408 665197 43414 665209
rect 43466 665197 43472 665249
rect 42160 664827 42166 664879
rect 42218 664867 42224 664879
rect 43024 664867 43030 664879
rect 42218 664839 43030 664867
rect 42218 664827 42224 664839
rect 43024 664827 43030 664839
rect 43082 664827 43088 664879
rect 42064 663939 42070 663991
rect 42122 663979 42128 663991
rect 42544 663979 42550 663991
rect 42122 663951 42550 663979
rect 42122 663939 42128 663951
rect 42544 663939 42550 663951
rect 42602 663939 42608 663991
rect 42160 663347 42166 663399
rect 42218 663387 42224 663399
rect 42544 663387 42550 663399
rect 42218 663359 42550 663387
rect 42218 663347 42224 663359
rect 42544 663347 42550 663359
rect 42602 663347 42608 663399
rect 42256 662385 42262 662437
rect 42314 662425 42320 662437
rect 42928 662425 42934 662437
rect 42314 662397 42934 662425
rect 42314 662385 42320 662397
rect 42928 662385 42934 662397
rect 42986 662385 42992 662437
rect 42928 662237 42934 662289
rect 42986 662277 42992 662289
rect 43600 662277 43606 662289
rect 42986 662249 43606 662277
rect 42986 662237 42992 662249
rect 43600 662237 43606 662249
rect 43658 662237 43664 662289
rect 672112 661349 672118 661401
rect 672170 661389 672176 661401
rect 674416 661389 674422 661401
rect 672170 661361 674422 661389
rect 672170 661349 672176 661361
rect 674416 661349 674422 661361
rect 674474 661349 674480 661401
rect 42064 661053 42070 661105
rect 42122 661093 42128 661105
rect 43120 661093 43126 661105
rect 42122 661065 43126 661093
rect 42122 661053 42128 661065
rect 43120 661053 43126 661065
rect 43178 661053 43184 661105
rect 42160 659869 42166 659921
rect 42218 659909 42224 659921
rect 42832 659909 42838 659921
rect 42218 659881 42838 659909
rect 42218 659869 42224 659881
rect 42832 659869 42838 659881
rect 42890 659869 42896 659921
rect 42064 659055 42070 659107
rect 42122 659095 42128 659107
rect 43024 659095 43030 659107
rect 42122 659067 43030 659095
rect 42122 659055 42128 659067
rect 43024 659055 43030 659067
rect 43082 659055 43088 659107
rect 42160 656835 42166 656887
rect 42218 656875 42224 656887
rect 42928 656875 42934 656887
rect 42218 656847 42934 656875
rect 42218 656835 42224 656847
rect 42928 656835 42934 656847
rect 42986 656835 42992 656887
rect 42832 656687 42838 656739
rect 42890 656727 42896 656739
rect 59536 656727 59542 656739
rect 42890 656699 59542 656727
rect 42890 656687 42896 656699
rect 59536 656687 59542 656699
rect 59594 656687 59600 656739
rect 649840 656687 649846 656739
rect 649898 656727 649904 656739
rect 679696 656727 679702 656739
rect 649898 656699 679702 656727
rect 649898 656687 649904 656699
rect 679696 656687 679702 656699
rect 679754 656687 679760 656739
rect 674416 656095 674422 656147
rect 674474 656135 674480 656147
rect 674896 656135 674902 656147
rect 674474 656107 674902 656135
rect 674474 656095 674480 656107
rect 674896 656095 674902 656107
rect 674954 656095 674960 656147
rect 672592 653727 672598 653779
rect 672650 653767 672656 653779
rect 674992 653767 674998 653779
rect 672650 653739 674998 653767
rect 672650 653727 672656 653739
rect 674992 653727 674998 653739
rect 675050 653727 675056 653779
rect 42448 649731 42454 649783
rect 42506 649771 42512 649783
rect 51856 649771 51862 649783
rect 42506 649743 51862 649771
rect 42506 649731 42512 649743
rect 51856 649731 51862 649743
rect 51914 649731 51920 649783
rect 42448 649509 42454 649561
rect 42506 649549 42512 649561
rect 53392 649549 53398 649561
rect 42506 649521 53398 649549
rect 42506 649509 42512 649521
rect 53392 649509 53398 649521
rect 53450 649509 53456 649561
rect 674896 649509 674902 649561
rect 674954 649549 674960 649561
rect 675184 649549 675190 649561
rect 674954 649521 675190 649549
rect 674954 649509 674960 649521
rect 675184 649509 675190 649521
rect 675242 649509 675248 649561
rect 671920 648251 671926 648303
rect 671978 648291 671984 648303
rect 675280 648291 675286 648303
rect 671978 648263 675286 648291
rect 671978 648251 671984 648263
rect 675280 648251 675286 648263
rect 675338 648251 675344 648303
rect 672880 648029 672886 648081
rect 672938 648069 672944 648081
rect 675280 648069 675286 648081
rect 672938 648041 675286 648069
rect 672938 648029 672944 648041
rect 675280 648029 675286 648041
rect 675338 648029 675344 648081
rect 675088 647807 675094 647859
rect 675146 647807 675152 647859
rect 675106 647563 675134 647807
rect 675088 647511 675094 647563
rect 675146 647511 675152 647563
rect 674512 646401 674518 646453
rect 674570 646441 674576 646453
rect 674896 646441 674902 646453
rect 674570 646413 674902 646441
rect 674570 646401 674576 646413
rect 674896 646401 674902 646413
rect 674954 646441 674960 646453
rect 675376 646441 675382 646453
rect 674954 646413 675382 646441
rect 674954 646401 674960 646413
rect 675376 646401 675382 646413
rect 675434 646401 675440 646453
rect 674608 645291 674614 645343
rect 674666 645331 674672 645343
rect 675184 645331 675190 645343
rect 674666 645303 675190 645331
rect 674666 645291 674672 645303
rect 675184 645291 675190 645303
rect 675242 645291 675248 645343
rect 654448 645217 654454 645269
rect 654506 645257 654512 645269
rect 666832 645257 666838 645269
rect 654506 645229 666838 645257
rect 654506 645217 654512 645229
rect 666832 645217 666838 645229
rect 666890 645217 666896 645269
rect 666736 645143 666742 645195
rect 666794 645183 666800 645195
rect 675184 645183 675190 645195
rect 666794 645155 675190 645183
rect 666794 645143 666800 645155
rect 675184 645143 675190 645155
rect 675242 645143 675248 645195
rect 671632 644773 671638 644825
rect 671690 644813 671696 644825
rect 675376 644813 675382 644825
rect 671690 644785 675382 644813
rect 671690 644773 671696 644785
rect 675376 644773 675382 644785
rect 675434 644773 675440 644825
rect 51856 644477 51862 644529
rect 51914 644517 51920 644529
rect 59248 644517 59254 644529
rect 51914 644489 59254 644517
rect 51914 644477 51920 644489
rect 59248 644477 59254 644489
rect 59306 644477 59312 644529
rect 672304 644033 672310 644085
rect 672362 644073 672368 644085
rect 675472 644073 675478 644085
rect 672362 644045 675478 644073
rect 672362 644033 672368 644045
rect 675472 644033 675478 644045
rect 675530 644033 675536 644085
rect 672592 643367 672598 643419
rect 672650 643407 672656 643419
rect 675376 643407 675382 643419
rect 672650 643379 675382 643407
rect 672650 643367 672656 643379
rect 675376 643367 675382 643379
rect 675434 643367 675440 643419
rect 671440 642257 671446 642309
rect 671498 642297 671504 642309
rect 675472 642297 675478 642309
rect 671498 642269 675478 642297
rect 671498 642257 671504 642269
rect 675472 642257 675478 642269
rect 675530 642257 675536 642309
rect 675184 641813 675190 641865
rect 675242 641853 675248 641865
rect 675376 641853 675382 641865
rect 675242 641825 675382 641853
rect 675242 641813 675248 641825
rect 675376 641813 675382 641825
rect 675434 641813 675440 641865
rect 669808 632489 669814 632541
rect 669866 632529 669872 632541
rect 674704 632529 674710 632541
rect 669866 632501 674710 632529
rect 669866 632489 669872 632501
rect 674704 632489 674710 632501
rect 674762 632489 674768 632541
rect 42448 632415 42454 632467
rect 42506 632455 42512 632467
rect 45040 632455 45046 632467
rect 42506 632427 45046 632455
rect 42506 632415 42512 632427
rect 45040 632415 45046 632427
rect 45098 632415 45104 632467
rect 43120 632119 43126 632171
rect 43178 632159 43184 632171
rect 43696 632159 43702 632171
rect 43178 632131 43702 632159
rect 43178 632119 43184 632131
rect 43696 632119 43702 632131
rect 43754 632119 43760 632171
rect 669712 631749 669718 631801
rect 669770 631789 669776 631801
rect 674704 631789 674710 631801
rect 669770 631761 674710 631789
rect 669770 631749 669776 631761
rect 674704 631749 674710 631761
rect 674762 631749 674768 631801
rect 661072 630565 661078 630617
rect 661130 630605 661136 630617
rect 674128 630605 674134 630617
rect 661130 630577 674134 630605
rect 661130 630565 661136 630577
rect 674128 630565 674134 630577
rect 674186 630565 674192 630617
rect 672496 630269 672502 630321
rect 672554 630309 672560 630321
rect 673840 630309 673846 630321
rect 672554 630281 673846 630309
rect 672554 630269 672560 630281
rect 673840 630269 673846 630281
rect 673898 630269 673904 630321
rect 671728 628419 671734 628471
rect 671786 628459 671792 628471
rect 673840 628459 673846 628471
rect 671786 628431 673846 628459
rect 671786 628419 671792 628431
rect 673840 628419 673846 628431
rect 673898 628419 673904 628471
rect 670960 628123 670966 628175
rect 671018 628163 671024 628175
rect 672688 628163 672694 628175
rect 671018 628135 672694 628163
rect 671018 628123 671024 628135
rect 672688 628123 672694 628135
rect 672746 628163 672752 628175
rect 673840 628163 673846 628175
rect 672746 628135 673846 628163
rect 672746 628123 672752 628135
rect 673840 628123 673846 628135
rect 673898 628123 673904 628175
rect 42448 627901 42454 627953
rect 42506 627941 42512 627953
rect 47824 627941 47830 627953
rect 42506 627913 47830 627941
rect 42506 627901 42512 627913
rect 47824 627901 47830 627913
rect 47882 627901 47888 627953
rect 40048 627827 40054 627879
rect 40106 627867 40112 627879
rect 42928 627867 42934 627879
rect 40106 627839 42934 627867
rect 40106 627827 40112 627839
rect 42928 627827 42934 627839
rect 42986 627827 42992 627879
rect 47632 627827 47638 627879
rect 47690 627867 47696 627879
rect 58000 627867 58006 627879
rect 47690 627839 58006 627867
rect 47690 627827 47696 627839
rect 58000 627827 58006 627839
rect 58058 627827 58064 627879
rect 670864 627753 670870 627805
rect 670922 627793 670928 627805
rect 675184 627793 675190 627805
rect 670922 627765 675190 627793
rect 670922 627753 670928 627765
rect 675184 627753 675190 627765
rect 675242 627753 675248 627805
rect 41488 627679 41494 627731
rect 41546 627719 41552 627731
rect 43120 627719 43126 627731
rect 41546 627691 43126 627719
rect 41546 627679 41552 627691
rect 43120 627679 43126 627691
rect 43178 627679 43184 627731
rect 42640 627605 42646 627657
rect 42698 627645 42704 627657
rect 43312 627645 43318 627657
rect 42698 627617 43318 627645
rect 42698 627605 42704 627617
rect 43312 627605 43318 627617
rect 43370 627605 43376 627657
rect 43024 627531 43030 627583
rect 43082 627571 43088 627583
rect 43408 627571 43414 627583
rect 43082 627543 43414 627571
rect 43082 627531 43088 627543
rect 43408 627531 43414 627543
rect 43466 627531 43472 627583
rect 41776 627383 41782 627435
rect 41834 627383 41840 627435
rect 41968 627383 41974 627435
rect 42026 627383 42032 627435
rect 42064 627383 42070 627435
rect 42122 627423 42128 627435
rect 43024 627423 43030 627435
rect 42122 627395 43030 627423
rect 42122 627383 42128 627395
rect 43024 627383 43030 627395
rect 43082 627383 43088 627435
rect 41794 627213 41822 627383
rect 41986 627349 42014 627383
rect 43504 627349 43510 627361
rect 41986 627321 43510 627349
rect 43504 627309 43510 627321
rect 43562 627309 43568 627361
rect 41776 627161 41782 627213
rect 41834 627161 41840 627213
rect 42160 625311 42166 625363
rect 42218 625351 42224 625363
rect 42928 625351 42934 625363
rect 42218 625323 42934 625351
rect 42218 625311 42224 625323
rect 42928 625311 42934 625323
rect 42986 625311 42992 625363
rect 42928 625163 42934 625215
rect 42986 625203 42992 625215
rect 43312 625203 43318 625215
rect 42986 625175 43318 625203
rect 42986 625163 42992 625175
rect 43312 625163 43318 625175
rect 43370 625163 43376 625215
rect 674608 624867 674614 624919
rect 674666 624907 674672 624919
rect 674896 624907 674902 624919
rect 674666 624879 674902 624907
rect 674666 624867 674672 624879
rect 674896 624867 674902 624879
rect 674954 624867 674960 624919
rect 42160 624645 42166 624697
rect 42218 624685 42224 624697
rect 42448 624685 42454 624697
rect 42218 624657 42454 624685
rect 42218 624645 42224 624657
rect 42448 624645 42454 624657
rect 42506 624645 42512 624697
rect 42448 623757 42454 623809
rect 42506 623797 42512 623809
rect 43696 623797 43702 623809
rect 42506 623769 43702 623797
rect 42506 623757 42512 623769
rect 43696 623757 43702 623769
rect 43754 623757 43760 623809
rect 42160 622203 42166 622255
rect 42218 622243 42224 622255
rect 43408 622243 43414 622255
rect 42218 622215 43414 622243
rect 42218 622203 42224 622215
rect 43408 622203 43414 622215
rect 43466 622203 43472 622255
rect 656368 622055 656374 622107
rect 656426 622095 656432 622107
rect 669712 622095 669718 622107
rect 656426 622067 669718 622095
rect 656426 622055 656432 622067
rect 669712 622055 669718 622067
rect 669770 622055 669776 622107
rect 42160 621611 42166 621663
rect 42218 621651 42224 621663
rect 43024 621651 43030 621663
rect 42218 621623 43030 621651
rect 42218 621611 42224 621623
rect 43024 621611 43030 621623
rect 43082 621611 43088 621663
rect 43024 621463 43030 621515
rect 43082 621503 43088 621515
rect 43504 621503 43510 621515
rect 43082 621475 43510 621503
rect 43082 621463 43088 621475
rect 43504 621463 43510 621475
rect 43562 621463 43568 621515
rect 42064 620871 42070 620923
rect 42122 620911 42128 620923
rect 42928 620911 42934 620923
rect 42122 620883 42934 620911
rect 42122 620871 42128 620883
rect 42928 620871 42934 620883
rect 42986 620871 42992 620923
rect 672208 619169 672214 619221
rect 672266 619209 672272 619221
rect 673840 619209 673846 619221
rect 672266 619181 673846 619209
rect 672266 619169 672272 619181
rect 673840 619169 673846 619181
rect 673898 619169 673904 619221
rect 672016 617837 672022 617889
rect 672074 617877 672080 617889
rect 673840 617877 673846 617889
rect 672074 617849 673846 617877
rect 672074 617837 672080 617849
rect 673840 617837 673846 617849
rect 673898 617837 673904 617889
rect 42064 617615 42070 617667
rect 42122 617655 42128 617667
rect 42928 617655 42934 617667
rect 42122 617627 42934 617655
rect 42122 617615 42128 617627
rect 42928 617615 42934 617627
rect 42986 617615 42992 617667
rect 42160 617319 42166 617371
rect 42218 617359 42224 617371
rect 43120 617359 43126 617371
rect 42218 617331 43126 617359
rect 42218 617319 42224 617331
rect 43120 617319 43126 617331
rect 43178 617319 43184 617371
rect 42160 616653 42166 616705
rect 42218 616693 42224 616705
rect 43024 616693 43030 616705
rect 42218 616665 43030 616693
rect 42218 616653 42224 616665
rect 43024 616653 43030 616665
rect 43082 616653 43088 616705
rect 42160 615987 42166 616039
rect 42218 616027 42224 616039
rect 42448 616027 42454 616039
rect 42218 615999 42454 616027
rect 42218 615987 42224 615999
rect 42448 615987 42454 615999
rect 42506 615987 42512 616039
rect 42160 613989 42166 614041
rect 42218 614029 42224 614041
rect 42448 614029 42454 614041
rect 42218 614001 42454 614029
rect 42218 613989 42224 614001
rect 42448 613989 42454 614001
rect 42506 613989 42512 614041
rect 42160 613619 42166 613671
rect 42218 613659 42224 613671
rect 42736 613659 42742 613671
rect 42218 613631 42742 613659
rect 42218 613619 42224 613631
rect 42736 613619 42742 613631
rect 42794 613619 42800 613671
rect 42448 613471 42454 613523
rect 42506 613511 42512 613523
rect 59440 613511 59446 613523
rect 42506 613483 59446 613511
rect 42506 613471 42512 613483
rect 59440 613471 59446 613483
rect 59498 613471 59504 613523
rect 649936 613471 649942 613523
rect 649994 613511 650000 613523
rect 679696 613511 679702 613523
rect 649994 613483 679702 613511
rect 649994 613471 650000 613483
rect 679696 613471 679702 613483
rect 679754 613471 679760 613523
rect 654448 613397 654454 613449
rect 654506 613437 654512 613449
rect 669520 613437 669526 613449
rect 654506 613409 669526 613437
rect 654506 613397 654512 613409
rect 669520 613397 669526 613409
rect 669578 613397 669584 613449
rect 42064 612805 42070 612857
rect 42122 612845 42128 612857
rect 42832 612845 42838 612857
rect 42122 612817 42838 612845
rect 42122 612805 42128 612817
rect 42832 612805 42838 612817
rect 42890 612805 42896 612857
rect 42736 607699 42742 607751
rect 42794 607739 42800 607751
rect 51856 607739 51862 607751
rect 42794 607711 51862 607739
rect 42794 607699 42800 607711
rect 51856 607699 51862 607711
rect 51914 607699 51920 607751
rect 42736 606811 42742 606863
rect 42794 606851 42800 606863
rect 53392 606851 53398 606863
rect 42794 606823 53398 606851
rect 42794 606811 42800 606823
rect 53392 606811 53398 606823
rect 53450 606811 53456 606863
rect 671824 603851 671830 603903
rect 671882 603891 671888 603903
rect 675088 603891 675094 603903
rect 671882 603863 675094 603891
rect 671882 603851 671888 603863
rect 675088 603851 675094 603863
rect 675146 603851 675152 603903
rect 672208 603629 672214 603681
rect 672266 603669 672272 603681
rect 674512 603669 674518 603681
rect 672266 603641 674518 603669
rect 672266 603629 672272 603641
rect 674512 603629 674518 603641
rect 674570 603669 674576 603681
rect 675280 603669 675286 603681
rect 674570 603641 675286 603669
rect 674570 603629 674576 603641
rect 675280 603629 675286 603641
rect 675338 603629 675344 603681
rect 673744 602815 673750 602867
rect 673802 602855 673808 602867
rect 674704 602855 674710 602867
rect 673802 602827 674710 602855
rect 673802 602815 673808 602827
rect 674704 602815 674710 602827
rect 674762 602855 674768 602867
rect 675472 602855 675478 602867
rect 674762 602827 675478 602855
rect 674762 602815 674768 602827
rect 675472 602815 675478 602827
rect 675530 602815 675536 602867
rect 673168 602667 673174 602719
rect 673226 602707 673232 602719
rect 675376 602707 675382 602719
rect 673226 602679 675382 602707
rect 673226 602667 673232 602679
rect 675376 602667 675382 602679
rect 675434 602667 675440 602719
rect 663760 602001 663766 602053
rect 663818 602041 663824 602053
rect 675184 602041 675190 602053
rect 663818 602013 675190 602041
rect 663818 602001 663824 602013
rect 675184 602001 675190 602013
rect 675242 602001 675248 602053
rect 672688 601927 672694 601979
rect 672746 601967 672752 601979
rect 675088 601967 675094 601979
rect 672746 601939 675094 601967
rect 672746 601927 672752 601939
rect 675088 601927 675094 601939
rect 675146 601927 675152 601979
rect 51856 601853 51862 601905
rect 51914 601893 51920 601905
rect 59536 601893 59542 601905
rect 51914 601865 59542 601893
rect 51914 601853 51920 601865
rect 59536 601853 59542 601865
rect 59594 601853 59600 601905
rect 672016 599559 672022 599611
rect 672074 599599 672080 599611
rect 675376 599599 675382 599611
rect 672074 599571 675382 599599
rect 672074 599559 672080 599571
rect 675376 599559 675382 599571
rect 675434 599559 675440 599611
rect 671536 599263 671542 599315
rect 671594 599303 671600 599315
rect 675376 599303 675382 599315
rect 671594 599275 675382 599303
rect 671594 599263 671600 599275
rect 675376 599263 675382 599275
rect 675434 599263 675440 599315
rect 654448 599041 654454 599093
rect 654506 599081 654512 599093
rect 669520 599081 669526 599093
rect 654506 599053 669526 599081
rect 654506 599041 654512 599053
rect 669520 599041 669526 599053
rect 669578 599041 669584 599093
rect 672112 598375 672118 598427
rect 672170 598415 672176 598427
rect 675472 598415 675478 598427
rect 672170 598387 675478 598415
rect 672170 598375 672176 598387
rect 675472 598375 675478 598387
rect 675530 598375 675536 598427
rect 672496 597117 672502 597169
rect 672554 597157 672560 597169
rect 675472 597157 675478 597169
rect 672554 597129 675478 597157
rect 672554 597117 672560 597129
rect 675472 597117 675478 597129
rect 675530 597117 675536 597169
rect 675184 596821 675190 596873
rect 675242 596861 675248 596873
rect 675376 596861 675382 596873
rect 675242 596833 675382 596861
rect 675242 596821 675248 596833
rect 675376 596821 675382 596833
rect 675434 596821 675440 596873
rect 42448 589199 42454 589251
rect 42506 589239 42512 589251
rect 45136 589239 45142 589251
rect 42506 589211 45142 589239
rect 42506 589199 42512 589211
rect 45136 589199 45142 589211
rect 45194 589199 45200 589251
rect 670864 587497 670870 587549
rect 670922 587537 670928 587549
rect 676816 587537 676822 587549
rect 670922 587509 676822 587537
rect 670922 587497 670928 587509
rect 676816 587497 676822 587509
rect 676874 587497 676880 587549
rect 53392 587423 53398 587475
rect 53450 587463 53456 587475
rect 59536 587463 59542 587475
rect 53450 587435 59542 587463
rect 53450 587423 53456 587435
rect 59536 587423 59542 587435
rect 59594 587423 59600 587475
rect 663952 586313 663958 586365
rect 664010 586353 664016 586365
rect 674416 586353 674422 586365
rect 664010 586325 674422 586353
rect 664010 586313 664016 586325
rect 674416 586313 674422 586325
rect 674474 586313 674480 586365
rect 40048 585943 40054 585995
rect 40106 585983 40112 585995
rect 42448 585983 42454 585995
rect 40106 585955 42454 585983
rect 40106 585943 40112 585955
rect 42448 585943 42454 585955
rect 42506 585943 42512 585995
rect 666928 585425 666934 585477
rect 666986 585465 666992 585477
rect 674416 585465 674422 585477
rect 666986 585437 674422 585465
rect 666986 585425 666992 585437
rect 674416 585425 674422 585437
rect 674474 585425 674480 585477
rect 43120 585351 43126 585403
rect 43178 585391 43184 585403
rect 43696 585391 43702 585403
rect 43178 585363 43702 585391
rect 43178 585351 43184 585363
rect 43696 585351 43702 585363
rect 43754 585351 43760 585403
rect 671728 584833 671734 584885
rect 671786 584873 671792 584885
rect 674608 584873 674614 584885
rect 671786 584845 674614 584873
rect 671786 584833 671792 584845
rect 674608 584833 674614 584845
rect 674666 584833 674672 584885
rect 42544 584759 42550 584811
rect 42602 584799 42608 584811
rect 43120 584799 43126 584811
rect 42602 584771 43126 584799
rect 42602 584759 42608 584771
rect 43120 584759 43126 584771
rect 43178 584759 43184 584811
rect 655216 584759 655222 584811
rect 655274 584799 655280 584811
rect 674704 584799 674710 584811
rect 655274 584771 674710 584799
rect 655274 584759 655280 584771
rect 674704 584759 674710 584771
rect 674762 584759 674768 584811
rect 42832 584685 42838 584737
rect 42890 584725 42896 584737
rect 50512 584725 50518 584737
rect 42890 584697 50518 584725
rect 42890 584685 42896 584697
rect 50512 584685 50518 584697
rect 50570 584685 50576 584737
rect 41968 584241 41974 584293
rect 42026 584281 42032 584293
rect 43216 584281 43222 584293
rect 42026 584253 43222 584281
rect 42026 584241 42032 584253
rect 43216 584241 43222 584253
rect 43274 584241 43280 584293
rect 41776 584167 41782 584219
rect 41834 584167 41840 584219
rect 42160 584167 42166 584219
rect 42218 584207 42224 584219
rect 42928 584207 42934 584219
rect 42218 584179 42934 584207
rect 42218 584167 42224 584179
rect 42928 584167 42934 584179
rect 42986 584167 42992 584219
rect 41794 583997 41822 584167
rect 41776 583945 41782 583997
rect 41834 583945 41840 583997
rect 672400 583575 672406 583627
rect 672458 583615 672464 583627
rect 674704 583615 674710 583627
rect 672458 583587 674710 583615
rect 672458 583575 672464 583587
rect 674704 583575 674710 583587
rect 674762 583575 674768 583627
rect 675184 582539 675190 582591
rect 675242 582579 675248 582591
rect 676816 582579 676822 582591
rect 675242 582551 676822 582579
rect 675242 582539 675248 582551
rect 676816 582539 676822 582551
rect 676874 582539 676880 582591
rect 42160 582095 42166 582147
rect 42218 582135 42224 582147
rect 42448 582135 42454 582147
rect 42218 582107 42454 582135
rect 42218 582095 42224 582107
rect 42448 582095 42454 582107
rect 42506 582095 42512 582147
rect 42064 581429 42070 581481
rect 42122 581469 42128 581481
rect 42832 581469 42838 581481
rect 42122 581441 42838 581469
rect 42122 581429 42128 581441
rect 42832 581429 42838 581441
rect 42890 581429 42896 581481
rect 42832 581281 42838 581333
rect 42890 581321 42896 581333
rect 43216 581321 43222 581333
rect 42890 581293 43222 581321
rect 42890 581281 42896 581293
rect 43216 581281 43222 581293
rect 43274 581281 43280 581333
rect 42064 580245 42070 580297
rect 42122 580285 42128 580297
rect 43024 580285 43030 580297
rect 42122 580257 43030 580285
rect 42122 580245 42128 580257
rect 43024 580245 43030 580257
rect 43082 580245 43088 580297
rect 42160 578987 42166 579039
rect 42218 579027 42224 579039
rect 43312 579027 43318 579039
rect 42218 578999 43318 579027
rect 42218 578987 42224 578999
rect 43312 578987 43318 578999
rect 43370 578987 43376 579039
rect 672400 578839 672406 578891
rect 672458 578879 672464 578891
rect 672784 578879 672790 578891
rect 672458 578851 672790 578879
rect 672458 578839 672464 578851
rect 672784 578839 672790 578851
rect 672842 578839 672848 578891
rect 42064 578395 42070 578447
rect 42122 578435 42128 578447
rect 42928 578435 42934 578447
rect 42122 578407 42934 578435
rect 42122 578395 42128 578407
rect 42928 578395 42934 578407
rect 42986 578395 42992 578447
rect 42160 577655 42166 577707
rect 42218 577695 42224 577707
rect 43120 577695 43126 577707
rect 42218 577667 43126 577695
rect 42218 577655 42224 577667
rect 43120 577655 43126 577667
rect 43178 577655 43184 577707
rect 43120 577507 43126 577559
rect 43178 577547 43184 577559
rect 43696 577547 43702 577559
rect 43178 577519 43702 577547
rect 43178 577507 43184 577519
rect 43696 577507 43702 577519
rect 43754 577507 43760 577559
rect 671920 575361 671926 575413
rect 671978 575401 671984 575413
rect 674704 575401 674710 575413
rect 671978 575373 674710 575401
rect 671978 575361 671984 575373
rect 674704 575361 674710 575373
rect 674762 575361 674768 575413
rect 671440 574473 671446 574525
rect 671498 574513 671504 574525
rect 674704 574513 674710 574525
rect 671498 574485 674710 574513
rect 671498 574473 671504 574485
rect 674704 574473 674710 574485
rect 674762 574473 674768 574525
rect 42160 574103 42166 574155
rect 42218 574143 42224 574155
rect 42832 574143 42838 574155
rect 42218 574115 42838 574143
rect 42218 574103 42224 574115
rect 42832 574103 42838 574115
rect 42890 574103 42896 574155
rect 672304 573585 672310 573637
rect 672362 573625 672368 573637
rect 674416 573625 674422 573637
rect 672362 573597 674422 573625
rect 672362 573585 672368 573597
rect 674416 573585 674422 573597
rect 674474 573585 674480 573637
rect 42064 573215 42070 573267
rect 42122 573255 42128 573267
rect 43024 573255 43030 573267
rect 42122 573227 43030 573255
rect 42122 573215 42128 573227
rect 43024 573215 43030 573227
rect 43082 573215 43088 573267
rect 654448 573141 654454 573193
rect 654506 573181 654512 573193
rect 661168 573181 661174 573193
rect 654506 573153 661174 573181
rect 654506 573141 654512 573153
rect 661168 573141 661174 573153
rect 661226 573141 661232 573193
rect 672880 572993 672886 573045
rect 672938 573033 672944 573045
rect 674704 573033 674710 573045
rect 672938 573005 674710 573033
rect 672938 572993 672944 573005
rect 674704 572993 674710 573005
rect 674762 572993 674768 573045
rect 42160 572623 42166 572675
rect 42218 572663 42224 572675
rect 42928 572663 42934 572675
rect 42218 572635 42934 572663
rect 42218 572623 42224 572635
rect 42928 572623 42934 572635
rect 42986 572623 42992 572675
rect 671632 571957 671638 572009
rect 671690 571997 671696 572009
rect 674416 571997 674422 572009
rect 671690 571969 674422 571997
rect 671690 571957 671696 571969
rect 674416 571957 674422 571969
rect 674474 571957 674480 572009
rect 672592 571365 672598 571417
rect 672650 571405 672656 571417
rect 674704 571405 674710 571417
rect 672650 571377 674710 571405
rect 672650 571365 672656 571377
rect 674704 571365 674710 571377
rect 674762 571365 674768 571417
rect 42160 570995 42166 571047
rect 42218 571035 42224 571047
rect 43120 571035 43126 571047
rect 42218 571007 43126 571035
rect 42218 570995 42224 571007
rect 43120 570995 43126 571007
rect 43178 570995 43184 571047
rect 42064 570403 42070 570455
rect 42122 570443 42128 570455
rect 42448 570443 42454 570455
rect 42122 570415 42454 570443
rect 42122 570403 42128 570415
rect 42448 570403 42454 570415
rect 42506 570403 42512 570455
rect 42352 570255 42358 570307
rect 42410 570295 42416 570307
rect 59536 570295 59542 570307
rect 42410 570267 59542 570295
rect 42410 570255 42416 570267
rect 59536 570255 59542 570267
rect 59594 570255 59600 570307
rect 42064 569663 42070 569715
rect 42122 569703 42128 569715
rect 42928 569703 42934 569715
rect 42122 569675 42934 569703
rect 42122 569663 42128 569675
rect 42928 569663 42934 569675
rect 42986 569663 42992 569715
rect 650032 567369 650038 567421
rect 650090 567409 650096 567421
rect 679792 567409 679798 567421
rect 650090 567381 679798 567409
rect 650090 567369 650096 567381
rect 679792 567369 679798 567381
rect 679850 567369 679856 567421
rect 34480 564483 34486 564535
rect 34538 564523 34544 564535
rect 53392 564523 53398 564535
rect 34538 564495 53398 564523
rect 34538 564483 34544 564495
rect 53392 564483 53398 564495
rect 53450 564483 53456 564535
rect 654448 564409 654454 564461
rect 654506 564449 654512 564461
rect 666640 564449 666646 564461
rect 654506 564421 666646 564449
rect 654506 564409 654512 564421
rect 666640 564409 666646 564421
rect 666698 564409 666704 564461
rect 672208 564409 672214 564461
rect 672266 564449 672272 564461
rect 674992 564449 674998 564461
rect 672266 564421 674998 564449
rect 672266 564409 672272 564421
rect 674992 564409 674998 564421
rect 675050 564409 675056 564461
rect 672208 564261 672214 564313
rect 672266 564301 672272 564313
rect 672784 564301 672790 564313
rect 672266 564273 672790 564301
rect 672266 564261 672272 564273
rect 672784 564261 672790 564273
rect 672842 564261 672848 564313
rect 42448 563447 42454 563499
rect 42506 563487 42512 563499
rect 50512 563487 50518 563499
rect 42506 563459 50518 563487
rect 42506 563447 42512 563459
rect 50512 563447 50518 563459
rect 50570 563447 50576 563499
rect 673744 561597 673750 561649
rect 673802 561637 673808 561649
rect 675088 561637 675094 561649
rect 673802 561609 675094 561637
rect 673802 561597 673808 561609
rect 675088 561597 675094 561609
rect 675146 561597 675152 561649
rect 674320 559525 674326 559577
rect 674378 559565 674384 559577
rect 675376 559565 675382 559577
rect 674378 559537 675382 559565
rect 674378 559525 674384 559537
rect 675376 559525 675382 559537
rect 675434 559525 675440 559577
rect 53392 558637 53398 558689
rect 53450 558677 53456 558689
rect 59536 558677 59542 558689
rect 53450 558649 59542 558677
rect 53450 558637 53456 558649
rect 59536 558637 59542 558649
rect 59594 558637 59600 558689
rect 673936 558045 673942 558097
rect 673994 558085 674000 558097
rect 675376 558085 675382 558097
rect 673994 558057 675382 558085
rect 673994 558045 674000 558057
rect 675376 558045 675382 558057
rect 675434 558045 675440 558097
rect 660880 555825 660886 555877
rect 660938 555865 660944 555877
rect 675184 555865 675190 555877
rect 660938 555837 675190 555865
rect 660938 555825 660944 555837
rect 675184 555825 675190 555837
rect 675242 555825 675248 555877
rect 674512 555011 674518 555063
rect 674570 555051 674576 555063
rect 675472 555051 675478 555063
rect 674570 555023 675478 555051
rect 674570 555011 674576 555023
rect 675472 555011 675478 555023
rect 675530 555011 675536 555063
rect 675088 554493 675094 554545
rect 675146 554533 675152 554545
rect 675376 554533 675382 554545
rect 675146 554505 675382 554533
rect 675146 554493 675152 554505
rect 675376 554493 675382 554505
rect 675434 554493 675440 554545
rect 674128 553901 674134 553953
rect 674186 553941 674192 553953
rect 675472 553941 675478 553953
rect 674186 553913 675478 553941
rect 674186 553901 674192 553913
rect 675472 553901 675478 553913
rect 675530 553901 675536 553953
rect 674800 553161 674806 553213
rect 674858 553201 674864 553213
rect 675376 553201 675382 553213
rect 674858 553173 675382 553201
rect 674858 553161 674864 553173
rect 675376 553161 675382 553173
rect 675434 553161 675440 553213
rect 674416 551903 674422 551955
rect 674474 551943 674480 551955
rect 675472 551943 675478 551955
rect 674474 551915 675478 551943
rect 674474 551903 674480 551915
rect 675472 551903 675478 551915
rect 675530 551903 675536 551955
rect 675184 551607 675190 551659
rect 675242 551647 675248 551659
rect 675376 551647 675382 551659
rect 675242 551619 675382 551647
rect 675242 551607 675248 551619
rect 675376 551607 675382 551619
rect 675434 551607 675440 551659
rect 654448 550127 654454 550179
rect 654506 550167 654512 550179
rect 663952 550167 663958 550179
rect 654506 550139 663958 550167
rect 654506 550127 654512 550139
rect 663952 550127 663958 550139
rect 664010 550127 664016 550179
rect 675184 550053 675190 550105
rect 675242 550093 675248 550105
rect 675472 550093 675478 550105
rect 675242 550065 675478 550093
rect 675242 550053 675248 550065
rect 675472 550053 675478 550065
rect 675530 550053 675536 550105
rect 674608 548203 674614 548255
rect 674666 548243 674672 548255
rect 675376 548243 675382 548255
rect 674666 548215 675382 548243
rect 674666 548203 674672 548215
rect 675376 548203 675382 548215
rect 675434 548203 675440 548255
rect 42640 546205 42646 546257
rect 42698 546245 42704 546257
rect 45232 546245 45238 546257
rect 42698 546217 45238 546245
rect 42698 546205 42704 546217
rect 45232 546205 45238 546217
rect 45290 546205 45296 546257
rect 42352 545539 42358 545591
rect 42410 545579 42416 545591
rect 42640 545579 42646 545591
rect 42410 545551 42646 545579
rect 42410 545539 42416 545551
rect 42640 545539 42646 545551
rect 42698 545539 42704 545591
rect 42832 544947 42838 544999
rect 42890 544947 42896 544999
rect 42850 544629 42878 544947
rect 42832 544577 42838 544629
rect 42890 544577 42896 544629
rect 40048 544281 40054 544333
rect 40106 544321 40112 544333
rect 42928 544321 42934 544333
rect 40106 544293 42934 544321
rect 40106 544281 40112 544293
rect 42928 544281 42934 544293
rect 42986 544281 42992 544333
rect 50512 543689 50518 543741
rect 50570 543729 50576 543741
rect 59536 543729 59542 543741
rect 50570 543701 59542 543729
rect 50570 543689 50576 543701
rect 59536 543689 59542 543701
rect 59594 543689 59600 543741
rect 43696 541469 43702 541521
rect 43754 541509 43760 541521
rect 53296 541509 53302 541521
rect 43754 541481 53302 541509
rect 43754 541469 43760 541481
rect 53296 541469 53302 541481
rect 53354 541469 53360 541521
rect 655408 541469 655414 541521
rect 655466 541509 655472 541521
rect 674704 541509 674710 541521
rect 655466 541481 674710 541509
rect 655466 541469 655472 541481
rect 674704 541469 674710 541481
rect 674762 541469 674768 541521
rect 672208 541395 672214 541447
rect 672266 541435 672272 541447
rect 673840 541435 673846 541447
rect 672266 541407 673846 541435
rect 672266 541395 672272 541407
rect 673840 541395 673846 541407
rect 673898 541395 673904 541447
rect 661264 541321 661270 541373
rect 661322 541361 661328 541373
rect 674224 541361 674230 541373
rect 661322 541333 674230 541361
rect 661322 541321 661328 541333
rect 674224 541321 674230 541333
rect 674282 541321 674288 541373
rect 674704 541321 674710 541373
rect 674762 541361 674768 541373
rect 675184 541361 675190 541373
rect 674762 541333 675190 541361
rect 674762 541321 674768 541333
rect 675184 541321 675190 541333
rect 675242 541321 675248 541373
rect 41968 541025 41974 541077
rect 42026 541065 42032 541077
rect 43504 541065 43510 541077
rect 42026 541037 43510 541065
rect 42026 541025 42032 541037
rect 43504 541025 43510 541037
rect 43562 541025 43568 541077
rect 41776 540951 41782 541003
rect 41834 540951 41840 541003
rect 42160 540951 42166 541003
rect 42218 540991 42224 541003
rect 43312 540991 43318 541003
rect 42218 540963 43318 540991
rect 42218 540951 42224 540963
rect 43312 540951 43318 540963
rect 43370 540951 43376 541003
rect 41794 540781 41822 540951
rect 41776 540729 41782 540781
rect 41834 540729 41840 540781
rect 664048 540433 664054 540485
rect 664106 540473 664112 540485
rect 674224 540473 674230 540485
rect 664106 540445 674230 540473
rect 664106 540433 664112 540445
rect 674224 540433 674230 540445
rect 674282 540433 674288 540485
rect 42928 540063 42934 540115
rect 42986 540063 42992 540115
rect 42946 539881 42974 540063
rect 43024 539881 43030 539893
rect 42946 539853 43030 539881
rect 43024 539841 43030 539853
rect 43082 539841 43088 539893
rect 42064 538879 42070 538931
rect 42122 538919 42128 538931
rect 43024 538919 43030 538931
rect 42122 538891 43030 538919
rect 42122 538879 42128 538891
rect 43024 538879 43030 538891
rect 43082 538879 43088 538931
rect 654448 538583 654454 538635
rect 654506 538623 654512 538635
rect 661072 538623 661078 538635
rect 654506 538595 661078 538623
rect 654506 538583 654512 538595
rect 661072 538583 661078 538595
rect 661130 538583 661136 538635
rect 674032 538583 674038 538635
rect 674090 538623 674096 538635
rect 675088 538623 675094 538635
rect 674090 538595 675094 538623
rect 674090 538583 674096 538595
rect 675088 538583 675094 538595
rect 675146 538583 675152 538635
rect 42160 538139 42166 538191
rect 42218 538179 42224 538191
rect 43696 538179 43702 538191
rect 42218 538151 43702 538179
rect 42218 538139 42224 538151
rect 43696 538139 43702 538151
rect 43754 538139 43760 538191
rect 42064 537029 42070 537081
rect 42122 537069 42128 537081
rect 42928 537069 42934 537081
rect 42122 537041 42934 537069
rect 42122 537029 42128 537041
rect 42928 537029 42934 537041
rect 42986 537029 42992 537081
rect 42064 535771 42070 535823
rect 42122 535811 42128 535823
rect 42832 535811 42838 535823
rect 42122 535783 42838 535811
rect 42122 535771 42128 535783
rect 42832 535771 42838 535783
rect 42890 535771 42896 535823
rect 42160 535031 42166 535083
rect 42218 535071 42224 535083
rect 42736 535071 42742 535083
rect 42218 535043 42742 535071
rect 42218 535031 42224 535043
rect 42736 535031 42742 535043
rect 42794 535031 42800 535083
rect 42160 534439 42166 534491
rect 42218 534479 42224 534491
rect 43120 534479 43126 534491
rect 42218 534451 43126 534479
rect 42218 534439 42224 534451
rect 43120 534439 43126 534451
rect 43178 534439 43184 534491
rect 43216 534439 43222 534491
rect 43274 534439 43280 534491
rect 43234 534269 43262 534439
rect 43216 534217 43222 534269
rect 43274 534217 43280 534269
rect 42064 533921 42070 533973
rect 42122 533961 42128 533973
rect 43024 533961 43030 533973
rect 42122 533933 43030 533961
rect 42122 533921 42128 533933
rect 43024 533921 43030 533933
rect 43082 533921 43088 533973
rect 43024 533773 43030 533825
rect 43082 533813 43088 533825
rect 43504 533813 43510 533825
rect 43082 533785 43510 533813
rect 43082 533773 43088 533785
rect 43504 533773 43510 533785
rect 43562 533773 43568 533825
rect 42256 532811 42262 532863
rect 42314 532851 42320 532863
rect 42640 532851 42646 532863
rect 42314 532823 42646 532851
rect 42314 532811 42320 532823
rect 42640 532811 42646 532823
rect 42698 532811 42704 532863
rect 672688 532737 672694 532789
rect 672746 532777 672752 532789
rect 673840 532777 673846 532789
rect 672746 532749 673846 532777
rect 672746 532737 672752 532749
rect 673840 532737 673846 532749
rect 673898 532737 673904 532789
rect 671824 532663 671830 532715
rect 671882 532703 671888 532715
rect 673744 532703 673750 532715
rect 671882 532675 673750 532703
rect 671882 532663 671888 532675
rect 673744 532663 673750 532675
rect 673802 532663 673808 532715
rect 42160 531331 42166 531383
rect 42218 531371 42224 531383
rect 43120 531371 43126 531383
rect 42218 531343 43126 531371
rect 42218 531331 42224 531343
rect 43120 531331 43126 531343
rect 43178 531331 43184 531383
rect 42256 530295 42262 530347
rect 42314 530335 42320 530347
rect 42928 530335 42934 530347
rect 42314 530307 42934 530335
rect 42314 530295 42320 530307
rect 42928 530295 42934 530307
rect 42986 530295 42992 530347
rect 42064 530147 42070 530199
rect 42122 530187 42128 530199
rect 42832 530187 42838 530199
rect 42122 530159 42838 530187
rect 42122 530147 42128 530159
rect 42832 530147 42838 530159
rect 42890 530147 42896 530199
rect 672496 529851 672502 529903
rect 672554 529891 672560 529903
rect 673840 529891 673846 529903
rect 672554 529863 673846 529891
rect 672554 529851 672560 529863
rect 673840 529851 673846 529863
rect 673898 529851 673904 529903
rect 671536 529185 671542 529237
rect 671594 529225 671600 529237
rect 673840 529225 673846 529237
rect 671594 529197 673846 529225
rect 671594 529185 671600 529197
rect 673840 529185 673846 529197
rect 673898 529185 673904 529237
rect 42160 527631 42166 527683
rect 42218 527671 42224 527683
rect 43024 527671 43030 527683
rect 42218 527643 43030 527671
rect 42218 527631 42224 527643
rect 43024 527631 43030 527643
rect 43082 527631 43088 527683
rect 42064 527187 42070 527239
rect 42122 527227 42128 527239
rect 42736 527227 42742 527239
rect 42122 527199 42742 527227
rect 42122 527187 42128 527199
rect 42736 527187 42742 527199
rect 42794 527187 42800 527239
rect 42352 527039 42358 527091
rect 42410 527079 42416 527091
rect 59536 527079 59542 527091
rect 42410 527051 59542 527079
rect 42410 527039 42416 527051
rect 59536 527039 59542 527051
rect 59594 527039 59600 527091
rect 654448 527039 654454 527091
rect 654506 527079 654512 527091
rect 669808 527079 669814 527091
rect 654506 527051 669814 527079
rect 654506 527039 654512 527051
rect 669808 527039 669814 527051
rect 669866 527039 669872 527091
rect 672016 526891 672022 526943
rect 672074 526931 672080 526943
rect 673840 526931 673846 526943
rect 672074 526903 673846 526931
rect 672074 526891 672080 526903
rect 673840 526891 673846 526903
rect 673898 526891 673904 526943
rect 672112 526743 672118 526795
rect 672170 526783 672176 526795
rect 673840 526783 673846 526795
rect 672170 526755 673846 526783
rect 672170 526743 672176 526755
rect 673840 526743 673846 526755
rect 673898 526743 673904 526795
rect 42160 526595 42166 526647
rect 42218 526635 42224 526647
rect 42640 526635 42646 526647
rect 42218 526607 42646 526635
rect 42218 526595 42224 526607
rect 42640 526595 42646 526607
rect 42698 526595 42704 526647
rect 650128 521267 650134 521319
rect 650186 521307 650192 521319
rect 679792 521307 679798 521319
rect 650186 521279 679798 521307
rect 650186 521267 650192 521279
rect 679792 521267 679798 521279
rect 679850 521267 679856 521319
rect 674512 518307 674518 518359
rect 674570 518347 674576 518359
rect 674896 518347 674902 518359
rect 674570 518319 674902 518347
rect 674570 518307 674576 518319
rect 674896 518307 674902 518319
rect 674954 518307 674960 518359
rect 654064 517271 654070 517323
rect 654122 517311 654128 517323
rect 663856 517311 663862 517323
rect 654122 517283 663862 517311
rect 654122 517271 654128 517283
rect 663856 517271 663862 517283
rect 663914 517271 663920 517323
rect 50512 512683 50518 512735
rect 50570 512723 50576 512735
rect 59344 512723 59350 512735
rect 50570 512695 59350 512723
rect 50570 512683 50576 512695
rect 59344 512683 59350 512695
rect 59402 512683 59408 512735
rect 673936 508317 673942 508369
rect 673994 508357 674000 508369
rect 674128 508357 674134 508369
rect 673994 508329 674134 508357
rect 673994 508317 674000 508329
rect 674128 508317 674134 508329
rect 674186 508317 674192 508369
rect 674320 508095 674326 508147
rect 674378 508095 674384 508147
rect 674338 507925 674366 508095
rect 674320 507873 674326 507925
rect 674378 507873 674384 507925
rect 674416 507873 674422 507925
rect 674474 507913 674480 507925
rect 674896 507913 674902 507925
rect 674474 507885 674902 507913
rect 674474 507873 674480 507885
rect 674896 507873 674902 507885
rect 674954 507873 674960 507925
rect 654928 504025 654934 504077
rect 654986 504065 654992 504077
rect 666640 504065 666646 504077
rect 654986 504037 666646 504065
rect 654986 504025 654992 504037
rect 666640 504025 666646 504037
rect 666698 504025 666704 504077
rect 53392 498253 53398 498305
rect 53450 498293 53456 498305
rect 57808 498293 57814 498305
rect 53450 498265 57814 498293
rect 53450 498253 53456 498265
rect 57808 498253 57814 498265
rect 57866 498253 57872 498305
rect 666832 497513 666838 497565
rect 666890 497553 666896 497565
rect 674512 497553 674518 497565
rect 666890 497525 674518 497553
rect 666890 497513 666896 497525
rect 674512 497513 674518 497525
rect 674570 497513 674576 497565
rect 669712 496625 669718 496677
rect 669770 496665 669776 496677
rect 674512 496665 674518 496677
rect 669770 496637 674518 496665
rect 669770 496625 669776 496637
rect 674512 496625 674518 496637
rect 674570 496625 674576 496677
rect 655312 495515 655318 495567
rect 655370 495555 655376 495567
rect 674704 495555 674710 495567
rect 655370 495527 674710 495555
rect 655370 495515 655376 495527
rect 674704 495515 674710 495527
rect 674762 495515 674768 495567
rect 53296 483823 53302 483875
rect 53354 483863 53360 483875
rect 59536 483863 59542 483875
rect 53354 483835 59542 483863
rect 53354 483823 53360 483835
rect 59536 483823 59542 483835
rect 59594 483823 59600 483875
rect 654448 480937 654454 480989
rect 654506 480977 654512 480989
rect 666832 480977 666838 480989
rect 654506 480949 666838 480977
rect 654506 480937 654512 480949
rect 666832 480937 666838 480949
rect 666890 480937 666896 480989
rect 650224 478125 650230 478177
rect 650282 478165 650288 478177
rect 679792 478165 679798 478177
rect 650282 478137 679798 478165
rect 650282 478125 650288 478137
rect 679792 478125 679798 478137
rect 679850 478125 679856 478177
rect 654448 470577 654454 470629
rect 654506 470617 654512 470629
rect 660976 470617 660982 470629
rect 654506 470589 660982 470617
rect 654506 470577 654512 470589
rect 660976 470577 660982 470589
rect 661034 470577 661040 470629
rect 50608 469467 50614 469519
rect 50666 469507 50672 469519
rect 59536 469507 59542 469519
rect 50666 469479 59542 469507
rect 50666 469467 50672 469479
rect 59536 469467 59542 469479
rect 59594 469467 59600 469519
rect 656368 457923 656374 457975
rect 656426 457963 656432 457975
rect 663856 457963 663862 457975
rect 656426 457935 663862 457963
rect 656426 457923 656432 457935
rect 663856 457923 663862 457935
rect 663914 457923 663920 457975
rect 45424 455037 45430 455089
rect 45482 455077 45488 455089
rect 59536 455077 59542 455089
rect 45482 455049 59542 455077
rect 45482 455037 45488 455049
rect 59536 455037 59542 455049
rect 59594 455037 59600 455089
rect 654448 446379 654454 446431
rect 654506 446419 654512 446431
rect 669712 446419 669718 446431
rect 654506 446391 669718 446419
rect 654506 446379 654512 446391
rect 669712 446379 669718 446391
rect 669770 446379 669776 446431
rect 45328 440681 45334 440733
rect 45386 440721 45392 440733
rect 57808 440721 57814 440733
rect 45386 440693 57814 440721
rect 45386 440681 45392 440693
rect 57808 440681 57814 440693
rect 57866 440681 57872 440733
rect 42640 436907 42646 436959
rect 42698 436947 42704 436959
rect 50512 436947 50518 436959
rect 42698 436919 50518 436947
rect 42698 436907 42704 436919
rect 50512 436907 50518 436919
rect 50570 436907 50576 436959
rect 42640 436093 42646 436145
rect 42698 436133 42704 436145
rect 53392 436133 53398 436145
rect 42698 436105 53398 436133
rect 42698 436093 42704 436105
rect 53392 436093 53398 436105
rect 53450 436093 53456 436145
rect 654448 434909 654454 434961
rect 654506 434949 654512 434961
rect 664048 434949 664054 434961
rect 654506 434921 664054 434949
rect 654506 434909 654512 434921
rect 664048 434909 664054 434921
rect 664106 434909 664112 434961
rect 53392 426251 53398 426303
rect 53450 426291 53456 426303
rect 59536 426291 59542 426303
rect 53450 426263 59542 426291
rect 53450 426251 53456 426263
rect 59536 426251 59542 426263
rect 59594 426251 59600 426303
rect 654448 423291 654454 423343
rect 654506 423331 654512 423343
rect 669616 423331 669622 423343
rect 654506 423303 669622 423331
rect 654506 423291 654512 423303
rect 669616 423291 669622 423303
rect 669674 423291 669680 423343
rect 42160 419961 42166 420013
rect 42218 420001 42224 420013
rect 42352 420001 42358 420013
rect 42218 419973 42358 420001
rect 42218 419961 42224 419973
rect 42352 419961 42358 419973
rect 42410 419961 42416 420013
rect 42640 418555 42646 418607
rect 42698 418595 42704 418607
rect 44656 418595 44662 418607
rect 42698 418567 44662 418595
rect 42698 418555 42704 418567
rect 44656 418555 44662 418567
rect 44714 418555 44720 418607
rect 37360 416927 37366 416979
rect 37418 416967 37424 416979
rect 42928 416967 42934 416979
rect 37418 416939 42934 416967
rect 37418 416927 37424 416939
rect 42928 416927 42934 416939
rect 42986 416927 42992 416979
rect 40144 416187 40150 416239
rect 40202 416227 40208 416239
rect 43120 416227 43126 416239
rect 40202 416199 43126 416227
rect 40202 416187 40208 416199
rect 43120 416187 43126 416199
rect 43178 416187 43184 416239
rect 40240 414781 40246 414833
rect 40298 414821 40304 414833
rect 42832 414821 42838 414833
rect 40298 414793 42838 414821
rect 40298 414781 40304 414793
rect 42832 414781 42838 414793
rect 42890 414781 42896 414833
rect 37264 414707 37270 414759
rect 37322 414747 37328 414759
rect 43312 414747 43318 414759
rect 37322 414719 43318 414747
rect 37322 414707 37328 414719
rect 43312 414707 43318 414719
rect 43370 414707 43376 414759
rect 41776 413375 41782 413427
rect 41834 413375 41840 413427
rect 41794 413205 41822 413375
rect 41776 413153 41782 413205
rect 41834 413153 41840 413205
rect 53488 411821 53494 411873
rect 53546 411861 53552 411873
rect 59536 411861 59542 411873
rect 53546 411833 59542 411861
rect 53546 411821 53552 411833
rect 59536 411821 59542 411833
rect 59594 411821 59600 411873
rect 42160 411303 42166 411355
rect 42218 411343 42224 411355
rect 42352 411343 42358 411355
rect 42218 411315 42358 411343
rect 42218 411303 42224 411315
rect 42352 411303 42358 411315
rect 42410 411303 42416 411355
rect 42064 410489 42070 410541
rect 42122 410529 42128 410541
rect 47440 410529 47446 410541
rect 42122 410501 47446 410529
rect 42122 410489 42128 410501
rect 47440 410489 47446 410501
rect 47498 410489 47504 410541
rect 42160 409453 42166 409505
rect 42218 409493 42224 409505
rect 42736 409493 42742 409505
rect 42218 409465 42742 409493
rect 42218 409453 42224 409465
rect 42736 409453 42742 409465
rect 42794 409453 42800 409505
rect 42832 409379 42838 409431
rect 42890 409379 42896 409431
rect 42850 409209 42878 409379
rect 43024 409231 43030 409283
rect 43082 409231 43088 409283
rect 42832 409157 42838 409209
rect 42890 409157 42896 409209
rect 43042 409061 43070 409231
rect 669520 409157 669526 409209
rect 669578 409197 669584 409209
rect 674416 409197 674422 409209
rect 669578 409169 674422 409197
rect 669578 409157 669584 409169
rect 674416 409157 674422 409169
rect 674474 409157 674480 409209
rect 655120 409083 655126 409135
rect 655178 409123 655184 409135
rect 674704 409123 674710 409135
rect 655178 409095 674710 409123
rect 655178 409083 655184 409095
rect 674704 409083 674710 409095
rect 674762 409083 674768 409135
rect 43024 409009 43030 409061
rect 43082 409009 43088 409061
rect 43120 409009 43126 409061
rect 43178 409049 43184 409061
rect 43312 409049 43318 409061
rect 43178 409021 43318 409049
rect 43178 409009 43184 409021
rect 43312 409009 43318 409021
rect 43370 409009 43376 409061
rect 654448 408935 654454 408987
rect 654506 408975 654512 408987
rect 669616 408975 669622 408987
rect 654506 408947 669622 408975
rect 654506 408935 654512 408947
rect 669616 408935 669622 408947
rect 669674 408935 669680 408987
rect 661168 408417 661174 408469
rect 661226 408457 661232 408469
rect 674704 408457 674710 408469
rect 661226 408429 674710 408457
rect 661226 408417 661232 408429
rect 674704 408417 674710 408429
rect 674762 408417 674768 408469
rect 42160 408195 42166 408247
rect 42218 408235 42224 408247
rect 42832 408235 42838 408247
rect 42218 408207 42838 408235
rect 42218 408195 42224 408207
rect 42832 408195 42838 408207
rect 42890 408195 42896 408247
rect 42064 407455 42070 407507
rect 42122 407495 42128 407507
rect 42928 407495 42934 407507
rect 42122 407467 42934 407495
rect 42122 407455 42128 407467
rect 42928 407455 42934 407467
rect 42986 407455 42992 407507
rect 42160 406863 42166 406915
rect 42218 406903 42224 406915
rect 43024 406903 43030 406915
rect 42218 406875 43030 406903
rect 42218 406863 42224 406875
rect 43024 406863 43030 406875
rect 43082 406863 43088 406915
rect 42160 403829 42166 403881
rect 42218 403869 42224 403881
rect 43120 403869 43126 403881
rect 42218 403841 43126 403869
rect 42218 403829 42224 403841
rect 43120 403829 43126 403841
rect 43178 403829 43184 403881
rect 42160 403311 42166 403363
rect 42218 403351 42224 403363
rect 42736 403351 42742 403363
rect 42218 403323 42742 403351
rect 42218 403311 42224 403323
rect 42736 403311 42742 403323
rect 42794 403311 42800 403363
rect 654640 397465 654646 397517
rect 654698 397505 654704 397517
rect 661168 397505 661174 397517
rect 654698 397477 661174 397505
rect 654698 397465 654704 397477
rect 661168 397465 661174 397477
rect 661226 397465 661232 397517
rect 42352 393913 42358 393965
rect 42410 393953 42416 393965
rect 50608 393953 50614 393965
rect 42410 393925 50614 393953
rect 42410 393913 42416 393925
rect 50608 393913 50614 393925
rect 50666 393913 50672 393965
rect 42352 393173 42358 393225
rect 42410 393213 42416 393225
rect 45424 393213 45430 393225
rect 42410 393185 45430 393213
rect 42410 393173 42416 393185
rect 45424 393173 45430 393185
rect 45482 393173 45488 393225
rect 42352 392285 42358 392337
rect 42410 392325 42416 392337
rect 53296 392325 53302 392337
rect 42410 392297 53302 392325
rect 42410 392285 42416 392297
rect 53296 392285 53302 392297
rect 53354 392285 53360 392337
rect 650320 391693 650326 391745
rect 650378 391733 650384 391745
rect 679696 391733 679702 391745
rect 650378 391705 679702 391733
rect 650378 391693 650384 391705
rect 679696 391693 679702 391705
rect 679754 391693 679760 391745
rect 654448 385921 654454 385973
rect 654506 385961 654512 385973
rect 669520 385961 669526 385973
rect 654506 385933 669526 385961
rect 654506 385921 654512 385933
rect 669520 385921 669526 385933
rect 669578 385921 669584 385973
rect 674896 384885 674902 384937
rect 674954 384925 674960 384937
rect 675280 384925 675286 384937
rect 674954 384897 675286 384925
rect 674954 384885 674960 384897
rect 675280 384885 675286 384897
rect 675338 384885 675344 384937
rect 674512 384293 674518 384345
rect 674570 384333 674576 384345
rect 675088 384333 675094 384345
rect 674570 384305 675094 384333
rect 674570 384293 674576 384305
rect 675088 384293 675094 384305
rect 675146 384293 675152 384345
rect 674032 383109 674038 383161
rect 674090 383149 674096 383161
rect 675376 383149 675382 383161
rect 674090 383121 675382 383149
rect 674090 383109 674096 383121
rect 675376 383109 675382 383121
rect 675434 383109 675440 383161
rect 45424 383035 45430 383087
rect 45482 383075 45488 383087
rect 59536 383075 59542 383087
rect 45482 383047 59542 383075
rect 45482 383035 45488 383047
rect 59536 383035 59542 383047
rect 59594 383035 59600 383087
rect 674704 378151 674710 378203
rect 674762 378191 674768 378203
rect 675376 378191 675382 378203
rect 674762 378163 675382 378191
rect 674762 378151 674768 378163
rect 675376 378151 675382 378163
rect 675434 378151 675440 378203
rect 674416 377559 674422 377611
rect 674474 377599 674480 377611
rect 675376 377599 675382 377611
rect 674474 377571 675382 377599
rect 674474 377559 674480 377571
rect 675376 377559 675382 377571
rect 675434 377559 675440 377611
rect 654448 377189 654454 377241
rect 654506 377229 654512 377241
rect 666736 377229 666742 377241
rect 654506 377201 666742 377229
rect 654506 377189 654512 377201
rect 666736 377189 666742 377201
rect 666794 377189 666800 377241
rect 674320 376819 674326 376871
rect 674378 376859 674384 376871
rect 675472 376859 675478 376871
rect 674378 376831 675478 376859
rect 674378 376819 674384 376831
rect 675472 376819 675478 376831
rect 675530 376819 675536 376871
rect 673936 375709 673942 375761
rect 673994 375749 674000 375761
rect 675472 375749 675478 375761
rect 673994 375721 675478 375749
rect 673994 375709 674000 375721
rect 675472 375709 675478 375721
rect 675530 375709 675536 375761
rect 42352 375191 42358 375243
rect 42410 375231 42416 375243
rect 47440 375231 47446 375243
rect 42410 375203 47446 375231
rect 42410 375191 42416 375203
rect 47440 375191 47446 375203
rect 47498 375191 47504 375243
rect 37168 371861 37174 371913
rect 37226 371901 37232 371913
rect 43312 371901 43318 371913
rect 37226 371873 43318 371901
rect 37226 371861 37232 371873
rect 43312 371861 43318 371873
rect 43370 371861 43376 371913
rect 37264 371787 37270 371839
rect 37322 371827 37328 371839
rect 43120 371827 43126 371839
rect 37322 371799 43126 371827
rect 37322 371787 37328 371799
rect 43120 371787 43126 371799
rect 43178 371787 43184 371839
rect 37360 371713 37366 371765
rect 37418 371753 37424 371765
rect 42832 371753 42838 371765
rect 37418 371725 42838 371753
rect 37418 371713 37424 371725
rect 42832 371713 42838 371725
rect 42890 371713 42896 371765
rect 40144 371639 40150 371691
rect 40202 371679 40208 371691
rect 42736 371679 42742 371691
rect 40202 371651 42742 371679
rect 40202 371639 40208 371651
rect 42736 371639 42742 371651
rect 42794 371639 42800 371691
rect 40048 371565 40054 371617
rect 40106 371605 40112 371617
rect 42352 371605 42358 371617
rect 40106 371577 42358 371605
rect 40106 371565 40112 371577
rect 42352 371565 42358 371577
rect 42410 371565 42416 371617
rect 41776 370159 41782 370211
rect 41834 370159 41840 370211
rect 41794 369989 41822 370159
rect 41776 369937 41782 369989
rect 41834 369937 41840 369989
rect 50512 368679 50518 368731
rect 50570 368719 50576 368731
rect 59536 368719 59542 368731
rect 50570 368691 59542 368719
rect 50570 368679 50576 368691
rect 59536 368679 59542 368691
rect 59594 368679 59600 368731
rect 42064 368087 42070 368139
rect 42122 368127 42128 368139
rect 43024 368127 43030 368139
rect 42122 368099 43030 368127
rect 42122 368087 42128 368099
rect 43024 368087 43030 368099
rect 43082 368087 43088 368139
rect 43024 367939 43030 367991
rect 43082 367979 43088 367991
rect 43312 367979 43318 367991
rect 43082 367951 43318 367979
rect 43082 367939 43088 367951
rect 43312 367939 43318 367951
rect 43370 367939 43376 367991
rect 42064 367347 42070 367399
rect 42122 367387 42128 367399
rect 50320 367387 50326 367399
rect 42122 367359 50326 367387
rect 42122 367347 42128 367359
rect 50320 367347 50326 367359
rect 50378 367347 50384 367399
rect 42064 366237 42070 366289
rect 42122 366277 42128 366289
rect 42352 366277 42358 366289
rect 42122 366249 42358 366277
rect 42122 366237 42128 366249
rect 42352 366237 42358 366249
rect 42410 366237 42416 366289
rect 42352 366089 42358 366141
rect 42410 366129 42416 366141
rect 43120 366129 43126 366141
rect 42410 366101 43126 366129
rect 42410 366089 42416 366101
rect 43120 366089 43126 366101
rect 43178 366089 43184 366141
rect 42160 364979 42166 365031
rect 42218 365019 42224 365031
rect 42736 365019 42742 365031
rect 42218 364991 42742 365019
rect 42218 364979 42224 364991
rect 42736 364979 42742 364991
rect 42794 364979 42800 365031
rect 661072 364905 661078 364957
rect 661130 364945 661136 364957
rect 674704 364945 674710 364957
rect 661130 364917 674710 364945
rect 661130 364905 661136 364917
rect 674704 364905 674710 364917
rect 674762 364905 674768 364957
rect 42064 364387 42070 364439
rect 42122 364427 42128 364439
rect 42928 364427 42934 364439
rect 42122 364399 42934 364427
rect 42122 364387 42128 364399
rect 42928 364387 42934 364399
rect 42986 364387 42992 364439
rect 663952 363869 663958 363921
rect 664010 363909 664016 363921
rect 674416 363909 674422 363921
rect 664010 363881 674422 363909
rect 664010 363869 664016 363881
rect 674416 363869 674422 363881
rect 674474 363869 674480 363921
rect 42160 363647 42166 363699
rect 42218 363687 42224 363699
rect 42832 363687 42838 363699
rect 42218 363659 42838 363687
rect 42218 363647 42224 363659
rect 42832 363647 42838 363659
rect 42890 363647 42896 363699
rect 654448 363499 654454 363551
rect 654506 363539 654512 363551
rect 660976 363539 660982 363551
rect 654506 363511 660982 363539
rect 654506 363499 654512 363511
rect 660976 363499 660982 363511
rect 661034 363499 661040 363551
rect 669808 363277 669814 363329
rect 669866 363317 669872 363329
rect 674704 363317 674710 363329
rect 669866 363289 674710 363317
rect 669866 363277 669872 363289
rect 674704 363277 674710 363289
rect 674762 363277 674768 363329
rect 42352 360095 42358 360147
rect 42410 360135 42416 360147
rect 43024 360135 43030 360147
rect 42410 360107 43030 360135
rect 42410 360095 42416 360107
rect 43024 360095 43030 360107
rect 43082 360095 43088 360147
rect 47824 354249 47830 354301
rect 47882 354289 47888 354301
rect 59536 354289 59542 354301
rect 47882 354261 59542 354289
rect 47882 354249 47888 354261
rect 59536 354249 59542 354261
rect 59594 354249 59600 354301
rect 42352 350697 42358 350749
rect 42410 350737 42416 350749
rect 53392 350737 53398 350749
rect 42410 350709 53398 350737
rect 42410 350697 42416 350709
rect 53392 350697 53398 350709
rect 53450 350697 53456 350749
rect 42640 349661 42646 349713
rect 42698 349701 42704 349713
rect 53488 349701 53494 349713
rect 42698 349673 53494 349701
rect 42698 349661 42704 349673
rect 53488 349661 53494 349673
rect 53546 349661 53552 349713
rect 42352 349069 42358 349121
rect 42410 349109 42416 349121
rect 45328 349109 45334 349121
rect 42410 349081 45334 349109
rect 42410 349069 42416 349081
rect 45328 349069 45334 349081
rect 45386 349069 45392 349121
rect 650416 345591 650422 345643
rect 650474 345631 650480 345643
rect 679792 345631 679798 345643
rect 650474 345603 679798 345631
rect 650474 345591 650480 345603
rect 679792 345591 679798 345603
rect 679850 345591 679856 345643
rect 674608 340929 674614 340981
rect 674666 340969 674672 340981
rect 675472 340969 675478 340981
rect 674666 340941 675478 340969
rect 674666 340929 674672 340941
rect 675472 340929 675478 340941
rect 675530 340929 675536 340981
rect 53296 339819 53302 339871
rect 53354 339859 53360 339871
rect 59536 339859 59542 339871
rect 53354 339831 59542 339859
rect 53354 339819 53360 339831
rect 59536 339819 59542 339831
rect 59594 339819 59600 339871
rect 654448 339819 654454 339871
rect 654506 339859 654512 339871
rect 666736 339859 666742 339871
rect 654506 339831 666742 339859
rect 654506 339819 654512 339831
rect 666736 339819 666742 339831
rect 666794 339819 666800 339871
rect 674032 339523 674038 339575
rect 674090 339563 674096 339575
rect 675376 339563 675382 339575
rect 674090 339535 675382 339563
rect 674090 339523 674096 339535
rect 675376 339523 675382 339535
rect 675434 339523 675440 339575
rect 674512 336563 674518 336615
rect 674570 336603 674576 336615
rect 675376 336603 675382 336615
rect 674570 336575 675382 336603
rect 674570 336563 674576 336575
rect 675376 336563 675382 336575
rect 675434 336563 675440 336615
rect 674320 332715 674326 332767
rect 674378 332755 674384 332767
rect 675376 332755 675382 332767
rect 674378 332727 675382 332755
rect 674378 332715 674384 332727
rect 675376 332715 675382 332727
rect 675434 332715 675440 332767
rect 674224 332197 674230 332249
rect 674282 332237 674288 332249
rect 675472 332237 675478 332249
rect 674282 332209 675478 332237
rect 674282 332197 674288 332209
rect 675472 332197 675478 332209
rect 675530 332197 675536 332249
rect 42160 331975 42166 332027
rect 42218 332015 42224 332027
rect 47920 332015 47926 332027
rect 42218 331987 47926 332015
rect 42218 331975 42224 331987
rect 47920 331975 47926 331987
rect 47978 331975 47984 332027
rect 674128 331531 674134 331583
rect 674186 331571 674192 331583
rect 675376 331571 675382 331583
rect 674186 331543 675382 331571
rect 674186 331531 674192 331543
rect 675376 331531 675382 331543
rect 675434 331531 675440 331583
rect 39952 331161 39958 331213
rect 40010 331201 40016 331213
rect 41776 331201 41782 331213
rect 40010 331173 41782 331201
rect 40010 331161 40016 331173
rect 41776 331161 41782 331173
rect 41834 331161 41840 331213
rect 37168 330421 37174 330473
rect 37226 330461 37232 330473
rect 40528 330461 40534 330473
rect 37226 330433 40534 330461
rect 37226 330421 37232 330433
rect 40528 330421 40534 330433
rect 40586 330421 40592 330473
rect 654064 329607 654070 329659
rect 654122 329647 654128 329659
rect 663760 329647 663766 329659
rect 654122 329619 663766 329647
rect 654122 329607 654128 329619
rect 663760 329607 663766 329619
rect 663818 329607 663824 329659
rect 40240 328497 40246 328549
rect 40298 328537 40304 328549
rect 43024 328537 43030 328549
rect 40298 328509 43030 328537
rect 40298 328497 40304 328509
rect 43024 328497 43030 328509
rect 43082 328497 43088 328549
rect 40048 328349 40054 328401
rect 40106 328389 40112 328401
rect 40106 328361 42494 328389
rect 40106 328349 40112 328361
rect 42466 328315 42494 328361
rect 42466 328287 42974 328315
rect 42946 328093 42974 328287
rect 43120 328275 43126 328327
rect 43178 328315 43184 328327
rect 43312 328315 43318 328327
rect 43178 328287 43318 328315
rect 43178 328275 43184 328287
rect 43312 328275 43318 328287
rect 43370 328275 43376 328327
rect 43024 328093 43030 328105
rect 42946 328065 43030 328093
rect 43024 328053 43030 328065
rect 43082 328053 43088 328105
rect 40528 327313 40534 327365
rect 40586 327353 40592 327365
rect 42352 327353 42358 327365
rect 40586 327325 42358 327353
rect 40586 327313 40592 327325
rect 42352 327313 42358 327325
rect 42410 327313 42416 327365
rect 41776 327017 41782 327069
rect 41834 327017 41840 327069
rect 41794 326773 41822 327017
rect 41776 326721 41782 326773
rect 41834 326721 41840 326773
rect 53392 325463 53398 325515
rect 53450 325503 53456 325515
rect 59536 325503 59542 325515
rect 53450 325475 59542 325503
rect 53450 325463 53456 325475
rect 59536 325463 59542 325475
rect 59594 325463 59600 325515
rect 42064 324871 42070 324923
rect 42122 324911 42128 324923
rect 42736 324911 42742 324923
rect 42122 324883 42742 324911
rect 42122 324871 42128 324883
rect 42736 324871 42742 324883
rect 42794 324871 42800 324923
rect 42448 324353 42454 324405
rect 42506 324393 42512 324405
rect 43312 324393 43318 324405
rect 42506 324365 43318 324393
rect 42506 324353 42512 324365
rect 43312 324353 43318 324365
rect 43370 324353 43376 324405
rect 42160 324131 42166 324183
rect 42218 324171 42224 324183
rect 53200 324171 53206 324183
rect 42218 324143 53206 324171
rect 42218 324131 42224 324143
rect 53200 324131 53206 324143
rect 53258 324131 53264 324183
rect 42160 323095 42166 323147
rect 42218 323135 42224 323147
rect 42352 323135 42358 323147
rect 42218 323107 42358 323135
rect 42218 323095 42224 323107
rect 42352 323095 42358 323107
rect 42410 323095 42416 323147
rect 42064 321763 42070 321815
rect 42122 321803 42128 321815
rect 43120 321803 43126 321815
rect 42122 321775 43126 321803
rect 42122 321763 42128 321775
rect 43120 321763 43126 321775
rect 43178 321763 43184 321815
rect 42160 321023 42166 321075
rect 42218 321063 42224 321075
rect 43024 321063 43030 321075
rect 42218 321035 43030 321063
rect 42218 321023 42224 321035
rect 43024 321023 43030 321035
rect 43082 321023 43088 321075
rect 42160 320579 42166 320631
rect 42218 320619 42224 320631
rect 42448 320619 42454 320631
rect 42218 320591 42454 320619
rect 42218 320579 42224 320591
rect 42448 320579 42454 320591
rect 42506 320579 42512 320631
rect 655216 319691 655222 319743
rect 655274 319731 655280 319743
rect 674416 319731 674422 319743
rect 655274 319703 674422 319731
rect 655274 319691 655280 319703
rect 674416 319691 674422 319703
rect 674474 319691 674480 319743
rect 666640 318877 666646 318929
rect 666698 318917 666704 318929
rect 674416 318917 674422 318929
rect 666698 318889 674422 318917
rect 666698 318877 666704 318889
rect 674416 318877 674422 318889
rect 674474 318877 674480 318929
rect 666832 318285 666838 318337
rect 666890 318325 666896 318337
rect 674704 318325 674710 318337
rect 666890 318297 674710 318325
rect 666890 318285 666896 318297
rect 674704 318285 674710 318297
rect 674762 318285 674768 318337
rect 45328 311033 45334 311085
rect 45386 311073 45392 311085
rect 59536 311073 59542 311085
rect 45386 311045 59542 311073
rect 45386 311033 45392 311045
rect 59536 311033 59542 311045
rect 59594 311033 59600 311085
rect 42256 307481 42262 307533
rect 42314 307521 42320 307533
rect 45424 307521 45430 307533
rect 42314 307493 45430 307521
rect 42314 307481 42320 307493
rect 45424 307481 45430 307493
rect 45482 307481 45488 307533
rect 42256 306741 42262 306793
rect 42314 306781 42320 306793
rect 50512 306781 50518 306793
rect 42314 306753 50518 306781
rect 42314 306741 42320 306753
rect 50512 306741 50518 306753
rect 50570 306741 50576 306793
rect 42832 305483 42838 305535
rect 42890 305523 42896 305535
rect 58960 305523 58966 305535
rect 42890 305495 58966 305523
rect 42890 305483 42896 305495
rect 58960 305483 58966 305495
rect 59018 305483 59024 305535
rect 650512 299563 650518 299615
rect 650570 299603 650576 299615
rect 679792 299603 679798 299615
rect 650570 299575 679798 299603
rect 650570 299563 650576 299575
rect 679792 299563 679798 299575
rect 679850 299563 679856 299615
rect 674800 299489 674806 299541
rect 674858 299529 674864 299541
rect 676816 299529 676822 299541
rect 674858 299501 676822 299529
rect 674858 299489 674864 299501
rect 676816 299489 676822 299501
rect 676874 299489 676880 299541
rect 674896 299415 674902 299467
rect 674954 299455 674960 299467
rect 676912 299455 676918 299467
rect 674954 299427 676918 299455
rect 674954 299415 674960 299427
rect 676912 299415 676918 299427
rect 676970 299415 676976 299467
rect 675280 299341 675286 299393
rect 675338 299381 675344 299393
rect 677104 299381 677110 299393
rect 675338 299353 677110 299381
rect 675338 299341 675344 299353
rect 677104 299341 677110 299353
rect 677162 299341 677168 299393
rect 45424 296677 45430 296729
rect 45482 296717 45488 296729
rect 59536 296717 59542 296729
rect 45482 296689 59542 296717
rect 45482 296677 45488 296689
rect 59536 296677 59542 296689
rect 59594 296677 59600 296729
rect 674320 295937 674326 295989
rect 674378 295977 674384 295989
rect 675376 295977 675382 295989
rect 674378 295949 675382 295977
rect 674378 295937 674384 295949
rect 675376 295937 675382 295949
rect 675434 295937 675440 295989
rect 674512 295345 674518 295397
rect 674570 295385 674576 295397
rect 675472 295385 675478 295397
rect 674570 295357 675478 295385
rect 674570 295345 674576 295357
rect 675472 295345 675478 295357
rect 675530 295345 675536 295397
rect 673936 294531 673942 294583
rect 673994 294571 674000 294583
rect 675376 294571 675382 294583
rect 673994 294543 675382 294571
rect 673994 294531 674000 294543
rect 675376 294531 675382 294543
rect 675434 294531 675440 294583
rect 674416 291053 674422 291105
rect 674474 291093 674480 291105
rect 675088 291093 675094 291105
rect 674474 291065 675094 291093
rect 674474 291053 674480 291065
rect 675088 291053 675094 291065
rect 675146 291053 675152 291105
rect 42640 289055 42646 289107
rect 42698 289095 42704 289107
rect 48016 289095 48022 289107
rect 42698 289067 48022 289095
rect 42698 289055 42704 289067
rect 48016 289055 48022 289067
rect 48074 289055 48080 289107
rect 41968 288907 41974 288959
rect 42026 288947 42032 288959
rect 42544 288947 42550 288959
rect 42026 288919 42550 288947
rect 42026 288907 42032 288919
rect 42544 288907 42550 288919
rect 42602 288907 42608 288959
rect 674896 288537 674902 288589
rect 674954 288577 674960 288589
rect 675472 288577 675478 288589
rect 674954 288549 675478 288577
rect 674954 288537 674960 288549
rect 675472 288537 675478 288549
rect 675530 288537 675536 288589
rect 39952 287945 39958 287997
rect 40010 287985 40016 287997
rect 41776 287985 41782 287997
rect 40010 287957 41782 287985
rect 40010 287945 40016 287957
rect 41776 287945 41782 287957
rect 41834 287945 41840 287997
rect 674224 287723 674230 287775
rect 674282 287763 674288 287775
rect 675376 287763 675382 287775
rect 674282 287735 675382 287763
rect 674282 287723 674288 287735
rect 675376 287723 675382 287735
rect 675434 287723 675440 287775
rect 674800 287353 674806 287405
rect 674858 287393 674864 287405
rect 675472 287393 675478 287405
rect 674858 287365 675478 287393
rect 674858 287353 674864 287365
rect 675472 287353 675478 287365
rect 675530 287353 675536 287405
rect 37360 286835 37366 286887
rect 37418 286875 37424 286887
rect 42736 286875 42742 286887
rect 37418 286847 42742 286875
rect 37418 286835 37424 286847
rect 42736 286835 42742 286847
rect 42794 286835 42800 286887
rect 674128 286539 674134 286591
rect 674186 286579 674192 286591
rect 675376 286579 675382 286591
rect 674186 286551 675382 286579
rect 674186 286539 674192 286551
rect 675376 286539 675382 286551
rect 675434 286539 675440 286591
rect 40144 285651 40150 285703
rect 40202 285691 40208 285703
rect 43120 285691 43126 285703
rect 40202 285663 43126 285691
rect 40202 285651 40208 285663
rect 43120 285651 43126 285663
rect 43178 285651 43184 285703
rect 40240 285133 40246 285185
rect 40298 285173 40304 285185
rect 42640 285173 42646 285185
rect 40298 285145 42646 285173
rect 40298 285133 40304 285145
rect 42640 285133 42646 285145
rect 42698 285133 42704 285185
rect 41776 283801 41782 283853
rect 41834 283801 41840 283853
rect 42160 283801 42166 283853
rect 42218 283841 42224 283853
rect 43312 283841 43318 283853
rect 42218 283813 43318 283841
rect 42218 283801 42224 283813
rect 43312 283801 43318 283813
rect 43370 283801 43376 283853
rect 41794 283409 41822 283801
rect 41776 283357 41782 283409
rect 41834 283357 41840 283409
rect 654448 282987 654454 283039
rect 654506 283027 654512 283039
rect 660880 283027 660886 283039
rect 654506 282999 660886 283027
rect 654506 282987 654512 282999
rect 660880 282987 660886 282999
rect 660938 282987 660944 283039
rect 45520 282247 45526 282299
rect 45578 282287 45584 282299
rect 59536 282287 59542 282299
rect 45578 282259 59542 282287
rect 45578 282247 45584 282259
rect 59536 282247 59542 282259
rect 59594 282247 59600 282299
rect 42160 281729 42166 281781
rect 42218 281769 42224 281781
rect 42544 281769 42550 281781
rect 42218 281741 42550 281769
rect 42218 281729 42224 281741
rect 42544 281729 42550 281741
rect 42602 281729 42608 281781
rect 42160 281063 42166 281115
rect 42218 281103 42224 281115
rect 47536 281103 47542 281115
rect 42218 281075 47542 281103
rect 42218 281063 42224 281075
rect 47536 281063 47542 281075
rect 47594 281063 47600 281115
rect 42160 279879 42166 279931
rect 42218 279919 42224 279931
rect 42736 279919 42742 279931
rect 42218 279891 42742 279919
rect 42218 279879 42224 279891
rect 42736 279879 42742 279891
rect 42794 279879 42800 279931
rect 42160 278547 42166 278599
rect 42218 278587 42224 278599
rect 42640 278587 42646 278599
rect 42218 278559 42646 278587
rect 42218 278547 42224 278559
rect 42640 278547 42646 278559
rect 42698 278547 42704 278599
rect 42160 277807 42166 277859
rect 42218 277847 42224 277859
rect 43120 277847 43126 277859
rect 42218 277819 43126 277847
rect 42218 277807 42224 277819
rect 43120 277807 43126 277819
rect 43178 277807 43184 277859
rect 43216 277807 43222 277859
rect 43274 277807 43280 277859
rect 43234 277637 43262 277807
rect 43216 277585 43222 277637
rect 43274 277585 43280 277637
rect 42064 277363 42070 277415
rect 42122 277403 42128 277415
rect 42832 277403 42838 277415
rect 42122 277375 42838 277403
rect 42122 277363 42128 277375
rect 42832 277363 42838 277375
rect 42890 277363 42896 277415
rect 303376 276327 303382 276379
rect 303434 276367 303440 276379
rect 435376 276367 435382 276379
rect 303434 276339 435382 276367
rect 303434 276327 303440 276339
rect 435376 276327 435382 276339
rect 435434 276327 435440 276379
rect 117232 276253 117238 276305
rect 117290 276293 117296 276305
rect 397552 276293 397558 276305
rect 117290 276265 397558 276293
rect 117290 276253 117296 276265
rect 397552 276253 397558 276265
rect 397610 276253 397616 276305
rect 120784 276179 120790 276231
rect 120842 276219 120848 276231
rect 398512 276219 398518 276231
rect 120842 276191 398518 276219
rect 120842 276179 120848 276191
rect 398512 276179 398518 276191
rect 398570 276179 398576 276231
rect 73264 276105 73270 276157
rect 73322 276145 73328 276157
rect 386320 276145 386326 276157
rect 73322 276117 386326 276145
rect 73322 276105 73328 276117
rect 386320 276105 386326 276117
rect 386378 276105 386384 276157
rect 113776 276031 113782 276083
rect 113834 276071 113840 276083
rect 396784 276071 396790 276083
rect 113834 276043 396790 276071
rect 113834 276031 113840 276043
rect 396784 276031 396790 276043
rect 396842 276031 396848 276083
rect 303568 275957 303574 276009
rect 303626 275997 303632 276009
rect 439024 275997 439030 276009
rect 303626 275969 439030 275997
rect 303626 275957 303632 275969
rect 439024 275957 439030 275969
rect 439082 275957 439088 276009
rect 303952 275883 303958 275935
rect 304010 275923 304016 275935
rect 442576 275923 442582 275935
rect 304010 275895 442582 275923
rect 304010 275883 304016 275895
rect 442576 275883 442582 275895
rect 442634 275883 442640 275935
rect 304432 275809 304438 275861
rect 304490 275849 304496 275861
rect 446320 275849 446326 275861
rect 304490 275821 446326 275849
rect 304490 275809 304496 275821
rect 446320 275809 446326 275821
rect 446378 275809 446384 275861
rect 305104 275735 305110 275787
rect 305162 275775 305168 275787
rect 449680 275775 449686 275787
rect 305162 275747 449686 275775
rect 305162 275735 305168 275747
rect 449680 275735 449686 275747
rect 449738 275735 449744 275787
rect 305200 275661 305206 275713
rect 305258 275701 305264 275713
rect 453232 275701 453238 275713
rect 305258 275673 453238 275701
rect 305258 275661 305264 275673
rect 453232 275661 453238 275673
rect 453290 275661 453296 275713
rect 421840 275587 421846 275639
rect 421898 275627 421904 275639
rect 649456 275627 649462 275639
rect 421898 275599 649462 275627
rect 421898 275587 421904 275599
rect 649456 275587 649462 275599
rect 649514 275587 649520 275639
rect 306640 275513 306646 275565
rect 306698 275553 306704 275565
rect 464368 275553 464374 275565
rect 306698 275525 464374 275553
rect 306698 275513 306704 275525
rect 464368 275513 464374 275525
rect 464426 275513 464432 275565
rect 307216 275439 307222 275491
rect 307274 275479 307280 275491
rect 467824 275479 467830 275491
rect 307274 275451 467830 275479
rect 307274 275439 307280 275451
rect 467824 275439 467830 275451
rect 467882 275439 467888 275491
rect 307696 275365 307702 275417
rect 307754 275405 307760 275417
rect 471376 275405 471382 275417
rect 307754 275377 471382 275405
rect 307754 275365 307760 275377
rect 471376 275365 471382 275377
rect 471434 275365 471440 275417
rect 307888 275291 307894 275343
rect 307946 275331 307952 275343
rect 475024 275331 475030 275343
rect 307946 275303 475030 275331
rect 307946 275291 307952 275303
rect 475024 275291 475030 275303
rect 475082 275291 475088 275343
rect 308368 275217 308374 275269
rect 308426 275257 308432 275269
rect 478576 275257 478582 275269
rect 308426 275229 478582 275257
rect 308426 275217 308432 275229
rect 478576 275217 478582 275229
rect 478634 275217 478640 275269
rect 308752 275143 308758 275195
rect 308810 275183 308816 275195
rect 481840 275183 481846 275195
rect 308810 275155 481846 275183
rect 308810 275143 308816 275155
rect 481840 275143 481846 275155
rect 481898 275143 481904 275195
rect 309424 275069 309430 275121
rect 309482 275109 309488 275121
rect 485680 275109 485686 275121
rect 309482 275081 485686 275109
rect 309482 275069 309488 275081
rect 485680 275069 485686 275081
rect 485738 275069 485744 275121
rect 64912 274995 64918 275047
rect 64970 275035 64976 275047
rect 181360 275035 181366 275047
rect 64970 275007 181366 275035
rect 64970 274995 64976 275007
rect 181360 274995 181366 275007
rect 181418 274995 181424 275047
rect 309904 274995 309910 275047
rect 309962 275035 309968 275047
rect 489232 275035 489238 275047
rect 309962 275007 489238 275035
rect 309962 274995 309968 275007
rect 489232 274995 489238 275007
rect 489290 274995 489296 275047
rect 573136 274995 573142 275047
rect 573194 275035 573200 275047
rect 649360 275035 649366 275047
rect 573194 275007 649366 275035
rect 573194 274995 573200 275007
rect 649360 274995 649366 275007
rect 649418 274995 649424 275047
rect 310096 274921 310102 274973
rect 310154 274961 310160 274973
rect 492880 274961 492886 274973
rect 310154 274933 492886 274961
rect 310154 274921 310160 274933
rect 492880 274921 492886 274933
rect 492938 274921 492944 274973
rect 669712 274921 669718 274973
rect 669770 274961 669776 274973
rect 674704 274961 674710 274973
rect 669770 274933 674710 274961
rect 669770 274921 669776 274933
rect 674704 274921 674710 274933
rect 674762 274921 674768 274973
rect 310480 274847 310486 274899
rect 310538 274887 310544 274899
rect 496432 274887 496438 274899
rect 310538 274859 496438 274887
rect 310538 274847 310544 274859
rect 496432 274847 496438 274859
rect 496490 274847 496496 274899
rect 311632 274773 311638 274825
rect 311690 274813 311696 274825
rect 503536 274813 503542 274825
rect 311690 274785 503542 274813
rect 311690 274773 311696 274785
rect 503536 274773 503542 274785
rect 503594 274773 503600 274825
rect 310960 274699 310966 274751
rect 311018 274739 311024 274751
rect 499888 274739 499894 274751
rect 311018 274711 499894 274739
rect 311018 274699 311024 274711
rect 499888 274699 499894 274711
rect 499946 274699 499952 274751
rect 42256 274625 42262 274677
rect 42314 274665 42320 274677
rect 42736 274665 42742 274677
rect 42314 274637 42742 274665
rect 42314 274625 42320 274637
rect 42736 274625 42742 274637
rect 42794 274625 42800 274677
rect 312112 274625 312118 274677
rect 312170 274665 312176 274677
rect 507088 274665 507094 274677
rect 312170 274637 507094 274665
rect 312170 274625 312176 274637
rect 507088 274625 507094 274637
rect 507146 274625 507152 274677
rect 312208 274551 312214 274603
rect 312266 274591 312272 274603
rect 510736 274591 510742 274603
rect 312266 274563 510742 274591
rect 312266 274551 312272 274563
rect 510736 274551 510742 274563
rect 510794 274551 510800 274603
rect 312688 274477 312694 274529
rect 312746 274517 312752 274529
rect 514288 274517 514294 274529
rect 312746 274489 514294 274517
rect 312746 274477 312752 274489
rect 514288 274477 514294 274489
rect 514346 274477 514352 274529
rect 313168 274403 313174 274455
rect 313226 274443 313232 274455
rect 517744 274443 517750 274455
rect 313226 274415 517750 274443
rect 313226 274403 313232 274415
rect 517744 274403 517750 274415
rect 517802 274403 517808 274455
rect 313744 274329 313750 274381
rect 313802 274369 313808 274381
rect 521392 274369 521398 274381
rect 313802 274341 521398 274369
rect 313802 274329 313808 274341
rect 521392 274329 521398 274341
rect 521450 274329 521456 274381
rect 314704 274255 314710 274307
rect 314762 274295 314768 274307
rect 528208 274295 528214 274307
rect 314762 274267 528214 274295
rect 314762 274255 314768 274267
rect 528208 274255 528214 274267
rect 528266 274255 528272 274307
rect 314896 274181 314902 274233
rect 314954 274221 314960 274233
rect 532144 274221 532150 274233
rect 314954 274193 532150 274221
rect 314954 274181 314960 274193
rect 532144 274181 532150 274193
rect 532202 274181 532208 274233
rect 42064 274107 42070 274159
rect 42122 274147 42128 274159
rect 43024 274147 43030 274159
rect 42122 274119 43030 274147
rect 42122 274107 42128 274119
rect 43024 274107 43030 274119
rect 43082 274107 43088 274159
rect 315280 274107 315286 274159
rect 315338 274147 315344 274159
rect 535600 274147 535606 274159
rect 315338 274119 535606 274147
rect 315338 274107 315344 274119
rect 535600 274107 535606 274119
rect 535658 274107 535664 274159
rect 315952 274033 315958 274085
rect 316010 274073 316016 274085
rect 539248 274073 539254 274085
rect 316010 274045 539254 274073
rect 316010 274033 316016 274045
rect 539248 274033 539254 274045
rect 539306 274033 539312 274085
rect 663856 274033 663862 274085
rect 663914 274073 663920 274085
rect 674704 274073 674710 274085
rect 663914 274045 674710 274073
rect 663914 274033 663920 274045
rect 674704 274033 674710 274045
rect 674762 274033 674768 274085
rect 316432 273959 316438 274011
rect 316490 273999 316496 274011
rect 542800 273999 542806 274011
rect 316490 273971 542806 273999
rect 316490 273959 316496 273971
rect 542800 273959 542806 273971
rect 542858 273959 542864 274011
rect 316624 273885 316630 273937
rect 316682 273925 316688 273937
rect 546352 273925 546358 273937
rect 316682 273897 546358 273925
rect 316682 273885 316688 273897
rect 546352 273885 546358 273897
rect 546410 273885 546416 273937
rect 358288 273811 358294 273863
rect 358346 273851 358352 273863
rect 429808 273851 429814 273863
rect 358346 273823 429814 273851
rect 358346 273811 358352 273823
rect 429808 273811 429814 273823
rect 429866 273811 429872 273863
rect 42256 273737 42262 273789
rect 42314 273777 42320 273789
rect 43120 273777 43126 273789
rect 42314 273749 43126 273777
rect 42314 273737 42320 273749
rect 43120 273737 43126 273749
rect 43178 273737 43184 273789
rect 302896 273737 302902 273789
rect 302954 273777 302960 273789
rect 432208 273777 432214 273789
rect 302954 273749 432214 273777
rect 302954 273737 302960 273749
rect 432208 273737 432214 273749
rect 432266 273737 432272 273789
rect 262096 273663 262102 273715
rect 262154 273703 262160 273715
rect 337552 273703 337558 273715
rect 262154 273675 337558 273703
rect 262154 273663 262160 273675
rect 337552 273663 337558 273675
rect 337610 273663 337616 273715
rect 358384 273663 358390 273715
rect 358442 273703 358448 273715
rect 433360 273703 433366 273715
rect 358442 273675 433366 273703
rect 358442 273663 358448 273675
rect 433360 273663 433366 273675
rect 433418 273663 433424 273715
rect 306160 273589 306166 273641
rect 306218 273629 306224 273641
rect 460720 273629 460726 273641
rect 306218 273601 460726 273629
rect 306218 273589 306224 273601
rect 460720 273589 460726 273601
rect 460778 273589 460784 273641
rect 239728 273515 239734 273567
rect 239786 273555 239792 273567
rect 370288 273555 370294 273567
rect 239786 273527 370294 273555
rect 239786 273515 239792 273527
rect 370288 273515 370294 273527
rect 370346 273515 370352 273567
rect 375664 273515 375670 273567
rect 375722 273555 375728 273567
rect 488080 273555 488086 273567
rect 375722 273527 488086 273555
rect 375722 273515 375728 273527
rect 488080 273515 488086 273527
rect 488138 273515 488144 273567
rect 240400 273441 240406 273493
rect 240458 273481 240464 273493
rect 377488 273481 377494 273493
rect 240458 273453 377494 273481
rect 240458 273441 240464 273453
rect 377488 273441 377494 273453
rect 377546 273441 377552 273493
rect 380656 273441 380662 273493
rect 380714 273481 380720 273493
rect 550096 273481 550102 273493
rect 380714 273453 550102 273481
rect 380714 273441 380720 273453
rect 550096 273441 550102 273453
rect 550154 273441 550160 273493
rect 241456 273367 241462 273419
rect 241514 273407 241520 273419
rect 384592 273407 384598 273419
rect 241514 273379 384598 273407
rect 241514 273367 241520 273379
rect 384592 273367 384598 273379
rect 384650 273367 384656 273419
rect 242128 273293 242134 273345
rect 242186 273333 242192 273345
rect 391696 273333 391702 273345
rect 242186 273305 391702 273333
rect 242186 273293 242192 273305
rect 391696 273293 391702 273305
rect 391754 273293 391760 273345
rect 664048 273293 664054 273345
rect 664106 273333 664112 273345
rect 674704 273333 674710 273345
rect 664106 273305 674710 273333
rect 664106 273293 664112 273305
rect 674704 273293 674710 273305
rect 674762 273293 674768 273345
rect 243184 273219 243190 273271
rect 243242 273259 243248 273271
rect 398896 273259 398902 273271
rect 243242 273231 398902 273259
rect 243242 273219 243248 273231
rect 398896 273219 398902 273231
rect 398954 273219 398960 273271
rect 243856 273145 243862 273197
rect 243914 273185 243920 273197
rect 406000 273185 406006 273197
rect 243914 273157 406006 273185
rect 243914 273145 243920 273157
rect 406000 273145 406006 273157
rect 406058 273145 406064 273197
rect 244720 273071 244726 273123
rect 244778 273111 244784 273123
rect 413200 273111 413206 273123
rect 244778 273083 413206 273111
rect 244778 273071 244784 273083
rect 413200 273071 413206 273083
rect 413258 273071 413264 273123
rect 245872 272997 245878 273049
rect 245930 273037 245936 273049
rect 419920 273037 419926 273049
rect 245930 273009 419926 273037
rect 245930 272997 245936 273009
rect 419920 272997 419926 273009
rect 419978 272997 419984 273049
rect 246448 272923 246454 272975
rect 246506 272963 246512 272975
rect 427408 272963 427414 272975
rect 246506 272935 427414 272963
rect 246506 272923 246512 272935
rect 427408 272923 427414 272935
rect 427466 272923 427472 272975
rect 247600 272849 247606 272901
rect 247658 272889 247664 272901
rect 434512 272889 434518 272901
rect 247658 272861 434518 272889
rect 247658 272849 247664 272861
rect 434512 272849 434518 272861
rect 434570 272849 434576 272901
rect 229072 272775 229078 272827
rect 229130 272815 229136 272827
rect 284656 272815 284662 272827
rect 229130 272787 284662 272815
rect 229130 272775 229136 272787
rect 284656 272775 284662 272787
rect 284714 272775 284720 272827
rect 322096 272775 322102 272827
rect 322154 272815 322160 272827
rect 322154 272787 327806 272815
rect 322154 272775 322160 272787
rect 230128 272701 230134 272753
rect 230186 272741 230192 272753
rect 291856 272741 291862 272753
rect 230186 272713 291862 272741
rect 230186 272701 230192 272713
rect 291856 272701 291862 272713
rect 291914 272701 291920 272753
rect 322960 272701 322966 272753
rect 323018 272741 323024 272753
rect 327778 272741 327806 272787
rect 327856 272775 327862 272827
rect 327914 272815 327920 272827
rect 582064 272815 582070 272827
rect 327914 272787 582070 272815
rect 327914 272775 327920 272787
rect 582064 272775 582070 272787
rect 582122 272775 582128 272827
rect 589168 272741 589174 272753
rect 323018 272713 327710 272741
rect 327778 272713 589174 272741
rect 323018 272701 323024 272713
rect 230800 272627 230806 272679
rect 230858 272667 230864 272679
rect 298960 272667 298966 272679
rect 230858 272639 298966 272667
rect 230858 272627 230864 272639
rect 298960 272627 298966 272639
rect 299018 272627 299024 272679
rect 323536 272627 323542 272679
rect 323594 272667 323600 272679
rect 327682 272667 327710 272713
rect 589168 272701 589174 272713
rect 589226 272701 589232 272753
rect 596368 272667 596374 272679
rect 323594 272639 327614 272667
rect 327682 272639 596374 272667
rect 323594 272627 323600 272639
rect 231856 272553 231862 272605
rect 231914 272593 231920 272605
rect 306064 272593 306070 272605
rect 231914 272565 306070 272593
rect 231914 272553 231920 272565
rect 306064 272553 306070 272565
rect 306122 272553 306128 272605
rect 324688 272553 324694 272605
rect 324746 272593 324752 272605
rect 327586 272593 327614 272639
rect 596368 272627 596374 272639
rect 596426 272627 596432 272679
rect 603472 272593 603478 272605
rect 324746 272565 327518 272593
rect 327586 272565 603478 272593
rect 324746 272553 324752 272565
rect 64816 272479 64822 272531
rect 64874 272519 64880 272531
rect 72016 272519 72022 272531
rect 64874 272491 72022 272519
rect 64874 272479 64880 272491
rect 72016 272479 72022 272491
rect 72074 272479 72080 272531
rect 261040 272479 261046 272531
rect 261098 272519 261104 272531
rect 327376 272519 327382 272531
rect 261098 272491 327382 272519
rect 261098 272479 261104 272491
rect 327376 272479 327382 272491
rect 327434 272479 327440 272531
rect 232720 272405 232726 272457
rect 232778 272445 232784 272457
rect 313264 272445 313270 272457
rect 232778 272417 313270 272445
rect 232778 272405 232784 272417
rect 313264 272405 313270 272417
rect 313322 272405 313328 272457
rect 325264 272405 325270 272457
rect 325322 272445 325328 272457
rect 327490 272445 327518 272565
rect 603472 272553 603478 272565
rect 603530 272553 603536 272605
rect 327568 272479 327574 272531
rect 327626 272519 327632 272531
rect 545200 272519 545206 272531
rect 327626 272491 545206 272519
rect 327626 272479 327632 272491
rect 545200 272479 545206 272491
rect 545258 272479 545264 272531
rect 610576 272445 610582 272457
rect 325322 272417 327422 272445
rect 327490 272417 610582 272445
rect 325322 272405 325328 272417
rect 233392 272331 233398 272383
rect 233450 272371 233456 272383
rect 320368 272371 320374 272383
rect 233450 272343 320374 272371
rect 233450 272331 233456 272343
rect 320368 272331 320374 272343
rect 320426 272331 320432 272383
rect 326224 272331 326230 272383
rect 326282 272371 326288 272383
rect 327394 272371 327422 272417
rect 610576 272405 610582 272417
rect 610634 272405 610640 272457
rect 617680 272371 617686 272383
rect 326282 272343 327326 272371
rect 327394 272343 617686 272371
rect 326282 272331 326288 272343
rect 64720 272257 64726 272309
rect 64778 272297 64784 272309
rect 66832 272297 66838 272309
rect 64778 272269 66838 272297
rect 64778 272257 64784 272269
rect 66832 272257 66838 272269
rect 66890 272257 66896 272309
rect 234448 272257 234454 272309
rect 234506 272297 234512 272309
rect 327184 272297 327190 272309
rect 234506 272269 327190 272297
rect 234506 272257 234512 272269
rect 327184 272257 327190 272269
rect 327242 272257 327248 272309
rect 327298 272297 327326 272343
rect 617680 272331 617686 272343
rect 617738 272331 617744 272383
rect 624880 272297 624886 272309
rect 327298 272269 624886 272297
rect 624880 272257 624886 272269
rect 624938 272257 624944 272309
rect 266512 272183 266518 272235
rect 266570 272223 266576 272235
rect 591568 272223 591574 272235
rect 266570 272195 591574 272223
rect 266570 272183 266576 272195
rect 591568 272183 591574 272195
rect 591626 272183 591632 272235
rect 267184 272109 267190 272161
rect 267242 272149 267248 272161
rect 595120 272149 595126 272161
rect 267242 272121 595126 272149
rect 267242 272109 267248 272121
rect 595120 272109 595126 272121
rect 595178 272109 595184 272161
rect 228112 272035 228118 272087
rect 228170 272075 228176 272087
rect 277552 272075 277558 272087
rect 228170 272047 277558 272075
rect 228170 272035 228176 272047
rect 277552 272035 277558 272047
rect 277610 272035 277616 272087
rect 302224 272035 302230 272087
rect 302282 272075 302288 272087
rect 428656 272075 428662 272087
rect 302282 272047 428662 272075
rect 302282 272035 302288 272047
rect 428656 272035 428662 272047
rect 428714 272035 428720 272087
rect 238864 271961 238870 272013
rect 238922 272001 238928 272013
rect 363184 272001 363190 272013
rect 238922 271973 363190 272001
rect 238922 271961 238928 271973
rect 363184 271961 363190 271973
rect 363242 271961 363248 272013
rect 364624 271961 364630 272013
rect 364682 272001 364688 272013
rect 393040 272001 393046 272013
rect 364682 271973 393046 272001
rect 364682 271961 364688 271973
rect 393040 271961 393046 271973
rect 393098 271961 393104 272013
rect 227920 271887 227926 271939
rect 227978 271927 227984 271939
rect 274000 271927 274006 271939
rect 227978 271899 274006 271927
rect 227978 271887 227984 271899
rect 274000 271887 274006 271899
rect 274058 271887 274064 271939
rect 301360 271887 301366 271939
rect 301418 271927 301424 271939
rect 387472 271927 387478 271939
rect 301418 271899 387478 271927
rect 301418 271887 301424 271899
rect 387472 271887 387478 271899
rect 387530 271887 387536 271939
rect 387664 271887 387670 271939
rect 387722 271927 387728 271939
rect 421456 271927 421462 271939
rect 387722 271899 421462 271927
rect 387722 271887 387728 271899
rect 421456 271887 421462 271899
rect 421514 271887 421520 271939
rect 237712 271813 237718 271865
rect 237770 271853 237776 271865
rect 356080 271853 356086 271865
rect 237770 271825 356086 271853
rect 237770 271813 237776 271825
rect 356080 271813 356086 271825
rect 356138 271813 356144 271865
rect 374128 271813 374134 271865
rect 374186 271853 374192 271865
rect 387376 271853 387382 271865
rect 374186 271825 387382 271853
rect 374186 271813 374192 271825
rect 387376 271813 387382 271825
rect 387434 271813 387440 271865
rect 393040 271813 393046 271865
rect 393098 271853 393104 271865
rect 426256 271853 426262 271865
rect 393098 271825 426262 271853
rect 393098 271813 393104 271825
rect 426256 271813 426262 271825
rect 426314 271813 426320 271865
rect 237136 271739 237142 271791
rect 237194 271779 237200 271791
rect 348976 271779 348982 271791
rect 237194 271751 348982 271779
rect 237194 271739 237200 271751
rect 348976 271739 348982 271751
rect 349034 271739 349040 271791
rect 356272 271739 356278 271791
rect 356330 271779 356336 271791
rect 415600 271779 415606 271791
rect 356330 271751 415606 271779
rect 356330 271739 356336 271751
rect 415600 271739 415606 271751
rect 415658 271739 415664 271791
rect 227440 271665 227446 271717
rect 227498 271705 227504 271717
rect 270352 271705 270358 271717
rect 227498 271677 270358 271705
rect 227498 271665 227504 271677
rect 270352 271665 270358 271677
rect 270410 271665 270416 271717
rect 300304 271665 300310 271717
rect 300362 271705 300368 271717
rect 410800 271705 410806 271717
rect 300362 271677 410806 271705
rect 300362 271665 300368 271677
rect 410800 271665 410806 271677
rect 410858 271665 410864 271717
rect 299152 271591 299158 271643
rect 299210 271631 299216 271643
rect 403600 271631 403606 271643
rect 299210 271603 403606 271631
rect 299210 271591 299216 271603
rect 403600 271591 403606 271603
rect 403658 271591 403664 271643
rect 235984 271517 235990 271569
rect 236042 271557 236048 271569
rect 341776 271557 341782 271569
rect 236042 271529 341782 271557
rect 236042 271517 236048 271529
rect 341776 271517 341782 271529
rect 341834 271517 341840 271569
rect 362800 271517 362806 271569
rect 362858 271557 362864 271569
rect 383344 271557 383350 271569
rect 362858 271529 383350 271557
rect 362858 271517 362864 271529
rect 383344 271517 383350 271529
rect 383402 271517 383408 271569
rect 387280 271517 387286 271569
rect 387338 271557 387344 271569
rect 394768 271557 394774 271569
rect 387338 271529 394774 271557
rect 387338 271517 387344 271529
rect 394768 271517 394774 271529
rect 394826 271517 394832 271569
rect 327280 271443 327286 271495
rect 327338 271483 327344 271495
rect 588880 271483 588886 271495
rect 327338 271455 588886 271483
rect 327338 271443 327344 271455
rect 588880 271443 588886 271455
rect 588938 271443 588944 271495
rect 235120 271369 235126 271421
rect 235178 271409 235184 271421
rect 334576 271409 334582 271421
rect 235178 271381 334582 271409
rect 235178 271369 235184 271381
rect 334576 271369 334582 271381
rect 334634 271369 334640 271421
rect 378448 271369 378454 271421
rect 378506 271409 378512 271421
rect 407344 271409 407350 271421
rect 378506 271381 407350 271409
rect 378506 271369 378512 271381
rect 407344 271369 407350 271381
rect 407402 271369 407408 271421
rect 298480 271295 298486 271347
rect 298538 271335 298544 271347
rect 396496 271335 396502 271347
rect 298538 271307 396502 271335
rect 298538 271295 298544 271307
rect 396496 271295 396502 271307
rect 396554 271295 396560 271347
rect 237424 271221 237430 271273
rect 237482 271261 237488 271273
rect 331024 271261 331030 271273
rect 237482 271233 331030 271261
rect 237482 271221 237488 271233
rect 331024 271221 331030 271233
rect 331082 271221 331088 271273
rect 376240 271221 376246 271273
rect 376298 271261 376304 271273
rect 459856 271261 459862 271273
rect 376298 271233 459862 271261
rect 376298 271221 376304 271233
rect 459856 271221 459862 271233
rect 459914 271221 459920 271273
rect 294832 271147 294838 271199
rect 294890 271187 294896 271199
rect 367888 271187 367894 271199
rect 294890 271159 367894 271187
rect 294890 271147 294896 271159
rect 367888 271147 367894 271159
rect 367946 271147 367952 271199
rect 377200 271147 377206 271199
rect 377258 271187 377264 271199
rect 387280 271187 387286 271199
rect 377258 271159 387286 271187
rect 377258 271147 377264 271159
rect 387280 271147 387286 271159
rect 387338 271147 387344 271199
rect 387376 271147 387382 271199
rect 387434 271187 387440 271199
rect 472336 271187 472342 271199
rect 387434 271159 472342 271187
rect 387434 271147 387440 271159
rect 472336 271147 472342 271159
rect 472394 271147 472400 271199
rect 296560 271073 296566 271125
rect 296618 271113 296624 271125
rect 382288 271113 382294 271125
rect 296618 271085 382294 271113
rect 296618 271073 296624 271085
rect 382288 271073 382294 271085
rect 382346 271073 382352 271125
rect 295888 270999 295894 271051
rect 295946 271039 295952 271051
rect 375088 271039 375094 271051
rect 295946 271011 375094 271039
rect 295946 270999 295952 271011
rect 375088 270999 375094 271011
rect 375146 270999 375152 271051
rect 379408 270999 379414 271051
rect 379466 271039 379472 271051
rect 394672 271039 394678 271051
rect 379466 271011 394678 271039
rect 379466 270999 379472 271011
rect 394672 270999 394678 271011
rect 394730 270999 394736 271051
rect 394768 270999 394774 271051
rect 394826 271039 394832 271051
rect 502672 271039 502678 271051
rect 394826 271011 502678 271039
rect 394826 270999 394832 271011
rect 502672 270999 502678 271011
rect 502730 270999 502736 271051
rect 297424 270925 297430 270977
rect 297482 270965 297488 270977
rect 389008 270965 389014 270977
rect 297482 270937 389014 270965
rect 297482 270925 297488 270937
rect 389008 270925 389014 270937
rect 389066 270925 389072 270977
rect 247888 270851 247894 270903
rect 247946 270891 247952 270903
rect 327760 270891 327766 270903
rect 247946 270863 327766 270891
rect 247946 270851 247952 270863
rect 327760 270851 327766 270863
rect 327818 270851 327824 270903
rect 328912 270851 328918 270903
rect 328970 270891 328976 270903
rect 562192 270891 562198 270903
rect 328970 270863 562198 270891
rect 328970 270851 328976 270863
rect 562192 270851 562198 270863
rect 562250 270851 562256 270903
rect 320944 270777 320950 270829
rect 321002 270817 321008 270829
rect 327856 270817 327862 270829
rect 321002 270789 327862 270817
rect 321002 270777 321008 270789
rect 327856 270777 327862 270789
rect 327914 270777 327920 270829
rect 327952 270777 327958 270829
rect 328010 270817 328016 270829
rect 570256 270817 570262 270829
rect 328010 270789 570262 270817
rect 328010 270777 328016 270789
rect 570256 270777 570262 270789
rect 570314 270777 570320 270829
rect 216784 270703 216790 270755
rect 216842 270743 216848 270755
rect 228880 270743 228886 270755
rect 216842 270715 228886 270743
rect 216842 270703 216848 270715
rect 228880 270703 228886 270715
rect 228938 270703 228944 270755
rect 230032 270703 230038 270755
rect 230090 270743 230096 270755
rect 333328 270743 333334 270755
rect 230090 270715 333334 270743
rect 230090 270703 230096 270715
rect 333328 270703 333334 270715
rect 333386 270703 333392 270755
rect 382192 270703 382198 270755
rect 382250 270743 382256 270755
rect 382250 270715 394622 270743
rect 382250 270703 382256 270715
rect 124144 270629 124150 270681
rect 124202 270669 124208 270681
rect 220624 270669 220630 270681
rect 124202 270641 220630 270669
rect 124202 270629 124208 270641
rect 220624 270629 220630 270641
rect 220682 270629 220688 270681
rect 220720 270629 220726 270681
rect 220778 270669 220784 270681
rect 327088 270669 327094 270681
rect 220778 270641 327094 270669
rect 220778 270629 220784 270641
rect 327088 270629 327094 270641
rect 327146 270629 327152 270681
rect 329872 270629 329878 270681
rect 329930 270669 329936 270681
rect 345808 270669 345814 270681
rect 329930 270641 345814 270669
rect 329930 270629 329936 270641
rect 345808 270629 345814 270641
rect 345866 270629 345872 270681
rect 351184 270629 351190 270681
rect 351242 270669 351248 270681
rect 372688 270669 372694 270681
rect 351242 270641 372694 270669
rect 351242 270629 351248 270641
rect 372688 270629 372694 270641
rect 372746 270629 372752 270681
rect 374416 270629 374422 270681
rect 374474 270669 374480 270681
rect 387280 270669 387286 270681
rect 374474 270641 387286 270669
rect 374474 270629 374480 270641
rect 387280 270629 387286 270641
rect 387338 270629 387344 270681
rect 387376 270629 387382 270681
rect 387434 270669 387440 270681
rect 390352 270669 390358 270681
rect 387434 270641 390358 270669
rect 387434 270629 387440 270641
rect 390352 270629 390358 270641
rect 390410 270629 390416 270681
rect 394594 270669 394622 270715
rect 394672 270703 394678 270755
rect 394730 270743 394736 270755
rect 403120 270743 403126 270755
rect 394730 270715 403126 270743
rect 394730 270703 394736 270715
rect 403120 270703 403126 270715
rect 403178 270703 403184 270755
rect 626032 270669 626038 270681
rect 394594 270641 626038 270669
rect 626032 270629 626038 270641
rect 626090 270629 626096 270681
rect 105040 270555 105046 270607
rect 105098 270595 105104 270607
rect 139792 270595 139798 270607
rect 105098 270567 139798 270595
rect 105098 270555 105104 270567
rect 139792 270555 139798 270567
rect 139850 270555 139856 270607
rect 160144 270555 160150 270607
rect 160202 270595 160208 270607
rect 160202 270567 168062 270595
rect 160202 270555 160208 270567
rect 101488 270481 101494 270533
rect 101546 270521 101552 270533
rect 139888 270521 139894 270533
rect 101546 270493 139894 270521
rect 101546 270481 101552 270493
rect 139888 270481 139894 270493
rect 139946 270481 139952 270533
rect 98320 270407 98326 270459
rect 98378 270447 98384 270459
rect 139984 270447 139990 270459
rect 98378 270419 139990 270447
rect 98378 270407 98384 270419
rect 139984 270407 139990 270419
rect 140042 270407 140048 270459
rect 94384 270333 94390 270385
rect 94442 270373 94448 270385
rect 140176 270373 140182 270385
rect 94442 270345 140182 270373
rect 94442 270333 94448 270345
rect 140176 270333 140182 270345
rect 140234 270333 140240 270385
rect 89584 270259 89590 270311
rect 89642 270299 89648 270311
rect 140080 270299 140086 270311
rect 89642 270271 140086 270299
rect 89642 270259 89648 270271
rect 140080 270259 140086 270271
rect 140138 270259 140144 270311
rect 168034 270299 168062 270567
rect 176464 270555 176470 270607
rect 176522 270595 176528 270607
rect 178480 270595 178486 270607
rect 176522 270567 178486 270595
rect 176522 270555 176528 270567
rect 178480 270555 178486 270567
rect 178538 270555 178544 270607
rect 180016 270555 180022 270607
rect 180074 270595 180080 270607
rect 181360 270595 181366 270607
rect 180074 270567 181366 270595
rect 180074 270555 180080 270567
rect 181360 270555 181366 270567
rect 181418 270555 181424 270607
rect 195856 270595 195862 270607
rect 181474 270567 195862 270595
rect 172912 270481 172918 270533
rect 172970 270521 172976 270533
rect 175600 270521 175606 270533
rect 172970 270493 175606 270521
rect 172970 270481 172976 270493
rect 175600 270481 175606 270493
rect 175658 270481 175664 270533
rect 174064 270407 174070 270459
rect 174122 270447 174128 270459
rect 181474 270447 181502 270567
rect 195856 270555 195862 270567
rect 195914 270555 195920 270607
rect 206512 270555 206518 270607
rect 206570 270595 206576 270607
rect 217456 270595 217462 270607
rect 206570 270567 217462 270595
rect 206570 270555 206576 270567
rect 217456 270555 217462 270567
rect 217514 270555 217520 270607
rect 337072 270595 337078 270607
rect 228802 270567 337078 270595
rect 187024 270481 187030 270533
rect 187082 270521 187088 270533
rect 216784 270521 216790 270533
rect 187082 270493 216790 270521
rect 187082 270481 187088 270493
rect 216784 270481 216790 270493
rect 216842 270481 216848 270533
rect 216880 270481 216886 270533
rect 216938 270521 216944 270533
rect 220528 270521 220534 270533
rect 216938 270493 220534 270521
rect 216938 270481 216944 270493
rect 220528 270481 220534 270493
rect 220586 270481 220592 270533
rect 174122 270419 181502 270447
rect 174122 270407 174128 270419
rect 182416 270407 182422 270459
rect 182474 270447 182480 270459
rect 195856 270447 195862 270459
rect 182474 270419 195862 270447
rect 182474 270407 182480 270419
rect 195856 270407 195862 270419
rect 195914 270407 195920 270459
rect 196048 270407 196054 270459
rect 196106 270447 196112 270459
rect 228802 270447 228830 270567
rect 337072 270555 337078 270567
rect 337130 270555 337136 270607
rect 357040 270555 357046 270607
rect 357098 270595 357104 270607
rect 397360 270595 397366 270607
rect 357098 270567 397366 270595
rect 357098 270555 357104 270567
rect 397360 270555 397366 270567
rect 397418 270555 397424 270607
rect 397456 270555 397462 270607
rect 397514 270595 397520 270607
rect 400336 270595 400342 270607
rect 397514 270567 400342 270595
rect 397514 270555 397520 270567
rect 400336 270555 400342 270567
rect 400394 270555 400400 270607
rect 403120 270555 403126 270607
rect 403178 270595 403184 270607
rect 604624 270595 604630 270607
rect 403178 270567 604630 270595
rect 403178 270555 403184 270567
rect 604624 270555 604630 270567
rect 604682 270555 604688 270607
rect 228880 270481 228886 270533
rect 228938 270521 228944 270533
rect 405904 270521 405910 270533
rect 228938 270493 405910 270521
rect 228938 270481 228944 270493
rect 405904 270481 405910 270493
rect 405962 270481 405968 270533
rect 407344 270481 407350 270533
rect 407402 270521 407408 270533
rect 597520 270521 597526 270533
rect 407402 270493 597526 270521
rect 407402 270481 407408 270493
rect 597520 270481 597526 270493
rect 597578 270481 597584 270533
rect 196106 270419 228830 270447
rect 196106 270407 196112 270419
rect 236080 270407 236086 270459
rect 236138 270447 236144 270459
rect 337072 270447 337078 270459
rect 236138 270419 337078 270447
rect 236138 270407 236144 270419
rect 337072 270407 337078 270419
rect 337130 270407 337136 270459
rect 357040 270407 357046 270459
rect 357098 270447 357104 270459
rect 387184 270447 387190 270459
rect 357098 270419 387190 270447
rect 357098 270407 357104 270419
rect 387184 270407 387190 270419
rect 387242 270407 387248 270459
rect 387280 270407 387286 270459
rect 387338 270447 387344 270459
rect 436912 270447 436918 270459
rect 387338 270419 436918 270447
rect 387338 270407 387344 270419
rect 436912 270407 436918 270419
rect 436970 270407 436976 270459
rect 459856 270407 459862 270459
rect 459914 270447 459920 270459
rect 579664 270447 579670 270459
rect 459914 270419 579670 270447
rect 459914 270407 459920 270419
rect 579664 270407 579670 270419
rect 579722 270407 579728 270459
rect 168112 270333 168118 270385
rect 168170 270373 168176 270385
rect 405712 270373 405718 270385
rect 168170 270345 220478 270373
rect 168170 270333 168176 270345
rect 195856 270299 195862 270311
rect 168034 270271 195862 270299
rect 195856 270259 195862 270271
rect 195914 270259 195920 270311
rect 195952 270259 195958 270311
rect 196010 270299 196016 270311
rect 213232 270299 213238 270311
rect 196010 270271 213238 270299
rect 196010 270259 196016 270271
rect 213232 270259 213238 270271
rect 213290 270259 213296 270311
rect 213328 270259 213334 270311
rect 213386 270299 213392 270311
rect 220336 270299 220342 270311
rect 213386 270271 220342 270299
rect 213386 270259 213392 270271
rect 220336 270259 220342 270271
rect 220394 270259 220400 270311
rect 220450 270299 220478 270345
rect 220642 270345 405718 270373
rect 220642 270299 220670 270345
rect 405712 270333 405718 270345
rect 405770 270333 405776 270385
rect 508240 270333 508246 270385
rect 508298 270373 508304 270385
rect 601072 270373 601078 270385
rect 508298 270345 601078 270373
rect 508298 270333 508304 270345
rect 601072 270333 601078 270345
rect 601130 270333 601136 270385
rect 220450 270271 220670 270299
rect 237616 270259 237622 270311
rect 237674 270299 237680 270311
rect 337072 270299 337078 270311
rect 237674 270271 337078 270299
rect 237674 270259 237680 270271
rect 337072 270259 337078 270271
rect 337130 270259 337136 270311
rect 357040 270259 357046 270311
rect 357098 270299 357104 270311
rect 380368 270299 380374 270311
rect 357098 270271 380374 270299
rect 357098 270259 357104 270271
rect 380368 270259 380374 270271
rect 380426 270259 380432 270311
rect 380464 270259 380470 270311
rect 380522 270299 380528 270311
rect 402160 270299 402166 270311
rect 380522 270271 402166 270299
rect 380522 270259 380528 270271
rect 402160 270259 402166 270271
rect 402218 270259 402224 270311
rect 402352 270259 402358 270311
rect 402410 270299 402416 270311
rect 554704 270299 554710 270311
rect 402410 270271 554710 270299
rect 402410 270259 402416 270271
rect 554704 270259 554710 270271
rect 554762 270259 554768 270311
rect 562192 270259 562198 270311
rect 562250 270299 562256 270311
rect 646288 270299 646294 270311
rect 562250 270271 646294 270299
rect 562250 270259 562256 270271
rect 646288 270259 646294 270271
rect 646346 270259 646352 270311
rect 84784 270185 84790 270237
rect 84842 270225 84848 270237
rect 140272 270225 140278 270237
rect 84842 270197 140278 270225
rect 84842 270185 84848 270197
rect 140272 270185 140278 270197
rect 140330 270185 140336 270237
rect 152656 270185 152662 270237
rect 152714 270225 152720 270237
rect 394864 270225 394870 270237
rect 152714 270197 394870 270225
rect 152714 270185 152720 270197
rect 394864 270185 394870 270197
rect 394922 270185 394928 270237
rect 400240 270185 400246 270237
rect 400298 270225 400304 270237
rect 568912 270225 568918 270237
rect 400298 270197 568918 270225
rect 400298 270185 400304 270197
rect 568912 270185 568918 270197
rect 568970 270185 568976 270237
rect 588880 270185 588886 270237
rect 588938 270225 588944 270237
rect 632080 270225 632086 270237
rect 588938 270197 632086 270225
rect 588938 270185 588944 270197
rect 632080 270185 632086 270197
rect 632138 270185 632144 270237
rect 80176 270111 80182 270163
rect 80234 270151 80240 270163
rect 140368 270151 140374 270163
rect 80234 270123 140374 270151
rect 80234 270111 80240 270123
rect 140368 270111 140374 270123
rect 140426 270111 140432 270163
rect 161008 270111 161014 270163
rect 161066 270151 161072 270163
rect 403888 270151 403894 270163
rect 161066 270123 403894 270151
rect 161066 270111 161072 270123
rect 403888 270111 403894 270123
rect 403946 270111 403952 270163
rect 408976 270111 408982 270163
rect 409034 270151 409040 270163
rect 422608 270151 422614 270163
rect 409034 270123 422614 270151
rect 409034 270111 409040 270123
rect 422608 270111 422614 270123
rect 422666 270111 422672 270163
rect 521776 270111 521782 270163
rect 521834 270151 521840 270163
rect 622480 270151 622486 270163
rect 521834 270123 622486 270151
rect 521834 270111 521840 270123
rect 622480 270111 622486 270123
rect 622538 270111 622544 270163
rect 75376 270037 75382 270089
rect 75434 270077 75440 270089
rect 139504 270077 139510 270089
rect 75434 270049 139510 270077
rect 75434 270037 75440 270049
rect 139504 270037 139510 270049
rect 139562 270037 139568 270089
rect 153808 270037 153814 270089
rect 153866 270077 153872 270089
rect 153866 270049 403166 270077
rect 153866 270037 153872 270049
rect 68176 269963 68182 270015
rect 68234 270003 68240 270015
rect 139312 270003 139318 270015
rect 68234 269975 139318 270003
rect 68234 269963 68240 269975
rect 139312 269963 139318 269975
rect 139370 269963 139376 270015
rect 142000 269963 142006 270015
rect 142058 270003 142064 270015
rect 380176 270003 380182 270015
rect 142058 269975 380182 270003
rect 142058 269963 142064 269975
rect 380176 269963 380182 269975
rect 380234 269963 380240 270015
rect 387088 270003 387094 270015
rect 380386 269975 387094 270003
rect 135280 269889 135286 269941
rect 135338 269929 135344 269941
rect 155536 269929 155542 269941
rect 135338 269901 155542 269929
rect 135338 269889 135344 269901
rect 155536 269889 155542 269901
rect 155594 269889 155600 269941
rect 166864 269889 166870 269941
rect 166922 269929 166928 269941
rect 182416 269929 182422 269941
rect 166922 269901 182422 269929
rect 166922 269889 166928 269901
rect 182416 269889 182422 269901
rect 182474 269889 182480 269941
rect 182512 269889 182518 269941
rect 182570 269929 182576 269941
rect 195856 269929 195862 269941
rect 182570 269901 195862 269929
rect 182570 269889 182576 269901
rect 195856 269889 195862 269901
rect 195914 269889 195920 269941
rect 195952 269889 195958 269941
rect 196010 269929 196016 269941
rect 209680 269929 209686 269941
rect 196010 269901 209686 269929
rect 196010 269889 196016 269901
rect 209680 269889 209686 269901
rect 209738 269889 209744 269941
rect 209776 269889 209782 269941
rect 209834 269929 209840 269941
rect 219856 269929 219862 269941
rect 209834 269901 219862 269929
rect 209834 269889 209840 269901
rect 219856 269889 219862 269901
rect 219914 269889 219920 269941
rect 219952 269889 219958 269941
rect 220010 269929 220016 269941
rect 236080 269929 236086 269941
rect 220010 269901 236086 269929
rect 220010 269889 220016 269901
rect 236080 269889 236086 269901
rect 236138 269889 236144 269941
rect 237520 269889 237526 269941
rect 237578 269929 237584 269941
rect 337072 269929 337078 269941
rect 237578 269901 337078 269929
rect 237578 269889 237584 269901
rect 337072 269889 337078 269901
rect 337130 269889 337136 269941
rect 337360 269889 337366 269941
rect 337418 269929 337424 269941
rect 356752 269929 356758 269941
rect 337418 269901 356758 269929
rect 337418 269889 337424 269901
rect 356752 269889 356758 269901
rect 356810 269889 356816 269941
rect 357040 269889 357046 269941
rect 357098 269929 357104 269941
rect 380080 269929 380086 269941
rect 357098 269901 380086 269929
rect 357098 269889 357104 269901
rect 380080 269889 380086 269901
rect 380138 269889 380144 269941
rect 127696 269815 127702 269867
rect 127754 269855 127760 269867
rect 380386 269855 380414 269975
rect 387088 269963 387094 269975
rect 387146 269963 387152 270015
rect 387280 269963 387286 270015
rect 387338 270003 387344 270015
rect 403024 270003 403030 270015
rect 387338 269975 403030 270003
rect 387338 269963 387344 269975
rect 403024 269963 403030 269975
rect 403082 269963 403088 270015
rect 403138 270003 403166 270049
rect 403216 270037 403222 270089
rect 403274 270077 403280 270089
rect 408400 270077 408406 270089
rect 403274 270049 408406 270077
rect 403274 270037 403280 270049
rect 408400 270037 408406 270049
rect 408458 270037 408464 270089
rect 411952 270077 411958 270089
rect 408994 270049 411958 270077
rect 405136 270003 405142 270015
rect 403138 269975 405142 270003
rect 405136 269963 405142 269975
rect 405194 269963 405200 270015
rect 406096 269963 406102 270015
rect 406154 270003 406160 270015
rect 408994 270003 409022 270049
rect 411952 270037 411958 270049
rect 412010 270037 412016 270089
rect 446224 270037 446230 270089
rect 446282 270077 446288 270089
rect 576112 270077 576118 270089
rect 446282 270049 576118 270077
rect 446282 270037 446288 270049
rect 576112 270037 576118 270049
rect 576170 270037 576176 270089
rect 406154 269975 409022 270003
rect 406154 269963 406160 269975
rect 409072 269963 409078 270015
rect 409130 270003 409136 270015
rect 583216 270003 583222 270015
rect 409130 269975 583222 270003
rect 409130 269963 409136 269975
rect 583216 269963 583222 269975
rect 583274 269963 583280 270015
rect 382288 269889 382294 269941
rect 382346 269929 382352 269941
rect 408976 269929 408982 269941
rect 382346 269901 408982 269929
rect 382346 269889 382352 269901
rect 408976 269889 408982 269901
rect 409034 269889 409040 269941
rect 409168 269889 409174 269941
rect 409226 269929 409232 269941
rect 593968 269929 593974 269941
rect 409226 269901 593974 269929
rect 409226 269889 409232 269901
rect 593968 269889 593974 269901
rect 594026 269889 594032 269941
rect 127754 269827 380414 269855
rect 127754 269815 127760 269827
rect 380560 269815 380566 269867
rect 380618 269855 380624 269867
rect 388816 269855 388822 269867
rect 380618 269827 388822 269855
rect 380618 269815 380624 269827
rect 388816 269815 388822 269827
rect 388874 269815 388880 269867
rect 391696 269815 391702 269867
rect 391754 269855 391760 269867
rect 590032 269855 590038 269867
rect 391754 269827 590038 269855
rect 391754 269815 391760 269827
rect 590032 269815 590038 269827
rect 590090 269815 590096 269867
rect 114640 269741 114646 269793
rect 114698 269781 114704 269793
rect 383152 269781 383158 269793
rect 114698 269753 383158 269781
rect 114698 269741 114704 269753
rect 383152 269741 383158 269753
rect 383210 269741 383216 269793
rect 383248 269741 383254 269793
rect 383306 269781 383312 269793
rect 407536 269781 407542 269793
rect 383306 269753 407542 269781
rect 383306 269741 383312 269753
rect 407536 269741 407542 269753
rect 407594 269741 407600 269793
rect 407632 269741 407638 269793
rect 407690 269781 407696 269793
rect 608176 269781 608182 269793
rect 407690 269753 608182 269781
rect 407690 269741 407696 269753
rect 608176 269741 608182 269753
rect 608234 269741 608240 269793
rect 74128 269667 74134 269719
rect 74186 269707 74192 269719
rect 367984 269707 367990 269719
rect 74186 269679 367990 269707
rect 74186 269667 74192 269679
rect 367984 269667 367990 269679
rect 368042 269667 368048 269719
rect 380080 269667 380086 269719
rect 380138 269707 380144 269719
rect 382768 269707 382774 269719
rect 380138 269679 382774 269707
rect 380138 269667 380144 269679
rect 382768 269667 382774 269679
rect 382826 269667 382832 269719
rect 382864 269667 382870 269719
rect 382922 269707 382928 269719
rect 633136 269707 633142 269719
rect 382922 269679 633142 269707
rect 382922 269667 382928 269679
rect 633136 269667 633142 269679
rect 633194 269667 633200 269719
rect 90832 269593 90838 269645
rect 90890 269633 90896 269645
rect 388624 269633 388630 269645
rect 90890 269605 388630 269633
rect 90890 269593 90896 269605
rect 388624 269593 388630 269605
rect 388682 269593 388688 269645
rect 388912 269593 388918 269645
rect 388970 269633 388976 269645
rect 611824 269633 611830 269645
rect 388970 269605 611830 269633
rect 388970 269593 388976 269605
rect 611824 269593 611830 269605
rect 611882 269593 611888 269645
rect 87184 269519 87190 269571
rect 87242 269559 87248 269571
rect 87242 269531 385982 269559
rect 87242 269519 87248 269531
rect 81328 269445 81334 269497
rect 81386 269485 81392 269497
rect 385648 269485 385654 269497
rect 81386 269457 385654 269485
rect 81386 269445 81392 269457
rect 385648 269445 385654 269457
rect 385706 269445 385712 269497
rect 385954 269485 385982 269531
rect 386032 269519 386038 269571
rect 386090 269559 386096 269571
rect 618928 269559 618934 269571
rect 386090 269531 618934 269559
rect 386090 269519 386096 269531
rect 618928 269519 618934 269531
rect 618986 269519 618992 269571
rect 388720 269485 388726 269497
rect 385954 269457 388726 269485
rect 388720 269445 388726 269457
rect 388778 269445 388784 269497
rect 388816 269445 388822 269497
rect 388874 269485 388880 269497
rect 394576 269485 394582 269497
rect 388874 269457 394582 269485
rect 388874 269445 388880 269457
rect 394576 269445 394582 269457
rect 394634 269445 394640 269497
rect 394672 269445 394678 269497
rect 394730 269485 394736 269497
rect 629680 269485 629686 269497
rect 394730 269457 629686 269485
rect 394730 269445 394736 269457
rect 629680 269445 629686 269457
rect 629738 269445 629744 269497
rect 78928 269371 78934 269423
rect 78986 269411 78992 269423
rect 382960 269411 382966 269423
rect 78986 269383 382966 269411
rect 78986 269371 78992 269383
rect 382960 269371 382966 269383
rect 383018 269371 383024 269423
rect 383632 269411 383638 269423
rect 383074 269383 383638 269411
rect 69328 269297 69334 269349
rect 69386 269337 69392 269349
rect 376048 269337 376054 269349
rect 69386 269309 376054 269337
rect 69386 269297 69392 269309
rect 376048 269297 376054 269309
rect 376106 269297 376112 269349
rect 380176 269297 380182 269349
rect 380234 269337 380240 269349
rect 383074 269337 383102 269383
rect 383632 269371 383638 269383
rect 383690 269371 383696 269423
rect 383728 269371 383734 269423
rect 383786 269411 383792 269423
rect 383786 269383 407486 269411
rect 383786 269371 383792 269383
rect 380234 269309 383102 269337
rect 380234 269297 380240 269309
rect 383152 269297 383158 269349
rect 383210 269337 383216 269349
rect 383210 269309 385886 269337
rect 383210 269297 383216 269309
rect 71728 269223 71734 269275
rect 71786 269263 71792 269275
rect 385744 269263 385750 269275
rect 71786 269235 385750 269263
rect 71786 269223 71792 269235
rect 385744 269223 385750 269235
rect 385802 269223 385808 269275
rect 385858 269263 385886 269309
rect 385936 269297 385942 269349
rect 385994 269337 386000 269349
rect 407458 269337 407486 269383
rect 407536 269371 407542 269423
rect 407594 269411 407600 269423
rect 636496 269411 636502 269423
rect 407594 269383 636502 269411
rect 407594 269371 407600 269383
rect 636496 269371 636502 269383
rect 636554 269371 636560 269423
rect 640336 269337 640342 269349
rect 385994 269309 407390 269337
rect 407458 269309 640342 269337
rect 385994 269297 386000 269309
rect 391408 269263 391414 269275
rect 385858 269235 391414 269263
rect 391408 269223 391414 269235
rect 391466 269223 391472 269275
rect 391792 269223 391798 269275
rect 391850 269263 391856 269275
rect 394480 269263 394486 269275
rect 391850 269235 394486 269263
rect 391850 269223 391856 269235
rect 394480 269223 394486 269235
rect 394538 269223 394544 269275
rect 394576 269223 394582 269275
rect 394634 269263 394640 269275
rect 407362 269263 407390 269309
rect 640336 269297 640342 269309
rect 640394 269297 640400 269349
rect 643888 269263 643894 269275
rect 394634 269235 407294 269263
rect 407362 269235 643894 269263
rect 394634 269223 394640 269235
rect 108688 269149 108694 269201
rect 108746 269189 108752 269201
rect 139696 269189 139702 269201
rect 108746 269161 139702 269189
rect 108746 269149 108752 269161
rect 139696 269149 139702 269161
rect 139754 269149 139760 269201
rect 155536 269149 155542 269201
rect 155594 269189 155600 269201
rect 182512 269189 182518 269201
rect 155594 269161 182518 269189
rect 155594 269149 155600 269161
rect 182512 269149 182518 269161
rect 182570 269149 182576 269201
rect 182704 269149 182710 269201
rect 182762 269189 182768 269201
rect 405616 269189 405622 269201
rect 182762 269161 405622 269189
rect 182762 269149 182768 269161
rect 405616 269149 405622 269161
rect 405674 269149 405680 269201
rect 407266 269189 407294 269235
rect 643888 269223 643894 269235
rect 643946 269223 643952 269275
rect 407266 269161 407774 269189
rect 112240 269075 112246 269127
rect 112298 269115 112304 269127
rect 139600 269115 139606 269127
rect 112298 269087 139606 269115
rect 112298 269075 112304 269087
rect 139600 269075 139606 269087
rect 139658 269075 139664 269127
rect 181264 269075 181270 269127
rect 181322 269115 181328 269127
rect 380464 269115 380470 269127
rect 181322 269087 380470 269115
rect 181322 269075 181328 269087
rect 380464 269075 380470 269087
rect 380522 269075 380528 269127
rect 382768 269075 382774 269127
rect 382826 269115 382832 269127
rect 388528 269115 388534 269127
rect 382826 269087 388534 269115
rect 382826 269075 382832 269087
rect 388528 269075 388534 269087
rect 388586 269075 388592 269127
rect 388816 269075 388822 269127
rect 388874 269115 388880 269127
rect 388874 269087 405758 269115
rect 388874 269075 388880 269087
rect 115792 269001 115798 269053
rect 115850 269041 115856 269053
rect 139408 269041 139414 269053
rect 115850 269013 139414 269041
rect 115850 269001 115856 269013
rect 139408 269001 139414 269013
rect 139466 269001 139472 269053
rect 185968 269001 185974 269053
rect 186026 269041 186032 269053
rect 405730 269041 405758 269087
rect 405808 269075 405814 269127
rect 405866 269115 405872 269127
rect 407632 269115 407638 269127
rect 405866 269087 407638 269115
rect 405866 269075 405872 269087
rect 407632 269075 407638 269087
rect 407690 269075 407696 269127
rect 407746 269115 407774 269161
rect 472336 269149 472342 269201
rect 472394 269189 472400 269201
rect 561808 269189 561814 269201
rect 472394 269161 561814 269189
rect 472394 269149 472400 269161
rect 561808 269149 561814 269161
rect 561866 269149 561872 269201
rect 570256 269149 570262 269201
rect 570314 269189 570320 269201
rect 639088 269189 639094 269201
rect 570314 269161 639094 269189
rect 570314 269149 570320 269161
rect 639088 269149 639094 269161
rect 639146 269149 639152 269201
rect 452368 269115 452374 269127
rect 407746 269087 452374 269115
rect 452368 269075 452374 269087
rect 452426 269075 452432 269127
rect 488080 269075 488086 269127
rect 488138 269115 488144 269127
rect 572560 269115 572566 269127
rect 488138 269087 572566 269115
rect 488138 269075 488144 269087
rect 572560 269075 572566 269087
rect 572618 269075 572624 269127
rect 186026 269013 403166 269041
rect 405730 269013 406814 269041
rect 186026 269001 186032 269013
rect 119344 268927 119350 268979
rect 119402 268967 119408 268979
rect 140944 268967 140950 268979
rect 119402 268939 140950 268967
rect 119402 268927 119408 268939
rect 140944 268927 140950 268939
rect 141002 268927 141008 268979
rect 184720 268927 184726 268979
rect 184778 268967 184784 268979
rect 387280 268967 387286 268979
rect 184778 268939 387286 268967
rect 184778 268927 184784 268939
rect 387280 268927 387286 268939
rect 387338 268927 387344 268979
rect 387376 268927 387382 268979
rect 387434 268967 387440 268979
rect 400144 268967 400150 268979
rect 387434 268939 400150 268967
rect 387434 268927 387440 268939
rect 400144 268927 400150 268939
rect 400202 268927 400208 268979
rect 403138 268967 403166 269013
rect 406672 268967 406678 268979
rect 403138 268939 406678 268967
rect 406672 268927 406678 268939
rect 406730 268927 406736 268979
rect 406786 268967 406814 269013
rect 502672 269001 502678 269053
rect 502730 269041 502736 269053
rect 586768 269041 586774 269053
rect 502730 269013 586774 269041
rect 502730 269001 502736 269013
rect 586768 269001 586774 269013
rect 586826 269001 586832 269053
rect 448912 268967 448918 268979
rect 406786 268939 448918 268967
rect 448912 268927 448918 268939
rect 448970 268927 448976 268979
rect 478768 268927 478774 268979
rect 478826 268967 478832 268979
rect 558256 268967 558262 268979
rect 478826 268939 558262 268967
rect 478826 268927 478832 268939
rect 558256 268927 558262 268939
rect 558314 268927 558320 268979
rect 135376 268853 135382 268905
rect 135434 268893 135440 268905
rect 259216 268893 259222 268905
rect 135434 268865 259222 268893
rect 135434 268853 135440 268865
rect 259216 268853 259222 268865
rect 259274 268853 259280 268905
rect 283792 268853 283798 268905
rect 283850 268893 283856 268905
rect 283850 268865 332126 268893
rect 283850 268853 283856 268865
rect 133552 268779 133558 268831
rect 133610 268819 133616 268831
rect 140560 268819 140566 268831
rect 133610 268791 140566 268819
rect 133610 268779 133616 268791
rect 140560 268779 140566 268791
rect 140618 268779 140624 268831
rect 175504 268779 175510 268831
rect 175562 268819 175568 268831
rect 187024 268819 187030 268831
rect 175562 268791 187030 268819
rect 175562 268779 175568 268791
rect 187024 268779 187030 268791
rect 187082 268779 187088 268831
rect 195856 268779 195862 268831
rect 195914 268819 195920 268831
rect 218800 268819 218806 268831
rect 195914 268791 218806 268819
rect 195914 268779 195920 268791
rect 218800 268779 218806 268791
rect 218858 268779 218864 268831
rect 219280 268779 219286 268831
rect 219338 268819 219344 268831
rect 219338 268791 324542 268819
rect 219338 268779 219344 268791
rect 122896 268705 122902 268757
rect 122954 268745 122960 268757
rect 140848 268745 140854 268757
rect 122954 268717 140854 268745
rect 122954 268705 122960 268717
rect 140848 268705 140854 268717
rect 140906 268705 140912 268757
rect 213232 268705 213238 268757
rect 213290 268745 213296 268757
rect 219952 268745 219958 268757
rect 213290 268717 219958 268745
rect 213290 268705 213296 268717
rect 219952 268705 219958 268717
rect 220010 268705 220016 268757
rect 226384 268705 226390 268757
rect 226442 268745 226448 268757
rect 324400 268745 324406 268757
rect 226442 268717 324406 268745
rect 226442 268705 226448 268717
rect 324400 268705 324406 268717
rect 324458 268705 324464 268757
rect 131248 268631 131254 268683
rect 131306 268671 131312 268683
rect 135376 268671 135382 268683
rect 131306 268643 135382 268671
rect 131306 268631 131312 268643
rect 135376 268631 135382 268643
rect 135434 268631 135440 268683
rect 212176 268631 212182 268683
rect 212234 268671 212240 268683
rect 313936 268671 313942 268683
rect 212234 268643 313942 268671
rect 212234 268631 212240 268643
rect 313936 268631 313942 268643
rect 313994 268631 314000 268683
rect 324514 268671 324542 268791
rect 331984 268671 331990 268683
rect 324514 268643 331990 268671
rect 331984 268631 331990 268643
rect 332042 268631 332048 268683
rect 332098 268671 332126 268865
rect 337072 268853 337078 268905
rect 337130 268893 337136 268905
rect 357040 268893 357046 268905
rect 337130 268865 357046 268893
rect 337130 268853 337136 268865
rect 357040 268853 357046 268865
rect 357098 268853 357104 268905
rect 371920 268853 371926 268905
rect 371978 268893 371984 268905
rect 543664 268893 543670 268905
rect 371978 268865 543670 268893
rect 371978 268853 371984 268865
rect 543664 268853 543670 268865
rect 543722 268853 543728 268905
rect 550096 268853 550102 268905
rect 550154 268893 550160 268905
rect 615376 268893 615382 268905
rect 550154 268865 615382 268893
rect 550154 268853 550160 268865
rect 615376 268853 615382 268865
rect 615434 268853 615440 268905
rect 349552 268779 349558 268831
rect 349610 268819 349616 268831
rect 358096 268819 358102 268831
rect 349610 268791 358102 268819
rect 349610 268779 349616 268791
rect 358096 268779 358102 268791
rect 358154 268779 358160 268831
rect 371344 268779 371350 268831
rect 371402 268819 371408 268831
rect 536848 268819 536854 268831
rect 371402 268791 536854 268819
rect 371402 268779 371408 268791
rect 536848 268779 536854 268791
rect 536906 268779 536912 268831
rect 337168 268705 337174 268757
rect 337226 268745 337232 268757
rect 337226 268717 339998 268745
rect 337226 268705 337232 268717
rect 339856 268671 339862 268683
rect 332098 268643 339862 268671
rect 339856 268631 339862 268643
rect 339914 268631 339920 268683
rect 339970 268671 339998 268717
rect 350128 268705 350134 268757
rect 350186 268745 350192 268757
rect 365584 268745 365590 268757
rect 350186 268717 365590 268745
rect 350186 268705 350192 268717
rect 365584 268705 365590 268717
rect 365642 268705 365648 268757
rect 370192 268705 370198 268757
rect 370250 268745 370256 268757
rect 529744 268745 529750 268757
rect 370250 268717 529750 268745
rect 370250 268705 370256 268717
rect 529744 268705 529750 268717
rect 529802 268705 529808 268757
rect 356944 268671 356950 268683
rect 339970 268643 356950 268671
rect 356944 268631 356950 268643
rect 357002 268631 357008 268683
rect 373168 268631 373174 268683
rect 373226 268671 373232 268683
rect 522544 268671 522550 268683
rect 373226 268643 522550 268671
rect 373226 268631 373232 268643
rect 522544 268631 522550 268643
rect 522602 268631 522608 268683
rect 217456 268557 217462 268609
rect 217514 268597 217520 268609
rect 219376 268597 219382 268609
rect 217514 268569 219382 268597
rect 217514 268557 217520 268569
rect 219376 268557 219382 268569
rect 219434 268557 219440 268609
rect 247696 268557 247702 268609
rect 247754 268597 247760 268609
rect 252208 268597 252214 268609
rect 247754 268569 252214 268597
rect 247754 268557 247760 268569
rect 252208 268557 252214 268569
rect 252266 268557 252272 268609
rect 269200 268557 269206 268609
rect 269258 268597 269264 268609
rect 331216 268597 331222 268609
rect 269258 268569 331222 268597
rect 269258 268557 269264 268569
rect 331216 268557 331222 268569
rect 331274 268557 331280 268609
rect 337264 268557 337270 268609
rect 337322 268597 337328 268609
rect 356848 268597 356854 268609
rect 337322 268569 356854 268597
rect 337322 268557 337328 268569
rect 356848 268557 356854 268569
rect 356906 268557 356912 268609
rect 368464 268557 368470 268609
rect 368522 268597 368528 268609
rect 515440 268597 515446 268609
rect 368522 268569 515446 268597
rect 368522 268557 368528 268569
rect 515440 268557 515446 268569
rect 515498 268557 515504 268609
rect 223600 268483 223606 268535
rect 223658 268523 223664 268535
rect 238288 268523 238294 268535
rect 223658 268495 238294 268523
rect 223658 268483 223664 268495
rect 238288 268483 238294 268495
rect 238346 268483 238352 268535
rect 240688 268483 240694 268535
rect 240746 268523 240752 268535
rect 267856 268523 267862 268535
rect 240746 268495 267862 268523
rect 240746 268483 240752 268495
rect 267856 268483 267862 268495
rect 267914 268483 267920 268535
rect 272752 268483 272758 268535
rect 272810 268523 272816 268535
rect 334096 268523 334102 268535
rect 272810 268495 334102 268523
rect 272810 268483 272816 268495
rect 334096 268483 334102 268495
rect 334154 268483 334160 268535
rect 367600 268483 367606 268535
rect 367658 268523 367664 268535
rect 508336 268523 508342 268535
rect 367658 268495 508342 268523
rect 367658 268483 367664 268495
rect 508336 268483 508342 268495
rect 508394 268483 508400 268535
rect 126544 268409 126550 268461
rect 126602 268449 126608 268461
rect 140752 268449 140758 268461
rect 126602 268421 140758 268449
rect 126602 268409 126608 268421
rect 140752 268409 140758 268421
rect 140810 268409 140816 268461
rect 218800 268409 218806 268461
rect 218858 268449 218864 268461
rect 237520 268449 237526 268461
rect 218858 268421 237526 268449
rect 218858 268409 218864 268421
rect 237520 268409 237526 268421
rect 237578 268409 237584 268461
rect 279952 268409 279958 268461
rect 280010 268449 280016 268461
rect 334192 268449 334198 268461
rect 280010 268421 334198 268449
rect 280010 268409 280016 268421
rect 334192 268409 334198 268421
rect 334250 268409 334256 268461
rect 336976 268409 336982 268461
rect 337034 268449 337040 268461
rect 346384 268449 346390 268461
rect 337034 268421 346390 268449
rect 337034 268409 337040 268421
rect 346384 268409 346390 268421
rect 346442 268409 346448 268461
rect 366928 268409 366934 268461
rect 366986 268449 366992 268461
rect 501136 268449 501142 268461
rect 366986 268421 501142 268449
rect 366986 268409 366992 268421
rect 501136 268409 501142 268421
rect 501194 268409 501200 268461
rect 130096 268335 130102 268387
rect 130154 268375 130160 268387
rect 140656 268375 140662 268387
rect 130154 268347 140662 268375
rect 130154 268335 130160 268347
rect 140656 268335 140662 268347
rect 140714 268335 140720 268387
rect 224176 268335 224182 268387
rect 224234 268375 224240 268387
rect 245488 268375 245494 268387
rect 224234 268347 245494 268375
rect 224234 268335 224240 268347
rect 245488 268335 245494 268347
rect 245546 268335 245552 268387
rect 264496 268335 264502 268387
rect 264554 268375 264560 268387
rect 282160 268375 282166 268387
rect 264554 268347 282166 268375
rect 264554 268335 264560 268347
rect 282160 268335 282166 268347
rect 282218 268335 282224 268387
rect 286096 268335 286102 268387
rect 286154 268375 286160 268387
rect 296752 268375 296758 268387
rect 286154 268347 296758 268375
rect 286154 268335 286160 268347
rect 296752 268335 296758 268347
rect 296810 268335 296816 268387
rect 298576 268335 298582 268387
rect 298634 268375 298640 268387
rect 338704 268375 338710 268387
rect 298634 268347 338710 268375
rect 298634 268335 298640 268347
rect 338704 268335 338710 268347
rect 338762 268335 338768 268387
rect 365872 268335 365878 268387
rect 365930 268375 365936 268387
rect 494032 268375 494038 268387
rect 365930 268347 494038 268375
rect 365930 268335 365936 268347
rect 494032 268335 494038 268347
rect 494090 268335 494096 268387
rect 209680 268261 209686 268313
rect 209738 268301 209744 268313
rect 237616 268301 237622 268313
rect 209738 268273 237622 268301
rect 209738 268261 209744 268273
rect 237616 268261 237622 268273
rect 237674 268261 237680 268313
rect 271600 268261 271606 268313
rect 271658 268301 271664 268313
rect 282832 268301 282838 268313
rect 271658 268273 282838 268301
rect 271658 268261 271664 268273
rect 282832 268261 282838 268273
rect 282890 268261 282896 268313
rect 339376 268301 339382 268313
rect 301186 268273 339382 268301
rect 259216 268187 259222 268239
rect 259274 268227 259280 268239
rect 279280 268227 279286 268239
rect 259274 268199 279286 268227
rect 259274 268187 259280 268199
rect 279280 268187 279286 268199
rect 279338 268187 279344 268239
rect 294256 268187 294262 268239
rect 294314 268227 294320 268239
rect 301186 268227 301214 268273
rect 339376 268261 339382 268273
rect 339434 268261 339440 268313
rect 365200 268261 365206 268313
rect 365258 268301 365264 268313
rect 486832 268301 486838 268313
rect 365258 268273 486838 268301
rect 365258 268261 365264 268273
rect 486832 268261 486838 268273
rect 486890 268261 486896 268313
rect 294314 268199 301214 268227
rect 294314 268187 294320 268199
rect 301264 268187 301270 268239
rect 301322 268227 301328 268239
rect 339664 268227 339670 268239
rect 301322 268199 339670 268227
rect 301322 268187 301328 268199
rect 339664 268187 339670 268199
rect 339722 268187 339728 268239
rect 364336 268187 364342 268239
rect 364394 268227 364400 268239
rect 479824 268227 479830 268239
rect 364394 268199 479830 268227
rect 364394 268187 364400 268199
rect 479824 268187 479830 268199
rect 479882 268187 479888 268239
rect 287056 268113 287062 268165
rect 287114 268153 287120 268165
rect 298576 268153 298582 268165
rect 287114 268125 298582 268153
rect 287114 268113 287120 268125
rect 298576 268113 298582 268125
rect 298634 268113 298640 268165
rect 308464 268113 308470 268165
rect 308522 268153 308528 268165
rect 343216 268153 343222 268165
rect 308522 268125 343222 268153
rect 308522 268113 308528 268125
rect 343216 268113 343222 268125
rect 343274 268113 343280 268165
rect 363184 268113 363190 268165
rect 363242 268153 363248 268165
rect 472624 268153 472630 268165
rect 363242 268125 472630 268153
rect 363242 268113 363248 268125
rect 472624 268113 472630 268125
rect 472682 268113 472688 268165
rect 287632 268039 287638 268091
rect 287690 268079 287696 268091
rect 307312 268079 307318 268091
rect 287690 268051 307318 268079
rect 287690 268039 287696 268051
rect 307312 268039 307318 268051
rect 307370 268039 307376 268091
rect 315664 268039 315670 268091
rect 315722 268079 315728 268091
rect 341968 268079 341974 268091
rect 315722 268051 341974 268079
rect 315722 268039 315728 268051
rect 341968 268039 341974 268051
rect 342026 268039 342032 268091
rect 362608 268039 362614 268091
rect 362666 268079 362672 268091
rect 465520 268079 465526 268091
rect 362666 268051 465526 268079
rect 362666 268039 362672 268051
rect 465520 268039 465526 268051
rect 465578 268039 465584 268091
rect 322768 267965 322774 268017
rect 322826 268005 322832 268017
rect 344656 268005 344662 268017
rect 322826 267977 344662 268005
rect 322826 267965 322832 267977
rect 344656 267965 344662 267977
rect 344714 267965 344720 268017
rect 361456 267965 361462 268017
rect 361514 268005 361520 268017
rect 458320 268005 458326 268017
rect 361514 267977 458326 268005
rect 361514 267965 361520 267977
rect 458320 267965 458326 267977
rect 458378 267965 458384 268017
rect 222544 267891 222550 267943
rect 222602 267931 222608 267943
rect 231184 267931 231190 267943
rect 222602 267903 231190 267931
rect 222602 267891 222608 267903
rect 231184 267891 231190 267903
rect 231242 267891 231248 267943
rect 319120 267891 319126 267943
rect 319178 267931 319184 267943
rect 341584 267931 341590 267943
rect 319178 267903 341590 267931
rect 319178 267891 319184 267903
rect 341584 267891 341590 267903
rect 341642 267891 341648 267943
rect 360592 267891 360598 267943
rect 360650 267931 360656 267943
rect 450832 267931 450838 267943
rect 360650 267903 450838 267931
rect 360650 267891 360656 267903
rect 450832 267891 450838 267903
rect 450890 267891 450896 267943
rect 66832 267817 66838 267869
rect 66890 267857 66896 267869
rect 66890 267829 69182 267857
rect 66890 267817 66896 267829
rect 69154 267783 69182 267829
rect 137200 267817 137206 267869
rect 137258 267857 137264 267869
rect 140464 267857 140470 267869
rect 137258 267829 140470 267857
rect 137258 267817 137264 267829
rect 140464 267817 140470 267829
rect 140522 267817 140528 267869
rect 147952 267817 147958 267869
rect 148010 267857 148016 267869
rect 149680 267857 149686 267869
rect 148010 267829 149686 267857
rect 148010 267817 148016 267829
rect 149680 267817 149686 267829
rect 149738 267817 149744 267869
rect 151408 267817 151414 267869
rect 151466 267857 151472 267869
rect 152560 267857 152566 267869
rect 151466 267829 152566 267857
rect 151466 267817 151472 267829
rect 152560 267817 152566 267829
rect 152618 267817 152624 267869
rect 158608 267817 158614 267869
rect 158666 267857 158672 267869
rect 161200 267857 161206 267869
rect 158666 267829 161206 267857
rect 158666 267817 158672 267829
rect 161200 267817 161206 267829
rect 161258 267817 161264 267869
rect 162160 267817 162166 267869
rect 162218 267857 162224 267869
rect 164080 267857 164086 267869
rect 162218 267829 164086 267857
rect 162218 267817 162224 267829
rect 164080 267817 164086 267829
rect 164138 267817 164144 267869
rect 165808 267817 165814 267869
rect 165866 267857 165872 267869
rect 166960 267857 166966 267869
rect 165866 267829 166966 267857
rect 165866 267817 165872 267829
rect 166960 267817 166966 267829
rect 167018 267817 167024 267869
rect 191056 267817 191062 267869
rect 191114 267857 191120 267869
rect 192880 267857 192886 267869
rect 191114 267829 192886 267857
rect 191114 267817 191120 267829
rect 192880 267817 192886 267829
rect 192938 267817 192944 267869
rect 222064 267817 222070 267869
rect 222122 267857 222128 267869
rect 227632 267857 227638 267869
rect 222122 267829 227638 267857
rect 222122 267817 222128 267829
rect 227632 267817 227638 267829
rect 227690 267817 227696 267869
rect 258544 267817 258550 267869
rect 258602 267857 258608 267869
rect 275920 267857 275926 267869
rect 258602 267829 275926 267857
rect 258602 267817 258608 267829
rect 275920 267817 275926 267829
rect 275978 267817 275984 267869
rect 278800 267817 278806 267869
rect 278858 267857 278864 267869
rect 283888 267857 283894 267869
rect 278858 267829 283894 267857
rect 278858 267817 278864 267829
rect 283888 267817 283894 267829
rect 283946 267817 283952 267869
rect 285616 267817 285622 267869
rect 285674 267857 285680 267869
rect 293008 267857 293014 267869
rect 285674 267829 293014 267857
rect 285674 267817 285680 267829
rect 293008 267817 293014 267829
rect 293066 267817 293072 267869
rect 324400 267817 324406 267869
rect 324458 267857 324464 267869
rect 330160 267857 330166 267869
rect 324458 267829 330166 267857
rect 324458 267817 324464 267829
rect 330160 267817 330166 267829
rect 330218 267817 330224 267869
rect 344176 267817 344182 267869
rect 344234 267857 344240 267869
rect 347536 267857 347542 267869
rect 344234 267829 347542 267857
rect 344234 267817 344240 267829
rect 347536 267817 347542 267829
rect 347594 267817 347600 267869
rect 359920 267817 359926 267869
rect 359978 267857 359984 267869
rect 444112 267857 444118 267869
rect 359978 267829 444118 267857
rect 359978 267817 359984 267829
rect 444112 267817 444118 267829
rect 444170 267817 444176 267869
rect 455632 267857 455638 267869
rect 447010 267829 447422 267857
rect 72112 267783 72118 267795
rect 69154 267755 72118 267783
rect 72112 267743 72118 267755
rect 72170 267743 72176 267795
rect 139120 267743 139126 267795
rect 139178 267783 139184 267795
rect 140272 267783 140278 267795
rect 139178 267755 140278 267783
rect 139178 267743 139184 267755
rect 140272 267743 140278 267755
rect 140330 267743 140336 267795
rect 181456 267743 181462 267795
rect 181514 267783 181520 267795
rect 191248 267783 191254 267795
rect 181514 267755 191254 267783
rect 181514 267743 181520 267755
rect 191248 267743 191254 267755
rect 191306 267743 191312 267795
rect 250480 267743 250486 267795
rect 250538 267783 250544 267795
rect 250538 267755 258974 267783
rect 250538 267743 250544 267755
rect 250768 267669 250774 267721
rect 250826 267709 250832 267721
rect 258832 267709 258838 267721
rect 250826 267681 258838 267709
rect 250826 267669 250832 267681
rect 258832 267669 258838 267681
rect 258890 267669 258896 267721
rect 258946 267709 258974 267755
rect 259120 267743 259126 267795
rect 259178 267783 259184 267795
rect 447010 267783 447038 267829
rect 259178 267755 447038 267783
rect 259178 267743 259184 267755
rect 447088 267743 447094 267795
rect 447146 267783 447152 267795
rect 447394 267783 447422 267829
rect 454978 267829 455638 267857
rect 454978 267783 455006 267829
rect 455632 267817 455638 267829
rect 455690 267817 455696 267869
rect 447146 267755 447326 267783
rect 447394 267755 455006 267783
rect 447146 267743 447152 267755
rect 447184 267709 447190 267721
rect 258946 267681 447190 267709
rect 447184 267669 447190 267681
rect 447242 267669 447248 267721
rect 447298 267709 447326 267755
rect 455056 267743 455062 267795
rect 455114 267783 455120 267795
rect 511888 267783 511894 267795
rect 455114 267755 511894 267783
rect 455114 267743 455120 267755
rect 511888 267743 511894 267755
rect 511946 267743 511952 267795
rect 463120 267709 463126 267721
rect 447298 267681 463126 267709
rect 463120 267669 463126 267681
rect 463178 267669 463184 267721
rect 210928 267595 210934 267647
rect 210986 267635 210992 267647
rect 275632 267635 275638 267647
rect 210986 267607 275638 267635
rect 210986 267595 210992 267607
rect 275632 267595 275638 267607
rect 275690 267595 275696 267647
rect 317488 267595 317494 267647
rect 317546 267635 317552 267647
rect 321808 267635 321814 267647
rect 317546 267607 321814 267635
rect 317546 267595 317552 267607
rect 321808 267595 321814 267607
rect 321866 267595 321872 267647
rect 321904 267595 321910 267647
rect 321962 267635 321968 267647
rect 524944 267635 524950 267647
rect 321962 267607 524950 267635
rect 321962 267595 321968 267607
rect 524944 267595 524950 267607
rect 525002 267595 525008 267647
rect 251248 267521 251254 267573
rect 251306 267561 251312 267573
rect 251306 267533 258782 267561
rect 251306 267521 251312 267533
rect 251920 267447 251926 267499
rect 251978 267487 251984 267499
rect 258754 267487 258782 267533
rect 258832 267521 258838 267573
rect 258890 267561 258896 267573
rect 447088 267561 447094 267573
rect 258890 267533 447094 267561
rect 258890 267521 258896 267533
rect 447088 267521 447094 267533
rect 447146 267521 447152 267573
rect 447184 267521 447190 267573
rect 447242 267561 447248 267573
rect 459568 267561 459574 267573
rect 447242 267533 459574 267561
rect 447242 267521 447248 267533
rect 459568 267521 459574 267533
rect 459626 267521 459632 267573
rect 466768 267487 466774 267499
rect 251978 267459 258686 267487
rect 258754 267459 466774 267487
rect 251978 267447 251984 267459
rect 252400 267373 252406 267425
rect 252458 267413 252464 267425
rect 258658 267413 258686 267459
rect 466768 267447 466774 267459
rect 466826 267447 466832 267499
rect 470224 267413 470230 267425
rect 252458 267385 258590 267413
rect 258658 267385 470230 267413
rect 252458 267373 252464 267385
rect 258562 267339 258590 267385
rect 470224 267373 470230 267385
rect 470282 267373 470288 267425
rect 473776 267339 473782 267351
rect 258562 267311 473782 267339
rect 473776 267299 473782 267311
rect 473834 267299 473840 267351
rect 207376 267225 207382 267277
rect 207434 267265 207440 267277
rect 258352 267265 258358 267277
rect 207434 267237 258358 267265
rect 207434 267225 207440 267237
rect 258352 267225 258358 267237
rect 258410 267225 258416 267277
rect 258544 267225 258550 267277
rect 258602 267265 258608 267277
rect 275248 267265 275254 267277
rect 258602 267237 275254 267265
rect 258602 267225 258608 267237
rect 275248 267225 275254 267237
rect 275306 267225 275312 267277
rect 289840 267225 289846 267277
rect 289898 267265 289904 267277
rect 325168 267265 325174 267277
rect 289898 267237 325174 267265
rect 289898 267225 289904 267237
rect 325168 267225 325174 267237
rect 325226 267225 325232 267277
rect 325456 267225 325462 267277
rect 325514 267265 325520 267277
rect 549904 267265 549910 267277
rect 325514 267237 549910 267265
rect 325514 267225 325520 267237
rect 549904 267225 549910 267237
rect 549962 267225 549968 267277
rect 225328 267151 225334 267203
rect 225386 267191 225392 267203
rect 247696 267191 247702 267203
rect 225386 267163 247702 267191
rect 225386 267151 225392 267163
rect 247696 267151 247702 267163
rect 247754 267151 247760 267203
rect 252976 267151 252982 267203
rect 253034 267191 253040 267203
rect 253034 267163 258398 267191
rect 253034 267151 253040 267163
rect 215728 267077 215734 267129
rect 215786 267117 215792 267129
rect 253648 267117 253654 267129
rect 215786 267089 253654 267117
rect 215786 267077 215792 267089
rect 253648 267077 253654 267089
rect 253706 267077 253712 267129
rect 253744 267077 253750 267129
rect 253802 267117 253808 267129
rect 258256 267117 258262 267129
rect 253802 267089 258262 267117
rect 253802 267077 253808 267089
rect 258256 267077 258262 267089
rect 258314 267077 258320 267129
rect 191920 267003 191926 267055
rect 191978 267043 191984 267055
rect 217648 267043 217654 267055
rect 191978 267015 217654 267043
rect 191978 267003 191984 267015
rect 217648 267003 217654 267015
rect 217706 267003 217712 267055
rect 222832 267003 222838 267055
rect 222890 267043 222896 267055
rect 253360 267043 253366 267055
rect 222890 267015 253366 267043
rect 222890 267003 222896 267015
rect 253360 267003 253366 267015
rect 253418 267003 253424 267055
rect 254128 267003 254134 267055
rect 254186 267043 254192 267055
rect 258370 267043 258398 267163
rect 258640 267151 258646 267203
rect 258698 267191 258704 267203
rect 477424 267191 477430 267203
rect 258698 267163 477430 267191
rect 258698 267151 258704 267163
rect 477424 267151 477430 267163
rect 477482 267151 477488 267203
rect 258448 267077 258454 267129
rect 258506 267117 258512 267129
rect 484432 267117 484438 267129
rect 258506 267089 484438 267117
rect 258506 267077 258512 267089
rect 484432 267077 484438 267089
rect 484490 267077 484496 267129
rect 480976 267043 480982 267055
rect 254186 267015 258302 267043
rect 258370 267015 480982 267043
rect 254186 267003 254192 267015
rect 189520 266929 189526 266981
rect 189578 266969 189584 266981
rect 223024 266969 223030 266981
rect 189578 266941 223030 266969
rect 189578 266929 189584 266941
rect 223024 266929 223030 266941
rect 223082 266929 223088 266981
rect 254512 266929 254518 266981
rect 254570 266969 254576 266981
rect 258274 266969 258302 267015
rect 480976 267003 480982 267015
rect 481034 267003 481040 267055
rect 487792 266969 487798 266981
rect 254570 266941 256478 266969
rect 258274 266941 487798 266969
rect 254570 266929 254576 266941
rect 203824 266855 203830 266907
rect 203882 266895 203888 266907
rect 252016 266895 252022 266907
rect 203882 266867 252022 266895
rect 203882 266855 203888 266867
rect 252016 266855 252022 266867
rect 252074 266855 252080 266907
rect 204976 266781 204982 266833
rect 205034 266821 205040 266833
rect 256240 266821 256246 266833
rect 205034 266793 256246 266821
rect 205034 266781 205040 266793
rect 256240 266781 256246 266793
rect 256298 266781 256304 266833
rect 256450 266821 256478 266941
rect 487792 266929 487798 266941
rect 487850 266929 487856 266981
rect 256528 266855 256534 266907
rect 256586 266895 256592 266907
rect 274768 266895 274774 266907
rect 256586 266867 274774 266895
rect 256586 266855 256592 266867
rect 274768 266855 274774 266867
rect 274826 266855 274832 266907
rect 276400 266855 276406 266907
rect 276458 266895 276464 266907
rect 294160 266895 294166 266907
rect 276458 266867 294166 266895
rect 276458 266855 276464 266867
rect 294160 266855 294166 266867
rect 294218 266855 294224 266907
rect 318064 266855 318070 266907
rect 318122 266895 318128 266907
rect 321712 266895 321718 266907
rect 318122 266867 321718 266895
rect 318122 266855 318128 266867
rect 321712 266855 321718 266867
rect 321770 266855 321776 266907
rect 321808 266855 321814 266907
rect 321866 266895 321872 266907
rect 553456 266895 553462 266907
rect 321866 266867 553462 266895
rect 321866 266855 321872 266867
rect 553456 266855 553462 266867
rect 553514 266855 553520 266907
rect 491632 266821 491638 266833
rect 256450 266793 491638 266821
rect 491632 266781 491638 266793
rect 491690 266781 491696 266833
rect 200176 266707 200182 266759
rect 200234 266747 200240 266759
rect 274192 266747 274198 266759
rect 200234 266719 274198 266747
rect 200234 266707 200240 266719
rect 274192 266707 274198 266719
rect 274250 266707 274256 266759
rect 288304 266707 288310 266759
rect 288362 266747 288368 266759
rect 314416 266747 314422 266759
rect 288362 266719 314422 266747
rect 288362 266707 288368 266719
rect 314416 266707 314422 266719
rect 314474 266707 314480 266759
rect 318640 266707 318646 266759
rect 318698 266747 318704 266759
rect 321616 266747 321622 266759
rect 318698 266719 321622 266747
rect 318698 266707 318704 266719
rect 321616 266707 321622 266719
rect 321674 266707 321680 266759
rect 321712 266707 321718 266759
rect 321770 266747 321776 266759
rect 557104 266747 557110 266759
rect 321770 266719 557110 266747
rect 321770 266707 321776 266719
rect 557104 266707 557110 266719
rect 557162 266707 557168 266759
rect 201424 266633 201430 266685
rect 201482 266673 201488 266685
rect 253840 266673 253846 266685
rect 201482 266645 253846 266673
rect 201482 266633 201488 266645
rect 253840 266633 253846 266645
rect 253898 266633 253904 266685
rect 254704 266633 254710 266685
rect 254762 266673 254768 266685
rect 495280 266673 495286 266685
rect 254762 266645 495286 266673
rect 254762 266633 254768 266645
rect 495280 266633 495286 266645
rect 495338 266633 495344 266685
rect 196720 266559 196726 266611
rect 196778 266599 196784 266611
rect 273616 266599 273622 266611
rect 196778 266571 273622 266599
rect 196778 266559 196784 266571
rect 273616 266559 273622 266571
rect 273674 266559 273680 266611
rect 289360 266559 289366 266611
rect 289418 266599 289424 266611
rect 321520 266599 321526 266611
rect 289418 266571 321526 266599
rect 289418 266559 289424 266571
rect 321520 266559 321526 266571
rect 321578 266559 321584 266611
rect 321616 266559 321622 266611
rect 321674 266599 321680 266611
rect 560656 266599 560662 266611
rect 321674 266571 560662 266599
rect 321674 266559 321680 266571
rect 560656 266559 560662 266571
rect 560714 266559 560720 266611
rect 197872 266485 197878 266537
rect 197930 266525 197936 266537
rect 255760 266525 255766 266537
rect 197930 266497 255766 266525
rect 197930 266485 197936 266497
rect 255760 266485 255766 266497
rect 255818 266485 255824 266537
rect 498832 266525 498838 266537
rect 255874 266497 498838 266525
rect 193072 266411 193078 266463
rect 193130 266451 193136 266463
rect 250000 266451 250006 266463
rect 193130 266423 250006 266451
rect 193130 266411 193136 266423
rect 250000 266411 250006 266423
rect 250058 266411 250064 266463
rect 250096 266411 250102 266463
rect 250154 266451 250160 266463
rect 250154 266423 254558 266451
rect 250154 266411 250160 266423
rect 138352 266337 138358 266389
rect 138410 266377 138416 266389
rect 254416 266377 254422 266389
rect 138410 266349 254422 266377
rect 138410 266337 138416 266349
rect 254416 266337 254422 266349
rect 254474 266337 254480 266389
rect 254530 266377 254558 266423
rect 255184 266411 255190 266463
rect 255242 266451 255248 266463
rect 255874 266451 255902 266497
rect 498832 266485 498838 266497
rect 498890 266485 498896 266537
rect 548560 266485 548566 266537
rect 548618 266525 548624 266537
rect 573136 266525 573142 266537
rect 548618 266497 573142 266525
rect 548618 266485 548624 266497
rect 573136 266485 573142 266497
rect 573194 266485 573200 266537
rect 255242 266423 255902 266451
rect 255242 266411 255248 266423
rect 266032 266411 266038 266463
rect 266090 266451 266096 266463
rect 299536 266451 299542 266463
rect 266090 266423 299542 266451
rect 266090 266411 266096 266423
rect 299536 266411 299542 266423
rect 299594 266411 299600 266463
rect 317968 266451 317974 266463
rect 299650 266423 317974 266451
rect 259120 266377 259126 266389
rect 254530 266349 259126 266377
rect 259120 266337 259126 266349
rect 259178 266337 259184 266389
rect 288688 266337 288694 266389
rect 288746 266377 288752 266389
rect 299650 266377 299678 266423
rect 317968 266411 317974 266423
rect 318026 266411 318032 266463
rect 318736 266411 318742 266463
rect 318794 266451 318800 266463
rect 564208 266451 564214 266463
rect 318794 266423 564214 266451
rect 318794 266411 318800 266423
rect 564208 266411 564214 266423
rect 564266 266411 564272 266463
rect 288746 266349 299678 266377
rect 288746 266337 288752 266349
rect 314224 266337 314230 266389
rect 314282 266377 314288 266389
rect 319600 266377 319606 266389
rect 314282 266349 319606 266377
rect 314282 266337 314288 266349
rect 319600 266337 319606 266349
rect 319658 266337 319664 266389
rect 319696 266337 319702 266389
rect 319754 266377 319760 266389
rect 571312 266377 571318 266389
rect 319754 266349 571318 266377
rect 319754 266337 319760 266349
rect 571312 266337 571318 266349
rect 571370 266337 571376 266389
rect 194320 266263 194326 266315
rect 194378 266303 194384 266315
rect 329008 266303 329014 266315
rect 194378 266275 329014 266303
rect 194378 266263 194384 266275
rect 329008 266263 329014 266275
rect 329066 266263 329072 266315
rect 372880 266263 372886 266315
rect 372938 266303 372944 266315
rect 551056 266303 551062 266315
rect 372938 266275 551062 266303
rect 372938 266263 372944 266275
rect 551056 266263 551062 266275
rect 551114 266263 551120 266315
rect 208528 266189 208534 266241
rect 208586 266229 208592 266241
rect 208586 266201 249950 266229
rect 208586 266189 208592 266201
rect 249922 266155 249950 266201
rect 250000 266189 250006 266241
rect 250058 266229 250064 266241
rect 250058 266201 272798 266229
rect 250058 266189 250064 266201
rect 257488 266155 257494 266167
rect 249922 266127 257494 266155
rect 257488 266115 257494 266127
rect 257546 266115 257552 266167
rect 257584 266115 257590 266167
rect 257642 266155 257648 266167
rect 272656 266155 272662 266167
rect 257642 266127 272662 266155
rect 257642 266115 257648 266127
rect 272656 266115 272662 266127
rect 272714 266115 272720 266167
rect 272770 266155 272798 266201
rect 272848 266189 272854 266241
rect 272906 266229 272912 266241
rect 445264 266229 445270 266241
rect 272906 266201 445270 266229
rect 272906 266189 272912 266201
rect 445264 266189 445270 266201
rect 445322 266189 445328 266241
rect 273520 266155 273526 266167
rect 272770 266127 273526 266155
rect 273520 266115 273526 266127
rect 273578 266115 273584 266167
rect 274096 266115 274102 266167
rect 274154 266155 274160 266167
rect 441712 266155 441718 266167
rect 274154 266127 441718 266155
rect 274154 266115 274160 266127
rect 441712 266115 441718 266127
rect 441770 266115 441776 266167
rect 254896 266041 254902 266093
rect 254954 266081 254960 266093
rect 256336 266081 256342 266093
rect 254954 266053 256342 266081
rect 254954 266041 254960 266053
rect 256336 266041 256342 266053
rect 256394 266041 256400 266093
rect 256432 266041 256438 266093
rect 256490 266081 256496 266093
rect 394576 266081 394582 266093
rect 256490 266053 394582 266081
rect 256490 266041 256496 266053
rect 394576 266041 394582 266053
rect 394634 266041 394640 266093
rect 394768 266041 394774 266093
rect 394826 266081 394832 266093
rect 394960 266081 394966 266093
rect 394826 266053 394966 266081
rect 394826 266041 394832 266053
rect 394960 266041 394966 266053
rect 395018 266041 395024 266093
rect 249328 265967 249334 266019
rect 249386 266007 249392 266019
rect 388816 266007 388822 266019
rect 249386 265979 388822 266007
rect 249386 265967 249392 265979
rect 388816 265967 388822 265979
rect 388874 265967 388880 266019
rect 218032 265893 218038 265945
rect 218090 265933 218096 265945
rect 276496 265933 276502 265945
rect 218090 265905 276502 265933
rect 218090 265893 218096 265905
rect 276496 265893 276502 265905
rect 276554 265893 276560 265945
rect 300688 265893 300694 265945
rect 300746 265933 300752 265945
rect 414352 265933 414358 265945
rect 300746 265905 414358 265933
rect 300746 265893 300752 265905
rect 414352 265893 414358 265905
rect 414410 265893 414416 265945
rect 249712 265819 249718 265871
rect 249770 265859 249776 265871
rect 256432 265859 256438 265871
rect 249770 265831 256438 265859
rect 249770 265819 249776 265831
rect 256432 265819 256438 265831
rect 256490 265819 256496 265871
rect 267856 265819 267862 265871
rect 267914 265859 267920 265871
rect 334960 265859 334966 265871
rect 267914 265831 334966 265859
rect 267914 265819 267920 265831
rect 334960 265819 334966 265831
rect 335018 265819 335024 265871
rect 356080 265819 356086 265871
rect 356138 265859 356144 265871
rect 406096 265859 406102 265871
rect 356138 265831 406102 265859
rect 356138 265819 356144 265831
rect 406096 265819 406102 265831
rect 406154 265819 406160 265871
rect 221488 265745 221494 265797
rect 221546 265785 221552 265797
rect 276976 265785 276982 265797
rect 221546 265757 276982 265785
rect 221546 265745 221552 265757
rect 276976 265745 276982 265757
rect 277034 265745 277040 265797
rect 294064 265745 294070 265797
rect 294122 265785 294128 265797
rect 360784 265785 360790 265797
rect 294122 265757 360790 265785
rect 294122 265745 294128 265757
rect 360784 265745 360790 265757
rect 360842 265745 360848 265797
rect 362128 265745 362134 265797
rect 362186 265785 362192 265797
rect 397744 265785 397750 265797
rect 362186 265757 397750 265785
rect 362186 265745 362192 265757
rect 397744 265745 397750 265757
rect 397802 265745 397808 265797
rect 225232 265671 225238 265723
rect 225290 265711 225296 265723
rect 277360 265711 277366 265723
rect 225290 265683 277366 265711
rect 225290 265671 225296 265683
rect 277360 265671 277366 265683
rect 277418 265671 277424 265723
rect 293680 265671 293686 265723
rect 293738 265711 293744 265723
rect 357232 265711 357238 265723
rect 293738 265683 357238 265711
rect 293738 265671 293744 265683
rect 357232 265671 357238 265683
rect 357290 265671 357296 265723
rect 373456 265671 373462 265723
rect 373514 265711 373520 265723
rect 402352 265711 402358 265723
rect 373514 265683 402358 265711
rect 373514 265671 373520 265683
rect 402352 265671 402358 265683
rect 402410 265671 402416 265723
rect 214576 265597 214582 265649
rect 214634 265637 214640 265649
rect 275824 265637 275830 265649
rect 214634 265609 275830 265637
rect 214634 265597 214640 265609
rect 275824 265597 275830 265609
rect 275882 265597 275888 265649
rect 275920 265597 275926 265649
rect 275978 265637 275984 265649
rect 337072 265637 337078 265649
rect 275978 265609 337078 265637
rect 275978 265597 275984 265609
rect 337072 265597 337078 265609
rect 337130 265597 337136 265649
rect 355600 265597 355606 265649
rect 355658 265637 355664 265649
rect 403216 265637 403222 265649
rect 355658 265609 403222 265637
rect 355658 265597 355664 265609
rect 403216 265597 403222 265609
rect 403274 265597 403280 265649
rect 228784 265523 228790 265575
rect 228842 265563 228848 265575
rect 228842 265535 257822 265563
rect 228842 265523 228848 265535
rect 232432 265449 232438 265501
rect 232490 265489 232496 265501
rect 257794 265489 257822 265535
rect 272656 265523 272662 265575
rect 272714 265563 272720 265575
rect 279568 265563 279574 265575
rect 272714 265535 279574 265563
rect 272714 265523 272720 265535
rect 279568 265523 279574 265535
rect 279626 265523 279632 265575
rect 293104 265523 293110 265575
rect 293162 265563 293168 265575
rect 353680 265563 353686 265575
rect 293162 265535 353686 265563
rect 293162 265523 293168 265535
rect 353680 265523 353686 265535
rect 353738 265523 353744 265575
rect 354928 265523 354934 265575
rect 354986 265563 354992 265575
rect 404464 265563 404470 265575
rect 354986 265535 404470 265563
rect 354986 265523 354992 265535
rect 404464 265523 404470 265535
rect 404522 265523 404528 265575
rect 277840 265489 277846 265501
rect 232490 265461 257726 265489
rect 257794 265461 277846 265489
rect 232490 265449 232496 265461
rect 243088 265375 243094 265427
rect 243146 265415 243152 265427
rect 257584 265415 257590 265427
rect 243146 265387 257590 265415
rect 243146 265375 243152 265387
rect 257584 265375 257590 265387
rect 257642 265375 257648 265427
rect 257698 265415 257726 265461
rect 277840 265449 277846 265461
rect 277898 265449 277904 265501
rect 292624 265449 292630 265501
rect 292682 265489 292688 265501
rect 350032 265489 350038 265501
rect 292682 265461 350038 265489
rect 292682 265449 292688 265461
rect 350032 265449 350038 265461
rect 350090 265449 350096 265501
rect 367216 265449 367222 265501
rect 367274 265489 367280 265501
rect 394096 265489 394102 265501
rect 367274 265461 394102 265489
rect 367274 265449 367280 265461
rect 394096 265449 394102 265461
rect 394154 265449 394160 265501
rect 278032 265415 278038 265427
rect 257698 265387 278038 265415
rect 278032 265375 278038 265387
rect 278090 265375 278096 265427
rect 292144 265375 292150 265427
rect 292202 265415 292208 265427
rect 346576 265415 346582 265427
rect 292202 265387 346582 265415
rect 292202 265375 292208 265387
rect 346576 265375 346582 265387
rect 346634 265375 346640 265427
rect 354544 265375 354550 265427
rect 354602 265415 354608 265427
rect 401200 265415 401206 265427
rect 354602 265387 401206 265415
rect 354602 265375 354608 265387
rect 401200 265375 401206 265387
rect 401258 265375 401264 265427
rect 235888 265301 235894 265353
rect 235946 265341 235952 265353
rect 278512 265341 278518 265353
rect 235946 265313 278518 265341
rect 235946 265301 235952 265313
rect 278512 265301 278518 265313
rect 278570 265301 278576 265353
rect 292048 265301 292054 265353
rect 292106 265341 292112 265353
rect 342736 265341 342742 265353
rect 292106 265313 342742 265341
rect 292106 265301 292112 265313
rect 342736 265301 342742 265313
rect 342794 265301 342800 265353
rect 357136 265301 357142 265353
rect 357194 265341 357200 265353
rect 382288 265341 382294 265353
rect 357194 265313 382294 265341
rect 357194 265301 357200 265313
rect 382288 265301 382294 265313
rect 382346 265301 382352 265353
rect 382384 265301 382390 265353
rect 382442 265341 382448 265353
rect 391696 265341 391702 265353
rect 382442 265313 391702 265341
rect 382442 265301 382448 265313
rect 391696 265301 391702 265313
rect 391754 265301 391760 265353
rect 239440 265227 239446 265279
rect 239498 265267 239504 265279
rect 279088 265267 279094 265279
rect 239498 265239 279094 265267
rect 239498 265227 239504 265239
rect 279088 265227 279094 265239
rect 279146 265227 279152 265279
rect 291568 265227 291574 265279
rect 291626 265267 291632 265279
rect 339088 265267 339094 265279
rect 291626 265239 339094 265267
rect 291626 265227 291632 265239
rect 339088 265227 339094 265239
rect 339146 265227 339152 265279
rect 358864 265227 358870 265279
rect 358922 265267 358928 265279
rect 374416 265267 374422 265279
rect 358922 265239 374422 265267
rect 358922 265227 358928 265239
rect 374416 265227 374422 265239
rect 374474 265227 374480 265279
rect 374992 265227 374998 265279
rect 375050 265267 375056 265279
rect 400240 265267 400246 265279
rect 375050 265239 400246 265267
rect 375050 265227 375056 265239
rect 400240 265227 400246 265239
rect 400298 265227 400304 265279
rect 246640 265153 246646 265205
rect 246698 265193 246704 265205
rect 280048 265193 280054 265205
rect 246698 265165 280054 265193
rect 246698 265153 246704 265165
rect 280048 265153 280054 265165
rect 280106 265153 280112 265205
rect 290416 265153 290422 265205
rect 290474 265193 290480 265205
rect 318160 265193 318166 265205
rect 290474 265165 318166 265193
rect 290474 265153 290480 265165
rect 318160 265153 318166 265165
rect 318218 265153 318224 265205
rect 335824 265193 335830 265205
rect 318274 265165 335830 265193
rect 141136 265079 141142 265131
rect 141194 265119 141200 265131
rect 151120 265119 151126 265131
rect 141194 265091 151126 265119
rect 141194 265079 141200 265091
rect 151120 265079 151126 265091
rect 151178 265079 151184 265131
rect 181456 265079 181462 265131
rect 181514 265119 181520 265131
rect 191536 265119 191542 265131
rect 181514 265091 191542 265119
rect 181514 265079 181520 265091
rect 191536 265079 191542 265091
rect 191594 265079 191600 265131
rect 250192 265079 250198 265131
rect 250250 265119 250256 265131
rect 280144 265119 280150 265131
rect 250250 265091 280150 265119
rect 250250 265079 250256 265091
rect 280144 265079 280150 265091
rect 280202 265079 280208 265131
rect 291184 265079 291190 265131
rect 291242 265119 291248 265131
rect 318274 265119 318302 265165
rect 335824 265153 335830 265165
rect 335882 265153 335888 265205
rect 367120 265153 367126 265205
rect 367178 265193 367184 265205
rect 390544 265193 390550 265205
rect 367178 265165 390550 265193
rect 367178 265153 367184 265165
rect 390544 265153 390550 265165
rect 390602 265153 390608 265205
rect 291242 265091 318302 265119
rect 291242 265079 291248 265091
rect 318352 265079 318358 265131
rect 318410 265119 318416 265131
rect 332272 265119 332278 265131
rect 318410 265091 332278 265119
rect 318410 265079 318416 265091
rect 332272 265079 332278 265091
rect 332330 265079 332336 265131
rect 369616 265079 369622 265131
rect 369674 265119 369680 265131
rect 373168 265119 373174 265131
rect 369674 265091 373174 265119
rect 369674 265079 369680 265091
rect 373168 265079 373174 265091
rect 373226 265079 373232 265131
rect 377872 265079 377878 265131
rect 377930 265119 377936 265131
rect 380080 265119 380086 265131
rect 377930 265091 380086 265119
rect 377930 265079 377936 265091
rect 380080 265079 380086 265091
rect 380138 265079 380144 265131
rect 380464 265079 380470 265131
rect 380522 265119 380528 265131
rect 388912 265119 388918 265131
rect 380522 265091 388918 265119
rect 380522 265079 380528 265091
rect 388912 265079 388918 265091
rect 388970 265079 388976 265131
rect 254032 265005 254038 265057
rect 254090 265045 254096 265057
rect 280624 265045 280630 265057
rect 254090 265017 280630 265045
rect 254090 265005 254096 265017
rect 280624 265005 280630 265017
rect 280682 265005 280688 265057
rect 290032 265005 290038 265057
rect 290090 265045 290096 265057
rect 328720 265045 328726 265057
rect 290090 265017 328726 265045
rect 290090 265005 290096 265017
rect 328720 265005 328726 265017
rect 328778 265005 328784 265057
rect 334018 265017 338942 265045
rect 87760 264931 87766 264983
rect 87818 264971 87824 264983
rect 106576 264971 106582 264983
rect 87818 264943 106582 264971
rect 87818 264931 87824 264943
rect 106576 264931 106582 264943
rect 106634 264931 106640 264983
rect 126736 264931 126742 264983
rect 126794 264971 126800 264983
rect 141136 264971 141142 264983
rect 126794 264943 141142 264971
rect 126794 264931 126800 264943
rect 141136 264931 141142 264943
rect 141194 264931 141200 264983
rect 151120 264931 151126 264983
rect 151178 264971 151184 264983
rect 168304 264971 168310 264983
rect 151178 264943 168310 264971
rect 151178 264931 151184 264943
rect 168304 264931 168310 264943
rect 168362 264931 168368 264983
rect 168400 264931 168406 264983
rect 168458 264971 168464 264983
rect 168458 264943 191486 264971
rect 168458 264931 168464 264943
rect 86434 264869 106526 264897
rect 66256 264783 66262 264835
rect 66314 264823 66320 264835
rect 86434 264823 86462 264869
rect 66314 264795 86462 264823
rect 106498 264823 106526 264869
rect 126754 264869 145790 264897
rect 126754 264823 126782 264869
rect 106498 264795 126782 264823
rect 145762 264823 145790 264869
rect 168400 264823 168406 264835
rect 145762 264795 168406 264823
rect 66314 264783 66320 264795
rect 168400 264783 168406 264795
rect 168458 264783 168464 264835
rect 168496 264783 168502 264835
rect 168554 264823 168560 264835
rect 181456 264823 181462 264835
rect 168554 264795 181462 264823
rect 168554 264783 168560 264795
rect 181456 264783 181462 264795
rect 181514 264783 181520 264835
rect 191458 264823 191486 264943
rect 202576 264931 202582 264983
rect 202634 264971 202640 264983
rect 218896 264971 218902 264983
rect 202634 264943 218902 264971
rect 202634 264931 202640 264943
rect 218896 264931 218902 264943
rect 218954 264931 218960 264983
rect 253360 264931 253366 264983
rect 253418 264971 253424 264983
rect 332752 264971 332758 264983
rect 253418 264943 332758 264971
rect 253418 264931 253424 264943
rect 332752 264931 332758 264943
rect 332810 264931 332816 264983
rect 333424 264931 333430 264983
rect 333482 264971 333488 264983
rect 334018 264971 334046 265017
rect 333482 264943 334046 264971
rect 333482 264931 333488 264943
rect 334096 264931 334102 264983
rect 334154 264971 334160 264983
rect 338800 264971 338806 264983
rect 334154 264943 338806 264971
rect 334154 264931 334160 264943
rect 338800 264931 338806 264943
rect 338858 264931 338864 264983
rect 338914 264971 338942 265017
rect 350896 265005 350902 265057
rect 350954 265045 350960 265057
rect 350954 265017 351422 265045
rect 350954 265005 350960 265017
rect 346288 264971 346294 264983
rect 338914 264943 346294 264971
rect 346288 264931 346294 264943
rect 346346 264931 346352 264983
rect 348400 264931 348406 264983
rect 348458 264971 348464 264983
rect 351280 264971 351286 264983
rect 348458 264943 351286 264971
rect 348458 264931 348464 264943
rect 351280 264931 351286 264943
rect 351338 264931 351344 264983
rect 351394 264971 351422 265017
rect 365680 265005 365686 265057
rect 365738 265045 365744 265057
rect 379888 265045 379894 265057
rect 365738 265017 379894 265045
rect 365738 265005 365744 265017
rect 379888 265005 379894 265017
rect 379946 265005 379952 265057
rect 381136 265005 381142 265057
rect 381194 265045 381200 265057
rect 386032 265045 386038 265057
rect 381194 265017 386038 265045
rect 381194 265005 381200 265017
rect 386032 265005 386038 265017
rect 386090 265005 386096 265057
rect 369136 264971 369142 264983
rect 351394 264943 369142 264971
rect 369136 264931 369142 264943
rect 369194 264931 369200 264983
rect 372400 264931 372406 264983
rect 372458 264971 372464 264983
rect 547600 264971 547606 264983
rect 372458 264943 547606 264971
rect 372458 264931 372464 264943
rect 547600 264931 547606 264943
rect 547658 264931 547664 264983
rect 191536 264857 191542 264909
rect 191594 264897 191600 264909
rect 216688 264897 216694 264909
rect 191594 264869 216694 264897
rect 191594 264857 191600 264869
rect 216688 264857 216694 264869
rect 216746 264857 216752 264909
rect 223024 264857 223030 264909
rect 223082 264897 223088 264909
rect 415312 264897 415318 264909
rect 223082 264869 415318 264897
rect 223082 264857 223088 264869
rect 415312 264857 415318 264869
rect 415370 264857 415376 264909
rect 216016 264823 216022 264835
rect 191458 264795 216022 264823
rect 216016 264783 216022 264795
rect 216074 264783 216080 264835
rect 227632 264783 227638 264835
rect 227690 264823 227696 264835
rect 249040 264823 249046 264835
rect 227690 264795 249046 264823
rect 227690 264783 227696 264795
rect 249040 264783 249046 264795
rect 249098 264783 249104 264835
rect 250384 264783 250390 264835
rect 250442 264823 250448 264835
rect 438064 264823 438070 264835
rect 250442 264795 438070 264823
rect 250442 264783 250448 264795
rect 438064 264783 438070 264795
rect 438122 264783 438128 264835
rect 106576 264709 106582 264761
rect 106634 264749 106640 264761
rect 126736 264749 126742 264761
rect 106634 264721 126742 264749
rect 106634 264709 106640 264721
rect 126736 264709 126742 264721
rect 126794 264709 126800 264761
rect 188368 264709 188374 264761
rect 188426 264749 188432 264761
rect 414832 264749 414838 264761
rect 188426 264721 414838 264749
rect 188426 264709 188432 264721
rect 414832 264709 414838 264721
rect 414890 264709 414896 264761
rect 178864 264635 178870 264687
rect 178922 264675 178928 264687
rect 412624 264675 412630 264687
rect 178922 264647 412630 264675
rect 178922 264635 178928 264647
rect 412624 264635 412630 264647
rect 412682 264635 412688 264687
rect 177616 264561 177622 264613
rect 177674 264601 177680 264613
rect 412528 264601 412534 264613
rect 177674 264573 412534 264601
rect 177674 264561 177680 264573
rect 412528 264561 412534 264573
rect 412586 264561 412592 264613
rect 67312 264487 67318 264539
rect 67370 264527 67376 264539
rect 87760 264527 87766 264539
rect 67370 264499 87766 264527
rect 67370 264487 67376 264499
rect 87760 264487 87766 264499
rect 87818 264487 87824 264539
rect 171664 264487 171670 264539
rect 171722 264527 171728 264539
rect 410896 264527 410902 264539
rect 171722 264499 410902 264527
rect 171722 264487 171728 264499
rect 410896 264487 410902 264499
rect 410954 264487 410960 264539
rect 170512 264413 170518 264465
rect 170570 264453 170576 264465
rect 410512 264453 410518 264465
rect 170570 264425 410518 264453
rect 170570 264413 170576 264425
rect 410512 264413 410518 264425
rect 410570 264413 410576 264465
rect 164560 264339 164566 264391
rect 164618 264379 164624 264391
rect 409360 264379 409366 264391
rect 164618 264351 409366 264379
rect 164618 264339 164624 264351
rect 409360 264339 409366 264351
rect 409418 264339 409424 264391
rect 42256 264265 42262 264317
rect 42314 264305 42320 264317
rect 53296 264305 53302 264317
rect 42314 264277 53302 264305
rect 42314 264265 42320 264277
rect 53296 264265 53302 264277
rect 53354 264265 53360 264317
rect 163408 264265 163414 264317
rect 163466 264305 163472 264317
rect 408976 264305 408982 264317
rect 163466 264277 408982 264305
rect 163466 264265 163472 264277
rect 408976 264265 408982 264277
rect 409034 264265 409040 264317
rect 156208 264191 156214 264243
rect 156266 264231 156272 264243
rect 407248 264231 407254 264243
rect 156266 264203 407254 264231
rect 156266 264191 156272 264203
rect 407248 264191 407254 264203
rect 407306 264191 407312 264243
rect 157456 264117 157462 264169
rect 157514 264157 157520 264169
rect 407728 264157 407734 264169
rect 157514 264129 407734 264157
rect 157514 264117 157520 264129
rect 407728 264117 407734 264129
rect 407786 264117 407792 264169
rect 150256 264043 150262 264095
rect 150314 264083 150320 264095
rect 406000 264083 406006 264095
rect 150314 264055 406006 264083
rect 150314 264043 150320 264055
rect 406000 264043 406006 264055
rect 406058 264043 406064 264095
rect 149104 263969 149110 264021
rect 149162 264009 149168 264021
rect 405520 264009 405526 264021
rect 149162 263981 405526 264009
rect 149162 263969 149168 263981
rect 405520 263969 405526 263981
rect 405578 263969 405584 264021
rect 405712 263969 405718 264021
rect 405770 264009 405776 264021
rect 410320 264009 410326 264021
rect 405770 263981 410326 264009
rect 405770 263969 405776 263981
rect 410320 263969 410326 263981
rect 410378 263969 410384 264021
rect 145552 263895 145558 263947
rect 145610 263935 145616 263947
rect 404368 263935 404374 263947
rect 145610 263907 404374 263935
rect 145610 263895 145616 263907
rect 404368 263895 404374 263907
rect 404426 263895 404432 263947
rect 405904 263895 405910 263947
rect 405962 263935 405968 263947
rect 412048 263935 412054 263947
rect 405962 263907 412054 263935
rect 405962 263895 405968 263907
rect 412048 263895 412054 263907
rect 412106 263895 412112 263947
rect 146992 263821 146998 263873
rect 147050 263861 147056 263873
rect 405040 263861 405046 263873
rect 147050 263833 405046 263861
rect 147050 263821 147056 263833
rect 405040 263821 405046 263833
rect 405098 263821 405104 263873
rect 405136 263821 405142 263873
rect 405194 263861 405200 263873
rect 406576 263861 406582 263873
rect 405194 263833 406582 263861
rect 405194 263821 405200 263833
rect 406576 263821 406582 263833
rect 406634 263821 406640 263873
rect 132496 263747 132502 263799
rect 132554 263787 132560 263799
rect 401584 263787 401590 263799
rect 132554 263759 401590 263787
rect 132554 263747 132560 263759
rect 401584 263747 401590 263759
rect 401642 263747 401648 263799
rect 403024 263747 403030 263799
rect 403082 263787 403088 263799
rect 414256 263787 414262 263799
rect 403082 263759 414262 263787
rect 403082 263747 403088 263759
rect 414256 263747 414262 263759
rect 414314 263747 414320 263799
rect 107440 263673 107446 263725
rect 107498 263713 107504 263725
rect 395248 263713 395254 263725
rect 107498 263685 395254 263713
rect 107498 263673 107504 263685
rect 395248 263673 395254 263685
rect 395306 263673 395312 263725
rect 395344 263673 395350 263725
rect 395402 263713 395408 263725
rect 396496 263713 396502 263725
rect 395402 263685 396502 263713
rect 395402 263673 395408 263685
rect 396496 263673 396502 263685
rect 396554 263673 396560 263725
rect 398608 263673 398614 263725
rect 398666 263713 398672 263725
rect 403984 263713 403990 263725
rect 398666 263685 403990 263713
rect 398666 263673 398672 263685
rect 403984 263673 403990 263685
rect 404042 263673 404048 263725
rect 405616 263673 405622 263725
rect 405674 263713 405680 263725
rect 413776 263713 413782 263725
rect 405674 263685 413782 263713
rect 405674 263673 405680 263685
rect 413776 263673 413782 263685
rect 413834 263673 413840 263725
rect 91984 263599 91990 263651
rect 92042 263639 92048 263651
rect 391504 263639 391510 263651
rect 92042 263611 391510 263639
rect 92042 263599 92048 263611
rect 391504 263599 391510 263611
rect 391562 263599 391568 263651
rect 394960 263599 394966 263651
rect 395018 263639 395024 263651
rect 408112 263639 408118 263651
rect 395018 263611 408118 263639
rect 395018 263599 395024 263611
rect 408112 263599 408118 263611
rect 408170 263599 408176 263651
rect 42256 263525 42262 263577
rect 42314 263565 42320 263577
rect 53392 263565 53398 263577
rect 42314 263537 53398 263565
rect 42314 263525 42320 263537
rect 53392 263525 53398 263537
rect 53450 263525 53456 263577
rect 76528 263525 76534 263577
rect 76586 263565 76592 263577
rect 387184 263565 387190 263577
rect 76586 263537 387190 263565
rect 76586 263525 76592 263537
rect 387184 263525 387190 263537
rect 387242 263525 387248 263577
rect 388720 263525 388726 263577
rect 388778 263565 388784 263577
rect 390256 263565 390262 263577
rect 388778 263537 390262 263565
rect 388778 263525 388784 263537
rect 390256 263525 390262 263537
rect 390314 263525 390320 263577
rect 390352 263525 390358 263577
rect 390410 263565 390416 263577
rect 394288 263565 394294 263577
rect 390410 263537 394294 263565
rect 390410 263525 390416 263537
rect 394288 263525 394294 263537
rect 394346 263525 394352 263577
rect 394864 263525 394870 263577
rect 394922 263565 394928 263577
rect 406096 263565 406102 263577
rect 394922 263537 406102 263565
rect 394922 263525 394928 263537
rect 406096 263525 406102 263537
rect 406154 263525 406160 263577
rect 195472 263451 195478 263503
rect 195530 263491 195536 263503
rect 218128 263491 218134 263503
rect 195530 263463 218134 263491
rect 195530 263451 195536 263463
rect 218128 263451 218134 263463
rect 218186 263451 218192 263503
rect 223792 263451 223798 263503
rect 223850 263491 223856 263503
rect 241840 263491 241846 263503
rect 223850 263463 241846 263491
rect 223850 263451 223856 263463
rect 241840 263451 241846 263463
rect 241898 263451 241904 263503
rect 256336 263451 256342 263503
rect 256394 263491 256400 263503
rect 336592 263491 336598 263503
rect 256394 263463 336598 263491
rect 256394 263451 256400 263463
rect 336592 263451 336598 263463
rect 336650 263451 336656 263503
rect 353392 263451 353398 263503
rect 353450 263491 353456 263503
rect 367120 263491 367126 263503
rect 353450 263463 367126 263491
rect 353450 263451 353456 263463
rect 367120 263451 367126 263463
rect 367178 263451 367184 263503
rect 371440 263451 371446 263503
rect 371498 263491 371504 263503
rect 540400 263491 540406 263503
rect 371498 263463 540406 263491
rect 371498 263451 371504 263463
rect 540400 263451 540406 263463
rect 540458 263451 540464 263503
rect 191248 263377 191254 263429
rect 191306 263417 191312 263429
rect 198736 263417 198742 263429
rect 191306 263389 198742 263417
rect 191306 263377 191312 263389
rect 198736 263377 198742 263389
rect 198794 263377 198800 263429
rect 224656 263377 224662 263429
rect 224714 263417 224720 263429
rect 227632 263417 227638 263429
rect 224714 263389 227638 263417
rect 224714 263377 224720 263389
rect 227632 263377 227638 263389
rect 227690 263377 227696 263429
rect 253648 263377 253654 263429
rect 253706 263417 253712 263429
rect 331600 263417 331606 263429
rect 253706 263389 331606 263417
rect 253706 263377 253712 263389
rect 331600 263377 331606 263389
rect 331658 263377 331664 263429
rect 334192 263377 334198 263429
rect 334250 263417 334256 263429
rect 339760 263417 339766 263429
rect 334250 263389 339766 263417
rect 334250 263377 334256 263389
rect 339760 263377 339766 263389
rect 339818 263377 339824 263429
rect 353872 263377 353878 263429
rect 353930 263417 353936 263429
rect 367216 263417 367222 263429
rect 353930 263389 367222 263417
rect 353930 263377 353936 263389
rect 367216 263377 367222 263389
rect 367274 263377 367280 263429
rect 370672 263377 370678 263429
rect 370730 263417 370736 263429
rect 533200 263417 533206 263429
rect 370730 263389 533206 263417
rect 370730 263377 370736 263389
rect 533200 263377 533206 263389
rect 533258 263377 533264 263429
rect 199120 263303 199126 263355
rect 199178 263343 199184 263355
rect 218320 263343 218326 263355
rect 199178 263315 218326 263343
rect 199178 263303 199184 263315
rect 218320 263303 218326 263315
rect 218378 263303 218384 263355
rect 255760 263303 255766 263355
rect 255818 263343 255824 263355
rect 329680 263343 329686 263355
rect 255818 263315 329686 263343
rect 255818 263303 255824 263315
rect 329680 263303 329686 263315
rect 329738 263303 329744 263355
rect 331216 263303 331222 263355
rect 331274 263343 331280 263355
rect 338128 263343 338134 263355
rect 331274 263315 338134 263343
rect 331274 263303 331280 263315
rect 338128 263303 338134 263315
rect 338186 263303 338192 263355
rect 340624 263303 340630 263355
rect 340682 263343 340688 263355
rect 346864 263343 346870 263355
rect 340682 263315 346870 263343
rect 340682 263303 340688 263315
rect 346864 263303 346870 263315
rect 346922 263303 346928 263355
rect 349072 263303 349078 263355
rect 349130 263343 349136 263355
rect 354832 263343 354838 263355
rect 349130 263315 354838 263343
rect 349130 263303 349136 263315
rect 354832 263303 354838 263315
rect 354890 263303 354896 263355
rect 355024 263303 355030 263355
rect 355082 263343 355088 263355
rect 365680 263343 365686 263355
rect 355082 263315 365686 263343
rect 355082 263303 355088 263315
rect 365680 263303 365686 263315
rect 365738 263303 365744 263355
rect 369712 263303 369718 263355
rect 369770 263343 369776 263355
rect 526192 263343 526198 263355
rect 369770 263315 526198 263343
rect 369770 263303 369776 263315
rect 526192 263303 526198 263315
rect 526250 263303 526256 263355
rect 252496 263229 252502 263281
rect 252554 263269 252560 263281
rect 258640 263269 258646 263281
rect 252554 263241 258646 263269
rect 252554 263229 252560 263241
rect 258640 263229 258646 263241
rect 258698 263229 258704 263281
rect 286576 263229 286582 263281
rect 286634 263269 286640 263281
rect 300112 263269 300118 263281
rect 286634 263241 300118 263269
rect 286634 263229 286640 263241
rect 300112 263229 300118 263241
rect 300170 263229 300176 263281
rect 327760 263229 327766 263281
rect 327818 263269 327824 263281
rect 335536 263269 335542 263281
rect 327818 263241 335542 263269
rect 327818 263229 327824 263241
rect 335536 263229 335542 263241
rect 335594 263229 335600 263281
rect 357808 263229 357814 263281
rect 357866 263269 357872 263281
rect 364624 263269 364630 263281
rect 357866 263241 364630 263269
rect 357866 263229 357872 263241
rect 364624 263229 364630 263241
rect 364682 263229 364688 263281
rect 369136 263229 369142 263281
rect 369194 263269 369200 263281
rect 518992 263269 518998 263281
rect 369194 263241 518998 263269
rect 369194 263229 369200 263241
rect 518992 263229 518998 263241
rect 519050 263229 519056 263281
rect 254416 263155 254422 263207
rect 254474 263195 254480 263207
rect 402832 263195 402838 263207
rect 254474 263167 402838 263195
rect 254474 263155 254480 263167
rect 402832 263155 402838 263167
rect 402890 263155 402896 263207
rect 406672 263155 406678 263207
rect 406730 263195 406736 263207
rect 414640 263195 414646 263207
rect 406730 263167 414646 263195
rect 406730 263155 406736 263167
rect 414640 263155 414646 263167
rect 414698 263155 414704 263207
rect 253840 263081 253846 263133
rect 253898 263121 253904 263133
rect 330064 263121 330070 263133
rect 253898 263093 330070 263121
rect 253898 263081 253904 263093
rect 330064 263081 330070 263093
rect 330122 263081 330128 263133
rect 330160 263081 330166 263133
rect 330218 263121 330224 263133
rect 332944 263121 332950 263133
rect 330218 263093 332950 263121
rect 330218 263081 330224 263093
rect 332944 263081 332950 263093
rect 333002 263081 333008 263133
rect 339664 263081 339670 263133
rect 339722 263121 339728 263133
rect 342064 263121 342070 263133
rect 339722 263093 342070 263121
rect 339722 263081 339728 263093
rect 342064 263081 342070 263093
rect 342122 263081 342128 263133
rect 349744 263081 349750 263133
rect 349802 263121 349808 263133
rect 362032 263121 362038 263133
rect 349802 263093 362038 263121
rect 349802 263081 349808 263093
rect 362032 263081 362038 263093
rect 362090 263081 362096 263133
rect 367408 263081 367414 263133
rect 367466 263121 367472 263133
rect 504688 263121 504694 263133
rect 367466 263093 504694 263121
rect 367466 263081 367472 263093
rect 504688 263081 504694 263093
rect 504746 263081 504752 263133
rect 223120 263007 223126 263059
rect 223178 263047 223184 263059
rect 234736 263047 234742 263059
rect 223178 263019 234742 263047
rect 223178 263007 223184 263019
rect 234736 263007 234742 263019
rect 234794 263007 234800 263059
rect 257488 263007 257494 263059
rect 257546 263047 257552 263059
rect 330736 263047 330742 263059
rect 257546 263019 330742 263047
rect 257546 263007 257552 263019
rect 330736 263007 330742 263019
rect 330794 263007 330800 263059
rect 331024 263007 331030 263059
rect 331082 263047 331088 263059
rect 334480 263047 334486 263059
rect 331082 263019 334486 263047
rect 331082 263007 331088 263019
rect 334480 263007 334486 263019
rect 334538 263007 334544 263059
rect 338704 263007 338710 263059
rect 338762 263047 338768 263059
rect 340336 263047 340342 263059
rect 338762 263019 340342 263047
rect 338762 263007 338768 263019
rect 340336 263007 340342 263019
rect 340394 263007 340400 263059
rect 354064 263007 354070 263059
rect 354122 263047 354128 263059
rect 362128 263047 362134 263059
rect 354122 263019 362134 263047
rect 354122 263007 354128 263019
rect 362128 263007 362134 263019
rect 362186 263007 362192 263059
rect 366544 263007 366550 263059
rect 366602 263047 366608 263059
rect 497296 263047 497302 263059
rect 366602 263019 497302 263047
rect 366602 263007 366608 263019
rect 497296 263007 497302 263019
rect 497354 263007 497360 263059
rect 261232 262933 261238 262985
rect 261290 262973 261296 262985
rect 326800 262973 326806 262985
rect 261290 262945 326806 262973
rect 261290 262933 261296 262945
rect 326800 262933 326806 262945
rect 326858 262933 326864 262985
rect 326992 262933 326998 262985
rect 327050 262973 327056 262985
rect 345328 262973 345334 262985
rect 327050 262945 345334 262973
rect 327050 262933 327056 262945
rect 345328 262933 345334 262945
rect 345386 262933 345392 262985
rect 351856 262933 351862 262985
rect 351914 262973 351920 262985
rect 355024 262973 355030 262985
rect 351914 262945 355030 262973
rect 351914 262933 351920 262945
rect 355024 262933 355030 262945
rect 355082 262933 355088 262985
rect 365392 262933 365398 262985
rect 365450 262973 365456 262985
rect 490480 262973 490486 262985
rect 365450 262945 490486 262973
rect 365450 262933 365456 262945
rect 490480 262933 490486 262945
rect 490538 262933 490544 262985
rect 248176 262859 248182 262911
rect 248234 262899 248240 262911
rect 274096 262899 274102 262911
rect 248234 262871 274102 262899
rect 248234 262859 248240 262871
rect 274096 262859 274102 262871
rect 274154 262859 274160 262911
rect 285520 262859 285526 262911
rect 285578 262899 285584 262911
rect 289456 262899 289462 262911
rect 285578 262871 289462 262899
rect 285578 262859 285584 262871
rect 289456 262859 289462 262871
rect 289514 262859 289520 262911
rect 290992 262859 290998 262911
rect 291050 262899 291056 262911
rect 341008 262899 341014 262911
rect 291050 262871 341014 262899
rect 291050 262859 291056 262871
rect 341008 262859 341014 262871
rect 341066 262859 341072 262911
rect 352336 262859 352342 262911
rect 352394 262899 352400 262911
rect 362800 262899 362806 262911
rect 352394 262871 362806 262899
rect 352394 262859 352400 262871
rect 362800 262859 362806 262871
rect 362858 262859 362864 262911
rect 364816 262859 364822 262911
rect 364874 262899 364880 262911
rect 483280 262899 483286 262911
rect 364874 262871 483286 262899
rect 364874 262859 364880 262871
rect 483280 262859 483286 262871
rect 483338 262859 483344 262911
rect 248656 262785 248662 262837
rect 248714 262825 248720 262837
rect 272848 262825 272854 262837
rect 248714 262797 272854 262825
rect 248714 262785 248720 262797
rect 272848 262785 272854 262797
rect 272906 262785 272912 262837
rect 294160 262785 294166 262837
rect 294218 262825 294224 262837
rect 339280 262825 339286 262837
rect 294218 262797 339286 262825
rect 294218 262785 294224 262797
rect 339280 262785 339286 262797
rect 339338 262785 339344 262837
rect 339376 262785 339382 262837
rect 339434 262825 339440 262837
rect 341488 262825 341494 262837
rect 339434 262797 341494 262825
rect 339434 262785 339440 262797
rect 341488 262785 341494 262797
rect 341546 262785 341552 262837
rect 341584 262785 341590 262837
rect 341642 262825 341648 262837
rect 344272 262825 344278 262837
rect 341642 262797 344278 262825
rect 341642 262785 341648 262797
rect 344272 262785 344278 262797
rect 344330 262785 344336 262837
rect 363664 262785 363670 262837
rect 363722 262825 363728 262837
rect 476176 262825 476182 262837
rect 363722 262797 476182 262825
rect 363722 262785 363728 262797
rect 476176 262785 476182 262797
rect 476234 262785 476240 262837
rect 257680 262711 257686 262763
rect 257738 262751 257744 262763
rect 281296 262751 281302 262763
rect 257738 262723 281302 262751
rect 257738 262711 257744 262723
rect 281296 262711 281302 262723
rect 281354 262711 281360 262763
rect 282352 262711 282358 262763
rect 282410 262751 282416 262763
rect 284368 262751 284374 262763
rect 282410 262723 284374 262751
rect 282410 262711 282416 262723
rect 284368 262711 284374 262723
rect 284426 262711 284432 262763
rect 297808 262711 297814 262763
rect 297866 262751 297872 262763
rect 341872 262751 341878 262763
rect 297866 262723 341878 262751
rect 297866 262711 297872 262723
rect 341872 262711 341878 262723
rect 341930 262711 341936 262763
rect 341968 262711 341974 262763
rect 342026 262751 342032 262763
rect 344080 262751 344086 262763
rect 342026 262723 344086 262751
rect 342026 262711 342032 262723
rect 344080 262711 344086 262723
rect 344138 262711 344144 262763
rect 362704 262711 362710 262763
rect 362762 262751 362768 262763
rect 468976 262751 468982 262763
rect 362762 262723 468982 262751
rect 362762 262711 362768 262723
rect 468976 262711 468982 262723
rect 469034 262711 469040 262763
rect 42256 262637 42262 262689
rect 42314 262677 42320 262689
rect 47824 262677 47830 262689
rect 42314 262649 47830 262677
rect 42314 262637 42320 262649
rect 47824 262637 47830 262649
rect 47882 262637 47888 262689
rect 260944 262637 260950 262689
rect 261002 262677 261008 262689
rect 261002 262649 268286 262677
rect 261002 262637 261008 262649
rect 268258 262455 268286 262649
rect 275152 262637 275158 262689
rect 275210 262677 275216 262689
rect 283504 262677 283510 262689
rect 275210 262649 283510 262677
rect 275210 262637 275216 262649
rect 283504 262637 283510 262649
rect 283562 262637 283568 262689
rect 287248 262637 287254 262689
rect 287306 262677 287312 262689
rect 303664 262677 303670 262689
rect 287306 262649 303670 262677
rect 287306 262637 287312 262649
rect 303664 262637 303670 262649
rect 303722 262637 303728 262689
rect 304912 262637 304918 262689
rect 304970 262677 304976 262689
rect 342736 262677 342742 262689
rect 304970 262649 342742 262677
rect 304970 262637 304976 262649
rect 342736 262637 342742 262649
rect 342794 262637 342800 262689
rect 362128 262637 362134 262689
rect 362186 262677 362192 262689
rect 461968 262677 461974 262689
rect 362186 262649 461974 262677
rect 362186 262637 362192 262649
rect 461968 262637 461974 262649
rect 462026 262637 462032 262689
rect 268336 262563 268342 262615
rect 268394 262603 268400 262615
rect 282352 262603 282358 262615
rect 268394 262575 282358 262603
rect 268394 262563 268400 262575
rect 282352 262563 282358 262575
rect 282410 262563 282416 262615
rect 285040 262563 285046 262615
rect 285098 262603 285104 262615
rect 285808 262603 285814 262615
rect 285098 262575 285814 262603
rect 285098 262563 285104 262575
rect 285808 262563 285814 262575
rect 285866 262563 285872 262615
rect 299536 262563 299542 262615
rect 299594 262603 299600 262615
rect 337744 262603 337750 262615
rect 299594 262575 337750 262603
rect 299594 262563 299600 262575
rect 337744 262563 337750 262575
rect 337802 262563 337808 262615
rect 361072 262563 361078 262615
rect 361130 262603 361136 262615
rect 454768 262603 454774 262615
rect 361130 262575 454774 262603
rect 361130 262563 361136 262575
rect 454768 262563 454774 262575
rect 454826 262563 454832 262615
rect 287824 262489 287830 262541
rect 287882 262529 287888 262541
rect 310864 262529 310870 262541
rect 287882 262501 310870 262529
rect 287882 262489 287888 262501
rect 310864 262489 310870 262501
rect 310922 262489 310928 262541
rect 312400 262489 312406 262541
rect 312458 262529 312464 262541
rect 343600 262529 343606 262541
rect 312458 262501 343606 262529
rect 312458 262489 312464 262501
rect 343600 262489 343606 262501
rect 343658 262489 343664 262541
rect 367984 262489 367990 262541
rect 368042 262529 368048 262541
rect 455056 262529 455062 262541
rect 368042 262501 455062 262529
rect 368042 262489 368048 262501
rect 455056 262489 455062 262501
rect 455114 262489 455120 262541
rect 281776 262455 281782 262467
rect 268258 262427 281782 262455
rect 281776 262415 281782 262427
rect 281834 262415 281840 262467
rect 313936 262415 313942 262467
rect 313994 262455 314000 262467
rect 331216 262455 331222 262467
rect 313994 262427 331222 262455
rect 313994 262415 314000 262427
rect 331216 262415 331222 262427
rect 331274 262415 331280 262467
rect 360400 262415 360406 262467
rect 360458 262455 360464 262467
rect 447664 262455 447670 262467
rect 360458 262427 447670 262455
rect 360458 262415 360464 262427
rect 447664 262415 447670 262427
rect 447722 262415 447728 262467
rect 317008 262341 317014 262393
rect 317066 262381 317072 262393
rect 325456 262381 325462 262393
rect 317066 262353 325462 262381
rect 317066 262341 317072 262353
rect 325456 262341 325462 262353
rect 325514 262341 325520 262393
rect 327088 262341 327094 262393
rect 327146 262381 327152 262393
rect 399184 262381 399190 262393
rect 327146 262353 399190 262381
rect 327146 262341 327152 262353
rect 399184 262341 399190 262353
rect 399242 262341 399248 262393
rect 400144 262341 400150 262393
rect 400202 262381 400208 262393
rect 409840 262381 409846 262393
rect 400202 262353 409846 262381
rect 400202 262341 400208 262353
rect 409840 262341 409846 262353
rect 409898 262341 409904 262393
rect 351760 262267 351766 262319
rect 351818 262307 351824 262319
rect 375952 262307 375958 262319
rect 351818 262279 375958 262307
rect 351818 262267 351824 262279
rect 375952 262267 375958 262279
rect 376010 262267 376016 262319
rect 376048 262267 376054 262319
rect 376106 262307 376112 262319
rect 384976 262307 384982 262319
rect 376106 262279 384982 262307
rect 376106 262267 376112 262279
rect 384976 262267 384982 262279
rect 385034 262267 385040 262319
rect 385648 262267 385654 262319
rect 385706 262307 385712 262319
rect 388240 262307 388246 262319
rect 385706 262279 388246 262307
rect 385706 262267 385712 262279
rect 388240 262267 388246 262279
rect 388298 262267 388304 262319
rect 388624 262267 388630 262319
rect 388682 262307 388688 262319
rect 390928 262307 390934 262319
rect 388682 262279 390934 262307
rect 388682 262267 388688 262279
rect 390928 262267 390934 262279
rect 390986 262267 390992 262319
rect 391408 262267 391414 262319
rect 391466 262307 391472 262319
rect 396976 262307 396982 262319
rect 391466 262279 396982 262307
rect 391466 262267 391472 262279
rect 396976 262267 396982 262279
rect 397034 262267 397040 262319
rect 397072 262267 397078 262319
rect 397130 262307 397136 262319
rect 401776 262307 401782 262319
rect 397130 262279 401782 262307
rect 397130 262267 397136 262279
rect 401776 262267 401782 262279
rect 401834 262267 401840 262319
rect 402160 262267 402166 262319
rect 402218 262307 402224 262319
rect 413104 262307 413110 262319
rect 402218 262279 413110 262307
rect 402218 262267 402224 262279
rect 413104 262267 413110 262279
rect 413162 262267 413168 262319
rect 336016 262233 336022 262245
rect 331042 262205 336022 262233
rect 144688 262119 144694 262171
rect 144746 262159 144752 262171
rect 146608 262159 146614 262171
rect 144746 262131 146614 262159
rect 144746 262119 144752 262131
rect 146608 262119 146614 262131
rect 146666 262119 146672 262171
rect 221584 262119 221590 262171
rect 221642 262159 221648 262171
rect 223984 262159 223990 262171
rect 221642 262131 223990 262159
rect 221642 262119 221648 262131
rect 223984 262119 223990 262131
rect 224042 262119 224048 262171
rect 247984 262119 247990 262171
rect 248042 262159 248048 262171
rect 250384 262159 250390 262171
rect 248042 262131 250390 262159
rect 248042 262119 248048 262131
rect 250384 262119 250390 262131
rect 250442 262119 250448 262171
rect 256240 262119 256246 262171
rect 256298 262159 256304 262171
rect 330544 262159 330550 262171
rect 256298 262131 330550 262159
rect 256298 262119 256304 262131
rect 330544 262119 330550 262131
rect 330602 262119 330608 262171
rect 251344 262045 251350 262097
rect 251402 262085 251408 262097
rect 331042 262085 331070 262205
rect 336016 262193 336022 262205
rect 336074 262193 336080 262245
rect 359344 262193 359350 262245
rect 359402 262233 359408 262245
rect 359402 262205 365822 262233
rect 359402 262193 359408 262205
rect 335344 262159 335350 262171
rect 251402 262057 331070 262085
rect 331138 262131 335350 262159
rect 251402 262045 251408 262057
rect 244240 261971 244246 262023
rect 244298 262011 244304 262023
rect 331138 262011 331166 262131
rect 335344 262119 335350 262131
rect 335402 262119 335408 262171
rect 352816 262119 352822 262171
rect 352874 262159 352880 262171
rect 362800 262159 362806 262171
rect 352874 262131 356990 262159
rect 352874 262119 352880 262131
rect 244298 261983 331166 262011
rect 356962 262011 356990 262131
rect 357250 262131 362806 262159
rect 357040 262045 357046 262097
rect 357098 262085 357104 262097
rect 357250 262085 357278 262131
rect 362800 262119 362806 262131
rect 362858 262119 362864 262171
rect 357098 262057 357278 262085
rect 365794 262085 365822 262205
rect 384400 262193 384406 262245
rect 384458 262233 384464 262245
rect 385840 262233 385846 262245
rect 384458 262205 385846 262233
rect 384458 262193 384464 262205
rect 385840 262193 385846 262205
rect 385898 262193 385904 262245
rect 386128 262193 386134 262245
rect 386186 262233 386192 262245
rect 390448 262233 390454 262245
rect 386186 262205 390454 262233
rect 386186 262193 386192 262205
rect 390448 262193 390454 262205
rect 390506 262193 390512 262245
rect 390640 262193 390646 262245
rect 390698 262233 390704 262245
rect 396304 262233 396310 262245
rect 390698 262205 396310 262233
rect 390698 262193 390704 262205
rect 396304 262193 396310 262205
rect 396362 262193 396368 262245
rect 400144 262233 400150 262245
rect 396418 262205 400150 262233
rect 382960 262119 382966 262171
rect 383018 262159 383024 262171
rect 388048 262159 388054 262171
rect 383018 262131 388054 262159
rect 383018 262119 383024 262131
rect 388048 262119 388054 262131
rect 388106 262119 388112 262171
rect 389008 262119 389014 262171
rect 389066 262159 389072 262171
rect 394192 262159 394198 262171
rect 389066 262131 394198 262159
rect 389066 262119 389072 262131
rect 394192 262119 394198 262131
rect 394250 262119 394256 262171
rect 394288 262119 394294 262171
rect 394346 262159 394352 262171
rect 396418 262159 396446 262205
rect 400144 262193 400150 262205
rect 400202 262193 400208 262245
rect 400336 262193 400342 262245
rect 400394 262233 400400 262245
rect 411568 262233 411574 262245
rect 400394 262205 411574 262233
rect 400394 262193 400400 262205
rect 411568 262193 411574 262205
rect 411626 262193 411632 262245
rect 394346 262131 396446 262159
rect 394346 262119 394352 262131
rect 396496 262119 396502 262171
rect 396554 262159 396560 262171
rect 403792 262159 403798 262171
rect 396554 262131 403798 262159
rect 396554 262119 396560 262131
rect 403792 262119 403798 262131
rect 403850 262119 403856 262171
rect 403888 262119 403894 262171
rect 403946 262159 403952 262171
rect 408304 262159 408310 262171
rect 403946 262131 408310 262159
rect 403946 262119 403952 262131
rect 408304 262119 408310 262131
rect 408362 262119 408368 262171
rect 440464 262085 440470 262097
rect 365794 262057 440470 262085
rect 357098 262045 357104 262057
rect 440464 262045 440470 262057
rect 440522 262045 440528 262097
rect 382576 262011 382582 262023
rect 356962 261983 382582 262011
rect 244298 261971 244304 261983
rect 382576 261971 382582 261983
rect 382634 261971 382640 262023
rect 382672 261971 382678 262023
rect 382730 262011 382736 262023
rect 394672 262011 394678 262023
rect 382730 261983 394678 262011
rect 382730 261971 382736 261983
rect 394672 261971 394678 261983
rect 394730 261971 394736 262023
rect 262096 261897 262102 261949
rect 262154 261937 262160 261949
rect 263344 261937 263350 261949
rect 262154 261909 263350 261937
rect 262154 261897 262160 261909
rect 263344 261897 263350 261909
rect 263402 261897 263408 261949
rect 324016 261897 324022 261949
rect 324074 261937 324080 261949
rect 346960 261937 346966 261949
rect 324074 261909 346966 261937
rect 324074 261897 324080 261909
rect 346960 261897 346966 261909
rect 347018 261897 347024 261949
rect 362800 261897 362806 261949
rect 362858 261937 362864 261949
rect 419056 261937 419062 261949
rect 362858 261909 419062 261937
rect 362858 261897 362864 261909
rect 419056 261897 419062 261909
rect 419114 261897 419120 261949
rect 243664 261823 243670 261875
rect 243722 261863 243728 261875
rect 402448 261863 402454 261875
rect 243722 261835 402454 261863
rect 243722 261823 243728 261835
rect 402448 261823 402454 261835
rect 402506 261823 402512 261875
rect 244240 261749 244246 261801
rect 244298 261789 244304 261801
rect 409552 261789 409558 261801
rect 244298 261761 409558 261789
rect 244298 261749 244304 261761
rect 409552 261749 409558 261761
rect 409610 261749 409616 261801
rect 245392 261675 245398 261727
rect 245450 261715 245456 261727
rect 416656 261715 416662 261727
rect 245450 261687 416662 261715
rect 245450 261675 245456 261687
rect 416656 261675 416662 261687
rect 416714 261675 416720 261727
rect 245968 261601 245974 261653
rect 246026 261641 246032 261653
rect 423856 261641 423862 261653
rect 246026 261613 423862 261641
rect 246026 261601 246032 261613
rect 423856 261601 423862 261613
rect 423914 261601 423920 261653
rect 246928 261527 246934 261579
rect 246986 261567 246992 261579
rect 431056 261567 431062 261579
rect 246986 261539 431062 261567
rect 246986 261527 246992 261539
rect 431056 261527 431062 261539
rect 431114 261527 431120 261579
rect 521296 261527 521302 261579
rect 521354 261567 521360 261579
rect 548560 261567 548566 261579
rect 521354 261539 548566 261567
rect 521354 261527 521360 261539
rect 548560 261527 548566 261539
rect 548618 261527 548624 261579
rect 239920 261453 239926 261505
rect 239978 261493 239984 261505
rect 373552 261493 373558 261505
rect 239978 261465 373558 261493
rect 239978 261453 239984 261465
rect 373552 261453 373558 261465
rect 373610 261453 373616 261505
rect 374608 261453 374614 261505
rect 374666 261493 374672 261505
rect 565456 261493 565462 261505
rect 374666 261465 565462 261493
rect 374666 261453 374672 261465
rect 565456 261453 565462 261465
rect 565514 261453 565520 261505
rect 320752 261379 320758 261431
rect 320810 261419 320816 261431
rect 578512 261419 578518 261431
rect 320810 261391 578518 261419
rect 320810 261379 320816 261391
rect 578512 261379 578518 261391
rect 578570 261379 578576 261431
rect 229648 261305 229654 261357
rect 229706 261345 229712 261357
rect 288208 261345 288214 261357
rect 229706 261317 288214 261345
rect 229706 261305 229712 261317
rect 288208 261305 288214 261317
rect 288266 261305 288272 261357
rect 321424 261305 321430 261357
rect 321482 261345 321488 261357
rect 585616 261345 585622 261357
rect 321482 261317 585622 261345
rect 321482 261305 321488 261317
rect 585616 261305 585622 261317
rect 585674 261305 585680 261357
rect 230320 261231 230326 261283
rect 230378 261271 230384 261283
rect 295408 261271 295414 261283
rect 230378 261243 295414 261271
rect 230378 261231 230384 261243
rect 295408 261231 295414 261243
rect 295466 261231 295472 261283
rect 302512 261271 302518 261283
rect 295522 261243 302518 261271
rect 231184 261157 231190 261209
rect 231242 261197 231248 261209
rect 295522 261197 295550 261243
rect 302512 261231 302518 261243
rect 302570 261231 302576 261283
rect 308176 261231 308182 261283
rect 308234 261271 308240 261283
rect 318352 261271 318358 261283
rect 308234 261243 318358 261271
rect 308234 261231 308240 261243
rect 318352 261231 318358 261243
rect 318410 261231 318416 261283
rect 322480 261231 322486 261283
rect 322538 261271 322544 261283
rect 592720 261271 592726 261283
rect 322538 261243 592726 261271
rect 322538 261231 322544 261243
rect 592720 261231 592726 261243
rect 592778 261231 592784 261283
rect 231242 261169 295550 261197
rect 231242 261157 231248 261169
rect 298000 261157 298006 261209
rect 298058 261197 298064 261209
rect 316720 261197 316726 261209
rect 298058 261169 316726 261197
rect 298058 261157 298064 261169
rect 316720 261157 316726 261169
rect 316778 261157 316784 261209
rect 323152 261157 323158 261209
rect 323210 261197 323216 261209
rect 599824 261197 599830 261209
rect 323210 261169 599830 261197
rect 323210 261157 323216 261169
rect 599824 261157 599830 261169
rect 599882 261157 599888 261209
rect 232336 261083 232342 261135
rect 232394 261123 232400 261135
rect 309712 261123 309718 261135
rect 232394 261095 309718 261123
rect 232394 261083 232400 261095
rect 309712 261083 309718 261095
rect 309770 261083 309776 261135
rect 318064 261083 318070 261135
rect 318122 261123 318128 261135
rect 338224 261123 338230 261135
rect 318122 261095 338230 261123
rect 318122 261083 318128 261095
rect 338224 261083 338230 261095
rect 338282 261083 338288 261135
rect 346960 261083 346966 261135
rect 347018 261123 347024 261135
rect 607024 261123 607030 261135
rect 347018 261095 607030 261123
rect 347018 261083 347024 261095
rect 607024 261083 607030 261095
rect 607082 261083 607088 261135
rect 225808 261009 225814 261061
rect 225866 261049 225872 261061
rect 255856 261049 255862 261061
rect 225866 261021 255862 261049
rect 225866 261009 225872 261021
rect 255856 261009 255862 261021
rect 255914 261009 255920 261061
rect 260656 261009 260662 261061
rect 260714 261049 260720 261061
rect 541648 261049 541654 261061
rect 260714 261021 541654 261049
rect 260714 261009 260720 261021
rect 541648 261009 541654 261021
rect 541706 261009 541712 261061
rect 225904 260935 225910 260987
rect 225962 260975 225968 260987
rect 259696 260975 259702 260987
rect 225962 260947 259702 260975
rect 225962 260935 225968 260947
rect 259696 260935 259702 260947
rect 259754 260935 259760 260987
rect 261712 260935 261718 260987
rect 261770 260975 261776 260987
rect 552304 260975 552310 260987
rect 261770 260947 552310 260975
rect 261770 260935 261776 260947
rect 552304 260935 552310 260947
rect 552362 260935 552368 260987
rect 232912 260861 232918 260913
rect 232970 260901 232976 260913
rect 298000 260901 298006 260913
rect 232970 260873 298006 260901
rect 232970 260861 232976 260873
rect 298000 260861 298006 260873
rect 298058 260861 298064 260913
rect 305680 260861 305686 260913
rect 305738 260901 305744 260913
rect 318256 260901 318262 260913
rect 305738 260873 318262 260901
rect 305738 260861 305744 260873
rect 318256 260861 318262 260873
rect 318314 260861 318320 260913
rect 325168 260861 325174 260913
rect 325226 260901 325232 260913
rect 614224 260901 614230 260913
rect 325226 260873 614230 260901
rect 325226 260861 325232 260873
rect 614224 260861 614230 260873
rect 614282 260861 614288 260913
rect 234064 260787 234070 260839
rect 234122 260827 234128 260839
rect 323920 260827 323926 260839
rect 234122 260799 323926 260827
rect 234122 260787 234128 260799
rect 323920 260787 323926 260799
rect 323978 260787 323984 260839
rect 325744 260787 325750 260839
rect 325802 260827 325808 260839
rect 620944 260827 620950 260839
rect 325802 260799 620950 260827
rect 325802 260787 325808 260799
rect 620944 260787 620950 260799
rect 621002 260787 621008 260839
rect 226384 260713 226390 260765
rect 226442 260753 226448 260765
rect 262096 260753 262102 260765
rect 226442 260725 262102 260753
rect 226442 260713 226448 260725
rect 262096 260713 262102 260725
rect 262154 260713 262160 260765
rect 262192 260713 262198 260765
rect 262250 260753 262256 260765
rect 555856 260753 555862 260765
rect 262250 260725 555862 260753
rect 262250 260713 262256 260725
rect 555856 260713 555862 260725
rect 555914 260713 555920 260765
rect 234928 260639 234934 260691
rect 234986 260679 234992 260691
rect 318160 260679 318166 260691
rect 234986 260651 318166 260679
rect 234986 260639 234992 260651
rect 318160 260639 318166 260651
rect 318218 260639 318224 260691
rect 318352 260639 318358 260691
rect 318410 260679 318416 260691
rect 328240 260679 328246 260691
rect 318410 260651 328246 260679
rect 318410 260639 318416 260651
rect 328240 260639 328246 260651
rect 328298 260639 328304 260691
rect 328336 260639 328342 260691
rect 328394 260679 328400 260691
rect 642736 260679 642742 260691
rect 328394 260651 642742 260679
rect 328394 260639 328400 260651
rect 642736 260639 642742 260651
rect 642794 260639 642800 260691
rect 240976 260565 240982 260617
rect 241034 260605 241040 260617
rect 381040 260605 381046 260617
rect 241034 260577 381046 260605
rect 241034 260565 241040 260577
rect 381040 260565 381046 260577
rect 381098 260565 381104 260617
rect 381520 260565 381526 260617
rect 381578 260605 381584 260617
rect 521776 260605 521782 260617
rect 381578 260577 521782 260605
rect 381578 260565 381584 260577
rect 521776 260565 521782 260577
rect 521834 260565 521840 260617
rect 239344 260491 239350 260543
rect 239402 260531 239408 260543
rect 366736 260531 366742 260543
rect 239402 260503 366742 260531
rect 239402 260491 239408 260503
rect 366736 260491 366742 260503
rect 366794 260491 366800 260543
rect 378928 260491 378934 260543
rect 378986 260531 378992 260543
rect 508240 260531 508246 260543
rect 378986 260503 508246 260531
rect 378986 260491 378992 260503
rect 508240 260491 508246 260503
rect 508298 260491 508304 260543
rect 228592 260417 228598 260469
rect 228650 260457 228656 260469
rect 280816 260457 280822 260469
rect 228650 260429 280822 260457
rect 228650 260417 228656 260429
rect 280816 260417 280822 260429
rect 280874 260417 280880 260469
rect 301840 260417 301846 260469
rect 301898 260457 301904 260469
rect 425008 260457 425014 260469
rect 301898 260429 425014 260457
rect 301898 260417 301904 260429
rect 425008 260417 425014 260429
rect 425066 260417 425072 260469
rect 238192 260343 238198 260395
rect 238250 260383 238256 260395
rect 359632 260383 359638 260395
rect 238250 260355 359638 260383
rect 238250 260343 238256 260355
rect 359632 260343 359638 260355
rect 359690 260343 359696 260395
rect 373936 260343 373942 260395
rect 373994 260383 374000 260395
rect 478768 260383 478774 260395
rect 373994 260355 478774 260383
rect 373994 260343 374000 260355
rect 478768 260343 478774 260355
rect 478826 260343 478832 260395
rect 226864 260269 226870 260321
rect 226922 260309 226928 260321
rect 266800 260309 266806 260321
rect 226922 260281 266806 260309
rect 226922 260269 226928 260281
rect 266800 260269 266806 260281
rect 266858 260269 266864 260321
rect 301168 260269 301174 260321
rect 301226 260309 301232 260321
rect 417904 260309 417910 260321
rect 301226 260281 417910 260309
rect 301226 260269 301232 260281
rect 417904 260269 417910 260281
rect 417962 260269 417968 260321
rect 237328 260195 237334 260247
rect 237386 260235 237392 260247
rect 352432 260235 352438 260247
rect 237386 260207 352438 260235
rect 237386 260195 237392 260207
rect 352432 260195 352438 260207
rect 352490 260195 352496 260247
rect 376144 260195 376150 260247
rect 376202 260235 376208 260247
rect 446224 260235 446230 260247
rect 376202 260207 446230 260235
rect 376202 260195 376208 260207
rect 446224 260195 446230 260207
rect 446282 260195 446288 260247
rect 236656 260121 236662 260173
rect 236714 260161 236720 260173
rect 345040 260161 345046 260173
rect 236714 260133 345046 260161
rect 236714 260121 236720 260133
rect 345040 260121 345046 260133
rect 345098 260121 345104 260173
rect 376720 260121 376726 260173
rect 376778 260161 376784 260173
rect 409072 260161 409078 260173
rect 376778 260133 409078 260161
rect 376778 260121 376784 260133
rect 409072 260121 409078 260133
rect 409130 260121 409136 260173
rect 299632 260047 299638 260099
rect 299690 260087 299696 260099
rect 407152 260087 407158 260099
rect 299690 260059 407158 260087
rect 299690 260047 299696 260059
rect 407152 260047 407158 260059
rect 407210 260047 407216 260099
rect 235600 259973 235606 260025
rect 235658 260013 235664 260025
rect 318064 260013 318070 260025
rect 235658 259985 318070 260013
rect 235658 259973 235664 259985
rect 318064 259973 318070 259985
rect 318122 259973 318128 260025
rect 318160 259973 318166 260025
rect 318218 260013 318224 260025
rect 331120 260013 331126 260025
rect 318218 259985 331126 260013
rect 318218 259973 318224 259985
rect 331120 259973 331126 259985
rect 331178 259973 331184 260025
rect 378256 259973 378262 260025
rect 378314 260013 378320 260025
rect 409168 260013 409174 260025
rect 378314 259985 409174 260013
rect 378314 259973 378320 259985
rect 409168 259973 409174 259985
rect 409226 259973 409232 260025
rect 233488 259899 233494 259951
rect 233546 259939 233552 259951
rect 233546 259911 288062 259939
rect 233546 259899 233552 259911
rect 72016 259529 72022 259581
rect 72074 259569 72080 259581
rect 77680 259569 77686 259581
rect 72074 259541 77686 259569
rect 72074 259529 72080 259541
rect 77680 259529 77686 259541
rect 77738 259529 77744 259581
rect 288034 259421 288062 259911
rect 298960 259899 298966 259951
rect 299018 259939 299024 259951
rect 400048 259939 400054 259951
rect 299018 259911 400054 259939
rect 299018 259899 299024 259911
rect 400048 259899 400054 259911
rect 400106 259899 400112 259951
rect 308080 259825 308086 259877
rect 308138 259865 308144 259877
rect 308176 259865 308182 259877
rect 308138 259837 308182 259865
rect 308138 259825 308144 259837
rect 308176 259825 308182 259837
rect 308234 259825 308240 259877
rect 328240 259825 328246 259877
rect 328298 259865 328304 259877
rect 334000 259865 334006 259877
rect 328298 259837 334006 259865
rect 328298 259825 328304 259837
rect 334000 259825 334006 259837
rect 334058 259825 334064 259877
rect 379984 259825 379990 259877
rect 380042 259865 380048 259877
rect 405808 259865 405814 259877
rect 380042 259837 405814 259865
rect 380042 259825 380048 259837
rect 405808 259825 405814 259837
rect 405866 259825 405872 259877
rect 298096 259751 298102 259803
rect 298154 259791 298160 259803
rect 392944 259791 392950 259803
rect 298154 259763 392950 259791
rect 298154 259751 298160 259763
rect 392944 259751 392950 259763
rect 393002 259751 393008 259803
rect 394672 259751 394678 259803
rect 394730 259791 394736 259803
rect 395056 259791 395062 259803
rect 394730 259763 395062 259791
rect 394730 259751 394736 259763
rect 395056 259751 395062 259763
rect 395114 259751 395120 259803
rect 296944 259677 296950 259729
rect 297002 259717 297008 259729
rect 385552 259717 385558 259729
rect 297002 259689 385558 259717
rect 297002 259677 297008 259689
rect 385552 259677 385558 259689
rect 385610 259677 385616 259729
rect 296368 259603 296374 259655
rect 296426 259643 296432 259655
rect 378640 259643 378646 259655
rect 296426 259615 378646 259643
rect 296426 259603 296432 259615
rect 378640 259603 378646 259615
rect 378698 259603 378704 259655
rect 295312 259529 295318 259581
rect 295370 259569 295376 259581
rect 371536 259569 371542 259581
rect 295370 259541 371542 259569
rect 295370 259529 295376 259541
rect 371536 259529 371542 259541
rect 371594 259529 371600 259581
rect 294352 259455 294358 259507
rect 294410 259495 294416 259507
rect 364432 259495 364438 259507
rect 294410 259467 364438 259495
rect 294410 259455 294416 259467
rect 364432 259455 364438 259467
rect 364490 259455 364496 259507
rect 308080 259421 308086 259433
rect 288034 259393 308086 259421
rect 308080 259381 308086 259393
rect 308138 259381 308144 259433
rect 318256 259381 318262 259433
rect 318314 259421 318320 259433
rect 457168 259421 457174 259433
rect 318314 259393 457174 259421
rect 318314 259381 318320 259393
rect 457168 259381 457174 259393
rect 457226 259381 457232 259433
rect 242512 259307 242518 259359
rect 242570 259347 242576 259359
rect 395152 259347 395158 259359
rect 242570 259319 395158 259347
rect 242570 259307 242576 259319
rect 395152 259307 395158 259319
rect 395210 259307 395216 259359
rect 241648 259233 241654 259285
rect 241706 259273 241712 259285
rect 388144 259273 388150 259285
rect 241706 259245 388150 259273
rect 241706 259233 241712 259245
rect 388144 259233 388150 259245
rect 388202 259233 388208 259285
rect 146512 259159 146518 259211
rect 146570 259199 146576 259211
rect 146608 259199 146614 259211
rect 146570 259171 146614 259199
rect 146570 259159 146576 259171
rect 146608 259159 146614 259171
rect 146666 259159 146672 259211
rect 639280 256347 639286 256399
rect 639338 256387 639344 256399
rect 679792 256387 679798 256399
rect 639338 256359 679798 256387
rect 639338 256347 639344 256359
rect 679792 256347 679798 256359
rect 679850 256347 679856 256399
rect 675088 253461 675094 253513
rect 675146 253501 675152 253513
rect 678256 253501 678262 253513
rect 675146 253473 678262 253501
rect 675146 253461 675152 253473
rect 678256 253461 678262 253473
rect 678314 253461 678320 253513
rect 72112 253387 72118 253439
rect 72170 253427 72176 253439
rect 77008 253427 77014 253439
rect 72170 253399 77014 253427
rect 72170 253387 72176 253399
rect 77008 253387 77014 253399
rect 77066 253387 77072 253439
rect 674800 251611 674806 251663
rect 674858 251651 674864 251663
rect 676912 251651 676918 251663
rect 674858 251623 676918 251651
rect 674858 251611 674864 251623
rect 676912 251611 676918 251623
rect 676970 251611 676976 251663
rect 674992 251537 674998 251589
rect 675050 251577 675056 251589
rect 676816 251577 676822 251589
rect 675050 251549 676822 251577
rect 675050 251537 675056 251549
rect 676816 251537 676822 251549
rect 676874 251537 676880 251589
rect 673936 250945 673942 250997
rect 673994 250985 674000 250997
rect 675376 250985 675382 250997
rect 673994 250957 675382 250985
rect 673994 250945 674000 250957
rect 675376 250945 675382 250957
rect 675434 250945 675440 250997
rect 198736 250575 198742 250627
rect 198794 250615 198800 250627
rect 198794 250587 201662 250615
rect 198794 250575 198800 250587
rect 201634 250541 201662 250587
rect 207280 250541 207286 250553
rect 201634 250513 207286 250541
rect 207280 250501 207286 250513
rect 207338 250501 207344 250553
rect 674608 250353 674614 250405
rect 674666 250393 674672 250405
rect 675472 250393 675478 250405
rect 674666 250365 675478 250393
rect 674666 250353 674672 250365
rect 675472 250353 675478 250365
rect 675530 250353 675536 250405
rect 674320 247023 674326 247075
rect 674378 247063 674384 247075
rect 675472 247063 675478 247075
rect 674378 247035 675478 247063
rect 674378 247023 674384 247035
rect 675472 247023 675478 247035
rect 675530 247023 675536 247075
rect 139504 246949 139510 247001
rect 139562 246989 139568 247001
rect 141424 246989 141430 247001
rect 139562 246961 141430 246989
rect 139562 246949 139568 246961
rect 141424 246949 141430 246961
rect 141482 246949 141488 247001
rect 674416 246949 674422 247001
rect 674474 246989 674480 247001
rect 675280 246989 675286 247001
rect 674474 246961 675286 246989
rect 674474 246949 674480 246961
rect 675280 246949 675286 246961
rect 675338 246949 675344 247001
rect 257008 246801 257014 246853
rect 257066 246841 257072 246853
rect 327952 246841 327958 246853
rect 257066 246813 327958 246841
rect 257066 246801 257072 246813
rect 327952 246801 327958 246813
rect 328010 246801 328016 246853
rect 262000 246727 262006 246779
rect 262058 246767 262064 246779
rect 331840 246767 331846 246779
rect 262058 246739 331846 246767
rect 262058 246727 262064 246739
rect 331840 246727 331846 246739
rect 331898 246727 331904 246779
rect 252880 246653 252886 246705
rect 252938 246693 252944 246705
rect 328768 246693 328774 246705
rect 252938 246665 328774 246693
rect 252938 246653 252944 246665
rect 328768 246653 328774 246665
rect 328826 246653 328832 246705
rect 258256 246579 258262 246631
rect 258314 246619 258320 246631
rect 332752 246619 332758 246631
rect 258314 246591 332758 246619
rect 258314 246579 258320 246591
rect 332752 246579 332758 246591
rect 332810 246579 332816 246631
rect 65104 246505 65110 246557
rect 65162 246545 65168 246557
rect 204976 246545 204982 246557
rect 65162 246517 204982 246545
rect 65162 246505 65168 246517
rect 204976 246505 204982 246517
rect 205034 246505 205040 246557
rect 257584 246505 257590 246557
rect 257642 246545 257648 246557
rect 334480 246545 334486 246557
rect 257642 246517 334486 246545
rect 257642 246505 257648 246517
rect 334480 246505 334486 246517
rect 334538 246505 334544 246557
rect 47920 246431 47926 246483
rect 47978 246471 47984 246483
rect 204880 246471 204886 246483
rect 47978 246443 204886 246471
rect 47978 246431 47984 246443
rect 204880 246431 204886 246443
rect 204938 246431 204944 246483
rect 256432 246431 256438 246483
rect 256490 246471 256496 246483
rect 336592 246471 336598 246483
rect 256490 246443 336598 246471
rect 256490 246431 256496 246443
rect 336592 246431 336598 246443
rect 336650 246431 336656 246483
rect 48016 246357 48022 246409
rect 48074 246397 48080 246409
rect 204496 246397 204502 246409
rect 48074 246369 204502 246397
rect 48074 246357 48080 246369
rect 204496 246357 204502 246369
rect 204554 246357 204560 246409
rect 255952 246357 255958 246409
rect 256010 246397 256016 246409
rect 338128 246397 338134 246409
rect 256010 246369 338134 246397
rect 256010 246357 256016 246369
rect 338128 246357 338134 246369
rect 338186 246357 338192 246409
rect 47440 246283 47446 246335
rect 47498 246323 47504 246335
rect 207184 246323 207190 246335
rect 47498 246295 207190 246323
rect 47498 246283 47504 246295
rect 207184 246283 207190 246295
rect 207242 246283 207248 246335
rect 255088 246283 255094 246335
rect 255146 246323 255152 246335
rect 339856 246323 339862 246335
rect 255146 246295 339862 246323
rect 255146 246283 255152 246295
rect 339856 246283 339862 246295
rect 339914 246283 339920 246335
rect 44656 246209 44662 246261
rect 44714 246249 44720 246261
rect 204784 246249 204790 246261
rect 44714 246221 204790 246249
rect 44714 246209 44720 246221
rect 204784 246209 204790 246221
rect 204842 246209 204848 246261
rect 254224 246209 254230 246261
rect 254282 246249 254288 246261
rect 341488 246249 341494 246261
rect 254282 246221 341494 246249
rect 254282 246209 254288 246221
rect 341488 246209 341494 246221
rect 341546 246209 341552 246261
rect 277552 246135 277558 246187
rect 277610 246175 277616 246187
rect 364336 246175 364342 246187
rect 277610 246147 364342 246175
rect 277610 246135 277616 246147
rect 364336 246135 364342 246147
rect 364394 246135 364400 246187
rect 139408 246061 139414 246113
rect 139466 246101 139472 246113
rect 141520 246101 141526 246113
rect 139466 246073 141526 246101
rect 139466 246061 139472 246073
rect 141520 246061 141526 246073
rect 141578 246061 141584 246113
rect 276400 246061 276406 246113
rect 276458 246101 276464 246113
rect 362800 246101 362806 246113
rect 276458 246073 362806 246101
rect 276458 246061 276464 246073
rect 362800 246061 362806 246073
rect 362858 246061 362864 246113
rect 674704 246061 674710 246113
rect 674762 246101 674768 246113
rect 675376 246101 675382 246113
rect 674762 246073 675382 246101
rect 674762 246061 674768 246073
rect 675376 246061 675382 246073
rect 675434 246061 675440 246113
rect 253744 245987 253750 246039
rect 253802 246027 253808 246039
rect 343216 246027 343222 246039
rect 253802 245999 343222 246027
rect 253802 245987 253808 245999
rect 343216 245987 343222 245999
rect 343274 245987 343280 246039
rect 273232 245913 273238 245965
rect 273290 245953 273296 245965
rect 360592 245953 360598 245965
rect 273290 245925 360598 245953
rect 273290 245913 273296 245925
rect 360592 245913 360598 245925
rect 360650 245913 360656 245965
rect 251536 245839 251542 245891
rect 251594 245879 251600 245891
rect 348016 245879 348022 245891
rect 251594 245851 348022 245879
rect 251594 245839 251600 245851
rect 348016 245839 348022 245851
rect 348074 245839 348080 245891
rect 139312 245765 139318 245817
rect 139370 245805 139376 245817
rect 143152 245805 143158 245817
rect 139370 245777 143158 245805
rect 139370 245765 139376 245777
rect 143152 245765 143158 245777
rect 143210 245765 143216 245817
rect 252016 245765 252022 245817
rect 252074 245805 252080 245817
rect 346288 245805 346294 245817
rect 252074 245777 346294 245805
rect 252074 245765 252080 245777
rect 346288 245765 346294 245777
rect 346346 245765 346352 245817
rect 250480 245691 250486 245743
rect 250538 245731 250544 245743
rect 349072 245731 349078 245743
rect 250538 245703 349078 245731
rect 250538 245691 250544 245703
rect 349072 245691 349078 245703
rect 349130 245691 349136 245743
rect 249808 245617 249814 245669
rect 249866 245657 249872 245669
rect 350800 245657 350806 245669
rect 249866 245629 350806 245657
rect 249866 245617 249872 245629
rect 350800 245617 350806 245629
rect 350858 245617 350864 245669
rect 248560 245543 248566 245595
rect 248618 245583 248624 245595
rect 354064 245583 354070 245595
rect 248618 245555 354070 245583
rect 248618 245543 248624 245555
rect 354064 245543 354070 245555
rect 354122 245543 354128 245595
rect 249328 245469 249334 245521
rect 249386 245509 249392 245521
rect 352816 245509 352822 245521
rect 249386 245481 352822 245509
rect 249386 245469 249392 245481
rect 352816 245469 352822 245481
rect 352874 245469 352880 245521
rect 263056 245395 263062 245447
rect 263114 245435 263120 245447
rect 372880 245435 372886 245447
rect 263114 245407 372886 245435
rect 263114 245395 263120 245407
rect 372880 245395 372886 245407
rect 372938 245395 372944 245447
rect 80656 245321 80662 245373
rect 80714 245361 80720 245373
rect 100720 245361 100726 245373
rect 80714 245333 100726 245361
rect 80714 245321 80720 245333
rect 100720 245321 100726 245333
rect 100778 245321 100784 245373
rect 247600 245321 247606 245373
rect 247658 245361 247664 245373
rect 355600 245361 355606 245373
rect 247658 245333 355606 245361
rect 247658 245321 247664 245333
rect 355600 245321 355606 245333
rect 355658 245321 355664 245373
rect 262672 245247 262678 245299
rect 262730 245287 262736 245299
rect 373456 245287 373462 245299
rect 262730 245259 373462 245287
rect 262730 245247 262736 245259
rect 373456 245247 373462 245259
rect 373514 245247 373520 245299
rect 246832 245173 246838 245225
rect 246890 245213 246896 245225
rect 357328 245213 357334 245225
rect 246890 245185 357334 245213
rect 246890 245173 246896 245185
rect 357328 245173 357334 245185
rect 357386 245173 357392 245225
rect 246352 245099 246358 245151
rect 246410 245139 246416 245151
rect 358864 245139 358870 245151
rect 246410 245111 358870 245139
rect 246410 245099 246416 245111
rect 358864 245099 358870 245111
rect 358922 245099 358928 245151
rect 158416 245025 158422 245077
rect 158474 245065 158480 245077
rect 168496 245065 168502 245077
rect 158474 245037 168502 245065
rect 158474 245025 158480 245037
rect 168496 245025 168502 245037
rect 168554 245025 168560 245077
rect 261424 245025 261430 245077
rect 261482 245065 261488 245077
rect 376720 245065 376726 245077
rect 261482 245037 376726 245065
rect 261482 245025 261488 245037
rect 376720 245025 376726 245037
rect 376778 245025 376784 245077
rect 260464 244951 260470 245003
rect 260522 244991 260528 245003
rect 378448 244991 378454 245003
rect 260522 244963 378454 244991
rect 260522 244951 260528 244963
rect 378448 244951 378454 244963
rect 378506 244951 378512 245003
rect 420496 244951 420502 245003
rect 420554 244991 420560 245003
rect 440560 244991 440566 245003
rect 420554 244963 440566 244991
rect 420554 244951 420560 244963
rect 440560 244951 440566 244963
rect 440618 244951 440624 245003
rect 204496 244877 204502 244929
rect 204554 244917 204560 244929
rect 205168 244917 205174 244929
rect 204554 244889 205174 244917
rect 204554 244877 204560 244889
rect 205168 244877 205174 244889
rect 205226 244917 205232 244929
rect 214096 244917 214102 244929
rect 205226 244889 214102 244917
rect 205226 244877 205232 244889
rect 214096 244877 214102 244889
rect 214154 244877 214160 244929
rect 259888 244877 259894 244929
rect 259946 244917 259952 244929
rect 379504 244917 379510 244929
rect 259946 244889 379510 244917
rect 259946 244877 259952 244889
rect 379504 244877 379510 244889
rect 379562 244877 379568 244929
rect 42352 244803 42358 244855
rect 42410 244843 42416 244855
rect 214480 244843 214486 244855
rect 42410 244815 214486 244843
rect 42410 244803 42416 244815
rect 214480 244803 214486 244815
rect 214538 244803 214544 244855
rect 259600 244803 259606 244855
rect 259658 244843 259664 244855
rect 380656 244843 380662 244855
rect 259658 244815 380662 244843
rect 259658 244803 259664 244815
rect 380656 244803 380662 244815
rect 380714 244803 380720 244855
rect 268720 244729 268726 244781
rect 268778 244769 268784 244781
rect 318256 244769 318262 244781
rect 268778 244741 318262 244769
rect 268778 244729 268784 244741
rect 318256 244729 318262 244741
rect 318314 244729 318320 244781
rect 217552 244655 217558 244707
rect 217610 244695 217616 244707
rect 257968 244695 257974 244707
rect 217610 244667 257974 244695
rect 217610 244655 217616 244667
rect 257968 244655 257974 244667
rect 258026 244655 258032 244707
rect 267568 244655 267574 244707
rect 267626 244695 267632 244707
rect 267626 244667 270398 244695
rect 267626 244655 267632 244667
rect 256336 244621 256342 244633
rect 236386 244593 256342 244621
rect 218416 244285 218422 244337
rect 218474 244325 218480 244337
rect 236386 244325 236414 244593
rect 256336 244581 256342 244593
rect 256394 244581 256400 244633
rect 236464 244507 236470 244559
rect 236522 244547 236528 244559
rect 268240 244547 268246 244559
rect 236522 244519 268246 244547
rect 236522 244507 236528 244519
rect 268240 244507 268246 244519
rect 268298 244507 268304 244559
rect 270370 244473 270398 244667
rect 278128 244655 278134 244707
rect 278186 244695 278192 244707
rect 318064 244695 318070 244707
rect 278186 244667 318070 244695
rect 278186 244655 278192 244667
rect 318064 244655 318070 244667
rect 318122 244655 318128 244707
rect 278032 244581 278038 244633
rect 278090 244621 278096 244633
rect 336400 244621 336406 244633
rect 278090 244593 336406 244621
rect 278090 244581 278096 244593
rect 336400 244581 336406 244593
rect 336458 244581 336464 244633
rect 270448 244507 270454 244559
rect 270506 244547 270512 244559
rect 318160 244547 318166 244559
rect 270506 244519 318166 244547
rect 270506 244507 270512 244519
rect 318160 244507 318166 244519
rect 318218 244507 318224 244559
rect 325456 244507 325462 244559
rect 325514 244547 325520 244559
rect 326800 244547 326806 244559
rect 325514 244519 326806 244547
rect 325514 244507 325520 244519
rect 326800 244507 326806 244519
rect 326858 244507 326864 244559
rect 338704 244473 338710 244485
rect 270370 244445 338710 244473
rect 338704 244433 338710 244445
rect 338762 244433 338768 244485
rect 398512 244473 398518 244485
rect 385570 244445 398518 244473
rect 261040 244359 261046 244411
rect 261098 244399 261104 244411
rect 335920 244399 335926 244411
rect 261098 244371 335926 244399
rect 261098 244359 261104 244371
rect 335920 244359 335926 244371
rect 335978 244359 335984 244411
rect 385570 244399 385598 244445
rect 398512 244433 398518 244445
rect 398570 244433 398576 244485
rect 337474 244371 385598 244399
rect 218474 244297 236414 244325
rect 218474 244285 218480 244297
rect 250192 244285 250198 244337
rect 250250 244325 250256 244337
rect 258832 244325 258838 244337
rect 250250 244297 258838 244325
rect 250250 244285 250256 244297
rect 258832 244285 258838 244297
rect 258890 244285 258896 244337
rect 277936 244285 277942 244337
rect 277994 244325 278000 244337
rect 337360 244325 337366 244337
rect 277994 244297 337366 244325
rect 277994 244285 278000 244297
rect 337360 244285 337366 244297
rect 337418 244285 337424 244337
rect 287632 244251 287638 244263
rect 251170 244223 287638 244251
rect 210160 244063 210166 244115
rect 210218 244103 210224 244115
rect 251170 244103 251198 244223
rect 287632 244211 287638 244223
rect 287690 244211 287696 244263
rect 294928 244211 294934 244263
rect 294986 244251 294992 244263
rect 306928 244251 306934 244263
rect 294986 244223 306934 244251
rect 294986 244211 294992 244223
rect 306928 244211 306934 244223
rect 306986 244211 306992 244263
rect 307024 244211 307030 244263
rect 307082 244251 307088 244263
rect 325360 244251 325366 244263
rect 307082 244223 325366 244251
rect 307082 244211 307088 244223
rect 325360 244211 325366 244223
rect 325418 244211 325424 244263
rect 325456 244211 325462 244263
rect 325514 244251 325520 244263
rect 337474 244251 337502 244371
rect 325514 244223 337502 244251
rect 325514 244211 325520 244223
rect 348496 244211 348502 244263
rect 348554 244251 348560 244263
rect 352816 244251 352822 244263
rect 348554 244223 352822 244251
rect 348554 244211 348560 244223
rect 352816 244211 352822 244223
rect 352874 244211 352880 244263
rect 254704 244137 254710 244189
rect 254762 244177 254768 244189
rect 356368 244177 356374 244189
rect 254762 244149 356374 244177
rect 254762 244137 254768 244149
rect 356368 244137 356374 244149
rect 356426 244137 356432 244189
rect 210218 244075 251198 244103
rect 210218 244063 210224 244075
rect 251248 244063 251254 244115
rect 251306 244103 251312 244115
rect 355024 244103 355030 244115
rect 251306 244075 355030 244103
rect 251306 244063 251312 244075
rect 355024 244063 355030 244075
rect 355082 244063 355088 244115
rect 77872 243989 77878 244041
rect 77930 244029 77936 244041
rect 149584 244029 149590 244041
rect 77930 244001 149590 244029
rect 77930 243989 77936 244001
rect 149584 243989 149590 244001
rect 149642 243989 149648 244041
rect 219472 243989 219478 244041
rect 219530 244029 219536 244041
rect 254032 244029 254038 244041
rect 219530 244001 254038 244029
rect 219530 243989 219536 244001
rect 254032 243989 254038 244001
rect 254090 243989 254096 244041
rect 256240 243989 256246 244041
rect 256298 244029 256304 244041
rect 357232 244029 357238 244041
rect 256298 244001 357238 244029
rect 256298 243989 256304 244001
rect 357232 243989 357238 244001
rect 357290 243989 357296 244041
rect 77008 243915 77014 243967
rect 77066 243955 77072 243967
rect 152464 243955 152470 243967
rect 77066 243927 152470 243955
rect 77066 243915 77072 243927
rect 152464 243915 152470 243927
rect 152522 243915 152528 243967
rect 248176 243915 248182 243967
rect 248234 243955 248240 243967
rect 353584 243955 353590 243967
rect 248234 243927 353590 243955
rect 248234 243915 248240 243927
rect 353584 243915 353590 243927
rect 353642 243915 353648 243967
rect 44944 243841 44950 243893
rect 45002 243881 45008 243893
rect 204688 243881 204694 243893
rect 45002 243853 204694 243881
rect 45002 243841 45008 243853
rect 204688 243841 204694 243853
rect 204746 243841 204752 243893
rect 220720 243841 220726 243893
rect 220778 243881 220784 243893
rect 250768 243881 250774 243893
rect 220778 243853 250774 243881
rect 220778 243841 220784 243853
rect 250768 243841 250774 243853
rect 250826 243841 250832 243893
rect 252976 243841 252982 243893
rect 253034 243881 253040 243893
rect 355792 243881 355798 243893
rect 253034 243853 355798 243881
rect 253034 243841 253040 243853
rect 355792 243841 355798 243853
rect 355850 243841 355856 243893
rect 45040 243767 45046 243819
rect 45098 243807 45104 243819
rect 204592 243807 204598 243819
rect 45098 243779 204598 243807
rect 45098 243767 45104 243779
rect 204592 243767 204598 243779
rect 204650 243767 204656 243819
rect 348496 243807 348502 243819
rect 247714 243779 348502 243807
rect 40240 243693 40246 243745
rect 40298 243733 40304 243745
rect 41776 243733 41782 243745
rect 40298 243705 41782 243733
rect 40298 243693 40304 243705
rect 41776 243693 41782 243705
rect 41834 243693 41840 243745
rect 45232 243693 45238 243745
rect 45290 243733 45296 243745
rect 206512 243733 206518 243745
rect 45290 243705 206518 243733
rect 45290 243693 45296 243705
rect 206512 243693 206518 243705
rect 206570 243693 206576 243745
rect 246928 243693 246934 243745
rect 246986 243733 246992 243745
rect 247714 243733 247742 243779
rect 348496 243767 348502 243779
rect 348554 243767 348560 243819
rect 360784 243767 360790 243819
rect 360842 243807 360848 243819
rect 397456 243807 397462 243819
rect 360842 243779 397462 243807
rect 360842 243767 360848 243779
rect 397456 243767 397462 243779
rect 397514 243767 397520 243819
rect 351856 243733 351862 243745
rect 246986 243705 247742 243733
rect 254242 243705 351862 243733
rect 246986 243693 246992 243705
rect 44560 243619 44566 243671
rect 44618 243659 44624 243671
rect 204496 243659 204502 243671
rect 44618 243631 204502 243659
rect 44618 243619 44624 243631
rect 204496 243619 204502 243631
rect 204554 243619 204560 243671
rect 41968 243545 41974 243597
rect 42026 243585 42032 243597
rect 42544 243585 42550 243597
rect 42026 243557 42550 243585
rect 42026 243545 42032 243557
rect 42544 243545 42550 243557
rect 42602 243545 42608 243597
rect 47728 243545 47734 243597
rect 47786 243585 47792 243597
rect 212368 243585 212374 243597
rect 47786 243557 212374 243585
rect 47786 243545 47792 243557
rect 212368 243545 212374 243557
rect 212426 243545 212432 243597
rect 245872 243545 245878 243597
rect 245930 243585 245936 243597
rect 254242 243585 254270 243705
rect 351856 243693 351862 243705
rect 351914 243693 351920 243745
rect 360208 243693 360214 243745
rect 360266 243733 360272 243745
rect 395920 243733 395926 243745
rect 360266 243705 395926 243733
rect 360266 243693 360272 243705
rect 395920 243693 395926 243705
rect 395978 243693 395984 243745
rect 254320 243619 254326 243671
rect 254378 243659 254384 243671
rect 254378 243631 257918 243659
rect 254378 243619 254384 243631
rect 245930 243557 254270 243585
rect 257890 243585 257918 243631
rect 258832 243619 258838 243671
rect 258890 243659 258896 243671
rect 354352 243659 354358 243671
rect 258890 243631 354358 243659
rect 258890 243619 258896 243631
rect 354352 243619 354358 243631
rect 354410 243619 354416 243671
rect 362032 243619 362038 243671
rect 362090 243659 362096 243671
rect 401776 243659 401782 243671
rect 362090 243631 401782 243659
rect 362090 243619 362096 243631
rect 401776 243619 401782 243631
rect 401834 243619 401840 243671
rect 350416 243585 350422 243597
rect 257890 243557 350422 243585
rect 245930 243545 245936 243557
rect 350416 243545 350422 243557
rect 350474 243545 350480 243597
rect 362416 243545 362422 243597
rect 362474 243585 362480 243597
rect 402832 243585 402838 243597
rect 362474 243557 402838 243585
rect 362474 243545 362480 243557
rect 402832 243545 402838 243557
rect 402890 243545 402896 243597
rect 45136 243471 45142 243523
rect 45194 243511 45200 243523
rect 212752 243511 212758 243523
rect 45194 243483 212758 243511
rect 45194 243471 45200 243483
rect 212752 243471 212758 243483
rect 212810 243471 212816 243523
rect 240976 243471 240982 243523
rect 241034 243511 241040 243523
rect 349648 243511 349654 243523
rect 241034 243483 349654 243511
rect 241034 243471 241040 243483
rect 349648 243471 349654 243483
rect 349706 243471 349712 243523
rect 363856 243471 363862 243523
rect 363914 243511 363920 243523
rect 405520 243511 405526 243523
rect 363914 243483 405526 243511
rect 363914 243471 363920 243483
rect 405520 243471 405526 243483
rect 405578 243471 405584 243523
rect 44752 243397 44758 243449
rect 44810 243437 44816 243449
rect 211888 243437 211894 243449
rect 44810 243409 211894 243437
rect 44810 243397 44816 243409
rect 211888 243397 211894 243409
rect 211946 243397 211952 243449
rect 239344 243397 239350 243449
rect 239402 243437 239408 243449
rect 349168 243437 349174 243449
rect 239402 243409 349174 243437
rect 239402 243397 239408 243409
rect 349168 243397 349174 243409
rect 349226 243397 349232 243449
rect 361936 243397 361942 243449
rect 361994 243437 362000 243449
rect 401104 243437 401110 243449
rect 361994 243409 401110 243437
rect 361994 243397 362000 243409
rect 401104 243397 401110 243409
rect 401162 243397 401168 243449
rect 44848 243323 44854 243375
rect 44906 243363 44912 243375
rect 212272 243363 212278 243375
rect 44906 243335 212278 243363
rect 44906 243323 44912 243335
rect 212272 243323 212278 243335
rect 212330 243323 212336 243375
rect 242128 243323 242134 243375
rect 242186 243363 242192 243375
rect 254320 243363 254326 243375
rect 242186 243335 254326 243363
rect 242186 243323 242192 243335
rect 254320 243323 254326 243335
rect 254378 243323 254384 243375
rect 351472 243363 351478 243375
rect 254434 243335 351478 243363
rect 243856 243249 243862 243301
rect 243914 243289 243920 243301
rect 254434 243289 254462 243335
rect 351472 243323 351478 243335
rect 351530 243323 351536 243375
rect 364624 243323 364630 243375
rect 364682 243363 364688 243375
rect 407248 243363 407254 243375
rect 364682 243335 407254 243363
rect 364682 243323 364688 243335
rect 407248 243323 407254 243335
rect 407306 243323 407312 243375
rect 243914 243261 254462 243289
rect 243914 243249 243920 243261
rect 264784 243249 264790 243301
rect 264842 243289 264848 243301
rect 313264 243289 313270 243301
rect 264842 243261 313270 243289
rect 264842 243249 264848 243261
rect 313264 243249 313270 243261
rect 313322 243249 313328 243301
rect 316528 243249 316534 243301
rect 316586 243289 316592 243301
rect 381136 243289 381142 243301
rect 316586 243261 381142 243289
rect 316586 243249 316592 243261
rect 381136 243249 381142 243261
rect 381194 243249 381200 243301
rect 265744 243175 265750 243227
rect 265802 243215 265808 243227
rect 311632 243215 311638 243227
rect 265802 243187 311638 243215
rect 265802 243175 265808 243187
rect 311632 243175 311638 243187
rect 311690 243175 311696 243227
rect 315568 243175 315574 243227
rect 315626 243215 315632 243227
rect 348496 243215 348502 243227
rect 315626 243187 348502 243215
rect 315626 243175 315632 243187
rect 348496 243175 348502 243187
rect 348554 243175 348560 243227
rect 368560 243175 368566 243227
rect 368618 243215 368624 243227
rect 378928 243215 378934 243227
rect 368618 243187 378934 243215
rect 368618 243175 368624 243187
rect 378928 243175 378934 243187
rect 378986 243175 378992 243227
rect 266608 243101 266614 243153
rect 266666 243141 266672 243153
rect 310480 243141 310486 243153
rect 266666 243113 310486 243141
rect 266666 243101 266672 243113
rect 310480 243101 310486 243113
rect 310538 243101 310544 243153
rect 326608 243101 326614 243153
rect 326666 243141 326672 243153
rect 374992 243141 374998 243153
rect 326666 243113 374998 243141
rect 326666 243101 326672 243113
rect 374992 243101 374998 243113
rect 375050 243101 375056 243153
rect 268048 243027 268054 243079
rect 268106 243067 268112 243079
rect 294928 243067 294934 243079
rect 268106 243039 294934 243067
rect 268106 243027 268112 243039
rect 294928 243027 294934 243039
rect 294986 243027 294992 243079
rect 305680 243067 305686 243079
rect 295042 243039 305686 243067
rect 268816 242953 268822 243005
rect 268874 242993 268880 243005
rect 295042 242993 295070 243039
rect 305680 243027 305686 243039
rect 305738 243027 305744 243079
rect 308002 243039 308318 243067
rect 268874 242965 295070 242993
rect 268874 242953 268880 242965
rect 295120 242953 295126 243005
rect 295178 242993 295184 243005
rect 302224 242993 302230 243005
rect 295178 242965 302230 242993
rect 295178 242953 295184 242965
rect 302224 242953 302230 242965
rect 302282 242953 302288 243005
rect 265840 242879 265846 242931
rect 265898 242919 265904 242931
rect 278128 242919 278134 242931
rect 265898 242891 278134 242919
rect 265898 242879 265904 242891
rect 278128 242879 278134 242891
rect 278186 242879 278192 242931
rect 282064 242879 282070 242931
rect 282122 242919 282128 242931
rect 308002 242919 308030 243039
rect 308290 242993 308318 243039
rect 312976 243027 312982 243079
rect 313034 243067 313040 243079
rect 326416 243067 326422 243079
rect 313034 243039 326422 243067
rect 313034 243027 313040 243039
rect 326416 243027 326422 243039
rect 326474 243027 326480 243079
rect 326704 243027 326710 243079
rect 326762 243067 326768 243079
rect 377200 243067 377206 243079
rect 326762 243039 377206 243067
rect 326762 243027 326768 243039
rect 377200 243027 377206 243039
rect 377258 243027 377264 243079
rect 326320 242993 326326 243005
rect 308290 242965 326326 242993
rect 326320 242953 326326 242965
rect 326378 242953 326384 243005
rect 326512 242953 326518 243005
rect 326570 242993 326576 243005
rect 372976 242993 372982 243005
rect 326570 242965 372982 242993
rect 326570 242953 326576 242965
rect 372976 242953 372982 242965
rect 373034 242953 373040 243005
rect 325744 242919 325750 242931
rect 282122 242891 308030 242919
rect 316834 242891 325750 242919
rect 282122 242879 282128 242891
rect 262768 242805 262774 242857
rect 262826 242845 262832 242857
rect 278032 242845 278038 242857
rect 262826 242817 278038 242845
rect 262826 242805 262832 242817
rect 278032 242805 278038 242817
rect 278090 242805 278096 242857
rect 283408 242805 283414 242857
rect 283466 242845 283472 242857
rect 283466 242817 298046 242845
rect 283466 242805 283472 242817
rect 263920 242731 263926 242783
rect 263978 242771 263984 242783
rect 277936 242771 277942 242783
rect 263978 242743 277942 242771
rect 263978 242731 263984 242743
rect 277936 242731 277942 242743
rect 277994 242731 278000 242783
rect 293584 242731 293590 242783
rect 293642 242771 293648 242783
rect 296656 242771 296662 242783
rect 293642 242743 296662 242771
rect 293642 242731 293648 242743
rect 296656 242731 296662 242743
rect 296714 242731 296720 242783
rect 270256 242657 270262 242709
rect 270314 242697 270320 242709
rect 295120 242697 295126 242709
rect 270314 242669 295126 242697
rect 270314 242657 270320 242669
rect 295120 242657 295126 242669
rect 295178 242657 295184 242709
rect 298018 242697 298046 242817
rect 298096 242805 298102 242857
rect 298154 242845 298160 242857
rect 316720 242845 316726 242857
rect 298154 242817 316726 242845
rect 298154 242805 298160 242817
rect 316720 242805 316726 242817
rect 316778 242805 316784 242857
rect 298192 242731 298198 242783
rect 298250 242771 298256 242783
rect 316834 242771 316862 242891
rect 325744 242879 325750 242891
rect 325802 242879 325808 242931
rect 330640 242879 330646 242931
rect 330698 242919 330704 242931
rect 361072 242919 361078 242931
rect 330698 242891 361078 242919
rect 330698 242879 330704 242891
rect 361072 242879 361078 242891
rect 361130 242879 361136 242931
rect 317200 242805 317206 242857
rect 317258 242845 317264 242857
rect 323536 242845 323542 242857
rect 317258 242817 323542 242845
rect 317258 242805 317264 242817
rect 323536 242805 323542 242817
rect 323594 242805 323600 242857
rect 331024 242805 331030 242857
rect 331082 242845 331088 242857
rect 362128 242845 362134 242857
rect 331082 242817 362134 242845
rect 331082 242805 331088 242817
rect 362128 242805 362134 242817
rect 362186 242805 362192 242857
rect 298250 242743 316862 242771
rect 298250 242731 298256 242743
rect 318256 242731 318262 242783
rect 318314 242771 318320 242783
rect 339568 242771 339574 242783
rect 318314 242743 339574 242771
rect 318314 242731 318320 242743
rect 339568 242731 339574 242743
rect 339626 242731 339632 242783
rect 348496 242731 348502 242783
rect 348554 242771 348560 242783
rect 368560 242771 368566 242783
rect 348554 242743 368566 242771
rect 348554 242731 348560 242743
rect 368560 242731 368566 242743
rect 368618 242731 368624 242783
rect 674896 242731 674902 242783
rect 674954 242771 674960 242783
rect 675376 242771 675382 242783
rect 674954 242743 675382 242771
rect 674954 242731 674960 242743
rect 675376 242731 675382 242743
rect 675434 242731 675440 242783
rect 324016 242697 324022 242709
rect 298018 242669 324022 242697
rect 324016 242657 324022 242669
rect 324074 242657 324080 242709
rect 330256 242657 330262 242709
rect 330314 242697 330320 242709
rect 360016 242697 360022 242709
rect 330314 242669 360022 242697
rect 330314 242657 330320 242669
rect 360016 242657 360022 242669
rect 360074 242657 360080 242709
rect 282928 242583 282934 242635
rect 282986 242623 282992 242635
rect 282986 242595 316574 242623
rect 282986 242583 282992 242595
rect 275248 242509 275254 242561
rect 275306 242549 275312 242561
rect 309424 242549 309430 242561
rect 275306 242521 309430 242549
rect 275306 242509 275312 242521
rect 309424 242509 309430 242521
rect 309482 242509 309488 242561
rect 316546 242549 316574 242595
rect 316720 242583 316726 242635
rect 316778 242623 316784 242635
rect 317200 242623 317206 242635
rect 316778 242595 317206 242623
rect 316778 242583 316784 242595
rect 317200 242583 317206 242595
rect 317258 242583 317264 242635
rect 318064 242583 318070 242635
rect 318122 242623 318128 242635
rect 337840 242623 337846 242635
rect 318122 242595 337846 242623
rect 318122 242583 318128 242595
rect 337840 242583 337846 242595
rect 337898 242583 337904 242635
rect 324688 242549 324694 242561
rect 316546 242521 324694 242549
rect 324688 242509 324694 242521
rect 324746 242509 324752 242561
rect 330736 242509 330742 242561
rect 330794 242549 330800 242561
rect 361648 242549 361654 242561
rect 330794 242521 361654 242549
rect 330794 242509 330800 242521
rect 361648 242509 361654 242521
rect 361706 242509 361712 242561
rect 139120 242435 139126 242487
rect 139178 242475 139184 242487
rect 140272 242475 140278 242487
rect 139178 242447 140278 242475
rect 139178 242435 139184 242447
rect 140272 242435 140278 242447
rect 140330 242435 140336 242487
rect 269872 242435 269878 242487
rect 269930 242475 269936 242487
rect 302992 242475 302998 242487
rect 269930 242447 302998 242475
rect 269930 242435 269936 242447
rect 302992 242435 302998 242447
rect 303050 242435 303056 242487
rect 326224 242475 326230 242487
rect 308194 242447 326230 242475
rect 293200 242361 293206 242413
rect 293258 242401 293264 242413
rect 293258 242373 308126 242401
rect 293258 242361 293264 242373
rect 140368 242287 140374 242339
rect 140426 242327 140432 242339
rect 141328 242327 141334 242339
rect 140426 242299 141334 242327
rect 140426 242287 140432 242299
rect 141328 242287 141334 242299
rect 141386 242287 141392 242339
rect 268912 242287 268918 242339
rect 268970 242327 268976 242339
rect 304624 242327 304630 242339
rect 268970 242299 304630 242327
rect 268970 242287 268976 242299
rect 304624 242287 304630 242299
rect 304682 242287 304688 242339
rect 308098 242327 308126 242373
rect 308194 242327 308222 242447
rect 326224 242435 326230 242447
rect 326282 242435 326288 242487
rect 318160 242361 318166 242413
rect 318218 242401 318224 242413
rect 340336 242401 340342 242413
rect 318218 242373 340342 242401
rect 318218 242361 318224 242373
rect 340336 242361 340342 242373
rect 340394 242361 340400 242413
rect 674992 242361 674998 242413
rect 675050 242401 675056 242413
rect 675376 242401 675382 242413
rect 675050 242373 675382 242401
rect 675050 242361 675056 242373
rect 675376 242361 675382 242373
rect 675434 242361 675440 242413
rect 308098 242299 308222 242327
rect 313456 242287 313462 242339
rect 313514 242327 313520 242339
rect 326608 242327 326614 242339
rect 313514 242299 326614 242327
rect 313514 242287 313520 242299
rect 326608 242287 326614 242299
rect 326666 242287 326672 242339
rect 283792 242213 283798 242265
rect 283850 242253 283856 242265
rect 298096 242253 298102 242265
rect 283850 242225 298102 242253
rect 283850 242213 283856 242225
rect 298096 242213 298102 242225
rect 298154 242213 298160 242265
rect 314800 242213 314806 242265
rect 314858 242253 314864 242265
rect 326704 242253 326710 242265
rect 314858 242225 326710 242253
rect 314858 242213 314864 242225
rect 326704 242213 326710 242225
rect 326762 242213 326768 242265
rect 37264 242139 37270 242191
rect 37322 242179 37328 242191
rect 42736 242179 42742 242191
rect 37322 242151 42742 242179
rect 37322 242139 37328 242151
rect 42736 242139 42742 242151
rect 42794 242139 42800 242191
rect 267874 242151 287006 242179
rect 40048 242065 40054 242117
rect 40106 242105 40112 242117
rect 42352 242105 42358 242117
rect 40106 242077 42358 242105
rect 40106 242065 40112 242077
rect 42352 242065 42358 242077
rect 42410 242065 42416 242117
rect 37360 241991 37366 242043
rect 37418 242031 37424 242043
rect 43120 242031 43126 242043
rect 37418 242003 43126 242031
rect 37418 241991 37424 242003
rect 43120 241991 43126 242003
rect 43178 241991 43184 242043
rect 140752 241991 140758 242043
rect 140810 242031 140816 242043
rect 141136 242031 141142 242043
rect 140810 242003 141142 242031
rect 140810 241991 140816 242003
rect 141136 241991 141142 242003
rect 141194 241991 141200 242043
rect 267874 242031 267902 242151
rect 286768 242031 286774 242043
rect 259234 242003 267902 242031
rect 286018 242003 286774 242031
rect 40144 241917 40150 241969
rect 40202 241957 40208 241969
rect 43024 241957 43030 241969
rect 40202 241929 43030 241957
rect 40202 241917 40208 241929
rect 43024 241917 43030 241929
rect 43082 241917 43088 241969
rect 44656 241917 44662 241969
rect 44714 241957 44720 241969
rect 206416 241957 206422 241969
rect 44714 241929 206422 241957
rect 44714 241917 44720 241929
rect 206416 241917 206422 241929
rect 206474 241917 206480 241969
rect 206512 241917 206518 241969
rect 206570 241957 206576 241969
rect 207088 241957 207094 241969
rect 206570 241929 207094 241957
rect 206570 241917 206576 241929
rect 207088 241917 207094 241929
rect 207146 241957 207152 241969
rect 213136 241957 213142 241969
rect 207146 241929 213142 241957
rect 207146 241917 207152 241929
rect 213136 241917 213142 241929
rect 213194 241917 213200 241969
rect 244624 241917 244630 241969
rect 244682 241957 244688 241969
rect 259234 241957 259262 242003
rect 244682 241929 259262 241957
rect 244682 241917 244688 241929
rect 43216 241843 43222 241895
rect 43274 241883 43280 241895
rect 43696 241883 43702 241895
rect 43274 241855 43702 241883
rect 43274 241843 43280 241855
rect 43696 241843 43702 241855
rect 43754 241883 43760 241895
rect 140752 241883 140758 241895
rect 43754 241855 140758 241883
rect 43754 241843 43760 241855
rect 140752 241843 140758 241855
rect 140810 241843 140816 241895
rect 152464 241843 152470 241895
rect 152522 241883 152528 241895
rect 152522 241855 167006 241883
rect 152522 241843 152528 241855
rect 41680 241769 41686 241821
rect 41738 241809 41744 241821
rect 43504 241809 43510 241821
rect 41738 241781 43510 241809
rect 41738 241769 41744 241781
rect 43504 241769 43510 241781
rect 43562 241809 43568 241821
rect 140656 241809 140662 241821
rect 43562 241781 140662 241809
rect 43562 241769 43568 241781
rect 140656 241769 140662 241781
rect 140714 241769 140720 241821
rect 166978 241735 167006 241855
rect 221392 241843 221398 241895
rect 221450 241883 221456 241895
rect 234544 241883 234550 241895
rect 221450 241855 234550 241883
rect 221450 241843 221456 241855
rect 234544 241843 234550 241855
rect 234602 241843 234608 241895
rect 240208 241843 240214 241895
rect 240266 241883 240272 241895
rect 259504 241883 259510 241895
rect 240266 241855 259510 241883
rect 240266 241843 240272 241855
rect 259504 241843 259510 241855
rect 259562 241843 259568 241895
rect 271888 241843 271894 241895
rect 271946 241883 271952 241895
rect 286018 241883 286046 242003
rect 286768 241991 286774 242003
rect 286826 241991 286832 242043
rect 286978 241957 287006 242151
rect 293008 242139 293014 242191
rect 293066 242179 293072 242191
rect 325264 242179 325270 242191
rect 293066 242151 325270 242179
rect 293066 242139 293072 242151
rect 325264 242139 325270 242151
rect 325322 242139 325328 242191
rect 287728 242065 287734 242117
rect 287786 242105 287792 242117
rect 298192 242105 298198 242117
rect 287786 242077 298198 242105
rect 287786 242065 287792 242077
rect 298192 242065 298198 242077
rect 298250 242065 298256 242117
rect 320464 242065 320470 242117
rect 320522 242105 320528 242117
rect 339472 242105 339478 242117
rect 320522 242077 339478 242105
rect 320522 242065 320528 242077
rect 339472 242065 339478 242077
rect 339530 242065 339536 242117
rect 292720 241991 292726 242043
rect 292778 242031 292784 242043
rect 324208 242031 324214 242043
rect 292778 242003 324214 242031
rect 292778 241991 292784 242003
rect 324208 241991 324214 242003
rect 324266 241991 324272 242043
rect 286978 241929 295934 241957
rect 271946 241855 286046 241883
rect 271946 241843 271952 241855
rect 286096 241843 286102 241895
rect 286154 241883 286160 241895
rect 289840 241883 289846 241895
rect 286154 241855 289846 241883
rect 286154 241843 286160 241855
rect 289840 241843 289846 241855
rect 289898 241843 289904 241895
rect 289936 241843 289942 241895
rect 289994 241883 290000 241895
rect 295792 241883 295798 241895
rect 289994 241855 295798 241883
rect 289994 241843 290000 241855
rect 295792 241843 295798 241855
rect 295850 241843 295856 241895
rect 295906 241883 295934 241929
rect 296656 241917 296662 241969
rect 296714 241957 296720 241969
rect 307024 241957 307030 241969
rect 296714 241929 307030 241957
rect 296714 241917 296720 241929
rect 307024 241917 307030 241929
rect 307082 241917 307088 241969
rect 338512 241957 338518 241969
rect 338146 241929 338518 241957
rect 330544 241883 330550 241895
rect 295906 241855 330550 241883
rect 330544 241843 330550 241855
rect 330602 241843 330608 241895
rect 331312 241843 331318 241895
rect 331370 241883 331376 241895
rect 338146 241883 338174 241929
rect 338512 241917 338518 241929
rect 338570 241917 338576 241969
rect 383536 241917 383542 241969
rect 383594 241957 383600 241969
rect 383594 241929 387326 241957
rect 383594 241917 383600 241929
rect 387298 241895 387326 241929
rect 331370 241855 338174 241883
rect 331370 241843 331376 241855
rect 338224 241843 338230 241895
rect 338282 241883 338288 241895
rect 352912 241883 352918 241895
rect 338282 241855 352918 241883
rect 338282 241843 338288 241855
rect 352912 241843 352918 241855
rect 352970 241843 352976 241895
rect 368272 241843 368278 241895
rect 368330 241883 368336 241895
rect 368330 241855 372638 241883
rect 368330 241843 368336 241855
rect 223120 241769 223126 241821
rect 223178 241809 223184 241821
rect 233968 241809 233974 241821
rect 223178 241781 233974 241809
rect 223178 241769 223184 241781
rect 233968 241769 233974 241781
rect 234026 241769 234032 241821
rect 239728 241769 239734 241821
rect 239786 241809 239792 241821
rect 239786 241781 242750 241809
rect 239786 241769 239792 241781
rect 216688 241735 216694 241747
rect 166978 241707 216694 241735
rect 216688 241695 216694 241707
rect 216746 241695 216752 241747
rect 228880 241695 228886 241747
rect 228938 241735 228944 241747
rect 241072 241735 241078 241747
rect 228938 241707 241078 241735
rect 228938 241695 228944 241707
rect 241072 241695 241078 241707
rect 241130 241695 241136 241747
rect 242722 241735 242750 241781
rect 245392 241769 245398 241821
rect 245450 241809 245456 241821
rect 273232 241809 273238 241821
rect 245450 241781 273238 241809
rect 245450 241769 245456 241781
rect 273232 241769 273238 241781
rect 273290 241769 273296 241821
rect 275440 241769 275446 241821
rect 275498 241809 275504 241821
rect 291088 241809 291094 241821
rect 275498 241781 291094 241809
rect 275498 241769 275504 241781
rect 291088 241769 291094 241781
rect 291146 241769 291152 241821
rect 291280 241769 291286 241821
rect 291338 241809 291344 241821
rect 298384 241809 298390 241821
rect 291338 241781 298390 241809
rect 291338 241769 291344 241781
rect 298384 241769 298390 241781
rect 298442 241769 298448 241821
rect 328912 241769 328918 241821
rect 328970 241809 328976 241821
rect 338128 241809 338134 241821
rect 328970 241781 338134 241809
rect 328970 241769 328976 241781
rect 338128 241769 338134 241781
rect 338186 241769 338192 241821
rect 338896 241769 338902 241821
rect 338954 241809 338960 241821
rect 353392 241809 353398 241821
rect 338954 241781 353398 241809
rect 338954 241769 338960 241781
rect 353392 241769 353398 241781
rect 353450 241769 353456 241821
rect 261232 241735 261238 241747
rect 242722 241707 261238 241735
rect 261232 241695 261238 241707
rect 261290 241695 261296 241747
rect 271024 241695 271030 241747
rect 271082 241735 271088 241747
rect 286480 241735 286486 241747
rect 271082 241707 286486 241735
rect 271082 241695 271088 241707
rect 286480 241695 286486 241707
rect 286538 241695 286544 241747
rect 289744 241695 289750 241747
rect 289802 241735 289808 241747
rect 296272 241735 296278 241747
rect 289802 241707 296278 241735
rect 289802 241695 289808 241707
rect 296272 241695 296278 241707
rect 296330 241695 296336 241747
rect 318256 241695 318262 241747
rect 318314 241735 318320 241747
rect 334960 241735 334966 241747
rect 318314 241707 334966 241735
rect 318314 241695 318320 241707
rect 334960 241695 334966 241707
rect 335018 241695 335024 241747
rect 337072 241695 337078 241747
rect 337130 241735 337136 241747
rect 345808 241735 345814 241747
rect 337130 241707 345814 241735
rect 337130 241695 337136 241707
rect 345808 241695 345814 241707
rect 345866 241695 345872 241747
rect 354544 241735 354550 241747
rect 345922 241707 354550 241735
rect 226864 241621 226870 241673
rect 226922 241661 226928 241673
rect 232144 241661 232150 241673
rect 226922 241633 232150 241661
rect 226922 241621 226928 241633
rect 232144 241621 232150 241633
rect 232202 241621 232208 241673
rect 244240 241661 244246 241673
rect 232258 241633 244246 241661
rect 227536 241547 227542 241599
rect 227594 241587 227600 241599
rect 232258 241587 232286 241633
rect 244240 241621 244246 241633
rect 244298 241621 244304 241673
rect 281296 241621 281302 241673
rect 281354 241661 281360 241673
rect 289936 241661 289942 241673
rect 281354 241633 289942 241661
rect 281354 241621 281360 241633
rect 289936 241621 289942 241633
rect 289994 241621 290000 241673
rect 290128 241621 290134 241673
rect 290186 241661 290192 241673
rect 290186 241633 301022 241661
rect 290186 241621 290192 241633
rect 227594 241559 232286 241587
rect 227594 241547 227600 241559
rect 236656 241547 236662 241599
rect 236714 241587 236720 241599
rect 248656 241587 248662 241599
rect 236714 241559 248662 241587
rect 236714 241547 236720 241559
rect 248656 241547 248662 241559
rect 248714 241547 248720 241599
rect 271984 241547 271990 241599
rect 272042 241587 272048 241599
rect 288112 241587 288118 241599
rect 272042 241559 288118 241587
rect 272042 241547 272048 241559
rect 288112 241547 288118 241559
rect 288170 241547 288176 241599
rect 228496 241473 228502 241525
rect 228554 241513 228560 241525
rect 238384 241513 238390 241525
rect 228554 241485 238390 241513
rect 228554 241473 228560 241485
rect 238384 241473 238390 241485
rect 238442 241473 238448 241525
rect 238768 241473 238774 241525
rect 238826 241513 238832 241525
rect 238826 241485 247262 241513
rect 238826 241473 238832 241485
rect 225904 241399 225910 241451
rect 225962 241439 225968 241451
rect 232336 241439 232342 241451
rect 225962 241411 232342 241439
rect 225962 241399 225968 241411
rect 232336 241399 232342 241411
rect 232394 241399 232400 241451
rect 236560 241439 236566 241451
rect 235234 241411 236566 241439
rect 225328 241325 225334 241377
rect 225386 241365 225392 241377
rect 232624 241365 232630 241377
rect 225386 241337 232630 241365
rect 225386 241325 225392 241337
rect 232624 241325 232630 241337
rect 232682 241325 232688 241377
rect 217264 241251 217270 241303
rect 217322 241291 217328 241303
rect 229168 241291 229174 241303
rect 217322 241263 229174 241291
rect 217322 241251 217328 241263
rect 229168 241251 229174 241263
rect 229226 241251 229232 241303
rect 235234 241291 235262 241411
rect 236560 241399 236566 241411
rect 236618 241399 236624 241451
rect 237232 241399 237238 241451
rect 237290 241439 237296 241451
rect 247120 241439 247126 241451
rect 237290 241411 247126 241439
rect 237290 241399 237296 241411
rect 247120 241399 247126 241411
rect 247178 241399 247184 241451
rect 235312 241325 235318 241377
rect 235370 241365 235376 241377
rect 245968 241365 245974 241377
rect 235370 241337 245974 241365
rect 235370 241325 235376 241337
rect 245968 241325 245974 241337
rect 246026 241325 246032 241377
rect 247234 241365 247262 241485
rect 247312 241473 247318 241525
rect 247370 241513 247376 241525
rect 262192 241513 262198 241525
rect 247370 241485 262198 241513
rect 247370 241473 247376 241485
rect 262192 241473 262198 241485
rect 262250 241473 262256 241525
rect 264400 241473 264406 241525
rect 264458 241513 264464 241525
rect 275632 241513 275638 241525
rect 264458 241485 275638 241513
rect 264458 241473 264464 241485
rect 275632 241473 275638 241485
rect 275690 241473 275696 241525
rect 283312 241473 283318 241525
rect 283370 241513 283376 241525
rect 289744 241513 289750 241525
rect 283370 241485 289750 241513
rect 283370 241473 283376 241485
rect 289744 241473 289750 241485
rect 289802 241473 289808 241525
rect 290704 241473 290710 241525
rect 290762 241513 290768 241525
rect 297616 241513 297622 241525
rect 290762 241485 297622 241513
rect 290762 241473 290768 241485
rect 297616 241473 297622 241485
rect 297674 241473 297680 241525
rect 273712 241399 273718 241451
rect 273770 241439 273776 241451
rect 286096 241439 286102 241451
rect 273770 241411 286102 241439
rect 273770 241399 273776 241411
rect 286096 241399 286102 241411
rect 286154 241399 286160 241451
rect 286672 241399 286678 241451
rect 286730 241439 286736 241451
rect 296944 241439 296950 241451
rect 286730 241411 296950 241439
rect 286730 241399 286736 241411
rect 296944 241399 296950 241411
rect 297002 241399 297008 241451
rect 262864 241365 262870 241377
rect 247234 241337 262870 241365
rect 262864 241325 262870 241337
rect 262922 241325 262928 241377
rect 271120 241325 271126 241377
rect 271178 241365 271184 241377
rect 286384 241365 286390 241377
rect 271178 241337 286390 241365
rect 271178 241325 271184 241337
rect 286384 241325 286390 241337
rect 286442 241325 286448 241377
rect 289456 241365 289462 241377
rect 286594 241337 289462 241365
rect 229858 241263 235262 241291
rect 220336 241103 220342 241155
rect 220394 241143 220400 241155
rect 229858 241143 229886 241263
rect 236272 241251 236278 241303
rect 236330 241291 236336 241303
rect 244912 241291 244918 241303
rect 236330 241263 244918 241291
rect 236330 241251 236336 241263
rect 244912 241251 244918 241263
rect 244970 241251 244976 241303
rect 272560 241251 272566 241303
rect 272618 241291 272624 241303
rect 286288 241291 286294 241303
rect 272618 241263 286294 241291
rect 272618 241251 272624 241263
rect 286288 241251 286294 241263
rect 286346 241251 286352 241303
rect 239344 241177 239350 241229
rect 239402 241217 239408 241229
rect 247312 241217 247318 241229
rect 239402 241189 247318 241217
rect 239402 241177 239408 241189
rect 247312 241177 247318 241189
rect 247370 241177 247376 241229
rect 273520 241177 273526 241229
rect 273578 241217 273584 241229
rect 286192 241217 286198 241229
rect 273578 241189 286198 241217
rect 273578 241177 273584 241189
rect 286192 241177 286198 241189
rect 286250 241177 286256 241229
rect 286594 241217 286622 241337
rect 289456 241325 289462 241337
rect 289514 241325 289520 241377
rect 289744 241325 289750 241377
rect 289802 241365 289808 241377
rect 300016 241365 300022 241377
rect 289802 241337 300022 241365
rect 289802 241325 289808 241337
rect 300016 241325 300022 241337
rect 300074 241325 300080 241377
rect 286768 241251 286774 241303
rect 286826 241291 286832 241303
rect 298288 241291 298294 241303
rect 286826 241263 298294 241291
rect 286826 241251 286832 241263
rect 298288 241251 298294 241263
rect 298346 241251 298352 241303
rect 286306 241189 286622 241217
rect 220394 241115 229886 241143
rect 220394 241103 220400 241115
rect 229936 241103 229942 241155
rect 229994 241143 230000 241155
rect 240400 241143 240406 241155
rect 229994 241115 240406 241143
rect 229994 241103 230000 241115
rect 240400 241103 240406 241115
rect 240458 241103 240464 241155
rect 240496 241103 240502 241155
rect 240554 241143 240560 241155
rect 264304 241143 264310 241155
rect 240554 241115 264310 241143
rect 240554 241103 240560 241115
rect 264304 241103 264310 241115
rect 264362 241103 264368 241155
rect 275920 241103 275926 241155
rect 275978 241143 275984 241155
rect 286306 241143 286334 241189
rect 287056 241177 287062 241229
rect 287114 241217 287120 241229
rect 291280 241217 291286 241229
rect 287114 241189 291286 241217
rect 287114 241177 287120 241189
rect 291280 241177 291286 241189
rect 291338 241177 291344 241229
rect 291376 241177 291382 241229
rect 291434 241217 291440 241229
rect 291434 241189 300926 241217
rect 291434 241177 291440 241189
rect 294352 241143 294358 241155
rect 275978 241115 286334 241143
rect 286402 241115 294358 241143
rect 275978 241103 275984 241115
rect 226480 241029 226486 241081
rect 226538 241069 226544 241081
rect 239440 241069 239446 241081
rect 226538 241041 239446 241069
rect 226538 241029 226544 241041
rect 239440 241029 239446 241041
rect 239498 241029 239504 241081
rect 247408 241029 247414 241081
rect 247466 241069 247472 241081
rect 267760 241069 267766 241081
rect 247466 241041 267766 241069
rect 247466 241029 247472 241041
rect 267760 241029 267766 241041
rect 267818 241029 267824 241081
rect 277360 241029 277366 241081
rect 277418 241069 277424 241081
rect 286000 241069 286006 241081
rect 277418 241041 286006 241069
rect 277418 241029 277424 241041
rect 286000 241029 286006 241041
rect 286058 241029 286064 241081
rect 286096 241029 286102 241081
rect 286154 241069 286160 241081
rect 286402 241069 286430 241115
rect 294352 241103 294358 241115
rect 294410 241103 294416 241155
rect 294448 241103 294454 241155
rect 294506 241143 294512 241155
rect 297712 241143 297718 241155
rect 294506 241115 297718 241143
rect 294506 241103 294512 241115
rect 297712 241103 297718 241115
rect 297770 241103 297776 241155
rect 286154 241041 286430 241069
rect 286154 241029 286160 241041
rect 286480 241029 286486 241081
rect 286538 241069 286544 241081
rect 300784 241069 300790 241081
rect 286538 241041 300790 241069
rect 286538 241029 286544 241041
rect 300784 241029 300790 241041
rect 300842 241029 300848 241081
rect 223312 240955 223318 241007
rect 223370 240995 223376 241007
rect 235312 240995 235318 241007
rect 223370 240967 235318 240995
rect 223370 240955 223376 240967
rect 235312 240955 235318 240967
rect 235370 240955 235376 241007
rect 243184 240995 243190 241007
rect 235474 240967 243190 240995
rect 42736 240881 42742 240933
rect 42794 240921 42800 240933
rect 43312 240921 43318 240933
rect 42794 240893 43318 240921
rect 42794 240881 42800 240893
rect 43312 240881 43318 240893
rect 43370 240881 43376 240933
rect 224560 240881 224566 240933
rect 224618 240921 224624 240933
rect 235474 240921 235502 240967
rect 243184 240955 243190 240967
rect 243242 240955 243248 241007
rect 243280 240955 243286 241007
rect 243338 240995 243344 241007
rect 264976 240995 264982 241007
rect 243338 240967 264982 240995
rect 243338 240955 243344 240967
rect 264976 240955 264982 240967
rect 265034 240955 265040 241007
rect 272848 240955 272854 241007
rect 272906 240995 272912 241007
rect 285424 240995 285430 241007
rect 272906 240967 285430 240995
rect 272906 240955 272912 240967
rect 285424 240955 285430 240967
rect 285482 240955 285488 241007
rect 285520 240955 285526 241007
rect 285578 240995 285584 241007
rect 290704 240995 290710 241007
rect 285578 240967 290710 240995
rect 285578 240955 285584 240967
rect 290704 240955 290710 240967
rect 290762 240955 290768 241007
rect 290800 240955 290806 241007
rect 290858 240995 290864 241007
rect 298480 240995 298486 241007
rect 290858 240967 298486 240995
rect 290858 240955 290864 240967
rect 298480 240955 298486 240967
rect 298538 240955 298544 241007
rect 249232 240921 249238 240933
rect 224618 240893 235502 240921
rect 237442 240893 249238 240921
rect 224618 240881 224624 240893
rect 223888 240807 223894 240859
rect 223946 240847 223952 240859
rect 236272 240847 236278 240859
rect 223946 240819 236278 240847
rect 223946 240807 223952 240819
rect 236272 240807 236278 240819
rect 236330 240807 236336 240859
rect 222544 240733 222550 240785
rect 222602 240773 222608 240785
rect 237232 240773 237238 240785
rect 222602 240745 237238 240773
rect 222602 240733 222608 240745
rect 237232 240733 237238 240745
rect 237290 240733 237296 240785
rect 221680 240659 221686 240711
rect 221738 240699 221744 240711
rect 237442 240699 237470 240893
rect 249232 240881 249238 240893
rect 249290 240881 249296 240933
rect 271504 240881 271510 240933
rect 271562 240921 271568 240933
rect 281680 240921 281686 240933
rect 271562 240893 281686 240921
rect 271562 240881 271568 240893
rect 281680 240881 281686 240893
rect 281738 240881 281744 240933
rect 283888 240881 283894 240933
rect 283946 240921 283952 240933
rect 296656 240921 296662 240933
rect 283946 240893 296662 240921
rect 283946 240881 283952 240893
rect 296656 240881 296662 240893
rect 296714 240881 296720 240933
rect 300898 240921 300926 241189
rect 300994 240995 301022 241633
rect 318832 241621 318838 241673
rect 318890 241661 318896 241673
rect 335536 241661 335542 241673
rect 318890 241633 335542 241661
rect 318890 241621 318896 241633
rect 335536 241621 335542 241633
rect 335594 241621 335600 241673
rect 338128 241621 338134 241673
rect 338186 241661 338192 241673
rect 345922 241661 345950 241707
rect 354544 241695 354550 241707
rect 354602 241695 354608 241747
rect 338186 241633 345950 241661
rect 338186 241621 338192 241633
rect 334576 241547 334582 241599
rect 334634 241587 334640 241599
rect 348112 241587 348118 241599
rect 334634 241559 348118 241587
rect 334634 241547 334640 241559
rect 348112 241547 348118 241559
rect 348170 241547 348176 241599
rect 348208 241547 348214 241599
rect 348266 241587 348272 241599
rect 358384 241587 358390 241599
rect 348266 241559 358390 241587
rect 348266 241547 348272 241559
rect 358384 241547 358390 241559
rect 358442 241547 358448 241599
rect 372610 241587 372638 241855
rect 378544 241843 378550 241895
rect 378602 241883 378608 241895
rect 385648 241883 385654 241895
rect 378602 241855 385654 241883
rect 378602 241843 378608 241855
rect 385648 241843 385654 241855
rect 385706 241843 385712 241895
rect 387280 241843 387286 241895
rect 387338 241843 387344 241895
rect 372688 241769 372694 241821
rect 372746 241809 372752 241821
rect 386128 241809 386134 241821
rect 372746 241781 386134 241809
rect 372746 241769 372752 241781
rect 386128 241769 386134 241781
rect 386186 241769 386192 241821
rect 377872 241695 377878 241747
rect 377930 241735 377936 241747
rect 387184 241735 387190 241747
rect 377930 241707 387190 241735
rect 377930 241695 377936 241707
rect 387184 241695 387190 241707
rect 387242 241695 387248 241747
rect 387280 241695 387286 241747
rect 387338 241735 387344 241747
rect 397840 241735 397846 241747
rect 387338 241707 397846 241735
rect 387338 241695 387344 241707
rect 397840 241695 397846 241707
rect 397898 241695 397904 241747
rect 373072 241621 373078 241673
rect 373130 241661 373136 241673
rect 384784 241661 384790 241673
rect 373130 241633 384790 241661
rect 373130 241621 373136 241633
rect 384784 241621 384790 241633
rect 384842 241621 384848 241673
rect 384880 241621 384886 241673
rect 384938 241661 384944 241673
rect 398992 241661 398998 241673
rect 384938 241633 398998 241661
rect 384938 241621 384944 241633
rect 398992 241621 398998 241633
rect 399050 241621 399056 241673
rect 389776 241587 389782 241599
rect 372610 241559 389782 241587
rect 389776 241547 389782 241559
rect 389834 241547 389840 241599
rect 674128 241547 674134 241599
rect 674186 241587 674192 241599
rect 675472 241587 675478 241599
rect 674186 241559 675478 241587
rect 674186 241547 674192 241559
rect 675472 241547 675478 241559
rect 675530 241547 675536 241599
rect 317872 241473 317878 241525
rect 317930 241513 317936 241525
rect 333808 241513 333814 241525
rect 317930 241485 333814 241513
rect 317930 241473 317936 241485
rect 333808 241473 333814 241485
rect 333866 241473 333872 241525
rect 338032 241473 338038 241525
rect 338090 241513 338096 241525
rect 355120 241513 355126 241525
rect 338090 241485 355126 241513
rect 338090 241473 338096 241485
rect 355120 241473 355126 241485
rect 355178 241473 355184 241525
rect 370480 241473 370486 241525
rect 370538 241513 370544 241525
rect 384976 241513 384982 241525
rect 370538 241485 384982 241513
rect 370538 241473 370544 241485
rect 384976 241473 384982 241485
rect 385034 241473 385040 241525
rect 385648 241473 385654 241525
rect 385706 241513 385712 241525
rect 388240 241513 388246 241525
rect 385706 241485 388246 241513
rect 385706 241473 385712 241485
rect 388240 241473 388246 241485
rect 388298 241473 388304 241525
rect 328528 241399 328534 241451
rect 328586 241439 328592 241451
rect 357136 241439 357142 241451
rect 328586 241411 357142 241439
rect 328586 241399 328592 241411
rect 357136 241399 357142 241411
rect 357194 241399 357200 241451
rect 385936 241439 385942 241451
rect 372130 241411 385942 241439
rect 329872 241325 329878 241377
rect 329930 241365 329936 241377
rect 359344 241365 359350 241377
rect 329930 241337 359350 241365
rect 329930 241325 329936 241337
rect 359344 241325 359350 241337
rect 359402 241325 359408 241377
rect 362800 241325 362806 241377
rect 362858 241365 362864 241377
rect 372130 241365 372158 241411
rect 385936 241399 385942 241411
rect 385994 241399 386000 241451
rect 386128 241399 386134 241451
rect 386186 241439 386192 241451
rect 399568 241439 399574 241451
rect 386186 241411 399574 241439
rect 386186 241399 386192 241411
rect 399568 241399 399574 241411
rect 399626 241399 399632 241451
rect 362858 241337 372158 241365
rect 362858 241325 362864 241337
rect 372208 241325 372214 241377
rect 372266 241365 372272 241377
rect 383536 241365 383542 241377
rect 372266 241337 383542 241365
rect 372266 241325 372272 241337
rect 383536 241325 383542 241337
rect 383594 241325 383600 241377
rect 383632 241325 383638 241377
rect 383690 241365 383696 241377
rect 389392 241365 389398 241377
rect 383690 241337 389398 241365
rect 383690 241325 383696 241337
rect 389392 241325 389398 241337
rect 389450 241325 389456 241377
rect 301168 241251 301174 241303
rect 301226 241291 301232 241303
rect 316624 241291 316630 241303
rect 301226 241263 316630 241291
rect 301226 241251 301232 241263
rect 316624 241251 316630 241263
rect 316682 241251 316688 241303
rect 327568 241251 327574 241303
rect 327626 241291 327632 241303
rect 338128 241291 338134 241303
rect 327626 241263 338134 241291
rect 327626 241251 327632 241263
rect 338128 241251 338134 241263
rect 338186 241251 338192 241303
rect 338512 241251 338518 241303
rect 338570 241291 338576 241303
rect 346384 241291 346390 241303
rect 338570 241263 346390 241291
rect 338570 241251 338576 241263
rect 346384 241251 346390 241263
rect 346442 241251 346448 241303
rect 381424 241251 381430 241303
rect 381482 241291 381488 241303
rect 392560 241291 392566 241303
rect 381482 241263 392566 241291
rect 381482 241251 381488 241263
rect 392560 241251 392566 241263
rect 392618 241251 392624 241303
rect 328048 241177 328054 241229
rect 328106 241217 328112 241229
rect 338032 241217 338038 241229
rect 328106 241189 338038 241217
rect 328106 241177 328112 241189
rect 338032 241177 338038 241189
rect 338090 241177 338096 241229
rect 338608 241177 338614 241229
rect 338666 241217 338672 241229
rect 344272 241217 344278 241229
rect 338666 241189 344278 241217
rect 338666 241177 338672 241189
rect 344272 241177 344278 241189
rect 344330 241177 344336 241229
rect 363184 241217 363190 241229
rect 348514 241189 363190 241217
rect 301072 241103 301078 241155
rect 301130 241143 301136 241155
rect 315472 241143 315478 241155
rect 301130 241115 315478 241143
rect 301130 241103 301136 241115
rect 315472 241103 315478 241115
rect 315530 241103 315536 241155
rect 332080 241103 332086 241155
rect 332138 241143 332144 241155
rect 332138 241115 338942 241143
rect 332138 241103 332144 241115
rect 302512 241029 302518 241081
rect 302570 241069 302576 241081
rect 315952 241069 315958 241081
rect 302570 241041 315958 241069
rect 302570 241029 302576 241041
rect 315952 241029 315958 241041
rect 316010 241029 316016 241081
rect 317776 241029 317782 241081
rect 317834 241069 317840 241081
rect 332944 241069 332950 241081
rect 317834 241041 332950 241069
rect 317834 241029 317840 241041
rect 332944 241029 332950 241041
rect 333002 241029 333008 241081
rect 333058 241041 338846 241069
rect 319216 240995 319222 241007
rect 300994 240967 319222 240995
rect 319216 240955 319222 240967
rect 319274 240955 319280 241007
rect 332464 240955 332470 241007
rect 332522 240995 332528 241007
rect 333058 240995 333086 241041
rect 332522 240967 333086 240995
rect 332522 240955 332528 240967
rect 333712 240955 333718 241007
rect 333770 240995 333776 241007
rect 333770 240967 338750 240995
rect 333770 240955 333776 240967
rect 322000 240921 322006 240933
rect 300898 240893 322006 240921
rect 322000 240881 322006 240893
rect 322058 240881 322064 240933
rect 335056 240881 335062 240933
rect 335114 240921 335120 240933
rect 335114 240893 338654 240921
rect 335114 240881 335120 240893
rect 250384 240847 250390 240859
rect 221738 240671 237470 240699
rect 237538 240819 250390 240847
rect 221738 240659 221744 240671
rect 41776 240585 41782 240637
rect 41834 240585 41840 240637
rect 221104 240585 221110 240637
rect 221162 240625 221168 240637
rect 237538 240625 237566 240819
rect 250384 240807 250390 240819
rect 250442 240807 250448 240859
rect 276880 240807 276886 240859
rect 276938 240847 276944 240859
rect 276938 240819 286046 240847
rect 276938 240807 276944 240819
rect 237616 240733 237622 240785
rect 237674 240773 237680 240785
rect 266032 240773 266038 240785
rect 237674 240745 266038 240773
rect 237674 240733 237680 240745
rect 266032 240733 266038 240745
rect 266090 240733 266096 240785
rect 276400 240773 276406 240785
rect 266818 240745 276406 240773
rect 238960 240659 238966 240711
rect 239018 240699 239024 240711
rect 266704 240699 266710 240711
rect 239018 240671 266710 240699
rect 239018 240659 239024 240671
rect 266704 240659 266710 240671
rect 266762 240659 266768 240711
rect 252496 240625 252502 240637
rect 221162 240597 237566 240625
rect 237634 240597 252502 240625
rect 221162 240585 221168 240597
rect 41794 240415 41822 240585
rect 225520 240511 225526 240563
rect 225578 240551 225584 240563
rect 228880 240551 228886 240563
rect 225578 240523 228886 240551
rect 225578 240511 225584 240523
rect 228880 240511 228886 240523
rect 228938 240511 228944 240563
rect 228976 240511 228982 240563
rect 229034 240551 229040 240563
rect 237424 240551 237430 240563
rect 229034 240523 237430 240551
rect 229034 240511 229040 240523
rect 237424 240511 237430 240523
rect 237482 240511 237488 240563
rect 226096 240437 226102 240489
rect 226154 240477 226160 240489
rect 229936 240477 229942 240489
rect 226154 240449 229942 240477
rect 226154 240437 226160 240449
rect 229936 240437 229942 240449
rect 229994 240437 230000 240489
rect 230032 240437 230038 240489
rect 230090 240477 230096 240489
rect 237328 240477 237334 240489
rect 230090 240449 237334 240477
rect 230090 240437 230096 240449
rect 237328 240437 237334 240449
rect 237386 240437 237392 240489
rect 41776 240363 41782 240415
rect 41834 240363 41840 240415
rect 224272 240363 224278 240415
rect 224330 240403 224336 240415
rect 227536 240403 227542 240415
rect 224330 240375 227542 240403
rect 224330 240363 224336 240375
rect 227536 240363 227542 240375
rect 227594 240363 227600 240415
rect 234352 240329 234358 240341
rect 228226 240301 234358 240329
rect 222064 240215 222070 240267
rect 222122 240255 222128 240267
rect 228226 240255 228254 240301
rect 234352 240289 234358 240301
rect 234410 240289 234416 240341
rect 222122 240227 228254 240255
rect 222122 240215 222128 240227
rect 228304 240215 228310 240267
rect 228362 240255 228368 240267
rect 235600 240255 235606 240267
rect 228362 240227 235606 240255
rect 228362 240215 228368 240227
rect 235600 240215 235606 240227
rect 235658 240215 235664 240267
rect 226864 240141 226870 240193
rect 226922 240181 226928 240193
rect 228496 240181 228502 240193
rect 226922 240153 228502 240181
rect 226922 240141 226928 240153
rect 228496 240141 228502 240153
rect 228554 240141 228560 240193
rect 228688 240141 228694 240193
rect 228746 240181 228752 240193
rect 234448 240181 234454 240193
rect 228746 240153 234454 240181
rect 228746 240141 228752 240153
rect 234448 240141 234454 240153
rect 234506 240141 234512 240193
rect 227920 240067 227926 240119
rect 227978 240107 227984 240119
rect 231760 240107 231766 240119
rect 227978 240079 231766 240107
rect 227978 240067 227984 240079
rect 231760 240067 231766 240079
rect 231818 240067 231824 240119
rect 226960 239993 226966 240045
rect 227018 240033 227024 240045
rect 228976 240033 228982 240045
rect 227018 240005 228982 240033
rect 227018 239993 227024 240005
rect 228976 239993 228982 240005
rect 229034 239993 229040 240045
rect 229072 239993 229078 240045
rect 229130 240033 229136 240045
rect 230800 240033 230806 240045
rect 229130 240005 230806 240033
rect 229130 239993 229136 240005
rect 230800 239993 230806 240005
rect 230858 239993 230864 240045
rect 218128 239919 218134 239971
rect 218186 239959 218192 239971
rect 225136 239959 225142 239971
rect 218186 239931 225142 239959
rect 218186 239919 218192 239931
rect 225136 239919 225142 239931
rect 225194 239919 225200 239971
rect 227344 239919 227350 239971
rect 227402 239959 227408 239971
rect 230032 239959 230038 239971
rect 227402 239931 230038 239959
rect 227402 239919 227408 239931
rect 230032 239919 230038 239931
rect 230090 239919 230096 239971
rect 230128 239919 230134 239971
rect 230186 239959 230192 239971
rect 230512 239959 230518 239971
rect 230186 239931 230518 239959
rect 230186 239919 230192 239931
rect 230512 239919 230518 239931
rect 230570 239919 230576 239971
rect 229552 239845 229558 239897
rect 229610 239885 229616 239897
rect 232240 239885 232246 239897
rect 229610 239857 232246 239885
rect 229610 239845 229616 239857
rect 232240 239845 232246 239857
rect 232298 239845 232304 239897
rect 229072 239771 229078 239823
rect 229130 239811 229136 239823
rect 233584 239811 233590 239823
rect 229130 239783 233590 239811
rect 229130 239771 229136 239783
rect 233584 239771 233590 239783
rect 233642 239771 233648 239823
rect 220240 239697 220246 239749
rect 220298 239737 220304 239749
rect 237634 239737 237662 240597
rect 252496 240585 252502 240597
rect 252554 240585 252560 240637
rect 266818 240625 266846 240745
rect 276400 240733 276406 240745
rect 276458 240733 276464 240785
rect 278512 240733 278518 240785
rect 278570 240773 278576 240785
rect 285904 240773 285910 240785
rect 278570 240745 285910 240773
rect 278570 240733 278576 240745
rect 285904 240733 285910 240745
rect 285962 240733 285968 240785
rect 280048 240659 280054 240711
rect 280106 240699 280112 240711
rect 285808 240699 285814 240711
rect 280106 240671 285814 240699
rect 280106 240659 280112 240671
rect 285808 240659 285814 240671
rect 285866 240659 285872 240711
rect 286018 240699 286046 240819
rect 287344 240807 287350 240859
rect 287402 240847 287408 240859
rect 315280 240847 315286 240859
rect 287402 240819 315286 240847
rect 287402 240807 287408 240819
rect 315280 240807 315286 240819
rect 315338 240807 315344 240859
rect 324496 240807 324502 240859
rect 324554 240847 324560 240859
rect 334576 240847 334582 240859
rect 324554 240819 334582 240847
rect 324554 240807 324560 240819
rect 334576 240807 334582 240819
rect 334634 240807 334640 240859
rect 334672 240807 334678 240859
rect 334730 240847 334736 240859
rect 334730 240819 338510 240847
rect 334730 240807 334736 240819
rect 287824 240733 287830 240785
rect 287882 240773 287888 240785
rect 290800 240773 290806 240785
rect 287882 240745 290806 240773
rect 287882 240733 287888 240745
rect 290800 240733 290806 240745
rect 290858 240733 290864 240785
rect 290992 240733 290998 240785
rect 291050 240773 291056 240785
rect 321424 240773 321430 240785
rect 291050 240745 321430 240773
rect 291050 240733 291056 240745
rect 321424 240733 321430 240745
rect 321482 240733 321488 240785
rect 327856 240773 327862 240785
rect 321634 240745 327862 240773
rect 288304 240699 288310 240711
rect 286018 240671 288310 240699
rect 288304 240659 288310 240671
rect 288362 240659 288368 240711
rect 289552 240659 289558 240711
rect 289610 240699 289616 240711
rect 289610 240671 299966 240699
rect 289610 240659 289616 240671
rect 252610 240597 266846 240625
rect 237904 240511 237910 240563
rect 237962 240551 237968 240563
rect 243280 240551 243286 240563
rect 237962 240523 243286 240551
rect 237962 240511 237968 240523
rect 243280 240511 243286 240523
rect 243338 240511 243344 240563
rect 244528 240511 244534 240563
rect 244586 240551 244592 240563
rect 252610 240551 252638 240597
rect 273232 240585 273238 240637
rect 273290 240625 273296 240637
rect 284656 240625 284662 240637
rect 273290 240597 284662 240625
rect 273290 240585 273296 240597
rect 284656 240585 284662 240597
rect 284714 240585 284720 240637
rect 286384 240585 286390 240637
rect 286442 240625 286448 240637
rect 299824 240625 299830 240637
rect 286442 240597 299830 240625
rect 286442 240585 286448 240597
rect 299824 240585 299830 240597
rect 299882 240585 299888 240637
rect 244586 240523 252638 240551
rect 244586 240511 244592 240523
rect 273328 240511 273334 240563
rect 273386 240551 273392 240563
rect 281584 240551 281590 240563
rect 273386 240523 281590 240551
rect 273386 240511 273392 240523
rect 281584 240511 281590 240523
rect 281642 240511 281648 240563
rect 281680 240511 281686 240563
rect 281738 240551 281744 240563
rect 285712 240551 285718 240563
rect 281738 240523 285718 240551
rect 281738 240511 281744 240523
rect 285712 240511 285718 240523
rect 285770 240511 285776 240563
rect 289264 240511 289270 240563
rect 289322 240551 289328 240563
rect 295312 240551 295318 240563
rect 289322 240523 295318 240551
rect 289322 240511 289328 240523
rect 295312 240511 295318 240523
rect 295370 240511 295376 240563
rect 299938 240551 299966 240671
rect 300016 240659 300022 240711
rect 300074 240699 300080 240711
rect 318352 240699 318358 240711
rect 300074 240671 318358 240699
rect 300074 240659 300080 240671
rect 318352 240659 318358 240671
rect 318410 240659 318416 240711
rect 315664 240585 315670 240637
rect 315722 240625 315728 240637
rect 321634 240625 321662 240745
rect 327856 240733 327862 240745
rect 327914 240733 327920 240785
rect 328240 240733 328246 240785
rect 328298 240773 328304 240785
rect 338128 240773 338134 240785
rect 328298 240745 338134 240773
rect 328298 240733 328304 240745
rect 338128 240733 338134 240745
rect 338186 240733 338192 240785
rect 326704 240659 326710 240711
rect 326762 240699 326768 240711
rect 338224 240699 338230 240711
rect 326762 240671 338230 240699
rect 326762 240659 326768 240671
rect 338224 240659 338230 240671
rect 338282 240659 338288 240711
rect 315722 240597 321662 240625
rect 315722 240585 315728 240597
rect 323632 240585 323638 240637
rect 323690 240625 323696 240637
rect 337072 240625 337078 240637
rect 323690 240597 337078 240625
rect 323690 240585 323696 240597
rect 337072 240585 337078 240597
rect 337130 240585 337136 240637
rect 338482 240625 338510 240819
rect 338626 240773 338654 240893
rect 338722 240847 338750 240967
rect 338818 240921 338846 241041
rect 338914 240995 338942 241115
rect 338992 241029 338998 241081
rect 339050 241069 339056 241081
rect 348514 241069 348542 241189
rect 363184 241177 363190 241189
rect 363242 241177 363248 241229
rect 373456 241177 373462 241229
rect 373514 241217 373520 241229
rect 384688 241217 384694 241229
rect 373514 241189 384694 241217
rect 373514 241177 373520 241189
rect 384688 241177 384694 241189
rect 384746 241177 384752 241229
rect 384784 241177 384790 241229
rect 384842 241217 384848 241229
rect 400720 241217 400726 241229
rect 384842 241189 400726 241217
rect 384842 241177 384848 241189
rect 400720 241177 400726 241189
rect 400778 241177 400784 241229
rect 374896 241103 374902 241155
rect 374954 241143 374960 241155
rect 403984 241143 403990 241155
rect 374954 241115 403990 241143
rect 374954 241103 374960 241115
rect 403984 241103 403990 241115
rect 404042 241103 404048 241155
rect 339050 241041 348542 241069
rect 339050 241029 339056 241041
rect 359824 241029 359830 241081
rect 359882 241069 359888 241081
rect 384496 241069 384502 241081
rect 359882 241041 384502 241069
rect 359882 241029 359888 241041
rect 384496 241029 384502 241041
rect 384554 241029 384560 241081
rect 406000 241069 406006 241081
rect 384610 241041 406006 241069
rect 363952 240995 363958 241007
rect 338914 240967 363958 240995
rect 363952 240955 363958 240967
rect 364010 240955 364016 241007
rect 375664 240955 375670 241007
rect 375722 240995 375728 241007
rect 384610 240995 384638 241041
rect 406000 241029 406006 241041
rect 406058 241029 406064 241081
rect 375722 240967 384638 240995
rect 375722 240955 375728 240967
rect 384688 240955 384694 241007
rect 384746 240995 384752 241007
rect 401584 240995 401590 241007
rect 384746 240967 401590 240995
rect 384746 240955 384752 240967
rect 401584 240955 401590 240967
rect 401642 240955 401648 241007
rect 364720 240921 364726 240933
rect 338818 240893 364726 240921
rect 364720 240881 364726 240893
rect 364778 240881 364784 240933
rect 374032 240881 374038 240933
rect 374090 240921 374096 240933
rect 402256 240921 402262 240933
rect 374090 240893 402262 240921
rect 374090 240881 374096 240893
rect 402256 240881 402262 240893
rect 402314 240881 402320 240933
rect 367984 240847 367990 240859
rect 338722 240819 367990 240847
rect 367984 240807 367990 240819
rect 368042 240807 368048 240859
rect 384112 240807 384118 240859
rect 384170 240847 384176 240859
rect 414256 240847 414262 240859
rect 384170 240819 414262 240847
rect 384170 240807 384176 240819
rect 414256 240807 414262 240819
rect 414314 240807 414320 240859
rect 370672 240773 370678 240785
rect 338626 240745 370678 240773
rect 370672 240733 370678 240745
rect 370730 240733 370736 240785
rect 375280 240733 375286 240785
rect 375338 240773 375344 240785
rect 405040 240773 405046 240785
rect 375338 240745 405046 240773
rect 375338 240733 375344 240745
rect 405040 240733 405046 240745
rect 405098 240733 405104 240785
rect 338608 240659 338614 240711
rect 338666 240699 338672 240711
rect 366928 240699 366934 240711
rect 338666 240671 366934 240699
rect 338666 240659 338672 240671
rect 366928 240659 366934 240671
rect 366986 240659 366992 240711
rect 372592 240659 372598 240711
rect 372650 240699 372656 240711
rect 384208 240699 384214 240711
rect 372650 240671 384214 240699
rect 372650 240659 372656 240671
rect 384208 240659 384214 240671
rect 384266 240659 384272 240711
rect 384304 240659 384310 240711
rect 384362 240699 384368 240711
rect 414640 240699 414646 240711
rect 384362 240671 414646 240699
rect 384362 240659 384368 240671
rect 414640 240659 414646 240671
rect 414698 240659 414704 240711
rect 369712 240625 369718 240637
rect 338482 240597 369718 240625
rect 369712 240585 369718 240597
rect 369770 240585 369776 240637
rect 376624 240585 376630 240637
rect 376682 240625 376688 240637
rect 407728 240625 407734 240637
rect 376682 240597 407734 240625
rect 376682 240585 376688 240597
rect 407728 240585 407734 240597
rect 407786 240585 407792 240637
rect 317488 240551 317494 240563
rect 299938 240523 317494 240551
rect 317488 240511 317494 240523
rect 317546 240511 317552 240563
rect 319216 240511 319222 240563
rect 319274 240551 319280 240563
rect 327760 240551 327766 240563
rect 319274 240523 327766 240551
rect 319274 240511 319280 240523
rect 327760 240511 327766 240523
rect 327818 240511 327824 240563
rect 327856 240511 327862 240563
rect 327914 240551 327920 240563
rect 332272 240551 332278 240563
rect 327914 240523 332278 240551
rect 327914 240511 327920 240523
rect 332272 240511 332278 240523
rect 332330 240511 332336 240563
rect 332848 240511 332854 240563
rect 332906 240551 332912 240563
rect 365872 240551 365878 240563
rect 332906 240523 365878 240551
rect 332906 240511 332912 240523
rect 365872 240511 365878 240523
rect 365930 240511 365936 240563
rect 374320 240511 374326 240563
rect 374378 240551 374384 240563
rect 403312 240551 403318 240563
rect 374378 240523 403318 240551
rect 374378 240511 374384 240523
rect 403312 240511 403318 240523
rect 403370 240511 403376 240563
rect 674800 240511 674806 240563
rect 674858 240551 674864 240563
rect 675472 240551 675478 240563
rect 674858 240523 675478 240551
rect 674858 240511 674864 240523
rect 675472 240511 675478 240523
rect 675530 240511 675536 240563
rect 238000 240437 238006 240489
rect 238058 240477 238064 240489
rect 240496 240477 240502 240489
rect 238058 240449 240502 240477
rect 238058 240437 238064 240449
rect 240496 240437 240502 240449
rect 240554 240437 240560 240489
rect 276784 240437 276790 240489
rect 276842 240477 276848 240489
rect 280336 240477 280342 240489
rect 276842 240449 280342 240477
rect 276842 240437 276848 240449
rect 280336 240437 280342 240449
rect 280394 240437 280400 240489
rect 280432 240437 280438 240489
rect 280490 240477 280496 240489
rect 295408 240477 295414 240489
rect 280490 240449 295414 240477
rect 280490 240437 280496 240449
rect 295408 240437 295414 240449
rect 295466 240437 295472 240489
rect 324112 240437 324118 240489
rect 324170 240477 324176 240489
rect 334192 240477 334198 240489
rect 324170 240449 334198 240477
rect 324170 240437 324176 240449
rect 334192 240437 334198 240449
rect 334250 240437 334256 240489
rect 334288 240437 334294 240489
rect 334346 240477 334352 240489
rect 368752 240477 368758 240489
rect 334346 240449 368758 240477
rect 334346 240437 334352 240449
rect 368752 240437 368758 240449
rect 368810 240437 368816 240489
rect 376240 240437 376246 240489
rect 376298 240477 376304 240489
rect 406576 240477 406582 240489
rect 376298 240449 406582 240477
rect 376298 240437 376304 240449
rect 406576 240437 406582 240449
rect 406634 240437 406640 240489
rect 549040 240437 549046 240489
rect 549098 240477 549104 240489
rect 650896 240477 650902 240489
rect 549098 240449 650902 240477
rect 549098 240437 549104 240449
rect 650896 240437 650902 240449
rect 650954 240437 650960 240489
rect 279088 240363 279094 240415
rect 279146 240403 279152 240415
rect 294448 240403 294454 240415
rect 279146 240375 294454 240403
rect 279146 240363 279152 240375
rect 294448 240363 294454 240375
rect 294506 240363 294512 240415
rect 321424 240363 321430 240415
rect 321482 240403 321488 240415
rect 327664 240403 327670 240415
rect 321482 240375 327670 240403
rect 321482 240363 321488 240375
rect 327664 240363 327670 240375
rect 327722 240363 327728 240415
rect 327760 240363 327766 240415
rect 327818 240403 327824 240415
rect 336016 240403 336022 240415
rect 327818 240375 336022 240403
rect 327818 240363 327824 240375
rect 336016 240363 336022 240375
rect 336074 240363 336080 240415
rect 338128 240363 338134 240415
rect 338186 240403 338192 240415
rect 356272 240403 356278 240415
rect 338186 240375 356278 240403
rect 338186 240363 338192 240375
rect 356272 240363 356278 240375
rect 356330 240363 356336 240415
rect 370000 240363 370006 240415
rect 370058 240403 370064 240415
rect 386608 240403 386614 240415
rect 370058 240375 386614 240403
rect 370058 240363 370064 240375
rect 386608 240363 386614 240375
rect 386666 240363 386672 240415
rect 275536 240289 275542 240341
rect 275594 240329 275600 240341
rect 275594 240301 285758 240329
rect 275594 240289 275600 240301
rect 240112 240215 240118 240267
rect 240170 240255 240176 240267
rect 260176 240255 260182 240267
rect 240170 240227 260182 240255
rect 240170 240215 240176 240227
rect 260176 240215 260182 240227
rect 260234 240215 260240 240267
rect 277744 240215 277750 240267
rect 277802 240255 277808 240267
rect 285616 240255 285622 240267
rect 277802 240227 285622 240255
rect 277802 240215 277808 240227
rect 285616 240215 285622 240227
rect 285674 240215 285680 240267
rect 278512 240141 278518 240193
rect 278570 240181 278576 240193
rect 284368 240181 284374 240193
rect 278570 240153 284374 240181
rect 278570 240141 278576 240153
rect 284368 240141 284374 240153
rect 284426 240141 284432 240193
rect 279088 240067 279094 240119
rect 279146 240107 279152 240119
rect 283504 240107 283510 240119
rect 279146 240079 283510 240107
rect 279146 240067 279152 240079
rect 283504 240067 283510 240079
rect 283562 240067 283568 240119
rect 272464 239993 272470 240045
rect 272522 240033 272528 240045
rect 273616 240033 273622 240045
rect 272522 240005 273622 240033
rect 272522 239993 272528 240005
rect 273616 239993 273622 240005
rect 273674 239993 273680 240045
rect 278992 239993 278998 240045
rect 279050 240033 279056 240045
rect 280816 240033 280822 240045
rect 279050 240005 280822 240033
rect 279050 239993 279056 240005
rect 280816 239993 280822 240005
rect 280874 239993 280880 240045
rect 273040 239919 273046 239971
rect 273098 239959 273104 239971
rect 276304 239959 276310 239971
rect 273098 239931 276310 239959
rect 273098 239919 273104 239931
rect 276304 239919 276310 239931
rect 276362 239919 276368 239971
rect 279856 239919 279862 239971
rect 279914 239959 279920 239971
rect 280624 239959 280630 239971
rect 279914 239931 280630 239959
rect 279914 239919 279920 239931
rect 280624 239919 280630 239931
rect 280682 239919 280688 239971
rect 268432 239845 268438 239897
rect 268490 239885 268496 239897
rect 274768 239885 274774 239897
rect 268490 239857 274774 239885
rect 268490 239845 268496 239857
rect 274768 239845 274774 239857
rect 274826 239845 274832 239897
rect 279280 239845 279286 239897
rect 279338 239885 279344 239897
rect 282352 239885 282358 239897
rect 279338 239857 282358 239885
rect 279338 239845 279344 239857
rect 282352 239845 282358 239857
rect 282410 239845 282416 239897
rect 285730 239885 285758 240301
rect 286192 240289 286198 240341
rect 286250 240329 286256 240341
rect 288496 240329 288502 240341
rect 286250 240301 288502 240329
rect 286250 240289 286256 240301
rect 288496 240289 288502 240301
rect 288554 240289 288560 240341
rect 288592 240289 288598 240341
rect 288650 240329 288656 240341
rect 294064 240329 294070 240341
rect 288650 240301 294070 240329
rect 288650 240289 288656 240301
rect 294064 240289 294070 240301
rect 294122 240289 294128 240341
rect 302320 240289 302326 240341
rect 302378 240289 302384 240341
rect 326224 240289 326230 240341
rect 326282 240329 326288 240341
rect 326282 240301 338750 240329
rect 326282 240289 326288 240301
rect 302338 240255 302366 240289
rect 302512 240255 302518 240267
rect 302338 240227 302518 240255
rect 302512 240215 302518 240227
rect 302570 240215 302576 240267
rect 324880 240215 324886 240267
rect 324938 240255 324944 240267
rect 329008 240255 329014 240267
rect 324938 240227 329014 240255
rect 324938 240215 324944 240227
rect 329008 240215 329014 240227
rect 329066 240215 329072 240267
rect 329200 240215 329206 240267
rect 329258 240255 329264 240267
rect 329776 240255 329782 240267
rect 329258 240227 329782 240255
rect 329258 240215 329264 240227
rect 329776 240215 329782 240227
rect 329834 240215 329840 240267
rect 333328 240215 333334 240267
rect 333386 240255 333392 240267
rect 338608 240255 338614 240267
rect 333386 240227 338614 240255
rect 333386 240215 333392 240227
rect 338608 240215 338614 240227
rect 338666 240215 338672 240267
rect 338722 240255 338750 240301
rect 342736 240289 342742 240341
rect 342794 240329 342800 240341
rect 343120 240329 343126 240341
rect 342794 240301 343126 240329
rect 342794 240289 342800 240301
rect 343120 240289 343126 240301
rect 343178 240289 343184 240341
rect 381520 240289 381526 240341
rect 381578 240329 381584 240341
rect 393712 240329 393718 240341
rect 381578 240301 393718 240329
rect 381578 240289 381584 240301
rect 393712 240289 393718 240301
rect 393770 240289 393776 240341
rect 342832 240255 342838 240267
rect 338722 240227 342838 240255
rect 342832 240215 342838 240227
rect 342890 240215 342896 240267
rect 381904 240215 381910 240267
rect 381962 240255 381968 240267
rect 394576 240255 394582 240267
rect 381962 240227 394582 240255
rect 381962 240215 381968 240227
rect 394576 240215 394582 240227
rect 394634 240215 394640 240267
rect 285904 240141 285910 240193
rect 285962 240181 285968 240193
rect 288592 240181 288598 240193
rect 285962 240153 288598 240181
rect 285962 240141 285968 240153
rect 288592 240141 288598 240153
rect 288650 240141 288656 240193
rect 288688 240141 288694 240193
rect 288746 240181 288752 240193
rect 298864 240181 298870 240193
rect 288746 240153 298870 240181
rect 288746 240141 288752 240153
rect 298864 240141 298870 240153
rect 298922 240141 298928 240193
rect 298960 240141 298966 240193
rect 299018 240181 299024 240193
rect 302416 240181 302422 240193
rect 299018 240153 302422 240181
rect 299018 240141 299024 240153
rect 302416 240141 302422 240153
rect 302474 240141 302480 240193
rect 325840 240141 325846 240193
rect 325898 240181 325904 240193
rect 325898 240153 338462 240181
rect 325898 240141 325904 240153
rect 286000 240067 286006 240119
rect 286058 240107 286064 240119
rect 286058 240079 291998 240107
rect 286058 240067 286064 240079
rect 286288 239993 286294 240045
rect 286346 240033 286352 240045
rect 291856 240033 291862 240045
rect 286346 240005 291862 240033
rect 286346 239993 286352 240005
rect 291856 239993 291862 240005
rect 291914 239993 291920 240045
rect 291970 240033 291998 240079
rect 292048 240067 292054 240119
rect 292106 240107 292112 240119
rect 300592 240107 300598 240119
rect 292106 240079 300598 240107
rect 292106 240067 292112 240079
rect 300592 240067 300598 240079
rect 300650 240067 300656 240119
rect 300688 240067 300694 240119
rect 300746 240107 300752 240119
rect 304624 240107 304630 240119
rect 300746 240079 304630 240107
rect 300746 240067 300752 240079
rect 304624 240067 304630 240079
rect 304682 240067 304688 240119
rect 324016 240067 324022 240119
rect 324074 240107 324080 240119
rect 331312 240107 331318 240119
rect 324074 240079 331318 240107
rect 324074 240067 324080 240079
rect 331312 240067 331318 240079
rect 331370 240067 331376 240119
rect 338224 240107 338230 240119
rect 331426 240079 338230 240107
rect 293968 240033 293974 240045
rect 291970 240005 293974 240033
rect 293968 239993 293974 240005
rect 294026 239993 294032 240045
rect 295888 239993 295894 240045
rect 295946 240033 295952 240045
rect 302512 240033 302518 240045
rect 295946 240005 302518 240033
rect 295946 239993 295952 240005
rect 302512 239993 302518 240005
rect 302570 239993 302576 240045
rect 303568 239993 303574 240045
rect 303626 240033 303632 240045
rect 305872 240033 305878 240045
rect 303626 240005 305878 240033
rect 303626 239993 303632 240005
rect 305872 239993 305878 240005
rect 305930 239993 305936 240045
rect 310864 239993 310870 240045
rect 310922 240033 310928 240045
rect 313936 240033 313942 240045
rect 310922 240005 313942 240033
rect 310922 239993 310928 240005
rect 313936 239993 313942 240005
rect 313994 239993 314000 240045
rect 323248 239993 323254 240045
rect 323306 240033 323312 240045
rect 331426 240033 331454 240079
rect 338224 240067 338230 240079
rect 338282 240067 338288 240119
rect 338434 240107 338462 240153
rect 338512 240141 338518 240193
rect 338570 240181 338576 240193
rect 338570 240153 342782 240181
rect 338570 240141 338576 240153
rect 342754 240107 342782 240153
rect 366832 240141 366838 240193
rect 366890 240181 366896 240193
rect 377872 240181 377878 240193
rect 366890 240153 377878 240181
rect 366890 240141 366896 240153
rect 377872 240141 377878 240153
rect 377930 240141 377936 240193
rect 380080 240141 380086 240193
rect 380138 240181 380144 240193
rect 390256 240181 390262 240193
rect 380138 240153 390262 240181
rect 380138 240141 380144 240153
rect 390256 240141 390262 240153
rect 390314 240141 390320 240193
rect 344656 240107 344662 240119
rect 338434 240079 339134 240107
rect 342754 240079 344662 240107
rect 323306 240005 331454 240033
rect 323306 239993 323312 240005
rect 331504 239993 331510 240045
rect 331562 240033 331568 240045
rect 338992 240033 338998 240045
rect 331562 240005 338998 240033
rect 331562 239993 331568 240005
rect 338992 239993 338998 240005
rect 339050 239993 339056 240045
rect 339106 240033 339134 240079
rect 344656 240067 344662 240079
rect 344714 240067 344720 240119
rect 368176 240067 368182 240119
rect 368234 240107 368240 240119
rect 378544 240107 378550 240119
rect 368234 240079 378550 240107
rect 368234 240067 368240 240079
rect 378544 240067 378550 240079
rect 378602 240067 378608 240119
rect 378832 240067 378838 240119
rect 378890 240107 378896 240119
rect 387664 240107 387670 240119
rect 378890 240079 387670 240107
rect 378890 240067 378896 240079
rect 387664 240067 387670 240079
rect 387722 240067 387728 240119
rect 388720 240067 388726 240119
rect 388778 240107 388784 240119
rect 396304 240107 396310 240119
rect 388778 240079 396310 240107
rect 388778 240067 388784 240079
rect 396304 240067 396310 240079
rect 396362 240067 396368 240119
rect 342736 240033 342742 240045
rect 339106 240005 342742 240033
rect 342736 239993 342742 240005
rect 342794 239993 342800 240045
rect 382864 239993 382870 240045
rect 382922 240033 382928 240045
rect 386512 240033 386518 240045
rect 382922 240005 386518 240033
rect 382922 239993 382928 240005
rect 386512 239993 386518 240005
rect 386570 239993 386576 240045
rect 386608 239993 386614 240045
rect 386666 240033 386672 240045
rect 393040 240033 393046 240045
rect 386666 240005 393046 240033
rect 386666 239993 386672 240005
rect 393040 239993 393046 240005
rect 393098 239993 393104 240045
rect 285808 239919 285814 239971
rect 285866 239959 285872 239971
rect 294928 239959 294934 239971
rect 285866 239931 294934 239959
rect 285866 239919 285872 239931
rect 294928 239919 294934 239931
rect 294986 239919 294992 239971
rect 296560 239919 296566 239971
rect 296618 239959 296624 239971
rect 302800 239959 302806 239971
rect 296618 239931 302806 239959
rect 296618 239919 296624 239931
rect 302800 239919 302806 239931
rect 302858 239919 302864 239971
rect 302896 239919 302902 239971
rect 302954 239959 302960 239971
rect 305488 239959 305494 239971
rect 302954 239931 305494 239959
rect 302954 239919 302960 239931
rect 305488 239919 305494 239931
rect 305546 239919 305552 239971
rect 309328 239919 309334 239971
rect 309386 239959 309392 239971
rect 309808 239959 309814 239971
rect 309386 239931 309814 239959
rect 309386 239919 309392 239931
rect 309808 239919 309814 239931
rect 309866 239919 309872 239971
rect 310000 239919 310006 239971
rect 310058 239959 310064 239971
rect 311152 239959 311158 239971
rect 310058 239931 311158 239959
rect 310058 239919 310064 239931
rect 311152 239919 311158 239931
rect 311210 239919 311216 239971
rect 311632 239919 311638 239971
rect 311690 239959 311696 239971
rect 327472 239959 327478 239971
rect 311690 239931 327478 239959
rect 311690 239919 311696 239931
rect 327472 239919 327478 239931
rect 327530 239919 327536 239971
rect 330928 239959 330934 239971
rect 327586 239931 330934 239959
rect 290416 239885 290422 239897
rect 285730 239857 290422 239885
rect 290416 239845 290422 239857
rect 290474 239845 290480 239897
rect 290512 239845 290518 239897
rect 290570 239885 290576 239897
rect 292240 239885 292246 239897
rect 290570 239857 292246 239885
rect 290570 239845 290576 239857
rect 292240 239845 292246 239857
rect 292298 239845 292304 239897
rect 292624 239845 292630 239897
rect 292682 239885 292688 239897
rect 300688 239885 300694 239897
rect 292682 239857 300694 239885
rect 292682 239845 292688 239857
rect 300688 239845 300694 239857
rect 300746 239845 300752 239897
rect 301360 239845 301366 239897
rect 301418 239885 301424 239897
rect 305008 239885 305014 239897
rect 301418 239857 305014 239885
rect 301418 239845 301424 239857
rect 305008 239845 305014 239857
rect 305066 239845 305072 239897
rect 321904 239845 321910 239897
rect 321962 239885 321968 239897
rect 327586 239885 327614 239931
rect 330928 239919 330934 239931
rect 330986 239919 330992 239971
rect 331120 239919 331126 239971
rect 331178 239959 331184 239971
rect 332944 239959 332950 239971
rect 331178 239931 332950 239959
rect 331178 239919 331184 239931
rect 332944 239919 332950 239931
rect 333002 239919 333008 239971
rect 334192 239919 334198 239971
rect 334250 239959 334256 239971
rect 347536 239959 347542 239971
rect 334250 239931 347542 239959
rect 334250 239919 334256 239931
rect 347536 239919 347542 239931
rect 347594 239919 347600 239971
rect 382288 239919 382294 239971
rect 382346 239959 382352 239971
rect 385456 239959 385462 239971
rect 382346 239931 385462 239959
rect 382346 239919 382352 239931
rect 385456 239919 385462 239931
rect 385514 239919 385520 239971
rect 321962 239857 327614 239885
rect 321962 239845 321968 239857
rect 327664 239845 327670 239897
rect 327722 239885 327728 239897
rect 341008 239885 341014 239897
rect 327722 239857 341014 239885
rect 327722 239845 327728 239857
rect 341008 239845 341014 239857
rect 341066 239845 341072 239897
rect 382960 239845 382966 239897
rect 383018 239885 383024 239897
rect 388048 239885 388054 239897
rect 383018 239857 388054 239885
rect 383018 239845 383024 239857
rect 388048 239845 388054 239857
rect 388106 239845 388112 239897
rect 279856 239771 279862 239823
rect 279914 239811 279920 239823
rect 281488 239811 281494 239823
rect 279914 239783 281494 239811
rect 279914 239771 279920 239783
rect 281488 239771 281494 239783
rect 281546 239771 281552 239823
rect 281584 239771 281590 239823
rect 281642 239811 281648 239823
rect 289264 239811 289270 239823
rect 281642 239783 289270 239811
rect 281642 239771 281648 239783
rect 289264 239771 289270 239783
rect 289322 239771 289328 239823
rect 289360 239771 289366 239823
rect 289418 239811 289424 239823
rect 299248 239811 299254 239823
rect 289418 239783 299254 239811
rect 289418 239771 289424 239783
rect 299248 239771 299254 239783
rect 299306 239771 299312 239823
rect 299632 239771 299638 239823
rect 299690 239811 299696 239823
rect 304240 239811 304246 239823
rect 299690 239783 304246 239811
rect 299690 239771 299696 239783
rect 304240 239771 304246 239783
rect 304298 239771 304304 239823
rect 311248 239771 311254 239823
rect 311306 239811 311312 239823
rect 314896 239811 314902 239823
rect 311306 239783 314902 239811
rect 311306 239771 311312 239783
rect 314896 239771 314902 239783
rect 314954 239771 314960 239823
rect 322288 239771 322294 239823
rect 322346 239811 322352 239823
rect 329104 239811 329110 239823
rect 322346 239783 329110 239811
rect 322346 239771 322352 239783
rect 329104 239771 329110 239783
rect 329162 239771 329168 239823
rect 329296 239771 329302 239823
rect 329354 239811 329360 239823
rect 348208 239811 348214 239823
rect 329354 239783 348214 239811
rect 329354 239771 329360 239783
rect 348208 239771 348214 239783
rect 348266 239771 348272 239823
rect 371248 239771 371254 239823
rect 371306 239811 371312 239823
rect 388720 239811 388726 239823
rect 371306 239783 388726 239811
rect 371306 239771 371312 239783
rect 388720 239771 388726 239783
rect 388778 239771 388784 239823
rect 277552 239737 277558 239749
rect 220298 239709 237662 239737
rect 262114 239709 277558 239737
rect 220298 239697 220304 239709
rect 222064 239623 222070 239675
rect 222122 239663 222128 239675
rect 236656 239663 236662 239675
rect 222122 239635 236662 239663
rect 222122 239623 222128 239635
rect 236656 239623 236662 239635
rect 236714 239623 236720 239675
rect 236752 239623 236758 239675
rect 236810 239663 236816 239675
rect 247408 239663 247414 239675
rect 236810 239635 247414 239663
rect 236810 239623 236816 239635
rect 247408 239623 247414 239635
rect 247466 239623 247472 239675
rect 224752 239549 224758 239601
rect 224810 239589 224816 239601
rect 242512 239589 242518 239601
rect 224810 239561 242518 239589
rect 224810 239549 224816 239561
rect 242512 239549 242518 239561
rect 242570 239549 242576 239601
rect 243760 239549 243766 239601
rect 243818 239589 243824 239601
rect 262114 239589 262142 239709
rect 277552 239697 277558 239709
rect 277610 239697 277616 239749
rect 278128 239697 278134 239749
rect 278186 239737 278192 239749
rect 284560 239737 284566 239749
rect 278186 239709 284566 239737
rect 278186 239697 278192 239709
rect 284560 239697 284566 239709
rect 284618 239697 284624 239749
rect 284656 239697 284662 239749
rect 284714 239737 284720 239749
rect 290800 239737 290806 239749
rect 284714 239709 290806 239737
rect 284714 239697 284720 239709
rect 290800 239697 290806 239709
rect 290858 239697 290864 239749
rect 290896 239697 290902 239749
rect 290954 239737 290960 239749
rect 300208 239737 300214 239749
rect 290954 239709 300214 239737
rect 290954 239697 290960 239709
rect 300208 239697 300214 239709
rect 300266 239697 300272 239749
rect 321808 239697 321814 239749
rect 321866 239737 321872 239749
rect 321866 239709 329150 239737
rect 321866 239697 321872 239709
rect 276208 239623 276214 239675
rect 276266 239663 276272 239675
rect 285232 239663 285238 239675
rect 276266 239635 285238 239663
rect 276266 239623 276272 239635
rect 285232 239623 285238 239635
rect 285290 239623 285296 239675
rect 296176 239663 296182 239675
rect 287266 239635 296182 239663
rect 243818 239561 262142 239589
rect 243818 239549 243824 239561
rect 277264 239549 277270 239601
rect 277322 239589 277328 239601
rect 287152 239589 287158 239601
rect 277322 239561 287158 239589
rect 277322 239549 277328 239561
rect 287152 239549 287158 239561
rect 287210 239549 287216 239601
rect 223792 239475 223798 239527
rect 223850 239515 223856 239527
rect 233584 239515 233590 239527
rect 223850 239487 233590 239515
rect 223850 239475 223856 239487
rect 233584 239475 233590 239487
rect 233642 239475 233648 239527
rect 246448 239515 246454 239527
rect 233698 239487 246454 239515
rect 233698 239441 233726 239487
rect 246448 239475 246454 239487
rect 246506 239475 246512 239527
rect 276976 239475 276982 239527
rect 277034 239515 277040 239527
rect 281584 239515 281590 239527
rect 277034 239487 281590 239515
rect 277034 239475 277040 239487
rect 281584 239475 281590 239487
rect 281642 239475 281648 239527
rect 282160 239475 282166 239527
rect 282218 239515 282224 239527
rect 287266 239515 287294 239635
rect 296176 239623 296182 239635
rect 296234 239623 296240 239675
rect 297424 239623 297430 239675
rect 297482 239663 297488 239675
rect 302896 239663 302902 239675
rect 297482 239635 302902 239663
rect 297482 239623 297488 239635
rect 302896 239623 302902 239635
rect 302954 239623 302960 239675
rect 305200 239623 305206 239675
rect 305258 239663 305264 239675
rect 306640 239663 306646 239675
rect 305258 239635 306646 239663
rect 305258 239623 305264 239635
rect 306640 239623 306646 239635
rect 306698 239623 306704 239675
rect 310768 239623 310774 239675
rect 310826 239663 310832 239675
rect 313168 239663 313174 239675
rect 310826 239635 313174 239663
rect 310826 239623 310832 239635
rect 313168 239623 313174 239635
rect 313226 239623 313232 239675
rect 321040 239623 321046 239675
rect 321098 239663 321104 239675
rect 328336 239663 328342 239675
rect 321098 239635 328342 239663
rect 321098 239623 321104 239635
rect 328336 239623 328342 239635
rect 328394 239623 328400 239675
rect 329122 239663 329150 239709
rect 330928 239697 330934 239749
rect 330986 239737 330992 239749
rect 343120 239737 343126 239749
rect 330986 239709 343126 239737
rect 330986 239697 330992 239709
rect 343120 239697 343126 239709
rect 343178 239697 343184 239749
rect 374800 239697 374806 239749
rect 374858 239737 374864 239749
rect 386032 239737 386038 239749
rect 374858 239709 386038 239737
rect 374858 239697 374864 239709
rect 386032 239697 386038 239709
rect 386090 239697 386096 239749
rect 341872 239663 341878 239675
rect 329122 239635 341878 239663
rect 341872 239623 341878 239635
rect 341930 239623 341936 239675
rect 370864 239623 370870 239675
rect 370922 239663 370928 239675
rect 383056 239663 383062 239675
rect 370922 239635 383062 239663
rect 370922 239623 370928 239635
rect 383056 239623 383062 239635
rect 383114 239623 383120 239675
rect 288688 239549 288694 239601
rect 288746 239589 288752 239601
rect 288746 239561 291854 239589
rect 288746 239549 288752 239561
rect 291664 239515 291670 239527
rect 282218 239487 287294 239515
rect 287362 239487 291670 239515
rect 282218 239475 282224 239487
rect 229762 239413 233726 239441
rect 222928 239253 222934 239305
rect 222986 239293 222992 239305
rect 229762 239293 229790 239413
rect 280432 239401 280438 239453
rect 280490 239441 280496 239453
rect 287362 239441 287390 239487
rect 291664 239475 291670 239487
rect 291722 239475 291728 239527
rect 291826 239515 291854 239561
rect 291952 239549 291958 239601
rect 292010 239589 292016 239601
rect 297040 239589 297046 239601
rect 292010 239561 297046 239589
rect 292010 239549 292016 239561
rect 297040 239549 297046 239561
rect 297098 239549 297104 239601
rect 301072 239589 301078 239601
rect 297154 239561 301078 239589
rect 297154 239515 297182 239561
rect 301072 239549 301078 239561
rect 301130 239549 301136 239601
rect 320080 239549 320086 239601
rect 320138 239589 320144 239601
rect 338800 239589 338806 239601
rect 320138 239561 338806 239589
rect 320138 239549 320144 239561
rect 338800 239549 338806 239561
rect 338858 239549 338864 239601
rect 380656 239549 380662 239601
rect 380714 239589 380720 239601
rect 390928 239589 390934 239601
rect 380714 239561 390934 239589
rect 380714 239549 380720 239561
rect 390928 239549 390934 239561
rect 390986 239549 390992 239601
rect 637552 239549 637558 239601
rect 637610 239589 637616 239601
rect 650128 239589 650134 239601
rect 637610 239561 650134 239589
rect 637610 239549 637616 239561
rect 650128 239549 650134 239561
rect 650186 239549 650192 239601
rect 291826 239487 297182 239515
rect 298000 239475 298006 239527
rect 298058 239515 298064 239527
rect 303280 239515 303286 239527
rect 298058 239487 303286 239515
rect 298058 239475 298064 239487
rect 303280 239475 303286 239487
rect 303338 239475 303344 239527
rect 310384 239475 310390 239527
rect 310442 239515 310448 239527
rect 312208 239515 312214 239527
rect 310442 239487 312214 239515
rect 310442 239475 310448 239487
rect 312208 239475 312214 239487
rect 312266 239475 312272 239527
rect 369616 239475 369622 239527
rect 369674 239515 369680 239527
rect 392464 239515 392470 239527
rect 369674 239487 392470 239515
rect 369674 239475 369680 239487
rect 392464 239475 392470 239487
rect 392522 239475 392528 239527
rect 638032 239475 638038 239527
rect 638090 239515 638096 239527
rect 650416 239515 650422 239527
rect 638090 239487 650422 239515
rect 638090 239475 638096 239487
rect 650416 239475 650422 239487
rect 650474 239475 650480 239527
rect 280490 239413 287390 239441
rect 280490 239401 280496 239413
rect 288784 239401 288790 239453
rect 288842 239441 288848 239453
rect 290512 239441 290518 239453
rect 288842 239413 290518 239441
rect 288842 239401 288848 239413
rect 290512 239401 290518 239413
rect 290570 239401 290576 239453
rect 290800 239401 290806 239453
rect 290858 239441 290864 239453
rect 295984 239441 295990 239453
rect 290858 239413 295990 239441
rect 290858 239401 290864 239413
rect 295984 239401 295990 239413
rect 296042 239401 296048 239453
rect 325360 239401 325366 239453
rect 325418 239441 325424 239453
rect 325418 239413 338462 239441
rect 325418 239401 325424 239413
rect 245008 239327 245014 239379
rect 245066 239367 245072 239379
rect 273520 239367 273526 239379
rect 245066 239339 273526 239367
rect 245066 239327 245072 239339
rect 273520 239327 273526 239339
rect 273578 239327 273584 239379
rect 274096 239327 274102 239379
rect 274154 239367 274160 239379
rect 285424 239367 285430 239379
rect 274154 239339 285430 239367
rect 274154 239327 274160 239339
rect 285424 239327 285430 239339
rect 285482 239327 285488 239379
rect 290032 239327 290038 239379
rect 290090 239367 290096 239379
rect 299824 239367 299830 239379
rect 290090 239339 299830 239367
rect 290090 239327 290096 239339
rect 299824 239327 299830 239339
rect 299882 239327 299888 239379
rect 304432 239327 304438 239379
rect 304490 239367 304496 239379
rect 306448 239367 306454 239379
rect 304490 239339 306454 239367
rect 304490 239327 304496 239339
rect 306448 239327 306454 239339
rect 306506 239327 306512 239379
rect 326320 239327 326326 239379
rect 326378 239367 326384 239379
rect 338434 239367 338462 239413
rect 368656 239401 368662 239453
rect 368714 239441 368720 239453
rect 390448 239441 390454 239453
rect 368714 239413 390454 239441
rect 368714 239401 368720 239413
rect 390448 239401 390454 239413
rect 390506 239401 390512 239453
rect 637648 239401 637654 239453
rect 637706 239441 637712 239453
rect 650224 239441 650230 239453
rect 637706 239413 650230 239441
rect 637706 239401 637712 239413
rect 650224 239401 650230 239413
rect 650282 239401 650288 239453
rect 349744 239367 349750 239379
rect 326378 239339 338366 239367
rect 338434 239339 349750 239367
rect 326378 239327 326384 239339
rect 222986 239265 229790 239293
rect 222986 239253 222992 239265
rect 229936 239253 229942 239305
rect 229994 239293 230000 239305
rect 231376 239293 231382 239305
rect 229994 239265 231382 239293
rect 229994 239253 230000 239265
rect 231376 239253 231382 239265
rect 231434 239253 231440 239305
rect 275056 239253 275062 239305
rect 275114 239293 275120 239305
rect 292144 239293 292150 239305
rect 275114 239265 292150 239293
rect 275114 239253 275120 239265
rect 292144 239253 292150 239265
rect 292202 239253 292208 239305
rect 292240 239253 292246 239305
rect 292298 239293 292304 239305
rect 301168 239293 301174 239305
rect 292298 239265 301174 239293
rect 292298 239253 292304 239265
rect 301168 239253 301174 239265
rect 301226 239253 301232 239305
rect 319600 239253 319606 239305
rect 319658 239293 319664 239305
rect 336976 239293 336982 239305
rect 319658 239265 336982 239293
rect 319658 239253 319664 239265
rect 336976 239253 336982 239265
rect 337034 239253 337040 239305
rect 338338 239293 338366 239339
rect 349744 239327 349750 239339
rect 349802 239327 349808 239379
rect 369040 239327 369046 239379
rect 369098 239367 369104 239379
rect 391504 239367 391510 239379
rect 369098 239339 391510 239367
rect 369098 239327 369104 239339
rect 391504 239327 391510 239339
rect 391562 239327 391568 239379
rect 494512 239327 494518 239379
rect 494570 239367 494576 239379
rect 497200 239367 497206 239379
rect 494570 239339 497206 239367
rect 494570 239327 494576 239339
rect 497200 239327 497206 239339
rect 497258 239327 497264 239379
rect 638800 239327 638806 239379
rect 638858 239367 638864 239379
rect 649552 239367 649558 239379
rect 638858 239339 649558 239367
rect 638858 239327 638864 239339
rect 649552 239327 649558 239339
rect 649610 239327 649616 239379
rect 352336 239293 352342 239305
rect 338338 239265 352342 239293
rect 352336 239253 352342 239265
rect 352394 239253 352400 239305
rect 370384 239253 370390 239305
rect 370442 239293 370448 239305
rect 394192 239293 394198 239305
rect 370442 239265 394198 239293
rect 370442 239253 370448 239265
rect 394192 239253 394198 239265
rect 394250 239253 394256 239305
rect 639376 239253 639382 239305
rect 639434 239293 639440 239305
rect 649744 239293 649750 239305
rect 639434 239265 649750 239293
rect 639434 239253 639440 239265
rect 649744 239253 649750 239265
rect 649802 239253 649808 239305
rect 140560 239179 140566 239231
rect 140618 239179 140624 239231
rect 216592 239179 216598 239231
rect 216650 239219 216656 239231
rect 233200 239219 233206 239231
rect 216650 239191 233206 239219
rect 216650 239179 216656 239191
rect 233200 239179 233206 239191
rect 233258 239179 233264 239231
rect 277840 239179 277846 239231
rect 277898 239219 277904 239231
rect 281200 239219 281206 239231
rect 277898 239191 281206 239219
rect 277898 239179 277904 239191
rect 281200 239179 281206 239191
rect 281258 239179 281264 239231
rect 282544 239179 282550 239231
rect 282602 239219 282608 239231
rect 287728 239219 287734 239231
rect 282602 239191 287734 239219
rect 282602 239179 282608 239191
rect 287728 239179 287734 239191
rect 287786 239179 287792 239231
rect 288016 239179 288022 239231
rect 288074 239219 288080 239231
rect 293104 239219 293110 239231
rect 288074 239191 293110 239219
rect 288074 239179 288080 239191
rect 293104 239179 293110 239191
rect 293162 239179 293168 239231
rect 294160 239179 294166 239231
rect 294218 239219 294224 239231
rect 301456 239219 301462 239231
rect 294218 239191 301462 239219
rect 294218 239179 294224 239191
rect 301456 239179 301462 239191
rect 301514 239179 301520 239231
rect 322672 239179 322678 239231
rect 322730 239219 322736 239231
rect 328912 239219 328918 239231
rect 322730 239191 328918 239219
rect 322730 239179 322736 239191
rect 328912 239179 328918 239191
rect 328970 239179 328976 239231
rect 329104 239179 329110 239231
rect 329162 239219 329168 239231
rect 343600 239219 343606 239231
rect 329162 239191 343606 239219
rect 329162 239179 329168 239191
rect 343600 239179 343606 239191
rect 343658 239179 343664 239231
rect 371824 239179 371830 239231
rect 371882 239219 371888 239231
rect 396976 239219 396982 239231
rect 371882 239191 396982 239219
rect 371882 239179 371888 239191
rect 396976 239179 396982 239191
rect 397034 239179 397040 239231
rect 505552 239179 505558 239231
rect 505610 239219 505616 239231
rect 674608 239219 674614 239231
rect 505610 239191 674614 239219
rect 505610 239179 505616 239191
rect 674608 239179 674614 239191
rect 674666 239219 674672 239231
rect 675088 239219 675094 239231
rect 674666 239191 675094 239219
rect 674666 239179 674672 239191
rect 675088 239179 675094 239191
rect 675146 239179 675152 239231
rect 140578 239009 140606 239179
rect 228592 239105 228598 239157
rect 228650 239145 228656 239157
rect 231376 239145 231382 239157
rect 228650 239117 231382 239145
rect 228650 239105 228656 239117
rect 231376 239105 231382 239117
rect 231434 239105 231440 239157
rect 237136 239105 237142 239157
rect 237194 239145 237200 239157
rect 238960 239145 238966 239157
rect 237194 239117 238966 239145
rect 237194 239105 237200 239117
rect 238960 239105 238966 239117
rect 239018 239105 239024 239157
rect 274672 239105 274678 239157
rect 274730 239145 274736 239157
rect 287920 239145 287926 239157
rect 274730 239117 287926 239145
rect 274730 239105 274736 239117
rect 287920 239105 287926 239117
rect 287978 239105 287984 239157
rect 288496 239105 288502 239157
rect 288554 239145 288560 239157
rect 301072 239145 301078 239157
rect 288554 239117 301078 239145
rect 288554 239105 288560 239117
rect 301072 239105 301078 239117
rect 301130 239105 301136 239157
rect 319696 239105 319702 239157
rect 319754 239145 319760 239157
rect 337744 239145 337750 239157
rect 319754 239117 337750 239145
rect 319754 239105 319760 239117
rect 337744 239105 337750 239117
rect 337802 239105 337808 239157
rect 381040 239105 381046 239157
rect 381098 239145 381104 239157
rect 391984 239145 391990 239157
rect 381098 239117 391990 239145
rect 381098 239105 381104 239117
rect 391984 239105 391990 239117
rect 392042 239105 392048 239157
rect 510352 239105 510358 239157
rect 510410 239145 510416 239157
rect 674992 239145 674998 239157
rect 510410 239117 674998 239145
rect 510410 239105 510416 239117
rect 674992 239105 674998 239117
rect 675050 239105 675056 239157
rect 144016 239031 144022 239083
rect 144074 239071 144080 239083
rect 174160 239071 174166 239083
rect 144074 239043 174166 239071
rect 144074 239031 144080 239043
rect 174160 239031 174166 239043
rect 174218 239031 174224 239083
rect 208720 239031 208726 239083
rect 208778 239071 208784 239083
rect 215632 239071 215638 239083
rect 208778 239043 215638 239071
rect 208778 239031 208784 239043
rect 215632 239031 215638 239043
rect 215690 239071 215696 239083
rect 222160 239071 222166 239083
rect 215690 239043 222166 239071
rect 215690 239031 215696 239043
rect 222160 239031 222166 239043
rect 222218 239031 222224 239083
rect 227728 239031 227734 239083
rect 227786 239071 227792 239083
rect 236176 239071 236182 239083
rect 227786 239043 236182 239071
rect 227786 239031 227792 239043
rect 236176 239031 236182 239043
rect 236234 239031 236240 239083
rect 236560 239031 236566 239083
rect 236618 239071 236624 239083
rect 238384 239071 238390 239083
rect 236618 239043 238390 239071
rect 236618 239031 236624 239043
rect 238384 239031 238390 239043
rect 238442 239031 238448 239083
rect 277648 239031 277654 239083
rect 277706 239071 277712 239083
rect 286576 239071 286582 239083
rect 277706 239043 286582 239071
rect 277706 239031 277712 239043
rect 286576 239031 286582 239043
rect 286634 239031 286640 239083
rect 294832 239031 294838 239083
rect 294890 239071 294896 239083
rect 302032 239071 302038 239083
rect 294890 239043 302038 239071
rect 294890 239031 294896 239043
rect 302032 239031 302038 239043
rect 302090 239031 302096 239083
rect 327088 239031 327094 239083
rect 327146 239071 327152 239083
rect 338896 239071 338902 239083
rect 327146 239043 338902 239071
rect 327146 239031 327152 239043
rect 338896 239031 338902 239043
rect 338954 239031 338960 239083
rect 379696 239031 379702 239083
rect 379754 239071 379760 239083
rect 388816 239071 388822 239083
rect 379754 239043 388822 239071
rect 379754 239031 379760 239043
rect 388816 239031 388822 239043
rect 388874 239031 388880 239083
rect 420592 239031 420598 239083
rect 420650 239071 420656 239083
rect 421840 239071 421846 239083
rect 420650 239043 421846 239071
rect 420650 239031 420656 239043
rect 421840 239031 421846 239043
rect 421898 239031 421904 239083
rect 541456 239031 541462 239083
rect 541514 239071 541520 239083
rect 549040 239071 549046 239083
rect 541514 239043 549046 239071
rect 541514 239031 541520 239043
rect 549040 239031 549046 239043
rect 549098 239031 549104 239083
rect 639760 239031 639766 239083
rect 639818 239071 639824 239083
rect 649936 239071 649942 239083
rect 639818 239043 649942 239071
rect 639818 239031 639824 239043
rect 649936 239031 649942 239043
rect 649994 239031 650000 239083
rect 140560 238957 140566 239009
rect 140618 238957 140624 239009
rect 264496 238957 264502 239009
rect 264554 238997 264560 239009
rect 314416 238997 314422 239009
rect 264554 238969 314422 238997
rect 264554 238957 264560 238969
rect 314416 238957 314422 238969
rect 314474 238957 314480 239009
rect 325456 238957 325462 239009
rect 325514 238997 325520 239009
rect 396784 238997 396790 239009
rect 325514 238969 396790 238997
rect 325514 238957 325520 238969
rect 396784 238957 396790 238969
rect 396842 238957 396848 239009
rect 140464 238883 140470 238935
rect 140522 238923 140528 238935
rect 141136 238923 141142 238935
rect 140522 238895 141142 238923
rect 140522 238883 140528 238895
rect 141136 238883 141142 238895
rect 141194 238883 141200 238935
rect 235312 238883 235318 238935
rect 235370 238923 235376 238935
rect 270832 238923 270838 238935
rect 235370 238895 270838 238923
rect 235370 238883 235376 238895
rect 270832 238883 270838 238895
rect 270890 238883 270896 238935
rect 271312 238883 271318 238935
rect 271370 238923 271376 238935
rect 340432 238923 340438 238935
rect 271370 238895 340438 238923
rect 271370 238883 271376 238895
rect 340432 238883 340438 238895
rect 340490 238883 340496 238935
rect 384016 238883 384022 238935
rect 384074 238923 384080 238935
rect 384592 238923 384598 238935
rect 384074 238895 384598 238923
rect 384074 238883 384080 238895
rect 384592 238883 384598 238895
rect 384650 238883 384656 238935
rect 266512 238809 266518 238861
rect 266570 238849 266576 238861
rect 338224 238849 338230 238861
rect 266570 238821 338230 238849
rect 266570 238809 266576 238821
rect 338224 238809 338230 238821
rect 338282 238809 338288 238861
rect 235792 238735 235798 238787
rect 235850 238775 235856 238787
rect 269104 238775 269110 238787
rect 235850 238747 269110 238775
rect 235850 238735 235856 238747
rect 269104 238735 269110 238747
rect 269162 238735 269168 238787
rect 277840 238775 277846 238787
rect 276418 238747 277846 238775
rect 256912 238661 256918 238713
rect 256970 238701 256976 238713
rect 276418 238701 276446 238747
rect 277840 238735 277846 238747
rect 277898 238735 277904 238787
rect 278704 238735 278710 238787
rect 278762 238775 278768 238787
rect 339952 238775 339958 238787
rect 278762 238747 339958 238775
rect 278762 238735 278768 238747
rect 339952 238735 339958 238747
rect 340010 238735 340016 238787
rect 256970 238673 276446 238701
rect 256970 238661 256976 238673
rect 276496 238661 276502 238713
rect 276554 238701 276560 238713
rect 336976 238701 336982 238713
rect 276554 238673 336982 238701
rect 276554 238661 276560 238673
rect 336976 238661 336982 238673
rect 337034 238661 337040 238713
rect 247984 238587 247990 238639
rect 248042 238627 248048 238639
rect 248042 238599 261662 238627
rect 248042 238587 248048 238599
rect 42160 238513 42166 238565
rect 42218 238553 42224 238565
rect 42544 238553 42550 238565
rect 42218 238525 42550 238553
rect 42218 238513 42224 238525
rect 42544 238513 42550 238525
rect 42602 238513 42608 238565
rect 217264 238513 217270 238565
rect 217322 238553 217328 238565
rect 259024 238553 259030 238565
rect 217322 238525 259030 238553
rect 217322 238513 217328 238525
rect 259024 238513 259030 238525
rect 259082 238513 259088 238565
rect 261634 238553 261662 238599
rect 261712 238587 261718 238639
rect 261770 238627 261776 238639
rect 336016 238627 336022 238639
rect 261770 238599 336022 238627
rect 261770 238587 261776 238599
rect 336016 238587 336022 238599
rect 336074 238587 336080 238639
rect 264208 238553 264214 238565
rect 261634 238525 264214 238553
rect 264208 238513 264214 238525
rect 264266 238513 264272 238565
rect 264880 238513 264886 238565
rect 264938 238553 264944 238565
rect 337744 238553 337750 238565
rect 264938 238525 337750 238553
rect 264938 238513 264944 238525
rect 337744 238513 337750 238525
rect 337802 238513 337808 238565
rect 237040 238439 237046 238491
rect 237098 238479 237104 238491
rect 257680 238479 257686 238491
rect 237098 238451 257686 238479
rect 237098 238439 237104 238451
rect 257680 238439 257686 238451
rect 257738 238439 257744 238491
rect 259984 238439 259990 238491
rect 260042 238479 260048 238491
rect 335536 238479 335542 238491
rect 260042 238451 335542 238479
rect 260042 238439 260048 238451
rect 335536 238439 335542 238451
rect 335594 238439 335600 238491
rect 219856 238365 219862 238417
rect 219914 238405 219920 238417
rect 253456 238405 253462 238417
rect 219914 238377 253462 238405
rect 219914 238365 219920 238377
rect 253456 238365 253462 238377
rect 253514 238365 253520 238417
rect 255184 238365 255190 238417
rect 255242 238405 255248 238417
rect 356656 238405 356662 238417
rect 255242 238377 356662 238405
rect 255242 238365 255248 238377
rect 356656 238365 356662 238377
rect 356714 238365 356720 238417
rect 218032 238291 218038 238343
rect 218090 238331 218096 238343
rect 257296 238331 257302 238343
rect 218090 238303 257302 238331
rect 218090 238291 218096 238303
rect 257296 238291 257302 238303
rect 257354 238291 257360 238343
rect 263440 238291 263446 238343
rect 263498 238331 263504 238343
rect 276496 238331 276502 238343
rect 263498 238303 276502 238331
rect 263498 238291 263504 238303
rect 276496 238291 276502 238303
rect 276554 238291 276560 238343
rect 277840 238291 277846 238343
rect 277898 238331 277904 238343
rect 357616 238331 357622 238343
rect 277898 238303 357622 238331
rect 277898 238291 277904 238303
rect 357616 238291 357622 238303
rect 357674 238291 357680 238343
rect 218512 238217 218518 238269
rect 218570 238257 218576 238269
rect 255664 238257 255670 238269
rect 218570 238229 255670 238257
rect 218570 238217 218576 238229
rect 255664 238217 255670 238229
rect 255722 238217 255728 238269
rect 355888 238257 355894 238269
rect 260866 238229 355894 238257
rect 220336 238143 220342 238195
rect 220394 238183 220400 238195
rect 251440 238183 251446 238195
rect 220394 238155 251446 238183
rect 220394 238143 220400 238155
rect 251440 238143 251446 238155
rect 251498 238143 251504 238195
rect 253936 238143 253942 238195
rect 253994 238183 254000 238195
rect 260866 238183 260894 238229
rect 355888 238217 355894 238229
rect 355946 238217 355952 238269
rect 355408 238183 355414 238195
rect 253994 238155 260894 238183
rect 264130 238155 355414 238183
rect 253994 238143 254000 238155
rect 252400 238069 252406 238121
rect 252458 238109 252464 238121
rect 264130 238109 264158 238155
rect 355408 238143 355414 238155
rect 355466 238143 355472 238195
rect 252458 238081 264158 238109
rect 252458 238069 252464 238081
rect 264208 238069 264214 238121
rect 264266 238109 264272 238121
rect 353200 238109 353206 238121
rect 264266 238081 353206 238109
rect 264266 238069 264272 238081
rect 353200 238069 353206 238081
rect 353258 238069 353264 238121
rect 249040 237995 249046 238047
rect 249098 238035 249104 238047
rect 353680 238035 353686 238047
rect 249098 238007 353686 238035
rect 249098 237995 249104 238007
rect 353680 237995 353686 238007
rect 353738 237995 353744 238047
rect 350992 237961 350998 237973
rect 257602 237933 350998 237961
rect 42160 237847 42166 237899
rect 42218 237887 42224 237899
rect 50416 237887 50422 237899
rect 42218 237859 50422 237887
rect 42218 237847 42224 237859
rect 50416 237847 50422 237859
rect 50474 237847 50480 237899
rect 243088 237847 243094 237899
rect 243146 237887 243152 237899
rect 257602 237887 257630 237933
rect 350992 237921 350998 237933
rect 351050 237921 351056 237973
rect 243146 237859 257630 237887
rect 243146 237847 243152 237859
rect 257680 237847 257686 237899
rect 257738 237887 257744 237899
rect 347824 237887 347830 237899
rect 257738 237859 347830 237887
rect 257738 237847 257744 237859
rect 347824 237847 347830 237859
rect 347882 237847 347888 237899
rect 361168 237847 361174 237899
rect 361226 237887 361232 237899
rect 399184 237887 399190 237899
rect 361226 237859 399190 237887
rect 361226 237847 361232 237859
rect 399184 237847 399190 237859
rect 399242 237847 399248 237899
rect 241648 237773 241654 237825
rect 241706 237813 241712 237825
rect 350032 237813 350038 237825
rect 241706 237785 350038 237813
rect 241706 237773 241712 237785
rect 350032 237773 350038 237785
rect 350090 237773 350096 237825
rect 361552 237773 361558 237825
rect 361610 237813 361616 237825
rect 400240 237813 400246 237825
rect 361610 237785 400246 237813
rect 361610 237773 361616 237785
rect 400240 237773 400246 237785
rect 400298 237773 400304 237825
rect 244720 237699 244726 237751
rect 244778 237739 244784 237751
rect 351472 237739 351478 237751
rect 244778 237711 351478 237739
rect 244778 237699 244784 237711
rect 351472 237699 351478 237711
rect 351530 237699 351536 237751
rect 363760 237699 363766 237751
rect 363818 237739 363824 237751
rect 404368 237739 404374 237751
rect 363818 237711 404374 237739
rect 363818 237699 363824 237711
rect 404368 237699 404374 237711
rect 404426 237699 404432 237751
rect 140368 237625 140374 237677
rect 140426 237665 140432 237677
rect 140656 237665 140662 237677
rect 140426 237637 140662 237665
rect 140426 237625 140432 237637
rect 140656 237625 140662 237637
rect 140714 237625 140720 237677
rect 239920 237625 239926 237677
rect 239978 237665 239984 237677
rect 349264 237665 349270 237677
rect 239978 237637 349270 237665
rect 239978 237625 239984 237637
rect 349264 237625 349270 237637
rect 349322 237625 349328 237677
rect 363376 237625 363382 237677
rect 363434 237665 363440 237677
rect 403792 237665 403798 237677
rect 363434 237637 403798 237665
rect 363434 237625 363440 237637
rect 403792 237625 403798 237637
rect 403850 237625 403856 237677
rect 233392 237551 233398 237603
rect 233450 237591 233456 237603
rect 346576 237591 346582 237603
rect 233450 237563 346582 237591
rect 233450 237551 233456 237563
rect 346576 237551 346582 237563
rect 346634 237551 346640 237603
rect 364240 237551 364246 237603
rect 364298 237591 364304 237603
rect 406096 237591 406102 237603
rect 364298 237563 406102 237591
rect 364298 237551 364304 237563
rect 406096 237551 406102 237563
rect 406154 237551 406160 237603
rect 277840 237477 277846 237529
rect 277898 237517 277904 237529
rect 312688 237517 312694 237529
rect 277898 237489 312694 237517
rect 277898 237477 277904 237489
rect 312688 237477 312694 237489
rect 312746 237477 312752 237529
rect 316048 237477 316054 237529
rect 316106 237517 316112 237529
rect 380176 237517 380182 237529
rect 316106 237489 380182 237517
rect 316106 237477 316112 237489
rect 380176 237477 380182 237489
rect 380234 237477 380240 237529
rect 266704 237403 266710 237455
rect 266762 237443 266768 237455
rect 309520 237443 309526 237455
rect 266762 237415 309526 237443
rect 266762 237403 266768 237415
rect 309520 237403 309526 237415
rect 309578 237403 309584 237455
rect 316816 237403 316822 237455
rect 316874 237443 316880 237455
rect 381712 237443 381718 237455
rect 316874 237415 381718 237443
rect 316874 237403 316880 237415
rect 381712 237403 381718 237415
rect 381770 237403 381776 237455
rect 140848 237329 140854 237381
rect 140906 237369 140912 237381
rect 141232 237369 141238 237381
rect 140906 237341 141238 237369
rect 140906 237329 140912 237341
rect 141232 237329 141238 237341
rect 141290 237329 141296 237381
rect 266224 237329 266230 237381
rect 266282 237369 266288 237381
rect 310960 237369 310966 237381
rect 266282 237341 310966 237369
rect 266282 237329 266288 237341
rect 310960 237329 310966 237341
rect 311018 237329 311024 237381
rect 315184 237329 315190 237381
rect 315242 237369 315248 237381
rect 377776 237369 377782 237381
rect 315242 237341 377782 237369
rect 315242 237329 315248 237341
rect 377776 237329 377782 237341
rect 377834 237329 377840 237381
rect 267088 237255 267094 237307
rect 267146 237295 267152 237307
rect 308752 237295 308758 237307
rect 267146 237267 308758 237295
rect 267146 237255 267152 237267
rect 308752 237255 308758 237267
rect 308810 237255 308816 237307
rect 313840 237255 313846 237307
rect 313898 237295 313904 237307
rect 375184 237295 375190 237307
rect 313898 237267 375190 237295
rect 313898 237255 313904 237267
rect 375184 237255 375190 237267
rect 375242 237255 375248 237307
rect 140848 237181 140854 237233
rect 140906 237221 140912 237233
rect 141328 237221 141334 237233
rect 140906 237193 141334 237221
rect 140906 237181 140912 237193
rect 141328 237181 141334 237193
rect 141386 237181 141392 237233
rect 267472 237181 267478 237233
rect 267530 237221 267536 237233
rect 307888 237221 307894 237233
rect 267530 237193 307894 237221
rect 267530 237181 267536 237193
rect 307888 237181 307894 237193
rect 307946 237181 307952 237233
rect 317392 237181 317398 237233
rect 317450 237221 317456 237233
rect 382576 237221 382582 237233
rect 317450 237193 382582 237221
rect 317450 237181 317456 237193
rect 382576 237181 382582 237193
rect 382634 237181 382640 237233
rect 269296 237107 269302 237159
rect 269354 237147 269360 237159
rect 303952 237147 303958 237159
rect 269354 237119 303958 237147
rect 269354 237107 269360 237119
rect 303952 237107 303958 237119
rect 304010 237107 304016 237159
rect 313072 237107 313078 237159
rect 313130 237147 313136 237159
rect 374128 237147 374134 237159
rect 313130 237119 374134 237147
rect 313130 237107 313136 237119
rect 374128 237107 374134 237119
rect 374186 237107 374192 237159
rect 269680 237033 269686 237085
rect 269738 237073 269744 237085
rect 278704 237073 278710 237085
rect 269738 237045 278710 237073
rect 269738 237033 269744 237045
rect 278704 237033 278710 237045
rect 278762 237033 278768 237085
rect 286960 237033 286966 237085
rect 287018 237073 287024 237085
rect 302128 237073 302134 237085
rect 287018 237045 302134 237073
rect 287018 237033 287024 237045
rect 302128 237033 302134 237045
rect 302186 237033 302192 237085
rect 314416 237033 314422 237085
rect 314474 237073 314480 237085
rect 376048 237073 376054 237085
rect 314474 237045 376054 237073
rect 314474 237033 314480 237045
rect 376048 237033 376054 237045
rect 376106 237033 376112 237085
rect 235696 236959 235702 237011
rect 235754 236999 235760 237011
rect 269776 236999 269782 237011
rect 235754 236971 269782 236999
rect 235754 236959 235760 236971
rect 269776 236959 269782 236971
rect 269834 236959 269840 237011
rect 274576 236959 274582 237011
rect 274634 236999 274640 237011
rect 305392 236999 305398 237011
rect 274634 236971 305398 236999
rect 274634 236959 274640 236971
rect 305392 236959 305398 236971
rect 305450 236959 305456 237011
rect 312592 236959 312598 237011
rect 312650 236999 312656 237011
rect 372400 236999 372406 237011
rect 312650 236971 372406 236999
rect 312650 236959 312656 236971
rect 372400 236959 372406 236971
rect 372458 236959 372464 237011
rect 265264 236885 265270 236937
rect 265322 236925 265328 236937
rect 277840 236925 277846 236937
rect 265322 236897 277846 236925
rect 265322 236885 265328 236897
rect 277840 236885 277846 236897
rect 277898 236885 277904 236937
rect 301840 236925 301846 236937
rect 277954 236897 301846 236925
rect 270640 236811 270646 236863
rect 270698 236851 270704 236863
rect 277954 236851 277982 236897
rect 301840 236885 301846 236897
rect 301898 236885 301904 236937
rect 302416 236885 302422 236937
rect 302474 236925 302480 236937
rect 303664 236925 303670 236937
rect 302474 236897 303670 236925
rect 302474 236885 302480 236897
rect 303664 236885 303670 236897
rect 303722 236885 303728 236937
rect 312208 236885 312214 236937
rect 312266 236925 312272 236937
rect 371344 236925 371350 236937
rect 312266 236897 371350 236925
rect 312266 236885 312272 236897
rect 371344 236885 371350 236897
rect 371402 236885 371408 236937
rect 270698 236823 277982 236851
rect 270698 236811 270704 236823
rect 284272 236811 284278 236863
rect 284330 236851 284336 236863
rect 322576 236851 322582 236863
rect 284330 236823 322582 236851
rect 284330 236811 284336 236823
rect 322576 236811 322582 236823
rect 322634 236811 322640 236863
rect 284752 236737 284758 236789
rect 284810 236777 284816 236789
rect 320944 236777 320950 236789
rect 284810 236749 320950 236777
rect 284810 236737 284816 236749
rect 320944 236737 320950 236749
rect 321002 236737 321008 236789
rect 42160 236663 42166 236715
rect 42218 236703 42224 236715
rect 43120 236703 43126 236715
rect 42218 236675 43126 236703
rect 42218 236663 42224 236675
rect 43120 236663 43126 236675
rect 43178 236663 43184 236715
rect 284368 236663 284374 236715
rect 284426 236703 284432 236715
rect 321520 236703 321526 236715
rect 284426 236675 321526 236703
rect 284426 236663 284432 236675
rect 321520 236663 321526 236675
rect 321578 236663 321584 236715
rect 285136 236589 285142 236641
rect 285194 236629 285200 236641
rect 319984 236629 319990 236641
rect 285194 236601 319990 236629
rect 285194 236589 285200 236601
rect 319984 236589 319990 236601
rect 320042 236589 320048 236641
rect 286096 236515 286102 236567
rect 286154 236555 286160 236567
rect 318736 236555 318742 236567
rect 286154 236527 318742 236555
rect 286154 236515 286160 236527
rect 318736 236515 318742 236527
rect 318794 236515 318800 236567
rect 43216 236441 43222 236493
rect 43274 236481 43280 236493
rect 43408 236481 43414 236493
rect 43274 236453 43414 236481
rect 43274 236441 43280 236453
rect 43408 236441 43414 236453
rect 43466 236441 43472 236493
rect 291760 236441 291766 236493
rect 291818 236481 291824 236493
rect 323152 236481 323158 236493
rect 291818 236453 323158 236481
rect 291818 236441 291824 236453
rect 323152 236441 323158 236453
rect 323210 236441 323216 236493
rect 43312 236367 43318 236419
rect 43370 236407 43376 236419
rect 43696 236407 43702 236419
rect 43370 236379 43702 236407
rect 43370 236367 43376 236379
rect 43696 236367 43702 236379
rect 43754 236367 43760 236419
rect 286576 236367 286582 236419
rect 286634 236407 286640 236419
rect 317008 236407 317014 236419
rect 286634 236379 317014 236407
rect 286634 236367 286640 236379
rect 317008 236367 317014 236379
rect 317066 236367 317072 236419
rect 290512 236293 290518 236345
rect 290570 236333 290576 236345
rect 319888 236333 319894 236345
rect 290570 236305 319894 236333
rect 290570 236293 290576 236305
rect 319888 236293 319894 236305
rect 319946 236293 319952 236345
rect 144016 236219 144022 236271
rect 144074 236259 144080 236271
rect 165520 236259 165526 236271
rect 144074 236231 165526 236259
rect 144074 236219 144080 236231
rect 165520 236219 165526 236231
rect 165578 236219 165584 236271
rect 286480 236219 286486 236271
rect 286538 236259 286544 236271
rect 317680 236259 317686 236271
rect 286538 236231 317686 236259
rect 286538 236219 286544 236231
rect 317680 236219 317686 236231
rect 317738 236219 317744 236271
rect 144112 236145 144118 236197
rect 144170 236185 144176 236197
rect 168400 236185 168406 236197
rect 144170 236157 168406 236185
rect 144170 236145 144176 236157
rect 168400 236145 168406 236157
rect 168458 236145 168464 236197
rect 290800 236145 290806 236197
rect 290858 236185 290864 236197
rect 320272 236185 320278 236197
rect 290858 236157 320278 236185
rect 290858 236145 290864 236157
rect 320272 236145 320278 236157
rect 320330 236145 320336 236197
rect 273520 236071 273526 236123
rect 273578 236111 273584 236123
rect 361456 236111 361462 236123
rect 273578 236083 361462 236111
rect 273578 236071 273584 236083
rect 361456 236071 361462 236083
rect 361514 236071 361520 236123
rect 257872 235775 257878 235827
rect 257930 235815 257936 235827
rect 333424 235815 333430 235827
rect 257930 235787 333430 235815
rect 257930 235775 257936 235787
rect 333424 235775 333430 235787
rect 333482 235775 333488 235827
rect 257392 235701 257398 235753
rect 257450 235741 257456 235753
rect 335344 235741 335350 235753
rect 257450 235713 335350 235741
rect 257450 235701 257456 235713
rect 335344 235701 335350 235713
rect 335402 235701 335408 235753
rect 248944 235627 248950 235679
rect 249002 235667 249008 235679
rect 329680 235667 329686 235679
rect 249002 235639 329686 235667
rect 249002 235627 249008 235639
rect 329680 235627 329686 235639
rect 329738 235627 329744 235679
rect 256048 235553 256054 235605
rect 256106 235593 256112 235605
rect 337552 235593 337558 235605
rect 256106 235565 337558 235593
rect 256106 235553 256112 235565
rect 337552 235553 337558 235565
rect 337610 235553 337616 235605
rect 255568 235479 255574 235531
rect 255626 235519 255632 235531
rect 339280 235519 339286 235531
rect 255626 235491 339286 235519
rect 255626 235479 255632 235491
rect 339280 235479 339286 235491
rect 339338 235479 339344 235531
rect 42160 235405 42166 235457
rect 42218 235445 42224 235457
rect 43024 235445 43030 235457
rect 42218 235417 43030 235445
rect 42218 235405 42224 235417
rect 43024 235405 43030 235417
rect 43082 235405 43088 235457
rect 254800 235405 254806 235457
rect 254858 235445 254864 235457
rect 340528 235445 340534 235457
rect 254858 235417 340534 235445
rect 254858 235405 254864 235417
rect 340528 235405 340534 235417
rect 340586 235405 340592 235457
rect 253840 235331 253846 235383
rect 253898 235371 253904 235383
rect 342064 235371 342070 235383
rect 253898 235343 342070 235371
rect 253898 235331 253904 235343
rect 342064 235331 342070 235343
rect 342122 235331 342128 235383
rect 253360 235257 253366 235309
rect 253418 235297 253424 235309
rect 344080 235297 344086 235309
rect 253418 235269 344086 235297
rect 253418 235257 253424 235269
rect 344080 235257 344086 235269
rect 344138 235257 344144 235309
rect 675088 235257 675094 235309
rect 675146 235297 675152 235309
rect 679792 235297 679798 235309
rect 675146 235269 679798 235297
rect 675146 235257 675152 235269
rect 679792 235257 679798 235269
rect 679850 235257 679856 235309
rect 252592 235183 252598 235235
rect 252650 235223 252656 235235
rect 345328 235223 345334 235235
rect 252650 235195 345334 235223
rect 252650 235183 252656 235195
rect 345328 235183 345334 235195
rect 345386 235183 345392 235235
rect 674992 235183 674998 235235
rect 675050 235223 675056 235235
rect 679984 235223 679990 235235
rect 675050 235195 679990 235223
rect 675050 235183 675056 235195
rect 679984 235183 679990 235195
rect 680042 235183 680048 235235
rect 251632 235109 251638 235161
rect 251690 235149 251696 235161
rect 346864 235149 346870 235161
rect 251690 235121 346870 235149
rect 251690 235109 251696 235121
rect 346864 235109 346870 235121
rect 346922 235109 346928 235161
rect 257776 235035 257782 235087
rect 257834 235075 257840 235087
rect 358000 235075 358006 235087
rect 257834 235047 358006 235075
rect 257834 235035 257840 235047
rect 358000 235035 358006 235047
rect 358058 235035 358064 235087
rect 251152 234961 251158 235013
rect 251210 235001 251216 235013
rect 348592 235001 348598 235013
rect 251210 234973 348598 235001
rect 251210 234961 251216 234973
rect 348592 234961 348598 234973
rect 348650 234961 348656 235013
rect 258928 234887 258934 234939
rect 258986 234927 258992 234939
rect 358096 234927 358102 234939
rect 258986 234899 358102 234927
rect 258986 234887 258992 234899
rect 358096 234887 358102 234899
rect 358154 234887 358160 234939
rect 42160 234813 42166 234865
rect 42218 234853 42224 234865
rect 42448 234853 42454 234865
rect 42218 234825 42454 234853
rect 42218 234813 42224 234825
rect 42448 234813 42454 234825
rect 42506 234813 42512 234865
rect 250384 234813 250390 234865
rect 250442 234853 250448 234865
rect 350128 234853 350134 234865
rect 250442 234825 350134 234853
rect 250442 234813 250448 234825
rect 350128 234813 350134 234825
rect 350186 234813 350192 234865
rect 210064 234739 210070 234791
rect 210122 234779 210128 234791
rect 383248 234779 383254 234791
rect 210122 234751 383254 234779
rect 210122 234739 210128 234751
rect 383248 234739 383254 234751
rect 383306 234739 383312 234791
rect 42448 234665 42454 234717
rect 42506 234705 42512 234717
rect 43120 234705 43126 234717
rect 42506 234677 43126 234705
rect 42506 234665 42512 234677
rect 43120 234665 43126 234677
rect 43178 234665 43184 234717
rect 249424 234665 249430 234717
rect 249482 234705 249488 234717
rect 351664 234705 351670 234717
rect 249482 234677 351670 234705
rect 249482 234665 249488 234677
rect 351664 234665 351670 234677
rect 351722 234665 351728 234717
rect 264016 234591 264022 234643
rect 264074 234631 264080 234643
rect 370960 234631 370966 234643
rect 264074 234603 370966 234631
rect 264074 234591 264080 234603
rect 370960 234591 370966 234603
rect 371018 234591 371024 234643
rect 248176 234517 248182 234569
rect 248234 234557 248240 234569
rect 354928 234557 354934 234569
rect 248234 234529 354934 234557
rect 248234 234517 248240 234529
rect 354928 234517 354934 234529
rect 354986 234517 354992 234569
rect 263632 234443 263638 234495
rect 263690 234483 263696 234495
rect 371920 234483 371926 234495
rect 263690 234455 371926 234483
rect 263690 234443 263696 234455
rect 371920 234443 371926 234455
rect 371978 234443 371984 234495
rect 247216 234369 247222 234421
rect 247274 234409 247280 234421
rect 356464 234409 356470 234421
rect 247274 234381 356470 234409
rect 247274 234369 247280 234381
rect 356464 234369 356470 234381
rect 356522 234369 356528 234421
rect 246736 234295 246742 234347
rect 246794 234335 246800 234347
rect 357808 234335 357814 234347
rect 246794 234307 357814 234335
rect 246794 234295 246800 234307
rect 357808 234295 357814 234307
rect 357866 234295 357872 234347
rect 245968 234221 245974 234273
rect 246026 234261 246032 234273
rect 359536 234261 359542 234273
rect 246026 234233 359542 234261
rect 246026 234221 246032 234233
rect 359536 234221 359542 234233
rect 359594 234221 359600 234273
rect 42064 234147 42070 234199
rect 42122 234187 42128 234199
rect 42352 234187 42358 234199
rect 42122 234159 42358 234187
rect 42122 234147 42128 234159
rect 42352 234147 42358 234159
rect 42410 234147 42416 234199
rect 262288 234147 262294 234199
rect 262346 234187 262352 234199
rect 374608 234187 374614 234199
rect 262346 234159 374614 234187
rect 262346 234147 262352 234159
rect 374608 234147 374614 234159
rect 374666 234147 374672 234199
rect 261808 234073 261814 234125
rect 261866 234113 261872 234125
rect 375760 234113 375766 234125
rect 261866 234085 375766 234113
rect 261866 234073 261872 234085
rect 375760 234073 375766 234085
rect 375818 234073 375824 234125
rect 260080 233999 260086 234051
rect 260138 234039 260144 234051
rect 379408 234039 379414 234051
rect 260138 234011 379414 234039
rect 260138 233999 260144 234011
rect 379408 233999 379414 234011
rect 379466 233999 379472 234051
rect 260848 233925 260854 233977
rect 260906 233965 260912 233977
rect 377392 233965 377398 233977
rect 260906 233937 377398 233965
rect 260906 233925 260912 233937
rect 377392 233925 377398 233937
rect 377450 233925 377456 233977
rect 243904 233851 243910 233903
rect 243962 233891 243968 233903
rect 363664 233891 363670 233903
rect 243962 233863 363670 233891
rect 243962 233851 243968 233863
rect 363664 233851 363670 233863
rect 363722 233851 363728 233903
rect 258976 233777 258982 233829
rect 259034 233817 259040 233829
rect 381232 233817 381238 233829
rect 259034 233789 381238 233817
rect 259034 233777 259040 233789
rect 381232 233777 381238 233789
rect 381290 233777 381296 233829
rect 207184 233703 207190 233755
rect 207242 233743 207248 233755
rect 213520 233743 213526 233755
rect 207242 233715 213526 233743
rect 207242 233703 207248 233715
rect 213520 233703 213526 233715
rect 213578 233703 213584 233755
rect 220144 233703 220150 233755
rect 220202 233703 220208 233755
rect 258832 233703 258838 233755
rect 258890 233743 258896 233755
rect 382384 233743 382390 233755
rect 258890 233715 382390 233743
rect 258890 233703 258896 233715
rect 382384 233703 382390 233715
rect 382442 233703 382448 233755
rect 210160 233629 210166 233681
rect 210218 233669 210224 233681
rect 212368 233669 212374 233681
rect 210218 233641 212374 233669
rect 210218 233629 210224 233641
rect 212368 233629 212374 233641
rect 212426 233629 212432 233681
rect 220162 233669 220190 233703
rect 358480 233669 358486 233681
rect 220162 233641 358486 233669
rect 358480 233629 358486 233641
rect 358538 233629 358544 233681
rect 210256 233555 210262 233607
rect 210314 233595 210320 233607
rect 212752 233595 212758 233607
rect 210314 233567 212758 233595
rect 210314 233555 210320 233567
rect 212752 233555 212758 233567
rect 212810 233555 212816 233607
rect 216496 233555 216502 233607
rect 216554 233595 216560 233607
rect 414832 233595 414838 233607
rect 216554 233567 414838 233595
rect 216554 233555 216560 233567
rect 414832 233555 414838 233567
rect 414890 233555 414896 233607
rect 144016 233259 144022 233311
rect 144074 233299 144080 233311
rect 171280 233299 171286 233311
rect 144074 233271 171286 233299
rect 144074 233259 144080 233271
rect 171280 233259 171286 233271
rect 171338 233259 171344 233311
rect 204976 233185 204982 233237
rect 205034 233225 205040 233237
rect 206800 233225 206806 233237
rect 205034 233197 206806 233225
rect 205034 233185 205040 233197
rect 206800 233185 206806 233197
rect 206858 233185 206864 233237
rect 645520 233185 645526 233237
rect 645578 233225 645584 233237
rect 649648 233225 649654 233237
rect 645578 233197 649654 233225
rect 645578 233185 645584 233197
rect 649648 233185 649654 233197
rect 649706 233185 649712 233237
rect 204496 233111 204502 233163
rect 204554 233151 204560 233163
rect 206896 233151 206902 233163
rect 204554 233123 206902 233151
rect 204554 233111 204560 233123
rect 206896 233111 206902 233123
rect 206954 233111 206960 233163
rect 645712 233111 645718 233163
rect 645770 233151 645776 233163
rect 649840 233151 649846 233163
rect 645770 233123 649846 233151
rect 645770 233111 645776 233123
rect 649840 233111 649846 233123
rect 649898 233111 649904 233163
rect 204688 233037 204694 233089
rect 204746 233077 204752 233089
rect 206704 233077 206710 233089
rect 204746 233049 206710 233077
rect 204746 233037 204752 233049
rect 206704 233037 206710 233049
rect 206762 233037 206768 233089
rect 645328 233037 645334 233089
rect 645386 233077 645392 233089
rect 650032 233077 650038 233089
rect 645386 233049 650038 233077
rect 645386 233037 645392 233049
rect 650032 233037 650038 233049
rect 650090 233037 650096 233089
rect 645136 232963 645142 233015
rect 645194 233003 645200 233015
rect 650320 233003 650326 233015
rect 645194 232975 650326 233003
rect 645194 232963 645200 232975
rect 650320 232963 650326 232975
rect 650378 232963 650384 233015
rect 645232 232889 645238 232941
rect 645290 232929 645296 232941
rect 650512 232929 650518 232941
rect 645290 232901 650518 232929
rect 645290 232889 645296 232901
rect 650512 232889 650518 232901
rect 650570 232889 650576 232941
rect 204592 232741 204598 232793
rect 204650 232781 204656 232793
rect 206608 232781 206614 232793
rect 204650 232753 206614 232781
rect 204650 232741 204656 232753
rect 206608 232741 206614 232753
rect 206666 232741 206672 232793
rect 144016 230521 144022 230573
rect 144074 230561 144080 230573
rect 151120 230561 151126 230573
rect 144074 230533 151126 230561
rect 144074 230521 144080 230533
rect 151120 230521 151126 230533
rect 151178 230521 151184 230573
rect 144112 230447 144118 230499
rect 144170 230487 144176 230499
rect 162640 230487 162646 230499
rect 144170 230459 162646 230487
rect 144170 230447 144176 230459
rect 162640 230447 162646 230459
rect 162698 230447 162704 230499
rect 141520 230373 141526 230425
rect 141578 230413 141584 230425
rect 201808 230413 201814 230425
rect 141578 230385 201814 230413
rect 141578 230373 141584 230385
rect 201808 230373 201814 230385
rect 201866 230373 201872 230425
rect 139984 230339 139990 230351
rect 139906 230311 139990 230339
rect 139906 229969 139934 230311
rect 139984 230299 139990 230311
rect 140042 230299 140048 230351
rect 141424 230299 141430 230351
rect 141482 230339 141488 230351
rect 201616 230339 201622 230351
rect 141482 230311 201622 230339
rect 141482 230299 141488 230311
rect 201616 230299 201622 230311
rect 201674 230299 201680 230351
rect 178576 230265 178582 230277
rect 175618 230237 178582 230265
rect 172720 230151 172726 230203
rect 172778 230191 172784 230203
rect 175618 230191 175646 230237
rect 178576 230225 178582 230237
rect 178634 230225 178640 230277
rect 172778 230163 175646 230191
rect 172778 230151 172784 230163
rect 178672 230151 178678 230203
rect 178730 230191 178736 230203
rect 201712 230191 201718 230203
rect 178730 230163 201718 230191
rect 178730 230151 178736 230163
rect 201712 230151 201718 230163
rect 201770 230151 201776 230203
rect 139984 230077 139990 230129
rect 140042 230117 140048 230129
rect 141328 230117 141334 230129
rect 140042 230089 141334 230117
rect 140042 230077 140048 230089
rect 141328 230077 141334 230089
rect 141386 230077 141392 230129
rect 143152 230077 143158 230129
rect 143210 230117 143216 230129
rect 146896 230117 146902 230129
rect 143210 230089 146902 230117
rect 143210 230077 143216 230089
rect 146896 230077 146902 230089
rect 146954 230077 146960 230129
rect 166864 230003 166870 230055
rect 166922 230043 166928 230055
rect 172720 230043 172726 230055
rect 166922 230015 172726 230043
rect 166922 230003 166928 230015
rect 172720 230003 172726 230015
rect 172778 230003 172784 230055
rect 139984 229969 139990 229981
rect 139906 229941 139990 229969
rect 139984 229929 139990 229941
rect 140042 229929 140048 229981
rect 661168 229485 661174 229537
rect 661226 229525 661232 229537
rect 674416 229525 674422 229537
rect 661226 229497 674422 229525
rect 661226 229485 661232 229497
rect 674416 229485 674422 229497
rect 674474 229485 674480 229537
rect 669616 228893 669622 228945
rect 669674 228933 669680 228945
rect 674704 228933 674710 228945
rect 669674 228905 674710 228933
rect 669674 228893 669680 228905
rect 674704 228893 674710 228905
rect 674762 228893 674768 228945
rect 141328 227897 141334 227909
rect 139906 227869 141334 227897
rect 139906 227613 139934 227869
rect 141328 227857 141334 227869
rect 141386 227857 141392 227909
rect 669520 227857 669526 227909
rect 669578 227897 669584 227909
rect 674416 227897 674422 227909
rect 669578 227869 674422 227897
rect 669578 227857 669584 227869
rect 674416 227857 674422 227869
rect 674474 227857 674480 227909
rect 140464 227783 140470 227835
rect 140522 227783 140528 227835
rect 140560 227783 140566 227835
rect 140618 227783 140624 227835
rect 140656 227783 140662 227835
rect 140714 227783 140720 227835
rect 140752 227783 140758 227835
rect 140810 227783 140816 227835
rect 140482 227613 140510 227783
rect 140578 227613 140606 227783
rect 140674 227613 140702 227783
rect 140770 227613 140798 227783
rect 144016 227709 144022 227761
rect 144074 227749 144080 227761
rect 188560 227749 188566 227761
rect 144074 227721 188566 227749
rect 144074 227709 144080 227721
rect 188560 227709 188566 227721
rect 188618 227709 188624 227761
rect 144208 227635 144214 227687
rect 144266 227675 144272 227687
rect 194320 227675 194326 227687
rect 144266 227647 194326 227675
rect 144266 227635 144272 227647
rect 194320 227635 194326 227647
rect 194378 227635 194384 227687
rect 139888 227561 139894 227613
rect 139946 227561 139952 227613
rect 140464 227561 140470 227613
rect 140522 227561 140528 227613
rect 140560 227561 140566 227613
rect 140618 227561 140624 227613
rect 140656 227561 140662 227613
rect 140714 227561 140720 227613
rect 140752 227561 140758 227613
rect 140810 227561 140816 227613
rect 144112 227561 144118 227613
rect 144170 227601 144176 227613
rect 197200 227601 197206 227613
rect 144170 227573 197206 227601
rect 144170 227561 144176 227573
rect 197200 227561 197206 227573
rect 197258 227561 197264 227613
rect 141232 227487 141238 227539
rect 141290 227527 141296 227539
rect 201808 227527 201814 227539
rect 141290 227499 201814 227527
rect 141290 227487 141296 227499
rect 201808 227487 201814 227499
rect 201866 227487 201872 227539
rect 140560 227413 140566 227465
rect 140618 227453 140624 227465
rect 197584 227453 197590 227465
rect 140618 227425 197590 227453
rect 140618 227413 140624 227425
rect 197584 227413 197590 227425
rect 197642 227413 197648 227465
rect 140944 227339 140950 227391
rect 141002 227379 141008 227391
rect 201712 227379 201718 227391
rect 141002 227351 201718 227379
rect 141002 227339 141008 227351
rect 201712 227339 201718 227351
rect 201770 227339 201776 227391
rect 140752 227265 140758 227317
rect 140810 227305 140816 227317
rect 201520 227305 201526 227317
rect 140810 227277 201526 227305
rect 140810 227265 140816 227277
rect 201520 227265 201526 227277
rect 201578 227265 201584 227317
rect 140464 227191 140470 227243
rect 140522 227231 140528 227243
rect 201616 227231 201622 227243
rect 140522 227203 201622 227231
rect 140522 227191 140528 227203
rect 201616 227191 201622 227203
rect 201674 227191 201680 227243
rect 144016 225637 144022 225689
rect 144074 225677 144080 225689
rect 156880 225677 156886 225689
rect 144074 225649 156886 225677
rect 144074 225637 144080 225649
rect 156880 225637 156886 225649
rect 156938 225637 156944 225689
rect 144016 224675 144022 224727
rect 144074 224715 144080 224727
rect 179920 224715 179926 224727
rect 144074 224687 179926 224715
rect 144074 224675 144080 224687
rect 179920 224675 179926 224687
rect 179978 224675 179984 224727
rect 140848 224601 140854 224653
rect 140906 224641 140912 224653
rect 201520 224641 201526 224653
rect 140906 224613 201526 224641
rect 140906 224601 140912 224613
rect 201520 224601 201526 224613
rect 201578 224601 201584 224653
rect 140656 224527 140662 224579
rect 140714 224567 140720 224579
rect 201712 224567 201718 224579
rect 140714 224539 201718 224567
rect 140714 224527 140720 224539
rect 201712 224527 201718 224539
rect 201770 224527 201776 224579
rect 141040 224453 141046 224505
rect 141098 224493 141104 224505
rect 201616 224493 201622 224505
rect 141098 224465 201622 224493
rect 141098 224453 141104 224465
rect 201616 224453 201622 224465
rect 201674 224453 201680 224505
rect 146800 224379 146806 224431
rect 146858 224419 146864 224431
rect 201712 224419 201718 224431
rect 146858 224391 201718 224419
rect 146858 224379 146864 224391
rect 201712 224379 201718 224391
rect 201770 224379 201776 224431
rect 149680 224305 149686 224357
rect 149738 224345 149744 224357
rect 201808 224345 201814 224357
rect 149738 224317 201814 224345
rect 149738 224305 149744 224317
rect 201808 224305 201814 224317
rect 201866 224305 201872 224357
rect 152560 224231 152566 224283
rect 152618 224271 152624 224283
rect 209968 224271 209974 224283
rect 152618 224243 209974 224271
rect 152618 224231 152624 224243
rect 209968 224231 209974 224243
rect 210026 224231 210032 224283
rect 209776 223195 209782 223247
rect 209834 223235 209840 223247
rect 210160 223235 210166 223247
rect 209834 223207 210166 223235
rect 209834 223195 209840 223207
rect 210160 223195 210166 223207
rect 210218 223195 210224 223247
rect 144016 221863 144022 221915
rect 144074 221903 144080 221915
rect 177040 221903 177046 221915
rect 144074 221875 177046 221903
rect 144074 221863 144080 221875
rect 177040 221863 177046 221875
rect 177098 221863 177104 221915
rect 144112 221789 144118 221841
rect 144170 221829 144176 221841
rect 202960 221829 202966 221841
rect 144170 221801 202966 221829
rect 144170 221789 144176 221801
rect 202960 221789 202966 221801
rect 203018 221789 203024 221841
rect 146416 221715 146422 221767
rect 146474 221755 146480 221767
rect 146704 221755 146710 221767
rect 146474 221727 146710 221755
rect 146474 221715 146480 221727
rect 146704 221715 146710 221727
rect 146762 221715 146768 221767
rect 155440 221715 155446 221767
rect 155498 221755 155504 221767
rect 198640 221755 198646 221767
rect 155498 221727 198646 221755
rect 155498 221715 155504 221727
rect 198640 221715 198646 221727
rect 198698 221715 198704 221767
rect 161200 221641 161206 221693
rect 161258 221681 161264 221693
rect 201712 221681 201718 221693
rect 161258 221653 201718 221681
rect 161258 221641 161264 221653
rect 201712 221641 201718 221653
rect 201770 221641 201776 221693
rect 164080 221567 164086 221619
rect 164138 221607 164144 221619
rect 209968 221607 209974 221619
rect 164138 221579 209974 221607
rect 164138 221567 164144 221579
rect 209968 221567 209974 221579
rect 210026 221567 210032 221619
rect 166960 221493 166966 221545
rect 167018 221533 167024 221545
rect 201616 221533 201622 221545
rect 167018 221505 201622 221533
rect 167018 221493 167024 221505
rect 201616 221493 201622 221505
rect 201674 221493 201680 221545
rect 169840 221419 169846 221471
rect 169898 221459 169904 221471
rect 201808 221459 201814 221471
rect 169898 221431 201814 221459
rect 169898 221419 169904 221431
rect 201808 221419 201814 221431
rect 201866 221419 201872 221471
rect 42352 221049 42358 221101
rect 42410 221089 42416 221101
rect 45424 221089 45430 221101
rect 42410 221061 45430 221089
rect 42410 221049 42416 221061
rect 45424 221049 45430 221061
rect 45482 221049 45488 221101
rect 42352 220309 42358 220361
rect 42410 220349 42416 220361
rect 45520 220349 45526 220361
rect 42410 220321 45526 220349
rect 42410 220309 42416 220321
rect 45520 220309 45526 220321
rect 45578 220309 45584 220361
rect 42352 219421 42358 219473
rect 42410 219461 42416 219473
rect 45328 219461 45334 219473
rect 42410 219433 45334 219461
rect 42410 219421 42416 219433
rect 45328 219421 45334 219433
rect 45386 219421 45392 219473
rect 144016 218903 144022 218955
rect 144074 218943 144080 218955
rect 174256 218943 174262 218955
rect 144074 218915 174262 218943
rect 144074 218903 144080 218915
rect 174256 218903 174262 218915
rect 174314 218903 174320 218955
rect 140272 218829 140278 218881
rect 140330 218869 140336 218881
rect 197584 218869 197590 218881
rect 140330 218841 197590 218869
rect 140330 218829 140336 218841
rect 197584 218829 197590 218841
rect 197642 218829 197648 218881
rect 175600 218755 175606 218807
rect 175658 218795 175664 218807
rect 209968 218795 209974 218807
rect 175658 218767 209974 218795
rect 175658 218755 175664 218767
rect 209968 218755 209974 218767
rect 210026 218755 210032 218807
rect 178480 218681 178486 218733
rect 178538 218721 178544 218733
rect 201712 218721 201718 218733
rect 178538 218693 201718 218721
rect 178538 218681 178544 218693
rect 201712 218681 201718 218693
rect 201770 218681 201776 218733
rect 181360 218607 181366 218659
rect 181418 218647 181424 218659
rect 198160 218647 198166 218659
rect 181418 218619 198166 218647
rect 181418 218607 181424 218619
rect 198160 218607 198166 218619
rect 198218 218607 198224 218659
rect 184240 218533 184246 218585
rect 184298 218573 184304 218585
rect 210160 218573 210166 218585
rect 184298 218545 210166 218573
rect 184298 218533 184304 218545
rect 210160 218533 210166 218545
rect 210218 218533 210224 218585
rect 144016 216683 144022 216735
rect 144074 216723 144080 216735
rect 154000 216723 154006 216735
rect 144074 216695 154006 216723
rect 144074 216683 144080 216695
rect 154000 216683 154006 216695
rect 154058 216683 154064 216735
rect 140080 215943 140086 215995
rect 140138 215983 140144 215995
rect 201616 215983 201622 215995
rect 140138 215955 201622 215983
rect 140138 215943 140144 215955
rect 201616 215943 201622 215955
rect 201674 215943 201680 215995
rect 139984 215869 139990 215921
rect 140042 215909 140048 215921
rect 210160 215909 210166 215921
rect 140042 215881 210166 215909
rect 140042 215869 140048 215881
rect 210160 215869 210166 215881
rect 210218 215869 210224 215921
rect 140080 215795 140086 215847
rect 140138 215835 140144 215847
rect 201808 215835 201814 215847
rect 140138 215807 201814 215835
rect 140138 215795 140144 215807
rect 201808 215795 201814 215807
rect 201866 215795 201872 215847
rect 140176 215721 140182 215773
rect 140234 215761 140240 215773
rect 201232 215761 201238 215773
rect 140234 215733 201238 215761
rect 140234 215721 140240 215733
rect 201232 215721 201238 215733
rect 201290 215721 201296 215773
rect 187120 215647 187126 215699
rect 187178 215687 187184 215699
rect 201712 215687 201718 215699
rect 187178 215659 201718 215687
rect 187178 215647 187184 215659
rect 201712 215647 201718 215659
rect 201770 215647 201776 215699
rect 192880 215573 192886 215625
rect 192938 215613 192944 215625
rect 209968 215613 209974 215625
rect 192938 215585 209974 215613
rect 192938 215573 192944 215585
rect 209968 215573 209974 215585
rect 210026 215573 210032 215625
rect 144016 213205 144022 213257
rect 144074 213245 144080 213257
rect 168496 213245 168502 213257
rect 144074 213217 168502 213245
rect 144074 213205 144080 213217
rect 168496 213205 168502 213217
rect 168554 213205 168560 213257
rect 144112 213131 144118 213183
rect 144170 213171 144176 213183
rect 171376 213171 171382 213183
rect 144170 213143 171382 213171
rect 144170 213131 144176 213143
rect 171376 213131 171382 213143
rect 171434 213131 171440 213183
rect 140080 213057 140086 213109
rect 140138 213097 140144 213109
rect 201616 213097 201622 213109
rect 140138 213069 201622 213097
rect 140138 213057 140144 213069
rect 201616 213057 201622 213069
rect 201674 213057 201680 213109
rect 139984 212983 139990 213035
rect 140042 212983 140048 213035
rect 140272 212983 140278 213035
rect 140330 213023 140336 213035
rect 201712 213023 201718 213035
rect 140330 212995 201718 213023
rect 140330 212983 140336 212995
rect 201712 212983 201718 212995
rect 201770 212983 201776 213035
rect 140002 212949 140030 212983
rect 209968 212949 209974 212961
rect 140002 212921 209974 212949
rect 209968 212909 209974 212921
rect 210026 212909 210032 212961
rect 144016 210245 144022 210297
rect 144074 210285 144080 210297
rect 148240 210285 148246 210297
rect 144074 210257 148246 210285
rect 144074 210245 144080 210257
rect 148240 210245 148246 210257
rect 148298 210245 148304 210297
rect 645616 210245 645622 210297
rect 645674 210285 645680 210297
rect 646096 210285 646102 210297
rect 645674 210257 646102 210285
rect 645674 210245 645680 210257
rect 646096 210245 646102 210257
rect 646154 210285 646160 210297
rect 679696 210285 679702 210297
rect 646154 210257 679702 210285
rect 646154 210245 646160 210257
rect 679696 210245 679702 210257
rect 679754 210245 679760 210297
rect 674608 210171 674614 210223
rect 674666 210211 674672 210223
rect 676816 210211 676822 210223
rect 674666 210183 676822 210211
rect 674666 210171 674672 210183
rect 676816 210171 676822 210183
rect 676874 210171 676880 210223
rect 209776 208469 209782 208521
rect 209834 208509 209840 208521
rect 210256 208509 210262 208521
rect 209834 208481 210262 208509
rect 209834 208469 209840 208481
rect 210256 208469 210262 208481
rect 210314 208469 210320 208521
rect 144016 207433 144022 207485
rect 144074 207473 144080 207485
rect 162736 207473 162742 207485
rect 144074 207445 162742 207473
rect 144074 207433 144080 207445
rect 162736 207433 162742 207445
rect 162794 207433 162800 207485
rect 144112 207359 144118 207411
rect 144170 207399 144176 207411
rect 165616 207399 165622 207411
rect 144170 207371 165622 207399
rect 144170 207359 144176 207371
rect 165616 207359 165622 207371
rect 165674 207359 165680 207411
rect 146416 207285 146422 207337
rect 146474 207325 146480 207337
rect 146704 207325 146710 207337
rect 146474 207297 146710 207325
rect 146474 207285 146480 207297
rect 146704 207285 146710 207297
rect 146762 207285 146768 207337
rect 674416 205731 674422 205783
rect 674474 205771 674480 205783
rect 675472 205771 675478 205783
rect 674474 205743 675478 205771
rect 674474 205731 674480 205743
rect 675472 205731 675478 205743
rect 675530 205731 675536 205783
rect 675184 205139 675190 205191
rect 675242 205179 675248 205191
rect 675472 205179 675478 205191
rect 675242 205151 675478 205179
rect 675242 205139 675248 205151
rect 675472 205139 675478 205151
rect 675530 205139 675536 205191
rect 675088 204883 675094 204895
rect 675010 204855 675094 204883
rect 675010 204673 675038 204855
rect 675088 204843 675094 204855
rect 675146 204843 675152 204895
rect 674992 204621 674998 204673
rect 675050 204621 675056 204673
rect 42160 204325 42166 204377
rect 42218 204365 42224 204377
rect 44656 204365 44662 204377
rect 42218 204337 44662 204365
rect 42218 204325 42224 204337
rect 44656 204325 44662 204337
rect 44714 204325 44720 204377
rect 146800 201661 146806 201713
rect 146858 201701 146864 201713
rect 185680 201701 185686 201713
rect 146858 201673 185686 201701
rect 146858 201661 146864 201673
rect 185680 201661 185686 201673
rect 185738 201661 185744 201713
rect 144208 201587 144214 201639
rect 144266 201627 144272 201639
rect 200080 201627 200086 201639
rect 144266 201599 200086 201627
rect 144266 201587 144272 201599
rect 200080 201587 200086 201599
rect 200138 201587 200144 201639
rect 40144 201513 40150 201565
rect 40202 201553 40208 201565
rect 42160 201553 42166 201565
rect 40202 201525 42166 201553
rect 40202 201513 40208 201525
rect 42160 201513 42166 201525
rect 42218 201513 42224 201565
rect 674320 201291 674326 201343
rect 674378 201331 674384 201343
rect 675376 201331 675382 201343
rect 674378 201303 675382 201331
rect 674378 201291 674384 201303
rect 675376 201291 675382 201303
rect 675434 201291 675440 201343
rect 37264 200181 37270 200233
rect 37322 200221 37328 200233
rect 43120 200221 43126 200233
rect 37322 200193 43126 200221
rect 37322 200181 37328 200193
rect 43120 200181 43126 200193
rect 43178 200181 43184 200233
rect 146800 198923 146806 198975
rect 146858 198963 146864 198975
rect 159760 198963 159766 198975
rect 146858 198935 159766 198963
rect 146858 198923 146864 198935
rect 159760 198923 159766 198935
rect 159818 198923 159824 198975
rect 37360 198849 37366 198901
rect 37418 198889 37424 198901
rect 43216 198889 43222 198901
rect 37418 198861 43222 198889
rect 37418 198849 37424 198861
rect 43216 198849 43222 198861
rect 43274 198849 43280 198901
rect 40240 198775 40246 198827
rect 40298 198815 40304 198827
rect 43024 198815 43030 198827
rect 40298 198787 43030 198815
rect 40298 198775 40304 198787
rect 43024 198775 43030 198787
rect 43082 198775 43088 198827
rect 146704 198701 146710 198753
rect 146762 198741 146768 198753
rect 191440 198741 191446 198753
rect 146762 198713 191446 198741
rect 146762 198701 146768 198713
rect 191440 198701 191446 198713
rect 191498 198701 191504 198753
rect 674800 197591 674806 197643
rect 674858 197631 674864 197643
rect 675376 197631 675382 197643
rect 674858 197603 675382 197631
rect 674858 197591 674864 197603
rect 675376 197591 675382 197603
rect 675434 197591 675440 197643
rect 42064 197443 42070 197495
rect 42122 197483 42128 197495
rect 42448 197483 42454 197495
rect 42122 197455 42454 197483
rect 42122 197443 42128 197455
rect 42448 197443 42454 197455
rect 42506 197443 42512 197495
rect 41872 197369 41878 197421
rect 41930 197369 41936 197421
rect 41968 197369 41974 197421
rect 42026 197369 42032 197421
rect 41890 197199 41918 197369
rect 41986 197261 42014 197369
rect 42352 197261 42358 197273
rect 41986 197233 42358 197261
rect 42352 197221 42358 197233
rect 42410 197221 42416 197273
rect 41872 197147 41878 197199
rect 41930 197147 41936 197199
rect 674608 196999 674614 197051
rect 674666 197039 674672 197051
rect 675472 197039 675478 197051
rect 674666 197011 675478 197039
rect 674666 196999 674672 197011
rect 675472 196999 675478 197011
rect 675530 196999 675536 197051
rect 674704 196555 674710 196607
rect 674762 196595 674768 196607
rect 675376 196595 675382 196607
rect 674762 196567 675382 196595
rect 674762 196555 674768 196567
rect 675376 196555 675382 196567
rect 675434 196555 675440 196607
rect 146800 195815 146806 195867
rect 146858 195855 146864 195867
rect 182800 195855 182806 195867
rect 146858 195827 182806 195855
rect 146858 195815 146864 195827
rect 182800 195815 182806 195827
rect 182858 195815 182864 195867
rect 42640 195741 42646 195793
rect 42698 195781 42704 195793
rect 43216 195781 43222 195793
rect 42698 195753 43222 195781
rect 42698 195741 42704 195753
rect 43216 195741 43222 195753
rect 43274 195741 43280 195793
rect 42160 195297 42166 195349
rect 42218 195337 42224 195349
rect 42352 195337 42358 195349
rect 42218 195309 42358 195337
rect 42218 195297 42224 195309
rect 42352 195297 42358 195309
rect 42410 195297 42416 195349
rect 42064 194483 42070 194535
rect 42122 194523 42128 194535
rect 47632 194523 47638 194535
rect 42122 194495 47638 194523
rect 42122 194483 42128 194495
rect 47632 194483 47638 194495
rect 47690 194483 47696 194535
rect 42064 193447 42070 193499
rect 42122 193487 42128 193499
rect 43120 193487 43126 193499
rect 42122 193459 43126 193487
rect 42122 193447 42128 193459
rect 43120 193447 43126 193459
rect 43178 193447 43184 193499
rect 146800 193003 146806 193055
rect 146858 193043 146864 193055
rect 148336 193043 148342 193055
rect 146858 193015 148342 193043
rect 146858 193003 146864 193015
rect 148336 193003 148342 193015
rect 148394 193003 148400 193055
rect 42160 192189 42166 192241
rect 42218 192229 42224 192241
rect 43024 192229 43030 192241
rect 42218 192201 43030 192229
rect 42218 192189 42224 192201
rect 43024 192189 43030 192201
rect 43082 192189 43088 192241
rect 42064 191449 42070 191501
rect 42122 191489 42128 191501
rect 42352 191489 42358 191501
rect 42122 191461 42358 191489
rect 42122 191449 42128 191461
rect 42352 191449 42358 191461
rect 42410 191449 42416 191501
rect 42352 191301 42358 191353
rect 42410 191341 42416 191353
rect 42640 191341 42646 191353
rect 42410 191313 42646 191341
rect 42410 191301 42416 191313
rect 42640 191301 42646 191313
rect 42698 191301 42704 191353
rect 146704 190191 146710 190243
rect 146762 190231 146768 190243
rect 148432 190231 148438 190243
rect 146762 190203 148438 190231
rect 146762 190191 146768 190203
rect 148432 190191 148438 190203
rect 148490 190191 148496 190243
rect 146800 190117 146806 190169
rect 146858 190157 146864 190169
rect 200176 190157 200182 190169
rect 146858 190129 200182 190157
rect 146858 190117 146864 190129
rect 200176 190117 200182 190129
rect 200234 190117 200240 190169
rect 42160 187823 42166 187875
rect 42218 187863 42224 187875
rect 42736 187863 42742 187875
rect 42218 187835 42742 187863
rect 42218 187823 42224 187835
rect 42736 187823 42742 187835
rect 42794 187823 42800 187875
rect 146704 187305 146710 187357
rect 146762 187345 146768 187357
rect 148528 187345 148534 187357
rect 146762 187317 148534 187345
rect 146762 187305 146768 187317
rect 148528 187305 148534 187317
rect 148586 187305 148592 187357
rect 146800 187231 146806 187283
rect 146858 187271 146864 187283
rect 194416 187271 194422 187283
rect 146858 187243 194422 187271
rect 146858 187231 146864 187243
rect 194416 187231 194422 187243
rect 194474 187231 194480 187283
rect 42160 187083 42166 187135
rect 42218 187123 42224 187135
rect 42448 187123 42454 187135
rect 42218 187095 42454 187123
rect 42218 187083 42224 187095
rect 42448 187083 42454 187095
rect 42506 187083 42512 187135
rect 42064 186491 42070 186543
rect 42122 186531 42128 186543
rect 42640 186531 42646 186543
rect 42122 186503 42646 186531
rect 42122 186491 42128 186503
rect 42640 186491 42646 186503
rect 42698 186491 42704 186543
rect 144016 184345 144022 184397
rect 144074 184385 144080 184397
rect 151216 184385 151222 184397
rect 144074 184357 151222 184385
rect 144074 184345 144080 184357
rect 151216 184345 151222 184357
rect 151274 184345 151280 184397
rect 655312 184345 655318 184397
rect 655370 184385 655376 184397
rect 674416 184385 674422 184397
rect 655370 184357 674422 184385
rect 655370 184345 655376 184357
rect 674416 184345 674422 184357
rect 674474 184345 674480 184397
rect 660976 183901 660982 183953
rect 661034 183941 661040 183953
rect 674704 183941 674710 183953
rect 661034 183913 674710 183941
rect 661034 183901 661040 183913
rect 674704 183901 674710 183913
rect 674762 183901 674768 183953
rect 666736 182865 666742 182917
rect 666794 182905 666800 182917
rect 674416 182905 674422 182917
rect 666794 182877 674422 182905
rect 666794 182865 666800 182877
rect 674416 182865 674422 182877
rect 674474 182865 674480 182917
rect 144016 181459 144022 181511
rect 144074 181499 144080 181511
rect 185776 181499 185782 181511
rect 144074 181471 185782 181499
rect 144074 181459 144080 181471
rect 185776 181459 185782 181471
rect 185834 181459 185840 181511
rect 144112 178647 144118 178699
rect 144170 178687 144176 178699
rect 148624 178687 148630 178699
rect 144170 178659 148630 178687
rect 144170 178647 144176 178659
rect 148624 178647 148630 178659
rect 148682 178647 148688 178699
rect 144016 178573 144022 178625
rect 144074 178613 144080 178625
rect 191536 178613 191542 178625
rect 144074 178585 191542 178613
rect 144074 178573 144080 178585
rect 191536 178573 191542 178585
rect 191594 178573 191600 178625
rect 144016 175687 144022 175739
rect 144074 175727 144080 175739
rect 188656 175727 188662 175739
rect 144074 175699 188662 175727
rect 144074 175687 144080 175699
rect 188656 175687 188662 175699
rect 188714 175687 188720 175739
rect 144016 172801 144022 172853
rect 144074 172841 144080 172853
rect 182896 172841 182902 172853
rect 144074 172813 182902 172841
rect 144074 172801 144080 172813
rect 182896 172801 182902 172813
rect 182954 172801 182960 172853
rect 144016 170359 144022 170411
rect 144074 170399 144080 170411
rect 159856 170399 159862 170411
rect 144074 170371 159862 170399
rect 144074 170359 144080 170371
rect 159856 170359 159862 170371
rect 159914 170359 159920 170411
rect 209968 169915 209974 169967
rect 210026 169955 210032 169967
rect 210160 169955 210166 169967
rect 210026 169927 210166 169955
rect 210026 169915 210032 169927
rect 210160 169915 210166 169927
rect 210218 169915 210224 169967
rect 209872 169841 209878 169893
rect 209930 169881 209936 169893
rect 209930 169853 210110 169881
rect 209930 169841 209936 169853
rect 209776 169767 209782 169819
rect 209834 169807 209840 169819
rect 209968 169807 209974 169819
rect 209834 169779 209974 169807
rect 209834 169767 209840 169779
rect 209968 169767 209974 169779
rect 210026 169767 210032 169819
rect 209872 169693 209878 169745
rect 209930 169733 209936 169745
rect 210082 169733 210110 169853
rect 209930 169705 210110 169733
rect 209930 169693 209936 169705
rect 647920 167177 647926 167229
rect 647978 167217 647984 167229
rect 674704 167217 674710 167229
rect 647978 167189 674710 167217
rect 647978 167177 647984 167189
rect 674704 167177 674710 167189
rect 674762 167177 674768 167229
rect 144016 167103 144022 167155
rect 144074 167143 144080 167155
rect 156976 167143 156982 167155
rect 144074 167115 156982 167143
rect 144074 167103 144080 167115
rect 156976 167103 156982 167115
rect 157034 167103 157040 167155
rect 144112 167029 144118 167081
rect 144170 167069 144176 167081
rect 148720 167069 148726 167081
rect 144170 167041 148726 167069
rect 144170 167029 144176 167041
rect 148720 167029 148726 167041
rect 148778 167029 148784 167081
rect 646192 164217 646198 164269
rect 646250 164257 646256 164269
rect 674608 164257 674614 164269
rect 646250 164229 674614 164257
rect 646250 164217 646256 164229
rect 674608 164217 674614 164229
rect 674666 164217 674672 164269
rect 144016 164143 144022 164195
rect 144074 164183 144080 164195
rect 148816 164183 148822 164195
rect 144074 164155 148822 164183
rect 144074 164143 144080 164155
rect 148816 164143 148822 164155
rect 148874 164143 148880 164195
rect 645904 164143 645910 164195
rect 645962 164183 645968 164195
rect 674704 164183 674710 164195
rect 645962 164155 674710 164183
rect 645962 164143 645968 164155
rect 674704 164143 674710 164155
rect 674762 164143 674768 164195
rect 675280 164069 675286 164121
rect 675338 164109 675344 164121
rect 677008 164109 677014 164121
rect 675338 164081 677014 164109
rect 675338 164069 675344 164081
rect 677008 164069 677014 164081
rect 677066 164069 677072 164121
rect 674800 163255 674806 163307
rect 674858 163295 674864 163307
rect 676816 163295 676822 163307
rect 674858 163267 676822 163295
rect 674858 163255 674864 163267
rect 676816 163255 676822 163267
rect 676874 163255 676880 163307
rect 144016 161331 144022 161383
rect 144074 161371 144080 161383
rect 148912 161371 148918 161383
rect 144074 161343 148918 161371
rect 144074 161331 144080 161343
rect 148912 161331 148918 161343
rect 148970 161331 148976 161383
rect 144112 161257 144118 161309
rect 144170 161297 144176 161309
rect 197296 161297 197302 161309
rect 144170 161269 197302 161297
rect 144170 161257 144176 161269
rect 197296 161257 197302 161269
rect 197354 161257 197360 161309
rect 674416 160739 674422 160791
rect 674474 160779 674480 160791
rect 675376 160779 675382 160791
rect 674474 160751 675382 160779
rect 674474 160739 674480 160751
rect 675376 160739 675382 160751
rect 675434 160739 675440 160791
rect 675184 159999 675190 160051
rect 675242 160039 675248 160051
rect 675472 160039 675478 160051
rect 675242 160011 675478 160039
rect 675242 159999 675248 160011
rect 675472 159999 675478 160011
rect 675530 159999 675536 160051
rect 674032 159407 674038 159459
rect 674090 159447 674096 159459
rect 675376 159447 675382 159459
rect 674090 159419 675382 159447
rect 674090 159407 674096 159419
rect 675376 159407 675382 159419
rect 675434 159407 675440 159459
rect 144016 158445 144022 158497
rect 144074 158485 144080 158497
rect 149200 158485 149206 158497
rect 144074 158457 149206 158485
rect 144074 158445 144080 158457
rect 149200 158445 149206 158457
rect 149258 158445 149264 158497
rect 144880 157113 144886 157165
rect 144938 157153 144944 157165
rect 146800 157153 146806 157165
rect 144938 157125 146806 157153
rect 144938 157113 144944 157125
rect 146800 157113 146806 157125
rect 146858 157113 146864 157165
rect 674992 157039 674998 157091
rect 675050 157079 675056 157091
rect 675184 157079 675190 157091
rect 675050 157051 675190 157079
rect 675050 157039 675056 157051
rect 675184 157039 675190 157051
rect 675242 157039 675248 157091
rect 144880 156965 144886 157017
rect 144938 157005 144944 157017
rect 146608 157005 146614 157017
rect 144938 156977 146614 157005
rect 144938 156965 144944 156977
rect 146608 156965 146614 156977
rect 146666 156965 146672 157017
rect 674896 156891 674902 156943
rect 674954 156931 674960 156943
rect 675472 156931 675478 156943
rect 674954 156903 675478 156931
rect 674954 156891 674960 156903
rect 675472 156891 675478 156903
rect 675530 156891 675536 156943
rect 144016 155559 144022 155611
rect 144074 155599 144080 155611
rect 149296 155599 149302 155611
rect 144074 155571 149302 155599
rect 144074 155559 144080 155571
rect 149296 155559 149302 155571
rect 149354 155559 149360 155611
rect 144016 152747 144022 152799
rect 144074 152787 144080 152799
rect 177136 152787 177142 152799
rect 144074 152759 177142 152787
rect 144074 152747 144080 152759
rect 177136 152747 177142 152759
rect 177194 152747 177200 152799
rect 144112 152673 144118 152725
rect 144170 152713 144176 152725
rect 180016 152713 180022 152725
rect 144170 152685 180022 152713
rect 144170 152673 144176 152685
rect 180016 152673 180022 152685
rect 180074 152673 180080 152725
rect 674320 152599 674326 152651
rect 674378 152639 674384 152651
rect 675376 152639 675382 152651
rect 674378 152611 675382 152639
rect 674378 152599 674384 152611
rect 675376 152599 675382 152611
rect 675434 152599 675440 152651
rect 674800 152155 674806 152207
rect 674858 152195 674864 152207
rect 675472 152195 675478 152207
rect 674858 152167 675478 152195
rect 674858 152155 674864 152167
rect 675472 152155 675478 152167
rect 675530 152155 675536 152207
rect 674512 151415 674518 151467
rect 674570 151455 674576 151467
rect 675376 151455 675382 151467
rect 674570 151427 675382 151455
rect 674570 151415 674576 151427
rect 675376 151415 675382 151427
rect 675434 151415 675440 151467
rect 144112 149861 144118 149913
rect 144170 149901 144176 149913
rect 149392 149901 149398 149913
rect 144170 149873 149398 149901
rect 144170 149861 144176 149873
rect 149392 149861 149398 149873
rect 149450 149861 149456 149913
rect 144016 149787 144022 149839
rect 144074 149827 144080 149839
rect 174352 149827 174358 149839
rect 144074 149799 174358 149827
rect 144074 149787 144080 149799
rect 174352 149787 174358 149799
rect 174410 149787 174416 149839
rect 209776 149787 209782 149839
rect 209834 149827 209840 149839
rect 209968 149827 209974 149839
rect 209834 149799 209974 149827
rect 209834 149787 209840 149799
rect 209968 149787 209974 149799
rect 210026 149787 210032 149839
rect 144016 149639 144022 149691
rect 144074 149679 144080 149691
rect 144304 149679 144310 149691
rect 144074 149651 144310 149679
rect 144074 149639 144080 149651
rect 144304 149639 144310 149651
rect 144362 149639 144368 149691
rect 144304 149491 144310 149543
rect 144362 149531 144368 149543
rect 144496 149531 144502 149543
rect 144362 149503 144502 149531
rect 144362 149491 144368 149503
rect 144496 149491 144502 149503
rect 144554 149491 144560 149543
rect 209968 148233 209974 148285
rect 210026 148273 210032 148285
rect 210160 148273 210166 148285
rect 210026 148245 210166 148273
rect 210026 148233 210032 148245
rect 210160 148233 210166 148245
rect 210218 148233 210224 148285
rect 144016 146975 144022 147027
rect 144074 147015 144080 147027
rect 149488 147015 149494 147027
rect 144074 146987 149494 147015
rect 144074 146975 144080 146987
rect 149488 146975 149494 146987
rect 149546 146975 149552 147027
rect 210064 147015 210070 147027
rect 209890 146987 210070 147015
rect 144208 146901 144214 146953
rect 144266 146941 144272 146953
rect 171472 146941 171478 146953
rect 144266 146913 171478 146941
rect 144266 146901 144272 146913
rect 171472 146901 171478 146913
rect 171530 146901 171536 146953
rect 209890 146719 209918 146987
rect 210064 146975 210070 146987
rect 210122 146975 210128 147027
rect 210256 146867 210262 146879
rect 209986 146839 210262 146867
rect 209986 146805 210014 146839
rect 210256 146827 210262 146839
rect 210314 146827 210320 146879
rect 209968 146753 209974 146805
rect 210026 146753 210032 146805
rect 210064 146719 210070 146731
rect 209890 146691 210070 146719
rect 210064 146679 210070 146691
rect 210122 146679 210128 146731
rect 144688 144311 144694 144363
rect 144746 144351 144752 144363
rect 144880 144351 144886 144363
rect 144746 144323 144886 144351
rect 144746 144311 144752 144323
rect 144880 144311 144886 144323
rect 144938 144311 144944 144363
rect 144208 144015 144214 144067
rect 144266 144055 144272 144067
rect 154096 144055 154102 144067
rect 144266 144027 154102 144055
rect 144266 144015 144272 144027
rect 154096 144015 154102 144027
rect 154154 144015 154160 144067
rect 144688 141391 144694 141403
rect 144130 141363 144694 141391
rect 144130 141021 144158 141363
rect 144688 141351 144694 141363
rect 144746 141351 144752 141403
rect 144400 141203 144406 141255
rect 144458 141243 144464 141255
rect 149584 141243 149590 141255
rect 144458 141215 149590 141243
rect 144458 141203 144464 141215
rect 149584 141203 149590 141215
rect 149642 141203 149648 141255
rect 144208 141129 144214 141181
rect 144266 141169 144272 141181
rect 168592 141169 168598 141181
rect 144266 141141 168598 141169
rect 144266 141129 144272 141141
rect 168592 141129 168598 141141
rect 168650 141129 168656 141181
rect 146512 141055 146518 141107
rect 146570 141055 146576 141107
rect 144208 141021 144214 141033
rect 144130 140993 144214 141021
rect 144208 140981 144214 140993
rect 144266 140981 144272 141033
rect 146530 141021 146558 141055
rect 147184 141021 147190 141033
rect 146530 140993 147190 141021
rect 147184 140981 147190 140993
rect 147242 140981 147248 141033
rect 146032 140463 146038 140515
rect 146090 140503 146096 140515
rect 146704 140503 146710 140515
rect 146090 140475 146710 140503
rect 146090 140463 146096 140475
rect 146704 140463 146710 140475
rect 146762 140463 146768 140515
rect 144208 138579 144214 138591
rect 144130 138551 144214 138579
rect 144130 138283 144158 138551
rect 144208 138539 144214 138551
rect 144266 138539 144272 138591
rect 655216 138539 655222 138591
rect 655274 138579 655280 138591
rect 674704 138579 674710 138591
rect 655274 138551 674710 138579
rect 655274 138539 655280 138551
rect 674704 138539 674710 138551
rect 674762 138539 674768 138591
rect 655120 138391 655126 138443
rect 655178 138431 655184 138443
rect 674416 138431 674422 138443
rect 655178 138403 674422 138431
rect 655178 138391 655184 138403
rect 674416 138391 674422 138403
rect 674474 138391 674480 138443
rect 144208 138317 144214 138369
rect 144266 138357 144272 138369
rect 149680 138357 149686 138369
rect 144266 138329 149686 138357
rect 144266 138317 144272 138329
rect 149680 138317 149686 138329
rect 149738 138317 149744 138369
rect 144130 138255 144254 138283
rect 144226 138135 144254 138255
rect 144400 138243 144406 138295
rect 144458 138283 144464 138295
rect 165712 138283 165718 138295
rect 144458 138255 165718 138283
rect 144458 138243 144464 138255
rect 165712 138243 165718 138255
rect 165770 138243 165776 138295
rect 144400 138135 144406 138147
rect 144226 138107 144406 138135
rect 144400 138095 144406 138107
rect 144458 138095 144464 138147
rect 144880 136911 144886 136963
rect 144938 136951 144944 136963
rect 144938 136923 145982 136951
rect 144938 136911 144944 136923
rect 144496 136763 144502 136815
rect 144554 136803 144560 136815
rect 144880 136803 144886 136815
rect 144554 136775 144886 136803
rect 144554 136763 144560 136775
rect 144880 136763 144886 136775
rect 144938 136763 144944 136815
rect 145954 136729 145982 136923
rect 145954 136701 146558 136729
rect 146530 136667 146558 136701
rect 146512 136615 146518 136667
rect 146570 136615 146576 136667
rect 144400 136245 144406 136297
rect 144458 136285 144464 136297
rect 144688 136285 144694 136297
rect 144458 136257 144694 136285
rect 144458 136245 144464 136257
rect 144688 136245 144694 136257
rect 144746 136245 144752 136297
rect 144592 136171 144598 136223
rect 144650 136171 144656 136223
rect 144610 136001 144638 136171
rect 144592 135949 144598 136001
rect 144650 135949 144656 136001
rect 655408 135579 655414 135631
rect 655466 135619 655472 135631
rect 674608 135619 674614 135631
rect 655466 135591 674614 135619
rect 655466 135579 655472 135591
rect 674608 135579 674614 135591
rect 674666 135579 674672 135631
rect 144496 135431 144502 135483
rect 144554 135471 144560 135483
rect 147088 135471 147094 135483
rect 144554 135443 147094 135471
rect 144554 135431 144560 135443
rect 147088 135431 147094 135443
rect 147146 135431 147152 135483
rect 646480 135357 646486 135409
rect 646538 135397 646544 135409
rect 674704 135397 674710 135409
rect 646538 135369 674710 135397
rect 646538 135357 646544 135369
rect 674704 135357 674710 135369
rect 674762 135357 674768 135409
rect 143920 134099 143926 134151
rect 143978 134139 143984 134151
rect 144400 134139 144406 134151
rect 143978 134111 144406 134139
rect 143978 134099 143984 134111
rect 144400 134099 144406 134111
rect 144458 134099 144464 134151
rect 146704 134099 146710 134151
rect 146762 134139 146768 134151
rect 146992 134139 146998 134151
rect 146762 134111 146998 134139
rect 146762 134099 146768 134111
rect 146992 134099 146998 134111
rect 147050 134099 147056 134151
rect 144496 132693 144502 132745
rect 144554 132733 144560 132745
rect 162928 132733 162934 132745
rect 144554 132705 162934 132733
rect 144554 132693 144560 132705
rect 162928 132693 162934 132705
rect 162986 132693 162992 132745
rect 144400 132545 144406 132597
rect 144458 132585 144464 132597
rect 208816 132585 208822 132597
rect 144458 132557 208822 132585
rect 144458 132545 144464 132557
rect 208816 132545 208822 132557
rect 208874 132545 208880 132597
rect 144208 132471 144214 132523
rect 144266 132511 144272 132523
rect 208912 132511 208918 132523
rect 144266 132483 208918 132511
rect 144266 132471 144272 132483
rect 208912 132471 208918 132483
rect 208970 132471 208976 132523
rect 143920 132397 143926 132449
rect 143978 132437 143984 132449
rect 144496 132437 144502 132449
rect 143978 132409 144502 132437
rect 143978 132397 143984 132409
rect 144496 132397 144502 132409
rect 144554 132397 144560 132449
rect 144208 130103 144214 130155
rect 144266 130143 144272 130155
rect 151312 130143 151318 130155
rect 144266 130115 151318 130143
rect 144266 130103 144272 130115
rect 151312 130103 151318 130115
rect 151370 130103 151376 130155
rect 144208 129585 144214 129637
rect 144266 129625 144272 129637
rect 209008 129625 209014 129637
rect 144266 129597 209014 129625
rect 144266 129585 144272 129597
rect 209008 129585 209014 129597
rect 209066 129585 209072 129637
rect 144208 129437 144214 129489
rect 144266 129477 144272 129489
rect 144688 129477 144694 129489
rect 144266 129449 144694 129477
rect 144266 129437 144272 129449
rect 144688 129437 144694 129449
rect 144746 129437 144752 129489
rect 146512 129403 146518 129415
rect 144706 129375 146518 129403
rect 144706 129341 144734 129375
rect 146512 129363 146518 129375
rect 146570 129363 146576 129415
rect 144688 129289 144694 129341
rect 144746 129289 144752 129341
rect 146896 126995 146902 127047
rect 146954 127035 146960 127047
rect 148144 127035 148150 127047
rect 146954 127007 148150 127035
rect 146954 126995 146960 127007
rect 148144 126995 148150 127007
rect 148202 126995 148208 127047
rect 209968 126995 209974 127047
rect 210026 127035 210032 127047
rect 210026 127007 210302 127035
rect 210026 126995 210032 127007
rect 146896 126773 146902 126825
rect 146954 126813 146960 126825
rect 148048 126813 148054 126825
rect 146954 126785 148054 126813
rect 146954 126773 146960 126785
rect 148048 126773 148054 126785
rect 148106 126773 148112 126825
rect 210274 126751 210302 127007
rect 146512 126699 146518 126751
rect 146570 126739 146576 126751
rect 200272 126739 200278 126751
rect 146570 126711 200278 126739
rect 146570 126699 146576 126711
rect 200272 126699 200278 126711
rect 200330 126699 200336 126751
rect 209968 126699 209974 126751
rect 210026 126739 210032 126751
rect 210160 126739 210166 126751
rect 210026 126711 210166 126739
rect 210026 126699 210032 126711
rect 210160 126699 210166 126711
rect 210218 126699 210224 126751
rect 210256 126699 210262 126751
rect 210314 126699 210320 126751
rect 146896 126625 146902 126677
rect 146954 126665 146960 126677
rect 147184 126665 147190 126677
rect 146954 126637 147190 126665
rect 146954 126625 146960 126637
rect 147184 126625 147190 126637
rect 147242 126625 147248 126677
rect 144784 125293 144790 125345
rect 144842 125333 144848 125345
rect 146608 125333 146614 125345
rect 144842 125305 146614 125333
rect 144842 125293 144848 125305
rect 146608 125293 146614 125305
rect 146666 125293 146672 125345
rect 144592 124479 144598 124531
rect 144650 124519 144656 124531
rect 146032 124519 146038 124531
rect 144650 124491 146038 124519
rect 144650 124479 144656 124491
rect 146032 124479 146038 124491
rect 146090 124479 146096 124531
rect 144592 123961 144598 124013
rect 144650 124001 144656 124013
rect 194512 124001 194518 124013
rect 144650 123973 194518 124001
rect 144650 123961 144656 123973
rect 194512 123961 194518 123973
rect 194570 123961 194576 124013
rect 144784 123887 144790 123939
rect 144842 123927 144848 123939
rect 197392 123927 197398 123939
rect 144842 123899 197398 123927
rect 144842 123887 144848 123899
rect 197392 123887 197398 123899
rect 197450 123887 197456 123939
rect 647824 121223 647830 121275
rect 647882 121263 647888 121275
rect 674704 121263 674710 121275
rect 647882 121235 674710 121263
rect 647882 121223 647888 121235
rect 674704 121223 674710 121235
rect 674762 121223 674768 121275
rect 144592 121149 144598 121201
rect 144650 121189 144656 121201
rect 203056 121189 203062 121201
rect 144650 121161 203062 121189
rect 144650 121149 144656 121161
rect 203056 121149 203062 121161
rect 203114 121149 203120 121201
rect 647920 121149 647926 121201
rect 647978 121189 647984 121201
rect 674800 121189 674806 121201
rect 647978 121161 674806 121189
rect 647978 121149 647984 121161
rect 674800 121149 674806 121161
rect 674858 121149 674864 121201
rect 647824 121075 647830 121127
rect 647882 121115 647888 121127
rect 674608 121115 674614 121127
rect 647882 121087 674614 121115
rect 647882 121075 647888 121087
rect 674608 121075 674614 121087
rect 674666 121075 674672 121127
rect 144784 121001 144790 121053
rect 144842 121041 144848 121053
rect 209104 121041 209110 121053
rect 144842 121013 209110 121041
rect 144842 121001 144848 121013
rect 209104 121001 209110 121013
rect 209162 121001 209168 121053
rect 674800 119965 674806 120017
rect 674858 120005 674864 120017
rect 675184 120005 675190 120017
rect 674858 119977 675190 120005
rect 674858 119965 674864 119977
rect 675184 119965 675190 119977
rect 675242 119965 675248 120017
rect 674128 118929 674134 118981
rect 674186 118969 674192 118981
rect 674416 118969 674422 118981
rect 674186 118941 674422 118969
rect 674186 118929 674192 118941
rect 674416 118929 674422 118941
rect 674474 118929 674480 118981
rect 144592 118559 144598 118611
rect 144650 118599 144656 118611
rect 191632 118599 191638 118611
rect 144650 118571 191638 118599
rect 144650 118559 144656 118571
rect 191632 118559 191638 118571
rect 191690 118559 191696 118611
rect 144592 118263 144598 118315
rect 144650 118303 144656 118315
rect 185872 118303 185878 118315
rect 144650 118275 185878 118303
rect 144650 118263 144656 118275
rect 185872 118263 185878 118275
rect 185930 118263 185936 118315
rect 144784 118115 144790 118167
rect 144842 118155 144848 118167
rect 209200 118155 209206 118167
rect 144842 118127 209206 118155
rect 144842 118115 144848 118127
rect 209200 118115 209206 118127
rect 209258 118115 209264 118167
rect 674608 118041 674614 118093
rect 674666 118081 674672 118093
rect 676816 118081 676822 118093
rect 674666 118053 676822 118081
rect 674666 118041 674672 118053
rect 676816 118041 676822 118053
rect 676874 118041 676880 118093
rect 144784 117967 144790 118019
rect 144842 118007 144848 118019
rect 146608 118007 146614 118019
rect 144842 117979 146614 118007
rect 144842 117967 144848 117979
rect 146608 117967 146614 117979
rect 146666 117967 146672 118019
rect 674416 117967 674422 118019
rect 674474 118007 674480 118019
rect 676912 118007 676918 118019
rect 674474 117979 676918 118007
rect 674474 117967 674480 117979
rect 676912 117967 676918 117979
rect 676970 117967 676976 118019
rect 146224 116635 146230 116687
rect 146282 116675 146288 116687
rect 146608 116675 146614 116687
rect 146282 116647 146614 116675
rect 146282 116635 146288 116647
rect 146608 116635 146614 116647
rect 146666 116635 146672 116687
rect 146224 115599 146230 115651
rect 146282 115639 146288 115651
rect 146282 115611 146846 115639
rect 146282 115599 146288 115611
rect 146818 115417 146846 115611
rect 146896 115417 146902 115429
rect 146818 115389 146902 115417
rect 146896 115377 146902 115389
rect 146954 115377 146960 115429
rect 146704 115303 146710 115355
rect 146762 115343 146768 115355
rect 209296 115343 209302 115355
rect 146762 115315 209302 115343
rect 146762 115303 146768 115315
rect 209296 115303 209302 115315
rect 209354 115303 209360 115355
rect 144592 115229 144598 115281
rect 144650 115269 144656 115281
rect 209392 115269 209398 115281
rect 144650 115241 209398 115269
rect 144650 115229 144656 115241
rect 209392 115229 209398 115241
rect 209450 115229 209456 115281
rect 146896 114899 146902 114911
rect 146434 114871 146902 114899
rect 146434 114159 146462 114871
rect 146896 114859 146902 114871
rect 146954 114859 146960 114911
rect 146512 114267 146518 114319
rect 146570 114307 146576 114319
rect 146992 114307 146998 114319
rect 146570 114279 146998 114307
rect 146570 114267 146576 114279
rect 146992 114267 146998 114279
rect 147050 114267 147056 114319
rect 146512 114159 146518 114171
rect 146434 114131 146518 114159
rect 146512 114119 146518 114131
rect 146570 114119 146576 114171
rect 674128 114119 674134 114171
rect 674186 114159 674192 114171
rect 675376 114159 675382 114171
rect 674186 114131 675382 114159
rect 674186 114119 674192 114131
rect 675376 114119 675382 114131
rect 675434 114119 675440 114171
rect 674032 113601 674038 113653
rect 674090 113641 674096 113653
rect 675184 113641 675190 113653
rect 674090 113613 675190 113641
rect 674090 113601 674096 113613
rect 675184 113601 675190 113613
rect 675242 113601 675248 113653
rect 674224 113305 674230 113357
rect 674282 113345 674288 113357
rect 675088 113345 675094 113357
rect 674282 113317 675094 113345
rect 674282 113305 674288 113317
rect 675088 113305 675094 113317
rect 675146 113305 675152 113357
rect 144784 113231 144790 113283
rect 144842 113271 144848 113283
rect 146896 113271 146902 113283
rect 144842 113243 146902 113271
rect 144842 113231 144848 113243
rect 146896 113231 146902 113243
rect 146954 113231 146960 113283
rect 647920 112861 647926 112913
rect 647978 112901 647984 112913
rect 665200 112901 665206 112913
rect 647978 112873 665206 112901
rect 647978 112861 647984 112873
rect 665200 112861 665206 112873
rect 665258 112861 665264 112913
rect 144592 112491 144598 112543
rect 144650 112531 144656 112543
rect 188752 112531 188758 112543
rect 144650 112503 188758 112531
rect 144650 112491 144656 112503
rect 188752 112491 188758 112503
rect 188810 112491 188816 112543
rect 144784 112417 144790 112469
rect 144842 112457 144848 112469
rect 203152 112457 203158 112469
rect 144842 112429 203158 112457
rect 144842 112417 144848 112429
rect 203152 112417 203158 112429
rect 203210 112417 203216 112469
rect 144592 112343 144598 112395
rect 144650 112383 144656 112395
rect 209488 112383 209494 112395
rect 144650 112355 209494 112383
rect 144650 112343 144656 112355
rect 209488 112343 209494 112355
rect 209546 112343 209552 112395
rect 674320 111159 674326 111211
rect 674378 111199 674384 111211
rect 675376 111199 675382 111211
rect 674378 111171 675382 111199
rect 674378 111159 674384 111171
rect 675376 111159 675382 111171
rect 675434 111159 675440 111211
rect 146512 111085 146518 111137
rect 146570 111125 146576 111137
rect 146570 111097 146654 111125
rect 146570 111085 146576 111097
rect 146224 110937 146230 110989
rect 146282 110977 146288 110989
rect 146512 110977 146518 110989
rect 146282 110949 146518 110977
rect 146282 110937 146288 110949
rect 146512 110937 146518 110949
rect 146570 110937 146576 110989
rect 146224 110789 146230 110841
rect 146282 110829 146288 110841
rect 146626 110829 146654 111097
rect 146282 110801 146654 110829
rect 146282 110789 146288 110801
rect 144784 109531 144790 109583
rect 144842 109571 144848 109583
rect 162832 109571 162838 109583
rect 144842 109543 162838 109571
rect 144842 109531 144848 109543
rect 162832 109531 162838 109543
rect 162890 109531 162896 109583
rect 144592 109457 144598 109509
rect 144650 109497 144656 109509
rect 182992 109497 182998 109509
rect 144650 109469 182998 109497
rect 144650 109457 144656 109469
rect 182992 109457 182998 109469
rect 183050 109457 183056 109509
rect 144784 109383 144790 109435
rect 144842 109423 144848 109435
rect 146032 109423 146038 109435
rect 144842 109395 146038 109423
rect 144842 109383 144848 109395
rect 146032 109383 146038 109395
rect 146090 109383 146096 109435
rect 144592 107459 144598 107511
rect 144650 107499 144656 107511
rect 160144 107499 160150 107511
rect 144650 107471 160150 107499
rect 144650 107459 144656 107471
rect 160144 107459 160150 107471
rect 160202 107459 160208 107511
rect 674512 107311 674518 107363
rect 674570 107351 674576 107363
rect 675376 107351 675382 107363
rect 674570 107323 675382 107351
rect 674570 107311 674576 107323
rect 675376 107311 675382 107323
rect 675434 107311 675440 107363
rect 674608 106941 674614 106993
rect 674666 106981 674672 106993
rect 675472 106981 675478 106993
rect 674666 106953 675478 106981
rect 674666 106941 674672 106953
rect 675472 106941 675478 106953
rect 675530 106941 675536 106993
rect 143920 106719 143926 106771
rect 143978 106759 143984 106771
rect 144784 106759 144790 106771
rect 143978 106731 144790 106759
rect 143978 106719 143984 106731
rect 144784 106719 144790 106731
rect 144842 106719 144848 106771
rect 146224 106685 146230 106697
rect 144802 106657 146230 106685
rect 144802 106623 144830 106657
rect 146224 106645 146230 106657
rect 146282 106645 146288 106697
rect 144784 106571 144790 106623
rect 144842 106571 144848 106623
rect 146032 106571 146038 106623
rect 146090 106611 146096 106623
rect 193936 106611 193942 106623
rect 146090 106583 193942 106611
rect 146090 106571 146096 106583
rect 193936 106571 193942 106583
rect 193994 106571 194000 106623
rect 144016 106497 144022 106549
rect 144074 106537 144080 106549
rect 146224 106537 146230 106549
rect 144074 106509 146230 106537
rect 144074 106497 144080 106509
rect 146224 106497 146230 106509
rect 146282 106497 146288 106549
rect 143920 106349 143926 106401
rect 143978 106389 143984 106401
rect 144304 106389 144310 106401
rect 143978 106361 144310 106389
rect 143978 106349 143984 106361
rect 144304 106349 144310 106361
rect 144362 106349 144368 106401
rect 673936 106127 673942 106179
rect 673994 106167 674000 106179
rect 675376 106167 675382 106179
rect 673994 106139 675382 106167
rect 673994 106127 674000 106139
rect 675376 106127 675382 106139
rect 675434 106127 675440 106179
rect 144112 105979 144118 106031
rect 144170 106019 144176 106031
rect 146032 106019 146038 106031
rect 144170 105991 146038 106019
rect 144170 105979 144176 105991
rect 146032 105979 146038 105991
rect 146090 105979 146096 106031
rect 674416 105165 674422 105217
rect 674474 105205 674480 105217
rect 675376 105205 675382 105217
rect 674474 105177 675382 105205
rect 674474 105165 674480 105177
rect 675376 105165 675382 105177
rect 675434 105165 675440 105217
rect 144016 104351 144022 104403
rect 144074 104391 144080 104403
rect 159952 104391 159958 104403
rect 144074 104363 159958 104391
rect 144074 104351 144080 104363
rect 159952 104351 159958 104363
rect 160010 104351 160016 104403
rect 144016 104203 144022 104255
rect 144074 104243 144080 104255
rect 157072 104243 157078 104255
rect 144074 104215 157078 104243
rect 144074 104203 144080 104215
rect 157072 104203 157078 104215
rect 157130 104203 157136 104255
rect 144112 103685 144118 103737
rect 144170 103725 144176 103737
rect 209584 103725 209590 103737
rect 144170 103697 209590 103725
rect 144170 103685 144176 103697
rect 209584 103685 209590 103697
rect 209642 103685 209648 103737
rect 146608 103611 146614 103663
rect 146666 103651 146672 103663
rect 201712 103651 201718 103663
rect 146666 103623 201718 103651
rect 146666 103611 146672 103623
rect 201712 103611 201718 103623
rect 201770 103611 201776 103663
rect 144784 103537 144790 103589
rect 144842 103577 144848 103589
rect 199984 103577 199990 103589
rect 144842 103549 199990 103577
rect 144842 103537 144848 103549
rect 199984 103537 199990 103549
rect 200042 103537 200048 103589
rect 146512 103463 146518 103515
rect 146570 103503 146576 103515
rect 210160 103503 210166 103515
rect 146570 103475 210166 103503
rect 146570 103463 146576 103475
rect 210160 103463 210166 103475
rect 210218 103463 210224 103515
rect 146704 103389 146710 103441
rect 146762 103429 146768 103441
rect 146992 103429 146998 103441
rect 146762 103401 146998 103429
rect 146762 103389 146768 103401
rect 146992 103389 146998 103401
rect 147050 103389 147056 103441
rect 144016 100873 144022 100925
rect 144074 100913 144080 100925
rect 149008 100913 149014 100925
rect 144074 100885 149014 100913
rect 144074 100873 144080 100885
rect 149008 100873 149014 100885
rect 149066 100873 149072 100925
rect 144112 100799 144118 100851
rect 144170 100839 144176 100851
rect 209680 100839 209686 100851
rect 144170 100811 209686 100839
rect 144170 100799 144176 100811
rect 209680 100799 209686 100811
rect 209738 100799 209744 100851
rect 201808 100765 201814 100777
rect 144322 100737 201814 100765
rect 144322 100703 144350 100737
rect 201808 100725 201814 100737
rect 201866 100725 201872 100777
rect 144304 100651 144310 100703
rect 144362 100651 144368 100703
rect 146896 100651 146902 100703
rect 146954 100691 146960 100703
rect 201616 100691 201622 100703
rect 146954 100663 201622 100691
rect 146954 100651 146960 100663
rect 201616 100651 201622 100663
rect 201674 100651 201680 100703
rect 151120 100577 151126 100629
rect 151178 100617 151184 100629
rect 201712 100617 201718 100629
rect 151178 100589 201718 100617
rect 151178 100577 151184 100589
rect 201712 100577 201718 100589
rect 201770 100577 201776 100629
rect 159760 100503 159766 100555
rect 159818 100543 159824 100555
rect 210160 100543 210166 100555
rect 159818 100515 210166 100543
rect 159818 100503 159824 100515
rect 210160 100503 210166 100515
rect 210218 100503 210224 100555
rect 185680 100429 185686 100481
rect 185738 100469 185744 100481
rect 201712 100469 201718 100481
rect 185738 100441 201718 100469
rect 185738 100429 185744 100441
rect 201712 100429 201718 100441
rect 201770 100429 201776 100481
rect 144016 98283 144022 98335
rect 144074 98323 144080 98335
rect 160048 98323 160054 98335
rect 144074 98295 160054 98323
rect 144074 98283 144080 98295
rect 160048 98283 160054 98295
rect 160106 98283 160112 98335
rect 144016 97987 144022 98039
rect 144074 98027 144080 98039
rect 177232 98027 177238 98039
rect 144074 97999 177238 98027
rect 144074 97987 144080 97999
rect 177232 97987 177238 97999
rect 177290 97987 177296 98039
rect 144112 97913 144118 97965
rect 144170 97953 144176 97965
rect 180112 97953 180118 97965
rect 144170 97925 180118 97953
rect 144170 97913 144176 97925
rect 180112 97913 180118 97925
rect 180170 97913 180176 97965
rect 156880 97765 156886 97817
rect 156938 97805 156944 97817
rect 210160 97805 210166 97817
rect 156938 97777 210166 97805
rect 156938 97765 156944 97777
rect 210160 97765 210166 97777
rect 210218 97765 210224 97817
rect 168496 97691 168502 97743
rect 168554 97731 168560 97743
rect 201808 97731 201814 97743
rect 168554 97703 201814 97731
rect 168554 97691 168560 97703
rect 201808 97691 201814 97703
rect 201866 97691 201872 97743
rect 171376 97617 171382 97669
rect 171434 97657 171440 97669
rect 201616 97657 201622 97669
rect 171434 97629 201622 97657
rect 171434 97617 171440 97629
rect 201616 97617 201622 97629
rect 201674 97617 201680 97669
rect 174256 97543 174262 97595
rect 174314 97583 174320 97595
rect 201712 97583 201718 97595
rect 174314 97555 201718 97583
rect 174314 97543 174320 97555
rect 201712 97543 201718 97555
rect 201770 97543 201776 97595
rect 154000 97469 154006 97521
rect 154058 97509 154064 97521
rect 210160 97509 210166 97521
rect 154058 97481 210166 97509
rect 154058 97469 154064 97481
rect 210160 97469 210166 97481
rect 210218 97469 210224 97521
rect 663184 96433 663190 96485
rect 663242 96473 663248 96485
rect 665200 96473 665206 96485
rect 663242 96445 665206 96473
rect 663242 96433 663248 96445
rect 665200 96433 665206 96445
rect 665258 96433 665264 96485
rect 144400 95397 144406 95449
rect 144458 95437 144464 95449
rect 146608 95437 146614 95449
rect 144458 95409 146614 95437
rect 144458 95397 144464 95409
rect 146608 95397 146614 95409
rect 146666 95397 146672 95449
rect 146512 95101 146518 95153
rect 146570 95141 146576 95153
rect 171568 95141 171574 95153
rect 146570 95113 171574 95141
rect 146570 95101 146576 95113
rect 171568 95101 171574 95113
rect 171626 95101 171632 95153
rect 144016 95027 144022 95079
rect 144074 95067 144080 95079
rect 174448 95067 174454 95079
rect 144074 95039 174454 95067
rect 144074 95027 144080 95039
rect 174448 95027 174454 95039
rect 174506 95027 174512 95079
rect 162736 94879 162742 94931
rect 162794 94919 162800 94931
rect 201712 94919 201718 94931
rect 162794 94891 201718 94919
rect 162794 94879 162800 94891
rect 201712 94879 201718 94891
rect 201770 94879 201776 94931
rect 165616 94805 165622 94857
rect 165674 94845 165680 94857
rect 210160 94845 210166 94857
rect 165674 94817 210166 94845
rect 165674 94805 165680 94817
rect 210160 94805 210166 94817
rect 210218 94805 210224 94857
rect 144592 94657 144598 94709
rect 144650 94697 144656 94709
rect 201616 94697 201622 94709
rect 144650 94669 201622 94697
rect 144650 94657 144656 94669
rect 201616 94657 201622 94669
rect 201674 94657 201680 94709
rect 193936 94065 193942 94117
rect 193994 94105 194000 94117
rect 209584 94105 209590 94117
rect 193994 94077 209590 94105
rect 193994 94065 194000 94077
rect 209584 94065 209590 94077
rect 209642 94065 209648 94117
rect 646480 92659 646486 92711
rect 646538 92699 646544 92711
rect 659824 92699 659830 92711
rect 646538 92671 659830 92699
rect 646538 92659 646544 92671
rect 659824 92659 659830 92671
rect 659882 92659 659888 92711
rect 647536 92585 647542 92637
rect 647594 92625 647600 92637
rect 661744 92625 661750 92637
rect 647594 92597 661750 92625
rect 647594 92585 647600 92597
rect 661744 92585 661750 92597
rect 661802 92585 661808 92637
rect 647344 92511 647350 92563
rect 647402 92551 647408 92563
rect 660688 92551 660694 92563
rect 647402 92523 660694 92551
rect 647402 92511 647408 92523
rect 660688 92511 660694 92523
rect 660746 92511 660752 92563
rect 646096 92437 646102 92489
rect 646154 92477 646160 92489
rect 663088 92477 663094 92489
rect 646154 92449 663094 92477
rect 646154 92437 646160 92449
rect 663088 92437 663094 92449
rect 663146 92437 663152 92489
rect 647824 92289 647830 92341
rect 647882 92329 647888 92341
rect 662512 92329 662518 92341
rect 647882 92301 662518 92329
rect 647882 92289 647888 92301
rect 662512 92289 662518 92301
rect 662570 92289 662576 92341
rect 144112 92215 144118 92267
rect 144170 92255 144176 92267
rect 154000 92255 154006 92267
rect 144170 92227 154006 92255
rect 144170 92215 144176 92227
rect 154000 92215 154006 92227
rect 154058 92215 154064 92267
rect 647248 92215 647254 92267
rect 647306 92255 647312 92267
rect 661168 92255 661174 92267
rect 647306 92227 661174 92255
rect 647306 92215 647312 92227
rect 661168 92215 661174 92227
rect 661226 92215 661232 92267
rect 144016 92141 144022 92193
rect 144074 92181 144080 92193
rect 168496 92181 168502 92193
rect 144074 92153 168502 92181
rect 144074 92141 144080 92153
rect 168496 92141 168502 92153
rect 168554 92141 168560 92193
rect 646576 92141 646582 92193
rect 646634 92181 646640 92193
rect 658864 92181 658870 92193
rect 646634 92153 658870 92181
rect 646634 92141 646640 92153
rect 658864 92141 658870 92153
rect 658922 92141 658928 92193
rect 146224 92067 146230 92119
rect 146282 92107 146288 92119
rect 201712 92107 201718 92119
rect 146282 92079 201718 92107
rect 146282 92067 146288 92079
rect 201712 92067 201718 92079
rect 201770 92067 201776 92119
rect 146032 91993 146038 92045
rect 146090 92033 146096 92045
rect 197680 92033 197686 92045
rect 146090 92005 197686 92033
rect 146090 91993 146096 92005
rect 197680 91993 197686 92005
rect 197738 91993 197744 92045
rect 151216 91919 151222 91971
rect 151274 91959 151280 91971
rect 201616 91959 201622 91971
rect 151274 91931 201622 91959
rect 151274 91919 151280 91931
rect 201616 91919 201622 91931
rect 201674 91919 201680 91971
rect 185776 91845 185782 91897
rect 185834 91885 185840 91897
rect 201808 91885 201814 91897
rect 185834 91857 201814 91885
rect 185834 91845 185840 91857
rect 201808 91845 201814 91857
rect 201866 91845 201872 91897
rect 144112 91179 144118 91231
rect 144170 91219 144176 91231
rect 144304 91219 144310 91231
rect 144170 91191 144310 91219
rect 144170 91179 144176 91191
rect 144304 91179 144310 91191
rect 144362 91179 144368 91231
rect 144016 89403 144022 89455
rect 144074 89443 144080 89455
rect 151120 89443 151126 89455
rect 144074 89415 151126 89443
rect 144074 89403 144080 89415
rect 151120 89403 151126 89415
rect 151178 89403 151184 89455
rect 144112 89329 144118 89381
rect 144170 89369 144176 89381
rect 163120 89369 163126 89381
rect 144170 89341 163126 89369
rect 144170 89329 144176 89341
rect 163120 89329 163126 89341
rect 163178 89329 163184 89381
rect 146224 89255 146230 89307
rect 146282 89295 146288 89307
rect 165808 89295 165814 89307
rect 146282 89267 165814 89295
rect 146282 89255 146288 89267
rect 165808 89255 165814 89267
rect 165866 89255 165872 89307
rect 144112 89181 144118 89233
rect 144170 89221 144176 89233
rect 144784 89221 144790 89233
rect 144170 89193 144790 89221
rect 144170 89181 144176 89193
rect 144784 89181 144790 89193
rect 144842 89181 144848 89233
rect 156976 89181 156982 89233
rect 157034 89221 157040 89233
rect 201808 89221 201814 89233
rect 157034 89193 201814 89221
rect 157034 89181 157040 89193
rect 201808 89181 201814 89193
rect 201866 89181 201872 89233
rect 159856 89107 159862 89159
rect 159914 89147 159920 89159
rect 201616 89147 201622 89159
rect 159914 89119 201622 89147
rect 159914 89107 159920 89119
rect 201616 89107 201622 89119
rect 201674 89107 201680 89159
rect 182896 89033 182902 89085
rect 182954 89073 182960 89085
rect 201520 89073 201526 89085
rect 182954 89045 201526 89073
rect 182954 89033 182960 89045
rect 201520 89033 201526 89045
rect 201578 89033 201584 89085
rect 188656 88959 188662 89011
rect 188714 88999 188720 89011
rect 198736 88999 198742 89011
rect 188714 88971 198742 88999
rect 188714 88959 188720 88971
rect 198736 88959 198742 88971
rect 198794 88959 198800 89011
rect 191536 88885 191542 88937
rect 191594 88925 191600 88937
rect 201712 88925 201718 88937
rect 191594 88897 201718 88925
rect 191594 88885 191600 88897
rect 201712 88885 201718 88897
rect 201770 88885 201776 88937
rect 646288 87553 646294 87605
rect 646346 87593 646352 87605
rect 650992 87593 650998 87605
rect 646346 87565 650998 87593
rect 646346 87553 646352 87565
rect 650992 87553 650998 87565
rect 651050 87553 651056 87605
rect 652336 87331 652342 87383
rect 652394 87371 652400 87383
rect 659344 87371 659350 87383
rect 652394 87343 659350 87371
rect 652394 87331 652400 87343
rect 659344 87331 659350 87343
rect 659402 87331 659408 87383
rect 658000 87297 658006 87309
rect 657058 87269 658006 87297
rect 657058 87161 657086 87269
rect 658000 87257 658006 87269
rect 658058 87257 658064 87309
rect 657040 87109 657046 87161
rect 657098 87109 657104 87161
rect 647920 87035 647926 87087
rect 647978 87075 647984 87087
rect 663280 87075 663286 87087
rect 647978 87047 663286 87075
rect 647978 87035 647984 87047
rect 663280 87035 663286 87047
rect 663338 87035 663344 87087
rect 646384 86739 646390 86791
rect 646442 86779 646448 86791
rect 651088 86779 651094 86791
rect 646442 86751 651094 86779
rect 646442 86739 646448 86751
rect 651088 86739 651094 86751
rect 651146 86739 651152 86791
rect 144016 86443 144022 86495
rect 144074 86483 144080 86495
rect 162736 86483 162742 86495
rect 144074 86455 162742 86483
rect 144074 86443 144080 86455
rect 162736 86443 162742 86455
rect 162794 86443 162800 86495
rect 144592 86369 144598 86421
rect 144650 86409 144656 86421
rect 144880 86409 144886 86421
rect 144650 86381 144886 86409
rect 144650 86369 144656 86381
rect 144880 86369 144886 86381
rect 144938 86369 144944 86421
rect 154096 86369 154102 86421
rect 154154 86409 154160 86421
rect 201904 86409 201910 86421
rect 154154 86381 201910 86409
rect 154154 86369 154160 86381
rect 201904 86369 201910 86381
rect 201962 86369 201968 86421
rect 171472 86295 171478 86347
rect 171530 86335 171536 86347
rect 201520 86335 201526 86347
rect 171530 86307 201526 86335
rect 171530 86295 171536 86307
rect 201520 86295 201526 86307
rect 201578 86295 201584 86347
rect 174352 86221 174358 86273
rect 174410 86261 174416 86273
rect 201808 86261 201814 86273
rect 174410 86233 201814 86261
rect 174410 86221 174416 86233
rect 201808 86221 201814 86233
rect 201866 86221 201872 86273
rect 177136 86147 177142 86199
rect 177194 86187 177200 86199
rect 201616 86187 201622 86199
rect 177194 86159 201622 86187
rect 177194 86147 177200 86159
rect 201616 86147 201622 86159
rect 201674 86147 201680 86199
rect 180016 86073 180022 86125
rect 180074 86113 180080 86125
rect 201712 86113 201718 86125
rect 180074 86085 201718 86113
rect 180074 86073 180080 86085
rect 201712 86073 201718 86085
rect 201770 86073 201776 86125
rect 144016 84963 144022 85015
rect 144074 85003 144080 85015
rect 201712 85003 201718 85015
rect 144074 84975 201718 85003
rect 144074 84963 144080 84975
rect 201712 84963 201718 84975
rect 201770 84963 201776 85015
rect 646480 84889 646486 84941
rect 646538 84929 646544 84941
rect 650896 84929 650902 84941
rect 646538 84901 650902 84929
rect 646538 84889 646544 84901
rect 650896 84889 650902 84901
rect 650954 84889 650960 84941
rect 145936 83631 145942 83683
rect 145994 83671 146000 83683
rect 146224 83671 146230 83683
rect 145994 83643 146230 83671
rect 145994 83631 146000 83643
rect 146224 83631 146230 83643
rect 146282 83631 146288 83683
rect 151312 83483 151318 83535
rect 151370 83523 151376 83535
rect 194608 83523 194614 83535
rect 151370 83495 194614 83523
rect 151370 83483 151376 83495
rect 194608 83483 194614 83495
rect 194666 83483 194672 83535
rect 162928 83409 162934 83461
rect 162986 83449 162992 83461
rect 201616 83449 201622 83461
rect 162986 83421 201622 83449
rect 162986 83409 162992 83421
rect 201616 83409 201622 83421
rect 201674 83409 201680 83461
rect 165712 83335 165718 83387
rect 165770 83375 165776 83387
rect 201712 83375 201718 83387
rect 165770 83347 201718 83375
rect 165770 83335 165776 83347
rect 201712 83335 201718 83347
rect 201770 83335 201776 83387
rect 168592 83261 168598 83313
rect 168650 83301 168656 83313
rect 201040 83301 201046 83313
rect 168650 83273 201046 83301
rect 168650 83261 168656 83273
rect 201040 83261 201046 83273
rect 201098 83261 201104 83313
rect 646288 83113 646294 83165
rect 646346 83153 646352 83165
rect 657040 83153 657046 83165
rect 646346 83125 657046 83153
rect 646346 83113 646352 83125
rect 657040 83113 657046 83125
rect 657098 83113 657104 83165
rect 144016 82077 144022 82129
rect 144074 82117 144080 82129
rect 197776 82117 197782 82129
rect 144074 82089 197782 82117
rect 144074 82077 144080 82089
rect 197776 82077 197782 82089
rect 197834 82077 197840 82129
rect 646096 81855 646102 81907
rect 646154 81895 646160 81907
rect 663280 81895 663286 81907
rect 646154 81867 663286 81895
rect 646154 81855 646160 81867
rect 663280 81855 663286 81867
rect 663338 81855 663344 81907
rect 646000 81781 646006 81833
rect 646058 81821 646064 81833
rect 663376 81821 663382 81833
rect 646058 81793 663382 81821
rect 646058 81781 646064 81793
rect 663376 81781 663382 81793
rect 663434 81781 663440 81833
rect 647632 81633 647638 81685
rect 647690 81673 647696 81685
rect 661072 81673 661078 81685
rect 647690 81645 661078 81673
rect 647690 81633 647696 81645
rect 661072 81633 661078 81645
rect 661130 81633 661136 81685
rect 647920 81411 647926 81463
rect 647978 81451 647984 81463
rect 657520 81451 657526 81463
rect 647978 81423 657526 81451
rect 647978 81411 647984 81423
rect 657520 81411 657526 81423
rect 657578 81411 657584 81463
rect 144016 80745 144022 80797
rect 144074 80785 144080 80797
rect 163024 80785 163030 80797
rect 144074 80757 163030 80785
rect 144074 80745 144080 80757
rect 163024 80745 163030 80757
rect 163082 80745 163088 80797
rect 144112 80671 144118 80723
rect 144170 80711 144176 80723
rect 144688 80711 144694 80723
rect 144170 80683 144694 80711
rect 144170 80671 144176 80683
rect 144688 80671 144694 80683
rect 144746 80671 144752 80723
rect 659440 80671 659446 80723
rect 659498 80711 659504 80723
rect 659536 80711 659542 80723
rect 659498 80683 659542 80711
rect 659498 80671 659504 80683
rect 659536 80671 659542 80683
rect 659594 80671 659600 80723
rect 185872 80597 185878 80649
rect 185930 80637 185936 80649
rect 201712 80637 201718 80649
rect 185930 80609 201718 80637
rect 185930 80597 185936 80609
rect 201712 80597 201718 80609
rect 201770 80597 201776 80649
rect 191632 80523 191638 80575
rect 191690 80563 191696 80575
rect 200368 80563 200374 80575
rect 191690 80535 200374 80563
rect 191690 80523 191696 80535
rect 200368 80523 200374 80535
rect 200426 80523 200432 80575
rect 646864 80227 646870 80279
rect 646922 80267 646928 80279
rect 656944 80267 656950 80279
rect 646922 80239 656950 80267
rect 646922 80227 646928 80239
rect 656944 80227 656950 80239
rect 657002 80227 657008 80279
rect 647920 79339 647926 79391
rect 647978 79379 647984 79391
rect 660688 79379 660694 79391
rect 647978 79351 660694 79379
rect 647978 79339 647984 79351
rect 660688 79339 660694 79351
rect 660746 79339 660752 79391
rect 640720 79191 640726 79243
rect 640778 79231 640784 79243
rect 663184 79231 663190 79243
rect 640778 79203 663190 79231
rect 640778 79191 640784 79203
rect 663184 79191 663190 79203
rect 663242 79191 663248 79243
rect 646864 78895 646870 78947
rect 646922 78935 646928 78947
rect 658864 78935 658870 78947
rect 646922 78907 658870 78935
rect 646922 78895 646928 78907
rect 658864 78895 658870 78907
rect 658922 78895 658928 78947
rect 646864 78303 646870 78355
rect 646922 78343 646928 78355
rect 651184 78343 651190 78355
rect 646922 78315 651190 78343
rect 646922 78303 646928 78315
rect 651184 78303 651190 78315
rect 651242 78303 651248 78355
rect 646480 78229 646486 78281
rect 646538 78269 646544 78281
rect 662512 78269 662518 78281
rect 646538 78241 662518 78269
rect 646538 78229 646544 78241
rect 662512 78229 662518 78241
rect 662570 78229 662576 78281
rect 144016 77859 144022 77911
rect 144074 77899 144080 77911
rect 165616 77899 165622 77911
rect 144074 77871 165622 77899
rect 144074 77859 144080 77871
rect 165616 77859 165622 77871
rect 165674 77859 165680 77911
rect 144112 77785 144118 77837
rect 144170 77825 144176 77837
rect 185680 77825 185686 77837
rect 144170 77797 185686 77825
rect 144170 77785 144176 77797
rect 185680 77785 185686 77797
rect 185738 77785 185744 77837
rect 149008 77711 149014 77763
rect 149066 77751 149072 77763
rect 201520 77751 201526 77763
rect 149066 77723 201526 77751
rect 149066 77711 149072 77723
rect 201520 77711 201526 77723
rect 201578 77711 201584 77763
rect 647920 77711 647926 77763
rect 647978 77751 647984 77763
rect 662896 77751 662902 77763
rect 647978 77723 662902 77751
rect 647978 77711 647984 77723
rect 662896 77711 662902 77723
rect 662954 77711 662960 77763
rect 157072 77637 157078 77689
rect 157130 77677 157136 77689
rect 201808 77677 201814 77689
rect 157130 77649 201814 77677
rect 157130 77637 157136 77649
rect 201808 77637 201814 77649
rect 201866 77637 201872 77689
rect 646672 77637 646678 77689
rect 646730 77677 646736 77689
rect 658288 77677 658294 77689
rect 646730 77649 658294 77677
rect 646730 77637 646736 77649
rect 658288 77637 658294 77649
rect 658346 77637 658352 77689
rect 160144 77563 160150 77615
rect 160202 77603 160208 77615
rect 195568 77603 195574 77615
rect 160202 77575 195574 77603
rect 160202 77563 160208 77575
rect 195568 77563 195574 77575
rect 195626 77563 195632 77615
rect 646288 77563 646294 77615
rect 646346 77603 646352 77615
rect 650896 77603 650902 77615
rect 646346 77575 650902 77603
rect 646346 77563 646352 77575
rect 650896 77563 650902 77575
rect 650954 77563 650960 77615
rect 182992 77489 182998 77541
rect 183050 77529 183056 77541
rect 201616 77529 201622 77541
rect 183050 77501 201622 77529
rect 183050 77489 183056 77501
rect 201616 77489 201622 77501
rect 201674 77489 201680 77541
rect 647824 77489 647830 77541
rect 647882 77529 647888 77541
rect 650992 77529 650998 77541
rect 647882 77501 650998 77529
rect 647882 77489 647888 77501
rect 650992 77489 650998 77501
rect 651050 77489 651056 77541
rect 185680 77415 185686 77467
rect 185738 77455 185744 77467
rect 201712 77455 201718 77467
rect 185738 77427 201718 77455
rect 185738 77415 185744 77427
rect 201712 77415 201718 77427
rect 201770 77415 201776 77467
rect 647440 77415 647446 77467
rect 647498 77455 647504 77467
rect 659440 77455 659446 77467
rect 647498 77427 659446 77455
rect 647498 77415 647504 77427
rect 659440 77415 659446 77427
rect 659498 77415 659504 77467
rect 188752 77341 188758 77393
rect 188810 77381 188816 77393
rect 210256 77381 210262 77393
rect 188810 77353 210262 77381
rect 188810 77341 188816 77353
rect 210256 77341 210262 77353
rect 210314 77341 210320 77393
rect 144112 76527 144118 76579
rect 144170 76567 144176 76579
rect 144592 76567 144598 76579
rect 144170 76539 144598 76567
rect 144170 76527 144176 76539
rect 144592 76527 144598 76539
rect 144650 76527 144656 76579
rect 144400 76453 144406 76505
rect 144458 76493 144464 76505
rect 144458 76465 144542 76493
rect 144458 76453 144464 76465
rect 144208 76305 144214 76357
rect 144266 76345 144272 76357
rect 144400 76345 144406 76357
rect 144266 76317 144406 76345
rect 144266 76305 144272 76317
rect 144400 76305 144406 76317
rect 144458 76305 144464 76357
rect 144514 76197 144542 76465
rect 144592 76305 144598 76357
rect 144650 76345 144656 76357
rect 145168 76345 145174 76357
rect 144650 76317 145174 76345
rect 144650 76305 144656 76317
rect 145168 76305 145174 76317
rect 145226 76305 145232 76357
rect 144784 76231 144790 76283
rect 144842 76271 144848 76283
rect 146032 76271 146038 76283
rect 144842 76243 146038 76271
rect 144842 76231 144848 76243
rect 146032 76231 146038 76243
rect 146090 76231 146096 76283
rect 145168 76197 145174 76209
rect 144514 76169 145174 76197
rect 145168 76157 145174 76169
rect 145226 76157 145232 76209
rect 647920 76083 647926 76135
rect 647978 76123 647984 76135
rect 661744 76123 661750 76135
rect 647978 76095 661750 76123
rect 647978 76083 647984 76095
rect 661744 76083 661750 76095
rect 661802 76083 661808 76135
rect 646480 75639 646486 75691
rect 646538 75679 646544 75691
rect 656848 75679 656854 75691
rect 646538 75651 656854 75679
rect 646538 75639 646544 75651
rect 656848 75639 656854 75651
rect 656906 75639 656912 75691
rect 144112 74973 144118 75025
rect 144170 75013 144176 75025
rect 160144 75013 160150 75025
rect 144170 74985 160150 75013
rect 144170 74973 144176 74985
rect 160144 74973 160150 74985
rect 160202 74973 160208 75025
rect 144016 74899 144022 74951
rect 144074 74939 144080 74951
rect 155536 74939 155542 74951
rect 144074 74911 155542 74939
rect 144074 74899 144080 74911
rect 155536 74899 155542 74911
rect 155594 74899 155600 74951
rect 144112 74825 144118 74877
rect 144170 74865 144176 74877
rect 208720 74865 208726 74877
rect 144170 74837 208726 74865
rect 144170 74825 144176 74837
rect 208720 74825 208726 74837
rect 208778 74825 208784 74877
rect 154000 74751 154006 74803
rect 154058 74791 154064 74803
rect 201712 74791 201718 74803
rect 154058 74763 201718 74791
rect 154058 74751 154064 74763
rect 201712 74751 201718 74763
rect 201770 74751 201776 74803
rect 171568 74677 171574 74729
rect 171626 74717 171632 74729
rect 200944 74717 200950 74729
rect 171626 74689 200950 74717
rect 171626 74677 171632 74689
rect 200944 74677 200950 74689
rect 201002 74677 201008 74729
rect 174448 74603 174454 74655
rect 174506 74643 174512 74655
rect 198352 74643 198358 74655
rect 174506 74615 198358 74643
rect 174506 74603 174512 74615
rect 198352 74603 198358 74615
rect 198410 74603 198416 74655
rect 177232 74529 177238 74581
rect 177290 74569 177296 74581
rect 201040 74569 201046 74581
rect 177290 74541 201046 74569
rect 177290 74529 177296 74541
rect 201040 74529 201046 74541
rect 201098 74529 201104 74581
rect 180112 74455 180118 74507
rect 180170 74495 180176 74507
rect 210256 74495 210262 74507
rect 180170 74467 210262 74495
rect 180170 74455 180176 74467
rect 210256 74455 210262 74467
rect 210314 74455 210320 74507
rect 144784 72679 144790 72731
rect 144842 72719 144848 72731
rect 145360 72719 145366 72731
rect 144842 72691 145366 72719
rect 144842 72679 144848 72691
rect 145360 72679 145366 72691
rect 145418 72679 145424 72731
rect 144112 72605 144118 72657
rect 144170 72645 144176 72657
rect 144304 72645 144310 72657
rect 144170 72617 144310 72645
rect 144170 72605 144176 72617
rect 144304 72605 144310 72617
rect 144362 72605 144368 72657
rect 145360 72531 145366 72583
rect 145418 72571 145424 72583
rect 146800 72571 146806 72583
rect 145418 72543 146806 72571
rect 145418 72531 145424 72543
rect 146800 72531 146806 72543
rect 146858 72531 146864 72583
rect 646288 72531 646294 72583
rect 646346 72571 646352 72583
rect 663280 72571 663286 72583
rect 646346 72543 663286 72571
rect 646346 72531 646352 72543
rect 663280 72531 663286 72543
rect 663338 72531 663344 72583
rect 144304 72457 144310 72509
rect 144362 72497 144368 72509
rect 146224 72497 146230 72509
rect 144362 72469 146230 72497
rect 144362 72457 144368 72469
rect 146224 72457 146230 72469
rect 146282 72457 146288 72509
rect 646096 72383 646102 72435
rect 646154 72423 646160 72435
rect 663472 72423 663478 72435
rect 646154 72395 663478 72423
rect 646154 72383 646160 72395
rect 663472 72383 663478 72395
rect 663530 72383 663536 72435
rect 146224 72309 146230 72361
rect 146282 72349 146288 72361
rect 146512 72349 146518 72361
rect 146282 72321 146518 72349
rect 146282 72309 146288 72321
rect 146512 72309 146518 72321
rect 146570 72309 146576 72361
rect 145168 72161 145174 72213
rect 145226 72201 145232 72213
rect 146512 72201 146518 72213
rect 145226 72173 146518 72201
rect 145226 72161 145232 72173
rect 146512 72161 146518 72173
rect 146570 72161 146576 72213
rect 647152 72161 647158 72213
rect 647210 72201 647216 72213
rect 660112 72201 660118 72213
rect 647210 72173 660118 72201
rect 647210 72161 647216 72173
rect 660112 72161 660118 72173
rect 660170 72161 660176 72213
rect 144016 72013 144022 72065
rect 144074 72053 144080 72065
rect 154096 72053 154102 72065
rect 144074 72025 154102 72053
rect 144074 72013 144080 72025
rect 154096 72013 154102 72025
rect 154154 72013 154160 72065
rect 146896 71939 146902 71991
rect 146954 71979 146960 71991
rect 200464 71979 200470 71991
rect 146954 71951 200470 71979
rect 146954 71939 146960 71951
rect 200464 71939 200470 71951
rect 200522 71939 200528 71991
rect 208624 71939 208630 71991
rect 208682 71979 208688 71991
rect 209200 71979 209206 71991
rect 208682 71951 209206 71979
rect 208682 71939 208688 71951
rect 209200 71939 209206 71951
rect 209258 71939 209264 71991
rect 151120 71865 151126 71917
rect 151178 71905 151184 71917
rect 201808 71905 201814 71917
rect 151178 71877 201814 71905
rect 151178 71865 151184 71877
rect 201808 71865 201814 71877
rect 201866 71865 201872 71917
rect 163120 71791 163126 71843
rect 163178 71831 163184 71843
rect 201616 71831 201622 71843
rect 163178 71803 201622 71831
rect 163178 71791 163184 71803
rect 201616 71791 201622 71803
rect 201674 71791 201680 71843
rect 165808 71717 165814 71769
rect 165866 71757 165872 71769
rect 209968 71757 209974 71769
rect 165866 71729 209974 71757
rect 165866 71717 165872 71729
rect 209968 71717 209974 71729
rect 210026 71717 210032 71769
rect 168496 71643 168502 71695
rect 168554 71683 168560 71695
rect 201712 71683 201718 71695
rect 168554 71655 201718 71683
rect 168554 71643 168560 71655
rect 201712 71643 201718 71655
rect 201770 71643 201776 71695
rect 144016 70237 144022 70289
rect 144074 70277 144080 70289
rect 149776 70277 149782 70289
rect 144074 70249 149782 70277
rect 144074 70237 144080 70249
rect 149776 70237 149782 70249
rect 149834 70237 149840 70289
rect 145168 69497 145174 69549
rect 145226 69537 145232 69549
rect 145552 69537 145558 69549
rect 145226 69509 145558 69537
rect 145226 69497 145232 69509
rect 145552 69497 145558 69509
rect 145610 69497 145616 69549
rect 144208 69349 144214 69401
rect 144266 69389 144272 69401
rect 145552 69389 145558 69401
rect 144266 69361 145558 69389
rect 144266 69349 144272 69361
rect 145552 69349 145558 69361
rect 145610 69349 145616 69401
rect 144016 69127 144022 69179
rect 144074 69167 144080 69179
rect 144074 69139 146942 69167
rect 144074 69127 144080 69139
rect 146914 69093 146942 69139
rect 201520 69093 201526 69105
rect 146914 69065 201526 69093
rect 201520 69053 201526 69065
rect 201578 69053 201584 69105
rect 149776 68979 149782 69031
rect 149834 69019 149840 69031
rect 201808 69019 201814 69031
rect 149834 68991 201814 69019
rect 149834 68979 149840 68991
rect 201808 68979 201814 68991
rect 201866 68979 201872 69031
rect 154096 68905 154102 68957
rect 154154 68945 154160 68957
rect 201616 68945 201622 68957
rect 154154 68917 201622 68945
rect 154154 68905 154160 68917
rect 201616 68905 201622 68917
rect 201674 68905 201680 68957
rect 155536 68831 155542 68883
rect 155594 68871 155600 68883
rect 201712 68871 201718 68883
rect 155594 68843 201718 68871
rect 155594 68831 155600 68843
rect 201712 68831 201718 68843
rect 201770 68831 201776 68883
rect 160144 68757 160150 68809
rect 160202 68797 160208 68809
rect 194704 68797 194710 68809
rect 160202 68769 194710 68797
rect 160202 68757 160208 68769
rect 194704 68757 194710 68769
rect 194762 68757 194768 68809
rect 144016 66981 144022 67033
rect 144074 67021 144080 67033
rect 152656 67021 152662 67033
rect 144074 66993 152662 67021
rect 144074 66981 144080 66993
rect 152656 66981 152662 66993
rect 152714 66981 152720 67033
rect 144208 66537 144214 66589
rect 144266 66577 144272 66589
rect 158320 66577 158326 66589
rect 144266 66549 158326 66577
rect 144266 66537 144272 66549
rect 158320 66537 158326 66549
rect 158378 66537 158384 66589
rect 144880 66315 144886 66367
rect 144938 66355 144944 66367
rect 145552 66355 145558 66367
rect 144938 66327 145558 66355
rect 144938 66315 144944 66327
rect 145552 66315 145558 66327
rect 145610 66315 145616 66367
rect 144016 66241 144022 66293
rect 144074 66281 144080 66293
rect 144074 66253 149822 66281
rect 144074 66241 144080 66253
rect 144208 66167 144214 66219
rect 144266 66207 144272 66219
rect 144688 66207 144694 66219
rect 144266 66179 144694 66207
rect 144266 66167 144272 66179
rect 144688 66167 144694 66179
rect 144746 66167 144752 66219
rect 149794 66207 149822 66253
rect 200176 66207 200182 66219
rect 149794 66179 200182 66207
rect 200176 66167 200182 66179
rect 200234 66167 200240 66219
rect 152656 66093 152662 66145
rect 152714 66133 152720 66145
rect 201712 66133 201718 66145
rect 152714 66105 201718 66133
rect 152714 66093 152720 66105
rect 201712 66093 201718 66105
rect 201770 66093 201776 66145
rect 145552 66019 145558 66071
rect 145610 66059 145616 66071
rect 145840 66059 145846 66071
rect 145610 66031 145846 66059
rect 145610 66019 145616 66031
rect 145840 66019 145846 66031
rect 145898 66019 145904 66071
rect 158320 66019 158326 66071
rect 158378 66059 158384 66071
rect 201616 66059 201622 66071
rect 158378 66031 201622 66059
rect 158378 66019 158384 66031
rect 201616 66019 201622 66031
rect 201674 66019 201680 66071
rect 146032 65575 146038 65627
rect 146090 65615 146096 65627
rect 146224 65615 146230 65627
rect 146090 65587 146230 65615
rect 146090 65575 146096 65587
rect 146224 65575 146230 65587
rect 146282 65575 146288 65627
rect 146224 64835 146230 64887
rect 146282 64875 146288 64887
rect 201712 64875 201718 64887
rect 146282 64847 201718 64875
rect 146282 64835 146288 64847
rect 201712 64835 201718 64847
rect 201770 64835 201776 64887
rect 144016 64761 144022 64813
rect 144074 64801 144080 64813
rect 193744 64801 193750 64813
rect 144074 64773 193750 64801
rect 144074 64761 144080 64773
rect 193744 64761 193750 64773
rect 193802 64761 193808 64813
rect 146896 63355 146902 63407
rect 146954 63395 146960 63407
rect 201712 63395 201718 63407
rect 146954 63367 201718 63395
rect 146954 63355 146960 63367
rect 201712 63355 201718 63367
rect 201770 63355 201776 63407
rect 208720 63059 208726 63111
rect 208778 63099 208784 63111
rect 209584 63099 209590 63111
rect 208778 63071 209590 63099
rect 208778 63059 208784 63071
rect 209584 63059 209590 63071
rect 209642 63059 209648 63111
rect 209680 62837 209686 62889
rect 209738 62877 209744 62889
rect 210160 62877 210166 62889
rect 209738 62849 210166 62877
rect 209738 62837 209744 62849
rect 210160 62837 210166 62849
rect 210218 62837 210224 62889
rect 144016 62171 144022 62223
rect 144074 62211 144080 62223
rect 151408 62211 151414 62223
rect 144074 62183 151414 62211
rect 144074 62171 144080 62183
rect 151408 62171 151414 62183
rect 151466 62171 151472 62223
rect 208240 61949 208246 62001
rect 208298 61989 208304 62001
rect 208912 61989 208918 62001
rect 208298 61961 208918 61989
rect 208298 61949 208304 61961
rect 208912 61949 208918 61961
rect 208970 61949 208976 62001
rect 208528 61875 208534 61927
rect 208586 61915 208592 61927
rect 209008 61915 209014 61927
rect 208586 61887 209014 61915
rect 208586 61875 208592 61887
rect 209008 61875 209014 61887
rect 209066 61875 209072 61927
rect 208144 61801 208150 61853
rect 208202 61841 208208 61853
rect 208816 61841 208822 61853
rect 208202 61813 208822 61841
rect 208202 61801 208208 61813
rect 208816 61801 208822 61813
rect 208874 61801 208880 61853
rect 147952 60765 147958 60817
rect 148010 60805 148016 60817
rect 148240 60805 148246 60817
rect 148010 60777 148246 60805
rect 148010 60765 148016 60777
rect 148240 60765 148246 60777
rect 148298 60765 148304 60817
rect 169936 60765 169942 60817
rect 169994 60805 170000 60817
rect 201712 60805 201718 60817
rect 169994 60777 201718 60805
rect 169994 60765 170000 60777
rect 201712 60765 201718 60777
rect 201770 60765 201776 60817
rect 167056 60691 167062 60743
rect 167114 60731 167120 60743
rect 194128 60731 194134 60743
rect 167114 60703 194134 60731
rect 167114 60691 167120 60703
rect 194128 60691 194134 60703
rect 194186 60691 194192 60743
rect 164176 60617 164182 60669
rect 164234 60657 164240 60669
rect 209968 60657 209974 60669
rect 164234 60629 209974 60657
rect 164234 60617 164240 60629
rect 209968 60617 209974 60629
rect 210026 60617 210032 60669
rect 152464 60543 152470 60595
rect 152522 60583 152528 60595
rect 201616 60583 201622 60595
rect 152522 60555 201622 60583
rect 152522 60543 152528 60555
rect 201616 60543 201622 60555
rect 201674 60543 201680 60595
rect 148432 60469 148438 60521
rect 148490 60509 148496 60521
rect 199312 60509 199318 60521
rect 148490 60481 199318 60509
rect 148490 60469 148496 60481
rect 199312 60469 199318 60481
rect 199370 60469 199376 60521
rect 146896 60395 146902 60447
rect 146954 60435 146960 60447
rect 201712 60435 201718 60447
rect 146954 60407 201718 60435
rect 146954 60395 146960 60407
rect 201712 60395 201718 60407
rect 201770 60395 201776 60447
rect 151408 60321 151414 60373
rect 151466 60361 151472 60373
rect 209968 60361 209974 60373
rect 151466 60333 209974 60361
rect 151466 60321 151472 60333
rect 209968 60321 209974 60333
rect 210026 60321 210032 60373
rect 146512 60247 146518 60299
rect 146570 60287 146576 60299
rect 169936 60287 169942 60299
rect 146570 60259 169942 60287
rect 146570 60247 146576 60259
rect 169936 60247 169942 60259
rect 169994 60247 170000 60299
rect 208624 59137 208630 59189
rect 208682 59177 208688 59189
rect 209008 59177 209014 59189
rect 208682 59149 209014 59177
rect 208682 59137 208688 59149
rect 209008 59137 209014 59149
rect 209066 59137 209072 59189
rect 144016 58989 144022 59041
rect 144074 59029 144080 59041
rect 201616 59029 201622 59041
rect 144074 59001 201622 59029
rect 144074 58989 144080 59001
rect 201616 58989 201622 59001
rect 201674 58989 201680 59041
rect 144112 58619 144118 58671
rect 144170 58659 144176 58671
rect 144170 58631 144254 58659
rect 144170 58619 144176 58631
rect 144226 58449 144254 58631
rect 144208 58397 144214 58449
rect 144266 58397 144272 58449
rect 144016 57509 144022 57561
rect 144074 57549 144080 57561
rect 167056 57549 167062 57561
rect 144074 57521 167062 57549
rect 144074 57509 144080 57521
rect 167056 57509 167062 57521
rect 167114 57509 167120 57561
rect 144112 57435 144118 57487
rect 144170 57475 144176 57487
rect 164176 57475 164182 57487
rect 144170 57447 164182 57475
rect 144170 57435 144176 57447
rect 164176 57435 164182 57447
rect 164234 57435 164240 57487
rect 144016 54623 144022 54675
rect 144074 54663 144080 54675
rect 152464 54663 152470 54675
rect 144074 54635 152470 54663
rect 144074 54623 144080 54635
rect 152464 54623 152470 54635
rect 152522 54623 152528 54675
rect 210064 54327 210070 54379
rect 210122 54367 210128 54379
rect 213808 54367 213814 54379
rect 210122 54339 213814 54367
rect 210122 54327 210128 54339
rect 213808 54327 213814 54339
rect 213866 54327 213872 54379
rect 214192 54327 214198 54379
rect 214250 54367 214256 54379
rect 216016 54367 216022 54379
rect 214250 54339 216022 54367
rect 214250 54327 214256 54339
rect 216016 54327 216022 54339
rect 216074 54327 216080 54379
rect 209776 54253 209782 54305
rect 209834 54293 209840 54305
rect 216400 54293 216406 54305
rect 209834 54265 216406 54293
rect 209834 54253 209840 54265
rect 216400 54253 216406 54265
rect 216458 54253 216464 54305
rect 206608 54179 206614 54231
rect 206666 54219 206672 54231
rect 218224 54219 218230 54231
rect 206666 54191 218230 54219
rect 206666 54179 206672 54191
rect 218224 54179 218230 54191
rect 218282 54179 218288 54231
rect 144016 54105 144022 54157
rect 144074 54145 144080 54157
rect 148432 54145 148438 54157
rect 144074 54117 148438 54145
rect 144074 54105 144080 54117
rect 148432 54105 148438 54117
rect 148490 54105 148496 54157
rect 206512 54105 206518 54157
rect 206570 54145 206576 54157
rect 220432 54145 220438 54157
rect 206570 54117 220438 54145
rect 206570 54105 206576 54117
rect 220432 54105 220438 54117
rect 220490 54105 220496 54157
rect 209488 54031 209494 54083
rect 209546 54071 209552 54083
rect 218224 54071 218230 54083
rect 209546 54043 218230 54071
rect 209546 54031 209552 54043
rect 218224 54031 218230 54043
rect 218282 54031 218288 54083
rect 206992 53957 206998 54009
rect 207050 53997 207056 54009
rect 218416 53997 218422 54009
rect 207050 53969 218422 53997
rect 207050 53957 207056 53969
rect 218416 53957 218422 53969
rect 218474 53957 218480 54009
rect 206896 53883 206902 53935
rect 206954 53923 206960 53935
rect 216208 53923 216214 53935
rect 206954 53895 216214 53923
rect 206954 53883 206960 53895
rect 216208 53883 216214 53895
rect 216266 53883 216272 53935
rect 210640 53809 210646 53861
rect 210698 53849 210704 53861
rect 210698 53821 246878 53849
rect 210698 53809 210704 53821
rect 206416 53735 206422 53787
rect 206474 53775 206480 53787
rect 206474 53747 221486 53775
rect 206474 53735 206480 53747
rect 209392 53661 209398 53713
rect 209450 53701 209456 53713
rect 209450 53673 219470 53701
rect 209450 53661 209456 53673
rect 219442 53639 219470 53673
rect 221458 53639 221486 53747
rect 246736 53701 246742 53713
rect 239074 53673 246742 53701
rect 210256 53587 210262 53639
rect 210314 53627 210320 53639
rect 210314 53599 217982 53627
rect 210314 53587 210320 53599
rect 210352 53513 210358 53565
rect 210410 53553 210416 53565
rect 217792 53553 217798 53565
rect 210410 53525 217798 53553
rect 210410 53513 210416 53525
rect 217792 53513 217798 53525
rect 217850 53513 217856 53565
rect 217954 53553 217982 53599
rect 219424 53587 219430 53639
rect 219482 53587 219488 53639
rect 221440 53587 221446 53639
rect 221498 53587 221504 53639
rect 231760 53587 231766 53639
rect 231818 53627 231824 53639
rect 239074 53627 239102 53673
rect 246736 53661 246742 53673
rect 246794 53661 246800 53713
rect 246850 53701 246878 53821
rect 282256 53735 282262 53787
rect 282314 53775 282320 53787
rect 282314 53747 299582 53775
rect 282314 53735 282320 53747
rect 282064 53701 282070 53713
rect 246850 53673 282070 53701
rect 282064 53661 282070 53673
rect 282122 53661 282128 53713
rect 299554 53701 299582 53747
rect 345616 53701 345622 53713
rect 299554 53673 345622 53701
rect 345616 53661 345622 53673
rect 345674 53661 345680 53713
rect 231818 53599 239102 53627
rect 231818 53587 231824 53599
rect 241840 53553 241846 53565
rect 217954 53525 241846 53553
rect 241840 53513 241846 53525
rect 241898 53513 241904 53565
rect 241936 53513 241942 53565
rect 241994 53553 242000 53565
rect 380176 53553 380182 53565
rect 241994 53525 380182 53553
rect 241994 53513 242000 53525
rect 380176 53513 380182 53525
rect 380234 53513 380240 53565
rect 443554 53525 443774 53553
rect 209584 53439 209590 53491
rect 209642 53479 209648 53491
rect 217264 53479 217270 53491
rect 209642 53451 217270 53479
rect 209642 53439 209648 53451
rect 217264 53439 217270 53451
rect 217322 53439 217328 53491
rect 218416 53439 218422 53491
rect 218474 53479 218480 53491
rect 219568 53479 219574 53491
rect 218474 53451 219574 53479
rect 218474 53439 218480 53451
rect 219568 53439 219574 53451
rect 219626 53439 219632 53491
rect 220624 53439 220630 53491
rect 220682 53479 220688 53491
rect 289168 53479 289174 53491
rect 220682 53451 289174 53479
rect 220682 53439 220688 53451
rect 289168 53439 289174 53451
rect 289226 53439 289232 53491
rect 417616 53439 417622 53491
rect 417674 53479 417680 53491
rect 440560 53479 440566 53491
rect 417674 53451 440566 53479
rect 417674 53439 417680 53451
rect 440560 53439 440566 53451
rect 440618 53439 440624 53491
rect 208720 53365 208726 53417
rect 208778 53405 208784 53417
rect 217552 53405 217558 53417
rect 208778 53377 217558 53405
rect 208778 53365 208784 53377
rect 217552 53365 217558 53377
rect 217610 53365 217616 53417
rect 262096 53405 262102 53417
rect 219970 53377 262102 53405
rect 206704 53291 206710 53343
rect 206762 53331 206768 53343
rect 217360 53331 217366 53343
rect 206762 53303 217366 53331
rect 206762 53291 206768 53303
rect 217360 53291 217366 53303
rect 217418 53291 217424 53343
rect 206800 53217 206806 53269
rect 206858 53257 206864 53269
rect 215536 53257 215542 53269
rect 206858 53229 215542 53257
rect 206858 53217 206864 53229
rect 215536 53217 215542 53229
rect 215594 53217 215600 53269
rect 210160 53143 210166 53195
rect 210218 53183 210224 53195
rect 219970 53183 219998 53377
rect 262096 53365 262102 53377
rect 262154 53365 262160 53417
rect 262192 53365 262198 53417
rect 262250 53405 262256 53417
rect 443554 53405 443582 53525
rect 262250 53377 443582 53405
rect 443746 53405 443774 53525
rect 463696 53405 463702 53417
rect 443746 53377 463702 53405
rect 262250 53365 262256 53377
rect 463696 53365 463702 53377
rect 463754 53365 463760 53417
rect 246736 53291 246742 53343
rect 246794 53331 246800 53343
rect 246794 53303 262142 53331
rect 246794 53291 246800 53303
rect 210218 53155 219998 53183
rect 210218 53143 210224 53155
rect 209968 53069 209974 53121
rect 210026 53109 210032 53121
rect 221776 53109 221782 53121
rect 210026 53081 221782 53109
rect 210026 53069 210032 53081
rect 221776 53069 221782 53081
rect 221834 53069 221840 53121
rect 262114 53109 262142 53303
rect 293698 53303 293822 53331
rect 262384 53217 262390 53269
rect 262442 53257 262448 53269
rect 282352 53257 282358 53269
rect 262442 53229 282358 53257
rect 262442 53217 262448 53229
rect 282352 53217 282358 53229
rect 282410 53217 282416 53269
rect 283600 53217 283606 53269
rect 283658 53257 283664 53269
rect 293698 53257 293726 53303
rect 293794 53269 293822 53303
rect 316912 53291 316918 53343
rect 316970 53331 316976 53343
rect 383152 53331 383158 53343
rect 316970 53303 383158 53331
rect 316970 53291 316976 53303
rect 383152 53291 383158 53303
rect 383210 53291 383216 53343
rect 383248 53291 383254 53343
rect 383306 53331 383312 53343
rect 423280 53331 423286 53343
rect 383306 53303 423286 53331
rect 383306 53291 383312 53303
rect 423280 53291 423286 53303
rect 423338 53291 423344 53343
rect 463600 53291 463606 53343
rect 463658 53331 463664 53343
rect 498736 53331 498742 53343
rect 463658 53303 498742 53331
rect 463658 53291 463664 53303
rect 498736 53291 498742 53303
rect 498794 53291 498800 53343
rect 283658 53229 293726 53257
rect 283658 53217 283664 53229
rect 293776 53217 293782 53269
rect 293834 53217 293840 53269
rect 348514 53229 362942 53257
rect 293680 53143 293686 53195
rect 293738 53183 293744 53195
rect 296560 53183 296566 53195
rect 293738 53155 296566 53183
rect 293738 53143 293744 53155
rect 296560 53143 296566 53155
rect 296618 53143 296624 53195
rect 296752 53143 296758 53195
rect 296810 53183 296816 53195
rect 328528 53183 328534 53195
rect 296810 53155 328534 53183
rect 296810 53143 296816 53155
rect 328528 53143 328534 53155
rect 328586 53143 328592 53195
rect 273616 53109 273622 53121
rect 262114 53081 273622 53109
rect 273616 53069 273622 53081
rect 273674 53069 273680 53121
rect 313840 53069 313846 53121
rect 313898 53109 313904 53121
rect 316720 53109 316726 53121
rect 313898 53081 316726 53109
rect 313898 53069 313904 53081
rect 316720 53069 316726 53081
rect 316778 53069 316784 53121
rect 328624 53069 328630 53121
rect 328682 53109 328688 53121
rect 348514 53109 348542 53229
rect 354256 53143 354262 53195
rect 354314 53143 354320 53195
rect 362914 53183 362942 53229
rect 391234 53229 403262 53257
rect 391234 53183 391262 53229
rect 362914 53155 391262 53183
rect 403234 53183 403262 53229
rect 417616 53217 417622 53269
rect 417674 53217 417680 53269
rect 440560 53217 440566 53269
rect 440618 53217 440624 53269
rect 509872 53217 509878 53269
rect 509930 53257 509936 53269
rect 525904 53257 525910 53269
rect 509930 53229 525910 53257
rect 509930 53217 509936 53229
rect 525904 53217 525910 53229
rect 525962 53217 525968 53269
rect 417634 53183 417662 53217
rect 403234 53155 417662 53183
rect 440578 53183 440606 53217
rect 509680 53183 509686 53195
rect 440578 53155 509686 53183
rect 509680 53143 509686 53155
rect 509738 53143 509744 53195
rect 328682 53081 348542 53109
rect 354274 53109 354302 53143
rect 374320 53109 374326 53121
rect 354274 53081 374326 53109
rect 328682 53069 328688 53081
rect 374320 53069 374326 53081
rect 374378 53069 374384 53121
rect 443536 53069 443542 53121
rect 443594 53109 443600 53121
rect 463600 53109 463606 53121
rect 443594 53081 463606 53109
rect 443594 53069 443600 53081
rect 463600 53069 463606 53081
rect 463658 53069 463664 53121
rect 211792 52995 211798 53047
rect 211850 53035 211856 53047
rect 261904 53035 261910 53047
rect 211850 53007 261910 53035
rect 211850 52995 211856 53007
rect 261904 52995 261910 53007
rect 261962 52995 261968 53047
rect 207088 52921 207094 52973
rect 207146 52961 207152 52973
rect 219280 52961 219286 52973
rect 207146 52933 219286 52961
rect 207146 52921 207152 52933
rect 219280 52921 219286 52933
rect 219338 52921 219344 52973
rect 221776 52921 221782 52973
rect 221834 52961 221840 52973
rect 231760 52961 231766 52973
rect 221834 52933 231766 52961
rect 221834 52921 221840 52933
rect 231760 52921 231766 52933
rect 231818 52921 231824 52973
rect 282352 52921 282358 52973
rect 282410 52961 282416 52973
rect 293680 52961 293686 52973
rect 282410 52933 293686 52961
rect 282410 52921 282416 52933
rect 293680 52921 293686 52933
rect 293738 52921 293744 52973
rect 293776 52921 293782 52973
rect 293834 52961 293840 52973
rect 313840 52961 313846 52973
rect 293834 52933 313846 52961
rect 293834 52921 293840 52933
rect 313840 52921 313846 52933
rect 313898 52921 313904 52973
rect 210064 52847 210070 52899
rect 210122 52887 210128 52899
rect 218800 52887 218806 52899
rect 210122 52859 218806 52887
rect 210122 52847 210128 52859
rect 218800 52847 218806 52859
rect 218858 52847 218864 52899
rect 273616 52847 273622 52899
rect 273674 52887 273680 52899
rect 283600 52887 283606 52899
rect 273674 52859 283606 52887
rect 273674 52847 273680 52859
rect 283600 52847 283606 52859
rect 283658 52847 283664 52899
rect 165616 52551 165622 52603
rect 165674 52591 165680 52603
rect 216112 52591 216118 52603
rect 165674 52563 216118 52591
rect 165674 52551 165680 52563
rect 216112 52551 216118 52563
rect 216170 52551 216176 52603
rect 162832 52403 162838 52455
rect 162890 52443 162896 52455
rect 217936 52443 217942 52455
rect 162890 52415 217942 52443
rect 162890 52403 162896 52415
rect 217936 52403 217942 52415
rect 217994 52403 218000 52455
rect 212272 52181 212278 52233
rect 212330 52221 212336 52233
rect 220432 52221 220438 52233
rect 212330 52193 220438 52221
rect 212330 52181 212336 52193
rect 220432 52181 220438 52193
rect 220490 52181 220496 52233
rect 160048 52107 160054 52159
rect 160106 52147 160112 52159
rect 215728 52147 215734 52159
rect 160106 52119 215734 52147
rect 160106 52107 160112 52119
rect 215728 52107 215734 52119
rect 215786 52107 215792 52159
rect 163024 52033 163030 52085
rect 163082 52073 163088 52085
rect 220912 52073 220918 52085
rect 163082 52045 220918 52073
rect 163082 52033 163088 52045
rect 220912 52033 220918 52045
rect 220970 52033 220976 52085
rect 159952 51959 159958 52011
rect 160010 51999 160016 52011
rect 216880 51999 216886 52011
rect 160010 51971 216886 51999
rect 160010 51959 160016 51971
rect 216880 51959 216886 51971
rect 216938 51959 216944 52011
rect 223600 51959 223606 52011
rect 223658 51999 223664 52011
rect 241168 51999 241174 52011
rect 223658 51971 241174 51999
rect 223658 51959 223664 51971
rect 241168 51959 241174 51971
rect 241226 51959 241232 52011
rect 162736 51885 162742 51937
rect 162794 51925 162800 51937
rect 227536 51925 227542 51937
rect 162794 51897 227542 51925
rect 162794 51885 162800 51897
rect 227536 51885 227542 51897
rect 227594 51885 227600 51937
rect 625744 51885 625750 51937
rect 625802 51925 625808 51937
rect 639664 51925 639670 51937
rect 625802 51897 639670 51925
rect 625802 51885 625808 51897
rect 639664 51885 639670 51897
rect 639722 51885 639728 51937
rect 209872 51811 209878 51863
rect 209930 51851 209936 51863
rect 214480 51851 214486 51863
rect 209930 51823 214486 51851
rect 209930 51811 209936 51823
rect 214480 51811 214486 51823
rect 214538 51811 214544 51863
rect 220432 51811 220438 51863
rect 220490 51851 220496 51863
rect 645520 51851 645526 51863
rect 220490 51823 645526 51851
rect 220490 51811 220496 51823
rect 645520 51811 645526 51823
rect 645578 51811 645584 51863
rect 208336 51737 208342 51789
rect 208394 51777 208400 51789
rect 213328 51777 213334 51789
rect 208394 51749 213334 51777
rect 208394 51737 208400 51749
rect 213328 51737 213334 51749
rect 213386 51737 213392 51789
rect 219472 51737 219478 51789
rect 219530 51777 219536 51789
rect 645712 51777 645718 51789
rect 219530 51749 645718 51777
rect 219530 51737 219536 51749
rect 645712 51737 645718 51749
rect 645770 51737 645776 51789
rect 208432 51663 208438 51715
rect 208490 51703 208496 51715
rect 214096 51703 214102 51715
rect 208490 51675 214102 51703
rect 208490 51663 208496 51675
rect 214096 51663 214102 51675
rect 214154 51663 214160 51715
rect 362896 51703 362902 51715
rect 241954 51675 291614 51703
rect 145744 51589 145750 51641
rect 145802 51629 145808 51641
rect 223600 51629 223606 51641
rect 145802 51601 223606 51629
rect 145802 51589 145808 51601
rect 223600 51589 223606 51601
rect 223658 51589 223664 51641
rect 241954 51629 241982 51675
rect 241906 51601 241982 51629
rect 211120 51515 211126 51567
rect 211178 51555 211184 51567
rect 241906 51555 241934 51601
rect 211178 51527 241934 51555
rect 291586 51555 291614 51675
rect 348610 51675 362902 51703
rect 348400 51629 348406 51641
rect 291778 51601 309470 51629
rect 291778 51555 291806 51601
rect 291586 51527 291806 51555
rect 309442 51555 309470 51601
rect 309634 51601 320894 51629
rect 309634 51555 309662 51601
rect 309442 51527 309662 51555
rect 320866 51555 320894 51601
rect 336898 51601 348406 51629
rect 336898 51555 336926 51601
rect 348400 51589 348406 51601
rect 348458 51589 348464 51641
rect 348496 51589 348502 51641
rect 348554 51629 348560 51641
rect 348610 51629 348638 51675
rect 362896 51663 362902 51675
rect 362954 51663 362960 51715
rect 403216 51703 403222 51715
rect 388834 51675 403222 51703
rect 348554 51601 348638 51629
rect 348554 51589 348560 51601
rect 320866 51527 336926 51555
rect 211178 51515 211184 51527
rect 383056 51515 383062 51567
rect 383114 51555 383120 51567
rect 388834 51555 388862 51675
rect 403216 51663 403222 51675
rect 403274 51663 403280 51715
rect 434896 51703 434902 51715
rect 429154 51675 434902 51703
rect 383114 51527 388862 51555
rect 383114 51515 383120 51527
rect 423376 51515 423382 51567
rect 423434 51555 423440 51567
rect 429154 51555 429182 51675
rect 434896 51663 434902 51675
rect 434954 51663 434960 51715
rect 509680 51663 509686 51715
rect 509738 51703 509744 51715
rect 520240 51703 520246 51715
rect 509738 51675 520246 51703
rect 509738 51663 509744 51675
rect 520240 51663 520246 51675
rect 520298 51663 520304 51715
rect 558832 51703 558838 51715
rect 550210 51675 558838 51703
rect 459280 51589 459286 51641
rect 459338 51629 459344 51641
rect 489616 51629 489622 51641
rect 459338 51601 489622 51629
rect 459338 51589 459344 51601
rect 489616 51589 489622 51601
rect 489674 51589 489680 51641
rect 550000 51629 550006 51641
rect 530050 51601 550006 51629
rect 423434 51527 429182 51555
rect 423434 51515 423440 51527
rect 520240 51515 520246 51567
rect 520298 51555 520304 51567
rect 530050 51555 530078 51601
rect 550000 51589 550006 51601
rect 550058 51589 550064 51641
rect 550096 51589 550102 51641
rect 550154 51629 550160 51641
rect 550210 51629 550238 51675
rect 558832 51663 558838 51675
rect 558890 51663 558896 51715
rect 601936 51703 601942 51715
rect 593986 51675 601942 51703
rect 550154 51601 550238 51629
rect 550154 51589 550160 51601
rect 520298 51527 530078 51555
rect 520298 51515 520304 51527
rect 558832 51515 558838 51567
rect 558890 51555 558896 51567
rect 593986 51555 594014 51675
rect 601936 51663 601942 51675
rect 601994 51663 602000 51715
rect 622000 51589 622006 51641
rect 622058 51629 622064 51641
rect 625744 51629 625750 51641
rect 622058 51601 625750 51629
rect 622058 51589 622064 51601
rect 625744 51589 625750 51601
rect 625802 51589 625808 51641
rect 558890 51527 594014 51555
rect 558890 51515 558896 51527
rect 211504 51441 211510 51493
rect 211562 51481 211568 51493
rect 219472 51481 219478 51493
rect 211562 51453 219478 51481
rect 211562 51441 211568 51453
rect 219472 51441 219478 51453
rect 219530 51441 219536 51493
rect 144976 51367 144982 51419
rect 145034 51407 145040 51419
rect 233776 51407 233782 51419
rect 145034 51379 233782 51407
rect 145034 51367 145040 51379
rect 233776 51367 233782 51379
rect 233834 51367 233840 51419
rect 145456 51293 145462 51345
rect 145514 51333 145520 51345
rect 235984 51333 235990 51345
rect 145514 51305 235990 51333
rect 145514 51293 145520 51305
rect 235984 51293 235990 51305
rect 236042 51293 236048 51345
rect 145648 51219 145654 51271
rect 145706 51259 145712 51271
rect 235024 51259 235030 51271
rect 145706 51231 235030 51259
rect 145706 51219 145712 51231
rect 235024 51219 235030 51231
rect 235082 51219 235088 51271
rect 146128 51145 146134 51197
rect 146186 51185 146192 51197
rect 231952 51185 231958 51197
rect 146186 51157 231958 51185
rect 146186 51145 146192 51157
rect 231952 51145 231958 51157
rect 232010 51145 232016 51197
rect 146416 51071 146422 51123
rect 146474 51111 146480 51123
rect 231184 51111 231190 51123
rect 146474 51083 231190 51111
rect 146474 51071 146480 51083
rect 231184 51071 231190 51083
rect 231242 51071 231248 51123
rect 146320 50997 146326 51049
rect 146378 51037 146384 51049
rect 231568 51037 231574 51049
rect 146378 51009 231574 51037
rect 146378 50997 146384 51009
rect 231568 50997 231574 51009
rect 231626 50997 231632 51049
rect 146800 50923 146806 50975
rect 146858 50963 146864 50975
rect 230512 50963 230518 50975
rect 146858 50935 230518 50963
rect 146858 50923 146864 50935
rect 230512 50923 230518 50935
rect 230570 50923 230576 50975
rect 498736 50923 498742 50975
rect 498794 50963 498800 50975
rect 504016 50963 504022 50975
rect 498794 50935 504022 50963
rect 498794 50923 498800 50935
rect 504016 50923 504022 50935
rect 504074 50923 504080 50975
rect 145072 50849 145078 50901
rect 145130 50889 145136 50901
rect 228976 50889 228982 50901
rect 145130 50861 228982 50889
rect 145130 50849 145136 50861
rect 228976 50849 228982 50861
rect 229034 50849 229040 50901
rect 289168 50849 289174 50901
rect 289226 50889 289232 50901
rect 302416 50889 302422 50901
rect 289226 50861 302422 50889
rect 289226 50849 289232 50861
rect 302416 50849 302422 50861
rect 302474 50849 302480 50901
rect 159376 50775 159382 50827
rect 159434 50815 159440 50827
rect 243856 50815 243862 50827
rect 159434 50787 243862 50815
rect 159434 50775 159440 50787
rect 243856 50775 243862 50787
rect 243914 50775 243920 50827
rect 145264 50701 145270 50753
rect 145322 50741 145328 50753
rect 228400 50741 228406 50753
rect 145322 50713 228406 50741
rect 145322 50701 145328 50713
rect 228400 50701 228406 50713
rect 228458 50701 228464 50753
rect 146704 50627 146710 50679
rect 146762 50667 146768 50679
rect 229744 50667 229750 50679
rect 146762 50639 229750 50667
rect 146762 50627 146768 50639
rect 229744 50627 229750 50639
rect 229802 50627 229808 50679
rect 145360 50553 145366 50605
rect 145418 50593 145424 50605
rect 229360 50593 229366 50605
rect 145418 50565 229366 50593
rect 145418 50553 145424 50565
rect 229360 50553 229366 50565
rect 229418 50553 229424 50605
rect 144112 50479 144118 50531
rect 144170 50519 144176 50531
rect 144170 50491 211166 50519
rect 144170 50479 144176 50491
rect 144880 50405 144886 50457
rect 144938 50445 144944 50457
rect 211138 50445 211166 50491
rect 224944 50445 224950 50457
rect 144938 50417 211070 50445
rect 211138 50417 224950 50445
rect 144938 50405 144944 50417
rect 145936 50331 145942 50383
rect 145994 50371 146000 50383
rect 211042 50371 211070 50417
rect 224944 50405 224950 50417
rect 225002 50405 225008 50457
rect 226096 50371 226102 50383
rect 145994 50343 210974 50371
rect 211042 50343 226102 50371
rect 145994 50331 146000 50343
rect 146032 50257 146038 50309
rect 146090 50297 146096 50309
rect 210832 50297 210838 50309
rect 146090 50269 210838 50297
rect 146090 50257 146096 50269
rect 210832 50257 210838 50269
rect 210890 50257 210896 50309
rect 210946 50297 210974 50343
rect 226096 50331 226102 50343
rect 226154 50331 226160 50383
rect 227152 50297 227158 50309
rect 210946 50269 227158 50297
rect 227152 50257 227158 50269
rect 227210 50257 227216 50309
rect 145840 50183 145846 50235
rect 145898 50223 145904 50235
rect 225712 50223 225718 50235
rect 145898 50195 225718 50223
rect 145898 50183 145904 50195
rect 225712 50183 225718 50195
rect 225770 50183 225776 50235
rect 144208 50109 144214 50161
rect 144266 50149 144272 50161
rect 223120 50149 223126 50161
rect 144266 50121 223126 50149
rect 144266 50109 144272 50121
rect 223120 50109 223126 50121
rect 223178 50109 223184 50161
rect 144400 50035 144406 50087
rect 144458 50075 144464 50087
rect 223504 50075 223510 50087
rect 144458 50047 223510 50075
rect 144458 50035 144464 50047
rect 223504 50035 223510 50047
rect 223562 50035 223568 50087
rect 144496 49961 144502 50013
rect 144554 50001 144560 50013
rect 224176 50001 224182 50013
rect 144554 49973 224182 50001
rect 144554 49961 144560 49973
rect 224176 49961 224182 49973
rect 224234 49961 224240 50013
rect 145168 49887 145174 49939
rect 145226 49927 145232 49939
rect 235600 49927 235606 49939
rect 145226 49899 235606 49927
rect 145226 49887 145232 49899
rect 235600 49887 235606 49899
rect 235658 49887 235664 49939
rect 145552 49813 145558 49865
rect 145610 49853 145616 49865
rect 234640 49853 234646 49865
rect 145610 49825 234646 49853
rect 145610 49813 145616 49825
rect 234640 49813 234646 49825
rect 234698 49813 234704 49865
rect 144304 49739 144310 49791
rect 144362 49779 144368 49791
rect 232432 49779 232438 49791
rect 144362 49751 232438 49779
rect 144362 49739 144368 49751
rect 232432 49739 232438 49751
rect 232490 49739 232496 49791
rect 210832 49665 210838 49717
rect 210890 49705 210896 49717
rect 226768 49705 226774 49717
rect 210890 49677 226774 49705
rect 210890 49665 210896 49677
rect 226768 49665 226774 49677
rect 226826 49665 226832 49717
rect 144592 49591 144598 49643
rect 144650 49631 144656 49643
rect 234544 49631 234550 49643
rect 144650 49603 234550 49631
rect 144650 49591 144656 49603
rect 234544 49591 234550 49603
rect 234602 49591 234608 49643
rect 144784 49517 144790 49569
rect 144842 49557 144848 49569
rect 236752 49557 236758 49569
rect 144842 49529 236758 49557
rect 144842 49517 144848 49529
rect 236752 49517 236758 49529
rect 236810 49517 236816 49569
rect 218608 49073 218614 49125
rect 218666 49113 218672 49125
rect 218666 49085 218942 49113
rect 218666 49073 218672 49085
rect 208624 48925 208630 48977
rect 208682 48965 208688 48977
rect 218914 48965 218942 49085
rect 345616 48999 345622 49051
rect 345674 49039 345680 49051
rect 353584 49039 353590 49051
rect 345674 49011 353590 49039
rect 345674 48999 345680 49011
rect 353584 48999 353590 49011
rect 353642 48999 353648 49051
rect 463696 48999 463702 49051
rect 463754 49039 463760 49051
rect 471376 49039 471382 49051
rect 463754 49011 471382 49039
rect 463754 48999 463760 49011
rect 471376 48999 471382 49011
rect 471434 48999 471440 49051
rect 625072 48999 625078 49051
rect 625130 49039 625136 49051
rect 640720 49039 640726 49051
rect 625130 49011 640726 49039
rect 625130 48999 625136 49011
rect 640720 48999 640726 49011
rect 640778 48999 640784 49051
rect 645616 48965 645622 48977
rect 208682 48937 218846 48965
rect 218914 48937 645622 48965
rect 208682 48925 208688 48937
rect 218818 48891 218846 48937
rect 645616 48925 645622 48937
rect 645674 48925 645680 48977
rect 218818 48863 219902 48891
rect 209296 48777 209302 48829
rect 209354 48817 209360 48829
rect 219088 48817 219094 48829
rect 209354 48789 219094 48817
rect 209354 48777 209360 48789
rect 219088 48777 219094 48789
rect 219146 48777 219152 48829
rect 209008 48629 209014 48681
rect 209066 48669 209072 48681
rect 219760 48669 219766 48681
rect 209066 48641 219766 48669
rect 209066 48629 209072 48641
rect 219760 48629 219766 48641
rect 219818 48629 219824 48681
rect 219874 48669 219902 48863
rect 224080 48851 224086 48903
rect 224138 48891 224144 48903
rect 645328 48891 645334 48903
rect 224138 48863 645334 48891
rect 224138 48851 224144 48863
rect 645328 48851 645334 48863
rect 645386 48851 645392 48903
rect 222928 48777 222934 48829
rect 222986 48817 222992 48829
rect 645136 48817 645142 48829
rect 222986 48789 645142 48817
rect 222986 48777 222992 48789
rect 645136 48777 645142 48789
rect 645194 48777 645200 48829
rect 222160 48703 222166 48755
rect 222218 48743 222224 48755
rect 645232 48743 645238 48755
rect 222218 48715 645238 48743
rect 222218 48703 222224 48715
rect 645232 48703 645238 48715
rect 645290 48703 645296 48755
rect 226384 48669 226390 48681
rect 219874 48641 226390 48669
rect 226384 48629 226390 48641
rect 226442 48629 226448 48681
rect 504016 48629 504022 48681
rect 504074 48669 504080 48681
rect 512560 48669 512566 48681
rect 504074 48641 512566 48669
rect 504074 48629 504080 48641
rect 512560 48629 512566 48641
rect 512618 48629 512624 48681
rect 203056 48555 203062 48607
rect 203114 48595 203120 48607
rect 208720 48595 208726 48607
rect 203114 48567 208726 48595
rect 203114 48555 203120 48567
rect 208720 48555 208726 48567
rect 208778 48555 208784 48607
rect 208816 48555 208822 48607
rect 208874 48595 208880 48607
rect 220528 48595 220534 48607
rect 208874 48567 220534 48595
rect 208874 48555 208880 48567
rect 220528 48555 220534 48567
rect 220586 48555 220592 48607
rect 191440 48481 191446 48533
rect 191498 48521 191504 48533
rect 240784 48521 240790 48533
rect 191498 48493 240790 48521
rect 191498 48481 191504 48493
rect 240784 48481 240790 48493
rect 240842 48481 240848 48533
rect 182800 48407 182806 48459
rect 182858 48447 182864 48459
rect 199216 48447 199222 48459
rect 182858 48419 199222 48447
rect 182858 48407 182864 48419
rect 199216 48407 199222 48419
rect 199274 48407 199280 48459
rect 200080 48407 200086 48459
rect 200138 48447 200144 48459
rect 241264 48447 241270 48459
rect 200138 48419 241270 48447
rect 200138 48407 200144 48419
rect 241264 48407 241270 48419
rect 241322 48407 241328 48459
rect 148816 48333 148822 48385
rect 148874 48373 148880 48385
rect 227920 48373 227926 48385
rect 148874 48345 227926 48373
rect 148874 48333 148880 48345
rect 227920 48333 227926 48345
rect 227978 48333 227984 48385
rect 149296 48259 149302 48311
rect 149354 48299 149360 48311
rect 230128 48299 230134 48311
rect 149354 48271 230134 48299
rect 149354 48259 149360 48271
rect 230128 48259 230134 48271
rect 230186 48259 230192 48311
rect 380176 48259 380182 48311
rect 380234 48299 380240 48311
rect 394576 48299 394582 48311
rect 380234 48271 394582 48299
rect 380234 48259 380240 48271
rect 394576 48259 394582 48271
rect 394634 48259 394640 48311
rect 149392 48185 149398 48237
rect 149450 48225 149456 48237
rect 208624 48225 208630 48237
rect 149450 48197 208630 48225
rect 149450 48185 149456 48197
rect 208624 48185 208630 48197
rect 208682 48185 208688 48237
rect 208720 48185 208726 48237
rect 208778 48225 208784 48237
rect 220144 48225 220150 48237
rect 208778 48197 220150 48225
rect 208778 48185 208784 48197
rect 220144 48185 220150 48197
rect 220202 48185 220208 48237
rect 149488 48111 149494 48163
rect 149546 48151 149552 48163
rect 208432 48151 208438 48163
rect 149546 48123 208438 48151
rect 149546 48111 149552 48123
rect 208432 48111 208438 48123
rect 208490 48111 208496 48163
rect 208528 48111 208534 48163
rect 208586 48151 208592 48163
rect 221968 48151 221974 48163
rect 208586 48123 221974 48151
rect 208586 48111 208592 48123
rect 221968 48111 221974 48123
rect 222026 48111 222032 48163
rect 149584 48037 149590 48089
rect 149642 48077 149648 48089
rect 208048 48077 208054 48089
rect 149642 48049 208054 48077
rect 149642 48037 149648 48049
rect 208048 48037 208054 48049
rect 208106 48037 208112 48089
rect 208240 48037 208246 48089
rect 208298 48077 208304 48089
rect 222352 48077 222358 48089
rect 208298 48049 222358 48077
rect 208298 48037 208304 48049
rect 222352 48037 222358 48049
rect 222410 48037 222416 48089
rect 149680 47963 149686 48015
rect 149738 48003 149744 48015
rect 149738 47975 208094 48003
rect 149738 47963 149744 47975
rect 208066 47929 208094 47975
rect 208144 47963 208150 48015
rect 208202 48003 208208 48015
rect 222736 48003 222742 48015
rect 208202 47975 222742 48003
rect 208202 47963 208208 47975
rect 222736 47963 222742 47975
rect 222794 47963 222800 48015
rect 223888 47929 223894 47941
rect 208066 47901 223894 47929
rect 223888 47889 223894 47901
rect 223946 47889 223952 47941
rect 199216 47815 199222 47867
rect 199274 47855 199280 47867
rect 240400 47855 240406 47867
rect 199274 47827 240406 47855
rect 199274 47815 199280 47827
rect 240400 47815 240406 47827
rect 240458 47815 240464 47867
rect 221680 47781 221686 47793
rect 151042 47753 221686 47781
rect 148144 47667 148150 47719
rect 148202 47707 148208 47719
rect 151042 47707 151070 47753
rect 221680 47741 221686 47753
rect 221738 47741 221744 47793
rect 221296 47707 221302 47719
rect 148202 47679 151070 47707
rect 151138 47679 221302 47707
rect 148202 47667 148208 47679
rect 148048 47593 148054 47645
rect 148106 47633 148112 47645
rect 151138 47633 151166 47679
rect 221296 47667 221302 47679
rect 221354 47667 221360 47719
rect 148106 47605 151166 47633
rect 148106 47593 148112 47605
rect 177040 47593 177046 47645
rect 177098 47633 177104 47645
rect 238576 47633 238582 47645
rect 177098 47605 238582 47633
rect 177098 47593 177104 47605
rect 238576 47593 238582 47605
rect 238634 47593 238640 47645
rect 208048 47519 208054 47571
rect 208106 47559 208112 47571
rect 224560 47559 224566 47571
rect 208106 47531 224566 47559
rect 208106 47519 208112 47531
rect 224560 47519 224566 47531
rect 224618 47519 224624 47571
rect 208432 47445 208438 47497
rect 208490 47485 208496 47497
rect 225328 47485 225334 47497
rect 208490 47457 225334 47485
rect 208490 47445 208496 47457
rect 225328 47445 225334 47457
rect 225386 47445 225392 47497
rect 149200 47371 149206 47423
rect 149258 47411 149264 47423
rect 233392 47411 233398 47423
rect 149258 47383 233398 47411
rect 149258 47371 149264 47383
rect 233392 47371 233398 47383
rect 233450 47371 233456 47423
rect 197200 46853 197206 46905
rect 197258 46893 197264 46905
rect 239056 46893 239062 46905
rect 197258 46865 239062 46893
rect 197258 46853 197264 46865
rect 239056 46853 239062 46865
rect 239114 46853 239120 46905
rect 148912 46779 148918 46831
rect 148970 46819 148976 46831
rect 234160 46819 234166 46831
rect 148970 46791 234166 46819
rect 148970 46779 148976 46791
rect 234160 46779 234166 46791
rect 234218 46779 234224 46831
rect 148624 46705 148630 46757
rect 148682 46745 148688 46757
rect 230608 46745 230614 46757
rect 148682 46717 230614 46745
rect 148682 46705 148688 46717
rect 230608 46705 230614 46717
rect 230666 46705 230672 46757
rect 148336 46631 148342 46683
rect 148394 46671 148400 46683
rect 232816 46671 232822 46683
rect 148394 46643 232822 46671
rect 148394 46631 148400 46643
rect 232816 46631 232822 46643
rect 232874 46631 232880 46683
rect 148528 46557 148534 46609
rect 148586 46597 148592 46609
rect 232336 46597 232342 46609
rect 148586 46569 232342 46597
rect 148586 46557 148592 46569
rect 232336 46557 232342 46569
rect 232394 46557 232400 46609
rect 148720 46483 148726 46535
rect 148778 46523 148784 46535
rect 228016 46523 228022 46535
rect 148778 46495 228022 46523
rect 148778 46483 148784 46495
rect 228016 46483 228022 46495
rect 228074 46483 228080 46535
rect 179920 46409 179926 46461
rect 179978 46449 179984 46461
rect 238960 46449 238966 46461
rect 179978 46421 238966 46449
rect 179978 46409 179984 46421
rect 238960 46409 238966 46421
rect 239018 46409 239024 46461
rect 148240 46335 148246 46387
rect 148298 46375 148304 46387
rect 236848 46375 236854 46387
rect 148298 46347 236854 46375
rect 148298 46335 148304 46347
rect 236848 46335 236854 46347
rect 236906 46335 236912 46387
rect 147952 46113 147958 46165
rect 148010 46153 148016 46165
rect 236368 46153 236374 46165
rect 148010 46125 236374 46153
rect 148010 46113 148016 46125
rect 236368 46113 236374 46125
rect 236426 46113 236432 46165
rect 212848 44781 212854 44833
rect 212906 44821 212912 44833
rect 408880 44821 408886 44833
rect 212906 44793 408886 44821
rect 212906 44781 212912 44793
rect 408880 44781 408886 44793
rect 408938 44781 408944 44833
rect 213904 44707 213910 44759
rect 213962 44747 213968 44759
rect 457744 44747 457750 44759
rect 213962 44719 457750 44747
rect 213962 44707 213968 44719
rect 457744 44707 457750 44719
rect 457802 44707 457808 44759
rect 141808 44633 141814 44685
rect 141866 44673 141872 44685
rect 155536 44673 155542 44685
rect 141866 44645 155542 44673
rect 141866 44633 141872 44645
rect 155536 44633 155542 44645
rect 155594 44633 155600 44685
rect 214672 44633 214678 44685
rect 214730 44673 214736 44685
rect 509776 44673 509782 44685
rect 214730 44645 509782 44673
rect 214730 44633 214736 44645
rect 509776 44633 509782 44645
rect 509834 44633 509840 44685
rect 509776 43227 509782 43279
rect 509834 43267 509840 43279
rect 509834 43239 521630 43267
rect 509834 43227 509840 43239
rect 521602 43205 521630 43239
rect 394576 43153 394582 43205
rect 394634 43193 394640 43205
rect 408976 43193 408982 43205
rect 394634 43165 408982 43193
rect 394634 43153 394640 43165
rect 408976 43153 408982 43165
rect 409034 43153 409040 43205
rect 521584 43153 521590 43205
rect 521642 43153 521648 43205
rect 212464 42339 212470 42391
rect 212522 42379 212528 42391
rect 310096 42379 310102 42391
rect 212522 42351 310102 42379
rect 212522 42339 212528 42351
rect 310096 42339 310102 42351
rect 310154 42339 310160 42391
rect 207280 42117 207286 42169
rect 207338 42157 207344 42169
rect 405232 42157 405238 42169
rect 207338 42129 405238 42157
rect 207338 42117 207344 42129
rect 405232 42117 405238 42129
rect 405290 42117 405296 42169
rect 512560 42117 512566 42169
rect 512618 42157 512624 42169
rect 520336 42157 520342 42169
rect 512618 42129 520342 42157
rect 512618 42117 512624 42129
rect 520336 42117 520342 42129
rect 520394 42117 520400 42169
rect 213520 42043 213526 42095
rect 213578 42083 213584 42095
rect 460048 42083 460054 42095
rect 213578 42055 460054 42083
rect 213578 42043 213584 42055
rect 460048 42043 460054 42055
rect 460106 42043 460112 42095
rect 514864 41747 514870 41799
rect 514922 41747 514928 41799
rect 214288 41673 214294 41725
rect 214346 41713 214352 41725
rect 514882 41713 514910 41747
rect 214346 41685 514910 41713
rect 214346 41673 214352 41685
<< via1 >>
rect 439222 1005745 439274 1005797
rect 466582 1005745 466634 1005797
rect 92374 1005523 92426 1005575
rect 371830 1005671 371882 1005723
rect 440662 1005671 440714 1005723
rect 446422 1005671 446474 1005723
rect 108598 1005449 108650 1005501
rect 357910 1005449 357962 1005501
rect 365014 1005449 365066 1005501
rect 383638 1005597 383690 1005649
rect 466486 1005523 466538 1005575
rect 93622 1005375 93674 1005427
rect 114166 1005375 114218 1005427
rect 298102 1005375 298154 1005427
rect 308758 1005375 308810 1005427
rect 364150 1005375 364202 1005427
rect 380566 1005449 380618 1005501
rect 430774 1005449 430826 1005501
rect 430870 1005449 430922 1005501
rect 446326 1005449 446378 1005501
rect 446422 1005449 446474 1005501
rect 471862 1005449 471914 1005501
rect 371062 1005375 371114 1005427
rect 380470 1005375 380522 1005427
rect 298390 1005301 298442 1005353
rect 309622 1005301 309674 1005353
rect 366742 1005301 366794 1005353
rect 380374 1005301 380426 1005353
rect 424534 1005301 424586 1005353
rect 439222 1005375 439274 1005427
rect 439414 1005375 439466 1005427
rect 470902 1005375 470954 1005427
rect 501142 1005375 501194 1005427
rect 518326 1005375 518378 1005427
rect 217270 1005227 217322 1005279
rect 218902 1005227 218954 1005279
rect 298294 1005227 298346 1005279
rect 307990 1005227 308042 1005279
rect 318646 1005227 318698 1005279
rect 331126 1005227 331178 1005279
rect 365782 1005227 365834 1005279
rect 380278 1005227 380330 1005279
rect 425302 1005227 425354 1005279
rect 460822 1005301 460874 1005353
rect 554518 1005301 554570 1005353
rect 572854 1005301 572906 1005353
rect 93718 1005153 93770 1005205
rect 115222 1005153 115274 1005205
rect 299926 1005153 299978 1005205
rect 315190 1005153 315242 1005205
rect 325462 1005153 325514 1005205
rect 331222 1005153 331274 1005205
rect 363478 1005153 363530 1005205
rect 371062 1005153 371114 1005205
rect 371830 1005153 371882 1005205
rect 380182 1005153 380234 1005205
rect 426070 1005153 426122 1005205
rect 437590 1005153 437642 1005205
rect 433174 1005079 433226 1005131
rect 439030 1005227 439082 1005279
rect 437878 1005153 437930 1005205
rect 471478 1005227 471530 1005279
rect 504598 1005227 504650 1005279
rect 521398 1005227 521450 1005279
rect 555766 1005227 555818 1005279
rect 573046 1005227 573098 1005279
rect 439222 1005153 439274 1005205
rect 471670 1005153 471722 1005205
rect 500758 1005153 500810 1005205
rect 512566 1005153 512618 1005205
rect 518326 1005153 518378 1005205
rect 521590 1005153 521642 1005205
rect 553750 1005153 553802 1005205
rect 572950 1005153 573002 1005205
rect 435574 1005005 435626 1005057
rect 440662 1005005 440714 1005057
rect 359926 1003969 359978 1004021
rect 380086 1003969 380138 1004021
rect 423382 1003895 423434 1003947
rect 453334 1003895 453386 1003947
rect 359062 1003821 359114 1003873
rect 377494 1003821 377546 1003873
rect 426454 1003821 426506 1003873
rect 463702 1003821 463754 1003873
rect 552598 1003821 552650 1003873
rect 572662 1003821 572714 1003873
rect 358390 1003747 358442 1003799
rect 377398 1003747 377450 1003799
rect 422518 1003747 422570 1003799
rect 461014 1003747 461066 1003799
rect 499990 1003747 500042 1003799
rect 515542 1003747 515594 1003799
rect 556534 1003747 556586 1003799
rect 574006 1003747 574058 1003799
rect 360694 1003673 360746 1003725
rect 377302 1003673 377354 1003725
rect 428086 1003673 428138 1003725
rect 472054 1003673 472106 1003725
rect 551734 1003673 551786 1003725
rect 572758 1003673 572810 1003725
rect 559222 1002637 559274 1002689
rect 566326 1002637 566378 1002689
rect 559990 1002563 560042 1002615
rect 566134 1002563 566186 1002615
rect 144022 1002489 144074 1002541
rect 150358 1002489 150410 1002541
rect 299638 1002489 299690 1002541
rect 307606 1002489 307658 1002541
rect 503446 1002489 503498 1002541
rect 515446 1002489 515498 1002541
rect 562198 1002489 562250 1002541
rect 567574 1002489 567626 1002541
rect 246550 1002415 246602 1002467
rect 254038 1002415 254090 1002467
rect 299542 1002415 299594 1002467
rect 305590 1002415 305642 1002467
rect 502774 1002415 502826 1002467
rect 513526 1002415 513578 1002467
rect 564598 1002415 564650 1002467
rect 568726 1002415 568778 1002467
rect 143926 1002341 143978 1002393
rect 153622 1002341 153674 1002393
rect 299830 1002341 299882 1002393
rect 306550 1002341 306602 1002393
rect 505078 1002341 505130 1002393
rect 521494 1002341 521546 1002393
rect 560470 1002341 560522 1002393
rect 564790 1002341 564842 1002393
rect 143734 1002267 143786 1002319
rect 178486 1002267 178538 1002319
rect 246742 1002267 246794 1002319
rect 253174 1002267 253226 1002319
rect 299734 1002267 299786 1002319
rect 304726 1002267 304778 1002319
rect 446326 1002267 446378 1002319
rect 489526 1002267 489578 1002319
rect 519190 1002267 519242 1002319
rect 561526 1002267 561578 1002319
rect 564694 1002267 564746 1002319
rect 460918 1002193 460970 1002245
rect 466582 1002193 466634 1002245
rect 471958 1002193 472010 1002245
rect 573046 1002193 573098 1002245
rect 573910 1002193 573962 1002245
rect 572950 1001823 573002 1001875
rect 573238 1001823 573290 1001875
rect 513526 1001601 513578 1001653
rect 518326 1001601 518378 1001653
rect 515446 1001527 515498 1001579
rect 516886 1001527 516938 1001579
rect 566134 1001453 566186 1001505
rect 567766 1001453 567818 1001505
rect 572854 1001305 572906 1001357
rect 574486 1001305 574538 1001357
rect 511030 1001231 511082 1001283
rect 516694 1001231 516746 1001283
rect 434134 1001083 434186 1001135
rect 472630 1001083 472682 1001135
rect 463702 1001009 463754 1001061
rect 471766 1001009 471818 1001061
rect 509398 1001009 509450 1001061
rect 516694 1001009 516746 1001061
rect 432502 1000935 432554 1000987
rect 472630 1000935 472682 1000987
rect 428950 1000861 429002 1000913
rect 472534 1000861 472586 1000913
rect 143830 1000787 143882 1000839
rect 160246 1000787 160298 1000839
rect 195094 1000787 195146 1000839
rect 208438 1000787 208490 1000839
rect 361558 1000787 361610 1000839
rect 383446 1000787 383498 1000839
rect 427318 1000787 427370 1000839
rect 472342 1000787 472394 1000839
rect 507766 1000713 507818 1000765
rect 516694 1000713 516746 1000765
rect 453334 1000417 453386 1000469
rect 463702 1000417 463754 1000469
rect 460822 1000343 460874 1000395
rect 472150 1000343 472202 1000395
rect 380470 999899 380522 999951
rect 383254 999899 383306 999951
rect 610582 999677 610634 999729
rect 625750 999677 625802 999729
rect 93046 999603 93098 999655
rect 127414 999603 127466 999655
rect 298102 999603 298154 999655
rect 298486 999603 298538 999655
rect 377302 999603 377354 999655
rect 383158 999603 383210 999655
rect 613462 999603 613514 999655
rect 625462 999603 625514 999655
rect 144214 999529 144266 999581
rect 158614 999529 158666 999581
rect 246646 999529 246698 999581
rect 262102 999529 262154 999581
rect 380182 999529 380234 999581
rect 383350 999529 383402 999581
rect 497590 999529 497642 999581
rect 516694 999529 516746 999581
rect 604726 999529 604778 999581
rect 625558 999529 625610 999581
rect 144118 999455 144170 999507
rect 155158 999455 155210 999507
rect 250486 999455 250538 999507
rect 263062 999455 263114 999507
rect 298102 999455 298154 999507
rect 311158 999455 311210 999507
rect 380374 999455 380426 999507
rect 382966 999455 383018 999507
rect 506326 999455 506378 999507
rect 516790 999455 516842 999507
rect 564694 999455 564746 999507
rect 143734 999381 143786 999433
rect 156886 999381 156938 999433
rect 246550 999381 246602 999433
rect 259606 999381 259658 999433
rect 299446 999381 299498 999433
rect 310294 999381 310346 999433
rect 380566 999381 380618 999433
rect 383542 999381 383594 999433
rect 399958 999381 400010 999433
rect 540310 999381 540362 999433
rect 561526 999381 561578 999433
rect 566326 999381 566378 999433
rect 593302 999455 593354 999507
rect 625846 999455 625898 999507
rect 460822 999307 460874 999359
rect 502390 999307 502442 999359
rect 516694 999307 516746 999359
rect 516886 999307 516938 999359
rect 520918 999307 520970 999359
rect 570454 999307 570506 999359
rect 590518 999381 590570 999433
rect 625654 999381 625706 999433
rect 570646 999307 570698 999359
rect 461014 999233 461066 999285
rect 471574 999233 471626 999285
rect 515542 999233 515594 999285
rect 523414 999233 523466 999285
rect 356278 998049 356330 998101
rect 368758 998049 368810 998101
rect 357046 997975 357098 998027
rect 368662 997975 368714 998027
rect 555286 997975 555338 998027
rect 570742 997975 570794 998027
rect 320950 997901 321002 997953
rect 367894 997901 367946 997953
rect 381718 997901 381770 997953
rect 561526 997901 561578 997953
rect 616342 997901 616394 997953
rect 331126 997827 331178 997879
rect 369046 997827 369098 997879
rect 557302 997827 557354 997879
rect 593302 997827 593354 997879
rect 574006 997753 574058 997805
rect 590518 997753 590570 997805
rect 567766 997679 567818 997731
rect 604726 997679 604778 997731
rect 573910 997605 573962 997657
rect 613462 997605 613514 997657
rect 564790 997531 564842 997583
rect 610582 997531 610634 997583
rect 460918 996939 460970 996991
rect 472246 996939 472298 996991
rect 377398 996865 377450 996917
rect 382870 996865 382922 996917
rect 201622 996643 201674 996695
rect 195766 996495 195818 996547
rect 205654 996495 205706 996547
rect 377494 996569 377546 996621
rect 382774 996569 382826 996621
rect 510262 996569 510314 996621
rect 521014 996569 521066 996621
rect 211702 996495 211754 996547
rect 298198 996495 298250 996547
rect 374518 996495 374570 996547
rect 508630 996495 508682 996547
rect 521206 996495 521258 996547
rect 320182 996421 320234 996473
rect 367126 996421 367178 996473
rect 144310 996273 144362 996325
rect 162262 996273 162314 996325
rect 115318 996125 115370 996177
rect 126742 996125 126794 996177
rect 115222 996051 115274 996103
rect 163126 996051 163178 996103
rect 177046 996051 177098 996103
rect 511126 996199 511178 996251
rect 198550 996125 198602 996177
rect 203638 996125 203690 996177
rect 214102 996125 214154 996177
rect 213334 996051 213386 996103
rect 266806 996125 266858 996177
rect 318646 996125 318698 996177
rect 371542 996125 371594 996177
rect 436342 996125 436394 996177
rect 436438 996125 436490 996177
rect 513430 996125 513482 996177
rect 562774 996125 562826 996177
rect 120982 995977 121034 996029
rect 164566 995977 164618 996029
rect 198646 995977 198698 996029
rect 202966 995977 203018 996029
rect 213046 995977 213098 996029
rect 216886 995977 216938 996029
rect 265942 996051 265994 996103
rect 317110 996051 317162 996103
rect 320950 996051 321002 996103
rect 381718 996051 381770 996103
rect 440662 996051 440714 996103
rect 265078 995977 265130 996029
rect 316342 995977 316394 996029
rect 320182 995977 320234 996029
rect 367126 995977 367178 996029
rect 434134 995977 434186 996029
rect 439414 995977 439466 996029
rect 470902 995977 470954 996029
rect 100630 995903 100682 995955
rect 94678 995829 94730 995881
rect 99958 995829 100010 995881
rect 82294 995755 82346 995807
rect 87862 995755 87914 995807
rect 102166 995755 102218 995807
rect 106486 995755 106538 995807
rect 113494 995829 113546 995881
rect 144118 995903 144170 995955
rect 152086 995903 152138 995955
rect 164182 995903 164234 995955
rect 215638 995903 215690 995955
rect 218902 995903 218954 995955
rect 266998 995903 267050 995955
rect 370582 995903 370634 995955
rect 374614 995903 374666 995955
rect 383350 995903 383402 995955
rect 177046 995829 177098 995881
rect 214102 995829 214154 995881
rect 246742 995829 246794 995881
rect 253366 995829 253418 995881
rect 259126 995829 259178 995881
rect 299446 995829 299498 995881
rect 382966 995829 383018 995881
rect 113302 995755 113354 995807
rect 118102 995755 118154 995807
rect 132406 995755 132458 995807
rect 133654 995755 133706 995807
rect 142966 995755 143018 995807
rect 143734 995755 143786 995807
rect 164086 995755 164138 995807
rect 165622 995755 165674 995807
rect 178486 995755 178538 995807
rect 185206 995755 185258 995807
rect 190582 995755 190634 995807
rect 204982 995755 205034 995807
rect 240886 995755 240938 995807
rect 245686 995755 245738 995807
rect 246550 995755 246602 995807
rect 283702 995755 283754 995807
rect 297334 995755 297386 995807
rect 298102 995755 298154 995807
rect 371350 995755 371402 995807
rect 374422 995755 374474 995807
rect 383638 995755 383690 995807
rect 384406 995755 384458 995807
rect 386038 995755 386090 995807
rect 471862 995903 471914 995955
rect 389398 995755 389450 995807
rect 396598 995755 396650 995807
rect 399958 995755 400010 995807
rect 438742 995755 438794 995807
rect 444886 995755 444938 995807
rect 472630 995755 472682 995807
rect 473302 995755 473354 995807
rect 91510 995681 91562 995733
rect 105334 995681 105386 995733
rect 127414 995681 127466 995733
rect 134326 995681 134378 995733
rect 141046 995681 141098 995733
rect 143830 995681 143882 995733
rect 163990 995681 164042 995733
rect 166294 995681 166346 995733
rect 194422 995681 194474 995733
rect 195094 995681 195146 995733
rect 198646 995681 198698 995733
rect 206614 995681 206666 995733
rect 243190 995681 243242 995733
rect 246646 995681 246698 995733
rect 294838 995681 294890 995733
rect 298198 995681 298250 995733
rect 383542 995681 383594 995733
rect 387478 995681 387530 995733
rect 472534 995681 472586 995733
rect 474070 995681 474122 995733
rect 511126 995903 511178 995955
rect 563542 996051 563594 996103
rect 513430 995977 513482 996029
rect 564790 995977 564842 996029
rect 521110 995903 521162 995955
rect 511894 995829 511946 995881
rect 523894 995829 523946 995881
rect 524086 995755 524138 995807
rect 528406 995755 528458 995807
rect 523990 995681 524042 995733
rect 528982 995681 529034 995733
rect 625462 995903 625514 995955
rect 625654 995829 625706 995881
rect 529846 995755 529898 995807
rect 537142 995755 537194 995807
rect 540310 995755 540362 995807
rect 625846 995755 625898 995807
rect 627094 995755 627146 995807
rect 630166 995755 630218 995807
rect 630934 995755 630986 995807
rect 532822 995681 532874 995733
rect 625750 995681 625802 995733
rect 626518 995681 626570 995733
rect 139318 995607 139370 995659
rect 143926 995607 143978 995659
rect 184342 995607 184394 995659
rect 195766 995607 195818 995659
rect 201718 995607 201770 995659
rect 206998 995607 207050 995659
rect 286774 995607 286826 995659
rect 298390 995607 298442 995659
rect 383446 995607 383498 995659
rect 384982 995607 385034 995659
rect 472342 995607 472394 995659
rect 477718 995607 477770 995659
rect 479446 995607 479498 995659
rect 137974 995533 138026 995585
rect 144022 995533 144074 995585
rect 287542 995533 287594 995585
rect 298486 995533 298538 995585
rect 383254 995533 383306 995585
rect 391702 995533 391754 995585
rect 472726 995533 472778 995585
rect 474646 995533 474698 995585
rect 81622 995459 81674 995511
rect 102166 995459 102218 995511
rect 236470 995459 236522 995511
rect 254806 995459 254858 995511
rect 287926 995459 287978 995511
rect 299830 995459 299882 995511
rect 383158 995459 383210 995511
rect 388054 995459 388106 995511
rect 471766 995459 471818 995511
rect 483862 995459 483914 995511
rect 523798 995607 523850 995659
rect 525430 995607 525482 995659
rect 563542 995607 563594 995659
rect 567382 995607 567434 995659
rect 625558 995607 625610 995659
rect 629590 995607 629642 995659
rect 523702 995533 523754 995585
rect 524758 995533 524810 995585
rect 562774 995533 562826 995585
rect 567478 995533 567530 995585
rect 629206 995459 629258 995511
rect 89782 995385 89834 995437
rect 92086 995385 92138 995437
rect 126742 995385 126794 995437
rect 144310 995385 144362 995437
rect 235798 995385 235850 995437
rect 247606 995385 247658 995437
rect 284374 995385 284426 995437
rect 299926 995385 299978 995437
rect 382870 995385 382922 995437
rect 393046 995385 393098 995437
rect 460822 995385 460874 995437
rect 630742 995385 630794 995437
rect 471574 995311 471626 995363
rect 479446 995311 479498 995363
rect 518518 995311 518570 995363
rect 533686 995311 533738 995363
rect 472150 995237 472202 995289
rect 478630 995237 478682 995289
rect 521014 995237 521066 995289
rect 537382 995237 537434 995289
rect 537526 995237 537578 995289
rect 645142 995237 645194 995289
rect 69142 995163 69194 995215
rect 343894 995163 343946 995215
rect 374518 995163 374570 995215
rect 649942 995163 649994 995215
rect 262198 995089 262250 995141
rect 645238 995089 645290 995141
rect 89014 995015 89066 995067
rect 570262 995015 570314 995067
rect 616342 995015 616394 995067
rect 640342 995015 640394 995067
rect 382774 994941 382826 994993
rect 395158 994941 395210 994993
rect 463702 994941 463754 994993
rect 482710 994941 482762 994993
rect 523414 994941 523466 994993
rect 537526 994941 537578 994993
rect 471670 994867 471722 994919
rect 481654 994867 481706 994919
rect 519190 994867 519242 994919
rect 530326 994867 530378 994919
rect 158422 994571 158474 994623
rect 178486 994571 178538 994623
rect 141238 994497 141290 994549
rect 146998 994497 147050 994549
rect 574486 994127 574538 994179
rect 635254 994127 635306 994179
rect 572758 993979 572810 994031
rect 636118 993979 636170 994031
rect 180502 993905 180554 993957
rect 201718 993905 201770 993957
rect 234934 993905 234986 993957
rect 250486 993905 250538 993957
rect 570646 993905 570698 993957
rect 639190 993905 639242 993957
rect 182998 993831 183050 993883
rect 207286 993831 207338 993883
rect 232150 993831 232202 993883
rect 253366 993831 253418 993883
rect 368662 993831 368714 993883
rect 392662 993831 392714 993883
rect 572662 993831 572714 993883
rect 634870 993831 634922 993883
rect 77686 993757 77738 993809
rect 100726 993757 100778 993809
rect 129334 993757 129386 993809
rect 152566 993757 152618 993809
rect 181366 993757 181418 993809
rect 212662 993757 212714 993809
rect 234358 993757 234410 993809
rect 261430 993757 261482 993809
rect 512758 993757 512810 993809
rect 534358 993757 534410 993809
rect 570742 993757 570794 993809
rect 637366 993757 637418 993809
rect 80182 993683 80234 993735
rect 107254 993683 107306 993735
rect 128470 993683 128522 993735
rect 159574 993683 159626 993735
rect 179830 993683 179882 993735
rect 211030 993683 211082 993735
rect 232534 993683 232586 993735
rect 264022 993683 264074 993735
rect 368758 993683 368810 993735
rect 393718 993683 393770 993735
rect 506614 993683 506666 993735
rect 538966 993683 539018 993735
rect 557974 993683 558026 993735
rect 641014 993683 641066 993735
rect 77302 993609 77354 993661
rect 108214 993609 108266 993661
rect 129718 993609 129770 993661
rect 161206 993609 161258 993661
rect 185398 993609 185450 993661
rect 236758 993609 236810 993661
rect 279286 993609 279338 993661
rect 282838 993609 282890 993661
rect 313846 993609 313898 993661
rect 362326 993609 362378 993661
rect 398806 993609 398858 993661
rect 429718 993609 429770 993661
rect 487798 993609 487850 993661
rect 530326 993609 530378 993661
rect 630838 993609 630890 993661
rect 632374 993609 632426 993661
rect 638902 993609 638954 993661
rect 643606 993609 643658 993661
rect 469462 993535 469514 993587
rect 479158 993535 479210 993587
rect 489526 993535 489578 993587
rect 331222 992129 331274 992181
rect 332566 992129 332618 992181
rect 285142 991611 285194 991663
rect 298582 991611 298634 991663
rect 241942 990871 241994 990923
rect 246454 990871 246506 990923
rect 629206 990871 629258 990923
rect 642166 990871 642218 990923
rect 640342 989465 640394 989517
rect 650230 989465 650282 989517
rect 645238 988503 645290 988555
rect 650038 988503 650090 988555
rect 604726 988207 604778 988259
rect 618550 988207 618602 988259
rect 64918 987763 64970 987815
rect 69142 987837 69194 987889
rect 223126 987763 223178 987815
rect 235606 987763 235658 987815
rect 236278 987763 236330 987815
rect 241942 987837 241994 987889
rect 518422 987763 518474 987815
rect 527638 987763 527690 987815
rect 570262 987763 570314 987815
rect 576310 987763 576362 987815
rect 645142 987763 645194 987815
rect 649366 987763 649418 987815
rect 219478 987171 219530 987223
rect 221878 987171 221930 987223
rect 374422 986505 374474 986557
rect 397846 986505 397898 986557
rect 570358 986505 570410 986557
rect 592438 986505 592490 986557
rect 630742 986505 630794 986557
rect 639382 986505 639434 986557
rect 326806 986431 326858 986483
rect 349174 986431 349226 986483
rect 377302 986431 377354 986483
rect 414070 986431 414122 986483
rect 445078 986431 445130 986483
rect 478966 986431 479018 986483
rect 521302 986431 521354 986483
rect 543766 986431 543818 986483
rect 573142 986431 573194 986483
rect 608758 986431 608810 986483
rect 622006 986431 622058 986483
rect 641110 986431 641162 986483
rect 73462 986357 73514 986409
rect 93622 986357 93674 986409
rect 138262 986357 138314 986409
rect 164086 986357 164138 986409
rect 273718 986357 273770 986409
rect 300502 986357 300554 986409
rect 323926 986357 323978 986409
rect 365398 986357 365450 986409
rect 374614 986357 374666 986409
rect 430294 986357 430346 986409
rect 440662 986357 440714 986409
rect 495190 986357 495242 986409
rect 518614 986357 518666 986409
rect 560086 986357 560138 986409
rect 570550 986357 570602 986409
rect 624982 986357 625034 986409
rect 630742 986357 630794 986409
rect 631030 986357 631082 986409
rect 203158 986283 203210 986335
rect 213046 986283 213098 986335
rect 273622 986135 273674 986187
rect 284278 986135 284330 986187
rect 154486 985987 154538 986039
rect 163990 985987 164042 986039
rect 89590 985839 89642 985891
rect 93718 985839 93770 985891
rect 45046 985469 45098 985521
rect 80758 985469 80810 985521
rect 100822 985469 100874 985521
rect 120886 985469 120938 985521
rect 146806 985469 146858 985521
rect 50518 985395 50570 985447
rect 122038 985395 122090 985447
rect 146998 985395 147050 985447
rect 201526 985469 201578 985521
rect 201622 985469 201674 985521
rect 218902 985469 218954 985521
rect 239158 985395 239210 985447
rect 251830 985395 251882 985447
rect 47830 985321 47882 985373
rect 186934 985321 186986 985373
rect 218998 985321 219050 985373
rect 80566 985247 80618 985299
rect 279382 985321 279434 985373
rect 285142 985321 285194 985373
rect 239158 985247 239210 985299
rect 45142 985173 45194 985225
rect 239062 985173 239114 985225
rect 239542 985173 239594 985225
rect 316726 985173 316778 985225
rect 44950 985099 45002 985151
rect 239158 985099 239210 985151
rect 239734 985099 239786 985151
rect 381622 985099 381674 985151
rect 444886 985099 444938 985151
rect 462742 985099 462794 985151
rect 44854 985025 44906 985077
rect 239062 985025 239114 985077
rect 239446 985025 239498 985077
rect 446518 985025 446570 985077
rect 42934 984951 42986 985003
rect 511414 984951 511466 985003
rect 642262 984951 642314 985003
rect 649462 984877 649514 984929
rect 65014 983841 65066 983893
rect 94966 983841 95018 983893
rect 47446 983767 47498 983819
rect 118102 983767 118154 983819
rect 618550 983767 618602 983819
rect 649654 983767 649706 983819
rect 44758 983693 44810 983745
rect 115222 983693 115274 983745
rect 568726 983693 568778 983745
rect 652246 983693 652298 983745
rect 44566 983619 44618 983671
rect 115318 983619 115370 983671
rect 567478 983619 567530 983671
rect 658006 983619 658058 983671
rect 65110 983545 65162 983597
rect 145270 983545 145322 983597
rect 567382 983545 567434 983597
rect 658102 983545 658154 983597
rect 65206 983471 65258 983523
rect 195382 983471 195434 983523
rect 217366 983471 217418 983523
rect 236278 983471 236330 983523
rect 544246 983471 544298 983523
rect 650902 983471 650954 983523
rect 273622 982287 273674 982339
rect 279382 982287 279434 982339
rect 643606 981769 643658 981821
rect 649846 981769 649898 981821
rect 639382 981325 639434 981377
rect 650134 981325 650186 981377
rect 130390 981029 130442 981081
rect 64726 980807 64778 980859
rect 106486 980955 106538 981007
rect 106582 980955 106634 981007
rect 130390 980881 130442 980933
rect 161302 980955 161354 981007
rect 64822 980659 64874 980711
rect 106486 980733 106538 980785
rect 106582 980733 106634 980785
rect 146902 980807 146954 980859
rect 178486 980881 178538 980933
rect 171286 980807 171338 980859
rect 146806 980733 146858 980785
rect 178486 980733 178538 980785
rect 238966 980807 239018 980859
rect 247606 980807 247658 980859
rect 247702 980807 247754 980859
rect 217366 980733 217418 980785
rect 217558 980733 217610 980785
rect 217654 980733 217706 980785
rect 218902 980733 218954 980785
rect 630838 980807 630890 980859
rect 273622 980733 273674 980785
rect 630934 980733 630986 980785
rect 675094 980733 675146 980785
rect 675286 980659 675338 980711
rect 53302 970595 53354 970647
rect 59542 970595 59594 970647
rect 42166 967265 42218 967317
rect 42934 967265 42986 967317
rect 42070 961345 42122 961397
rect 42550 961345 42602 961397
rect 42166 960679 42218 960731
rect 42358 960679 42410 960731
rect 673942 958977 673994 959029
rect 675478 958977 675530 959029
rect 675094 958385 675146 958437
rect 675382 958385 675434 958437
rect 675190 956979 675242 957031
rect 675478 956979 675530 957031
rect 43126 956165 43178 956217
rect 59542 956165 59594 956217
rect 42070 955277 42122 955329
rect 42934 955277 42986 955329
rect 669526 954685 669578 954737
rect 675382 954685 675434 954737
rect 42166 954611 42218 954663
rect 42838 954611 42890 954663
rect 674134 953871 674186 953923
rect 675478 953871 675530 953923
rect 674038 952021 674090 952073
rect 675478 952021 675530 952073
rect 649558 951799 649610 951851
rect 653782 951799 653834 951851
rect 42358 948543 42410 948595
rect 42646 948543 42698 948595
rect 42358 947729 42410 947781
rect 47542 947729 47594 947781
rect 42166 947655 42218 947707
rect 50326 947655 50378 947707
rect 655222 944843 655274 944895
rect 674710 944843 674762 944895
rect 655126 944621 655178 944673
rect 674710 944621 674762 944673
rect 50326 944547 50378 944599
rect 59542 944547 59594 944599
rect 672310 942327 672362 942379
rect 674710 942327 674762 942379
rect 658102 942179 658154 942231
rect 674710 942179 674762 942231
rect 654358 942031 654410 942083
rect 674614 942031 674666 942083
rect 652246 941883 652298 941935
rect 674806 941883 674858 941935
rect 658006 939071 658058 939123
rect 674710 939071 674762 939123
rect 42358 930931 42410 930983
rect 44566 930931 44618 930983
rect 47542 930191 47594 930243
rect 59542 930191 59594 930243
rect 654454 927453 654506 927505
rect 666742 927453 666794 927505
rect 649558 927379 649610 927431
rect 679798 927379 679850 927431
rect 654454 915835 654506 915887
rect 660982 915835 661034 915887
rect 47446 912949 47498 913001
rect 59542 912949 59594 913001
rect 53206 901479 53258 901531
rect 58198 901479 58250 901531
rect 654454 901479 654506 901531
rect 663958 901479 664010 901531
rect 50422 884163 50474 884215
rect 59542 884163 59594 884215
rect 654454 878391 654506 878443
rect 660886 878391 660938 878443
rect 674998 872101 675050 872153
rect 675478 872101 675530 872153
rect 674518 871657 674570 871709
rect 675190 871657 675242 871709
rect 675382 871657 675434 871709
rect 674326 868993 674378 869045
rect 675478 868993 675530 869045
rect 674230 868327 674282 868379
rect 675382 868327 675434 868379
rect 673654 867809 673706 867861
rect 675382 867809 675434 867861
rect 654454 866921 654506 866973
rect 669622 866921 669674 866973
rect 666646 865293 666698 865345
rect 675382 865293 675434 865345
rect 674902 863961 674954 864013
rect 674998 863961 675050 864013
rect 50326 858263 50378 858315
rect 59542 858263 59594 858315
rect 654454 855377 654506 855429
rect 661174 855377 661226 855429
rect 675190 846645 675242 846697
rect 675382 846645 675434 846697
rect 53398 843833 53450 843885
rect 59542 843833 59594 843885
rect 674806 843833 674858 843885
rect 674902 843833 674954 843885
rect 654454 832363 654506 832415
rect 666838 832363 666890 832415
rect 50614 829477 50666 829529
rect 59542 829477 59594 829529
rect 675382 826591 675434 826643
rect 675574 826591 675626 826643
rect 42358 823853 42410 823905
rect 50422 823853 50474 823905
rect 42358 822225 42410 822277
rect 53206 822225 53258 822277
rect 42454 821855 42506 821907
rect 58966 821855 59018 821907
rect 654454 820819 654506 820871
rect 663766 820819 663818 820871
rect 47542 815047 47594 815099
rect 59542 815047 59594 815099
rect 654454 809275 654506 809327
rect 664054 809275 664106 809327
rect 650134 809201 650186 809253
rect 653782 809201 653834 809253
rect 42262 805131 42314 805183
rect 44758 805131 44810 805183
rect 42358 804391 42410 804443
rect 42934 804391 42986 804443
rect 42454 804095 42506 804147
rect 42742 804095 42794 804147
rect 40150 803429 40202 803481
rect 42454 803429 42506 803481
rect 41974 802393 42026 802445
rect 42838 802393 42890 802445
rect 43030 801579 43082 801631
rect 43414 801579 43466 801631
rect 43030 801431 43082 801483
rect 44854 801431 44906 801483
rect 53206 800617 53258 800669
rect 59542 800617 59594 800669
rect 41686 800543 41738 800595
rect 43510 800543 43562 800595
rect 41590 800469 41642 800521
rect 43318 800469 43370 800521
rect 41878 800173 41930 800225
rect 41878 799729 41930 799781
rect 42166 798027 42218 798079
rect 42454 798027 42506 798079
rect 42070 797287 42122 797339
rect 43030 797287 43082 797339
rect 43030 797139 43082 797191
rect 43318 797139 43370 797191
rect 42166 796251 42218 796303
rect 43126 796251 43178 796303
rect 43126 796103 43178 796155
rect 43414 796103 43466 796155
rect 42166 794993 42218 795045
rect 42742 794993 42794 795045
rect 42166 793809 42218 793861
rect 42454 793809 42506 793861
rect 42166 793143 42218 793195
rect 42838 793143 42890 793195
rect 43030 793069 43082 793121
rect 42838 792995 42890 793047
rect 42742 792921 42794 792973
rect 43030 792921 43082 792973
rect 42262 792107 42314 792159
rect 43126 792107 43178 792159
rect 42166 791959 42218 792011
rect 42454 791959 42506 792011
rect 43126 791959 43178 792011
rect 43510 791959 43562 792011
rect 674710 791959 674762 792011
rect 674902 791959 674954 792011
rect 42262 790109 42314 790161
rect 42838 790109 42890 790161
rect 42166 789887 42218 789939
rect 43030 789887 43082 789939
rect 42166 789443 42218 789495
rect 42934 789443 42986 789495
rect 42166 787001 42218 787053
rect 43126 787001 43178 787053
rect 42166 786409 42218 786461
rect 42742 786409 42794 786461
rect 654454 786261 654506 786313
rect 669718 786261 669770 786313
rect 42070 785743 42122 785795
rect 42454 785743 42506 785795
rect 674518 784929 674570 784981
rect 675382 784929 675434 784981
rect 672886 783449 672938 783501
rect 675286 783449 675338 783501
rect 674998 782857 675050 782909
rect 675286 782857 675338 782909
rect 672790 782191 672842 782243
rect 674614 782191 674666 782243
rect 675286 782191 675338 782243
rect 663862 780563 663914 780615
rect 675094 780563 675146 780615
rect 42742 780415 42794 780467
rect 50614 780415 50666 780467
rect 674902 780415 674954 780467
rect 675478 780415 675530 780467
rect 42454 779897 42506 779949
rect 47542 779897 47594 779949
rect 672502 779749 672554 779801
rect 675382 779749 675434 779801
rect 672214 779305 672266 779357
rect 675478 779305 675530 779357
rect 42742 778861 42794 778913
rect 53398 778861 53450 778913
rect 672598 778565 672650 778617
rect 675382 778565 675434 778617
rect 672022 777603 672074 777655
rect 675478 777603 675530 777655
rect 675094 777011 675146 777063
rect 675382 777011 675434 777063
rect 674230 775457 674282 775509
rect 675382 775457 675434 775509
rect 654454 774717 654506 774769
rect 669814 774717 669866 774769
rect 674326 773607 674378 773659
rect 675382 773607 675434 773659
rect 53398 771831 53450 771883
rect 59542 771831 59594 771883
rect 660982 767465 661034 767517
rect 674422 767465 674474 767517
rect 666742 766873 666794 766925
rect 674710 766873 674762 766925
rect 663958 765837 664010 765889
rect 674422 765837 674474 765889
rect 672310 765245 672362 765297
rect 674710 765245 674762 765297
rect 654454 763247 654506 763299
rect 661078 763247 661130 763299
rect 672694 763247 672746 763299
rect 674710 763247 674762 763299
rect 672406 762507 672458 762559
rect 674710 762507 674762 762559
rect 42742 762211 42794 762263
rect 44854 762211 44906 762263
rect 38998 760287 39050 760339
rect 42742 760287 42794 760339
rect 43126 759325 43178 759377
rect 43414 759325 43466 759377
rect 43030 757771 43082 757823
rect 44950 757771 45002 757823
rect 50422 757475 50474 757527
rect 59542 757475 59594 757527
rect 42454 757253 42506 757305
rect 43606 757253 43658 757305
rect 41974 757105 42026 757157
rect 43798 757105 43850 757157
rect 42070 757031 42122 757083
rect 43510 757031 43562 757083
rect 41782 756957 41834 757009
rect 41878 756957 41930 757009
rect 43702 756883 43754 756935
rect 41782 756735 41834 756787
rect 42070 754885 42122 754937
rect 42742 754885 42794 754937
rect 42454 754293 42506 754345
rect 42934 754293 42986 754345
rect 42166 754071 42218 754123
rect 43030 754071 43082 754123
rect 42070 753035 42122 753087
rect 43414 753035 43466 753087
rect 43222 752221 43274 752273
rect 43606 752221 43658 752273
rect 43126 751851 43178 751903
rect 42934 751777 42986 751829
rect 43126 751629 43178 751681
rect 43414 751629 43466 751681
rect 42070 751185 42122 751237
rect 42934 751185 42986 751237
rect 42742 750963 42794 751015
rect 43606 750963 43658 751015
rect 42166 750371 42218 750423
rect 43126 750371 43178 750423
rect 43126 750223 43178 750275
rect 43510 750223 43562 750275
rect 42070 749927 42122 749979
rect 43030 749927 43082 749979
rect 42262 748891 42314 748943
rect 42742 748891 42794 748943
rect 649654 748817 649706 748869
rect 679702 748817 679754 748869
rect 42070 746079 42122 746131
rect 43126 746079 43178 746131
rect 672790 745931 672842 745983
rect 674998 745931 675050 745983
rect 674710 745857 674762 745909
rect 674902 745857 674954 745909
rect 42166 745635 42218 745687
rect 42454 745635 42506 745687
rect 42166 743785 42218 743837
rect 42838 743785 42890 743837
rect 42070 743045 42122 743097
rect 42934 743045 42986 743097
rect 47542 743045 47594 743097
rect 59542 743045 59594 743097
rect 42166 742601 42218 742653
rect 42742 742601 42794 742653
rect 674038 741565 674090 741617
rect 674422 741565 674474 741617
rect 672310 738087 672362 738139
rect 674998 738087 675050 738139
rect 675478 738087 675530 738139
rect 674902 738013 674954 738065
rect 674998 737939 675050 737991
rect 674902 737865 674954 737917
rect 675382 737865 675434 737917
rect 660982 737347 661034 737399
rect 675190 737347 675242 737399
rect 654454 737273 654506 737325
rect 663958 737273 664010 737325
rect 42646 737199 42698 737251
rect 53398 737199 53450 737251
rect 42358 736681 42410 736733
rect 50422 736681 50474 736733
rect 674518 735645 674570 735697
rect 675478 735645 675530 735697
rect 42358 735423 42410 735475
rect 58966 735423 59018 735475
rect 672118 733573 672170 733625
rect 675478 733573 675530 733625
rect 674134 732315 674186 732367
rect 675478 732315 675530 732367
rect 675190 732019 675242 732071
rect 675382 732019 675434 732071
rect 674710 730465 674762 730517
rect 675478 730465 675530 730517
rect 50422 728615 50474 728667
rect 58390 728615 58442 728667
rect 674614 728615 674666 728667
rect 675478 728615 675530 728667
rect 669622 722473 669674 722525
rect 674422 722473 674474 722525
rect 660886 721733 660938 721785
rect 674422 721733 674474 721785
rect 661174 720845 661226 720897
rect 674422 720845 674474 720897
rect 671926 719143 671978 719195
rect 674422 719143 674474 719195
rect 672406 717663 672458 717715
rect 674422 717663 674474 717715
rect 43318 717219 43370 717271
rect 44950 717219 45002 717271
rect 40150 715887 40202 715939
rect 41878 715887 41930 715939
rect 672694 715295 672746 715347
rect 673654 715295 673706 715347
rect 53398 714259 53450 714311
rect 58390 714259 58442 714311
rect 654454 714259 654506 714311
rect 666934 714259 666986 714311
rect 41590 714037 41642 714089
rect 41686 714037 41738 714089
rect 43510 714037 43562 714089
rect 41782 713963 41834 714015
rect 43606 713963 43658 714015
rect 41782 713519 41834 713571
rect 42934 711743 42986 711795
rect 43510 711373 43562 711425
rect 43222 711225 43274 711277
rect 43702 711225 43754 711277
rect 42166 710781 42218 710833
rect 45142 710781 45194 710833
rect 672886 710485 672938 710537
rect 674422 710485 674474 710537
rect 42166 709893 42218 709945
rect 42358 709893 42410 709945
rect 672022 709893 672074 709945
rect 674806 709893 674858 709945
rect 672214 709005 672266 709057
rect 674422 709005 674474 709057
rect 42550 707895 42602 707947
rect 43414 707895 43466 707947
rect 42166 707377 42218 707429
rect 43030 707377 43082 707429
rect 672502 707377 672554 707429
rect 674422 707377 674474 707429
rect 43030 707229 43082 707281
rect 43606 707229 43658 707281
rect 672598 706785 672650 706837
rect 674806 706785 674858 706837
rect 42934 706415 42986 706467
rect 43510 706415 43562 706467
rect 42166 705823 42218 705875
rect 42262 705601 42314 705653
rect 42838 703603 42890 703655
rect 42070 703529 42122 703581
rect 42166 702863 42218 702915
rect 43030 702863 43082 702915
rect 649750 702715 649802 702767
rect 679702 702715 679754 702767
rect 42166 702271 42218 702323
rect 42550 702271 42602 702323
rect 42070 700569 42122 700621
rect 42934 700569 42986 700621
rect 42166 700051 42218 700103
rect 42838 700051 42890 700103
rect 42358 699829 42410 699881
rect 57814 699829 57866 699881
rect 672310 699829 672362 699881
rect 672598 699829 672650 699881
rect 42646 693983 42698 694035
rect 53398 693983 53450 694035
rect 672214 692873 672266 692925
rect 675382 692873 675434 692925
rect 672598 692651 672650 692703
rect 675478 692651 675530 692703
rect 42646 692429 42698 692481
rect 50422 692429 50474 692481
rect 654454 691245 654506 691297
rect 661270 691245 661322 691297
rect 674326 690653 674378 690705
rect 675478 690653 675530 690705
rect 675094 689765 675146 689817
rect 675382 689765 675434 689817
rect 674422 689321 674474 689373
rect 675382 689321 675434 689373
rect 672022 688581 672074 688633
rect 675478 688581 675530 688633
rect 674230 687323 674282 687375
rect 675478 687323 675530 687375
rect 669622 686213 669674 686265
rect 675382 686213 675434 686265
rect 50422 685473 50474 685525
rect 59542 685473 59594 685525
rect 674806 685473 674858 685525
rect 675478 685473 675530 685525
rect 674902 683623 674954 683675
rect 675478 683623 675530 683675
rect 663766 677333 663818 677385
rect 674422 677333 674474 677385
rect 666838 676445 666890 676497
rect 674422 676445 674474 676497
rect 42742 676297 42794 676349
rect 42646 676001 42698 676053
rect 664054 675705 664106 675757
rect 674422 675705 674474 675757
rect 42358 675631 42410 675683
rect 47734 675631 47786 675683
rect 671926 674817 671978 674869
rect 674422 674817 674474 674869
rect 41878 674521 41930 674573
rect 43126 674521 43178 674573
rect 672502 674003 672554 674055
rect 674422 674003 674474 674055
rect 43318 673781 43370 673833
rect 45046 673781 45098 673833
rect 40246 672375 40298 672427
rect 41878 672375 41930 672427
rect 42070 671931 42122 671983
rect 42454 671931 42506 671983
rect 53398 671043 53450 671095
rect 59446 671043 59498 671095
rect 672406 670969 672458 671021
rect 675190 670969 675242 671021
rect 41302 670895 41354 670947
rect 42934 670895 42986 670947
rect 43222 670895 43274 670947
rect 43606 670895 43658 670947
rect 42262 670747 42314 670799
rect 43414 670747 43466 670799
rect 41974 670673 42026 670725
rect 43126 670673 43178 670725
rect 41782 670599 41834 670651
rect 41878 670599 41930 670651
rect 42934 670525 42986 670577
rect 41782 670303 41834 670355
rect 42166 668527 42218 668579
rect 42934 668527 42986 668579
rect 42934 668379 42986 668431
rect 43222 668379 43274 668431
rect 654454 668157 654506 668209
rect 664054 668157 664106 668209
rect 649846 668083 649898 668135
rect 652246 668083 652298 668135
rect 42166 667861 42218 667913
rect 43318 667861 43370 667913
rect 42166 665345 42218 665397
rect 42934 665345 42986 665397
rect 42934 665197 42986 665249
rect 43414 665197 43466 665249
rect 42166 664827 42218 664879
rect 43030 664827 43082 664879
rect 42070 663939 42122 663991
rect 42550 663939 42602 663991
rect 42166 663347 42218 663399
rect 42550 663347 42602 663399
rect 42262 662385 42314 662437
rect 42934 662385 42986 662437
rect 42934 662237 42986 662289
rect 43606 662237 43658 662289
rect 672118 661349 672170 661401
rect 674422 661349 674474 661401
rect 42070 661053 42122 661105
rect 43126 661053 43178 661105
rect 42166 659869 42218 659921
rect 42838 659869 42890 659921
rect 42070 659055 42122 659107
rect 43030 659055 43082 659107
rect 42166 656835 42218 656887
rect 42934 656835 42986 656887
rect 42838 656687 42890 656739
rect 59542 656687 59594 656739
rect 649846 656687 649898 656739
rect 679702 656687 679754 656739
rect 674422 656095 674474 656147
rect 674902 656095 674954 656147
rect 672598 653727 672650 653779
rect 674998 653727 675050 653779
rect 42454 649731 42506 649783
rect 51862 649731 51914 649783
rect 42454 649509 42506 649561
rect 53398 649509 53450 649561
rect 674902 649509 674954 649561
rect 675190 649509 675242 649561
rect 671926 648251 671978 648303
rect 675286 648251 675338 648303
rect 672886 648029 672938 648081
rect 675286 648029 675338 648081
rect 675094 647807 675146 647859
rect 675094 647511 675146 647563
rect 674518 646401 674570 646453
rect 674902 646401 674954 646453
rect 675382 646401 675434 646453
rect 674614 645291 674666 645343
rect 675190 645291 675242 645343
rect 654454 645217 654506 645269
rect 666838 645217 666890 645269
rect 666742 645143 666794 645195
rect 675190 645143 675242 645195
rect 671638 644773 671690 644825
rect 675382 644773 675434 644825
rect 51862 644477 51914 644529
rect 59254 644477 59306 644529
rect 672310 644033 672362 644085
rect 675478 644033 675530 644085
rect 672598 643367 672650 643419
rect 675382 643367 675434 643419
rect 671446 642257 671498 642309
rect 675478 642257 675530 642309
rect 675190 641813 675242 641865
rect 675382 641813 675434 641865
rect 669814 632489 669866 632541
rect 674710 632489 674762 632541
rect 42454 632415 42506 632467
rect 45046 632415 45098 632467
rect 43126 632119 43178 632171
rect 43702 632119 43754 632171
rect 669718 631749 669770 631801
rect 674710 631749 674762 631801
rect 661078 630565 661130 630617
rect 674134 630565 674186 630617
rect 672502 630269 672554 630321
rect 673846 630269 673898 630321
rect 671734 628419 671786 628471
rect 673846 628419 673898 628471
rect 670966 628123 671018 628175
rect 672694 628123 672746 628175
rect 673846 628123 673898 628175
rect 42454 627901 42506 627953
rect 47830 627901 47882 627953
rect 40054 627827 40106 627879
rect 42934 627827 42986 627879
rect 47638 627827 47690 627879
rect 58006 627827 58058 627879
rect 670870 627753 670922 627805
rect 675190 627753 675242 627805
rect 41494 627679 41546 627731
rect 43126 627679 43178 627731
rect 42646 627605 42698 627657
rect 43318 627605 43370 627657
rect 43030 627531 43082 627583
rect 43414 627531 43466 627583
rect 41782 627383 41834 627435
rect 41974 627383 42026 627435
rect 42070 627383 42122 627435
rect 43030 627383 43082 627435
rect 43510 627309 43562 627361
rect 41782 627161 41834 627213
rect 42166 625311 42218 625363
rect 42934 625311 42986 625363
rect 42934 625163 42986 625215
rect 43318 625163 43370 625215
rect 674614 624867 674666 624919
rect 674902 624867 674954 624919
rect 42166 624645 42218 624697
rect 42454 624645 42506 624697
rect 42454 623757 42506 623809
rect 43702 623757 43754 623809
rect 42166 622203 42218 622255
rect 43414 622203 43466 622255
rect 656374 622055 656426 622107
rect 669718 622055 669770 622107
rect 42166 621611 42218 621663
rect 43030 621611 43082 621663
rect 43030 621463 43082 621515
rect 43510 621463 43562 621515
rect 42070 620871 42122 620923
rect 42934 620871 42986 620923
rect 672214 619169 672266 619221
rect 673846 619169 673898 619221
rect 672022 617837 672074 617889
rect 673846 617837 673898 617889
rect 42070 617615 42122 617667
rect 42934 617615 42986 617667
rect 42166 617319 42218 617371
rect 43126 617319 43178 617371
rect 42166 616653 42218 616705
rect 43030 616653 43082 616705
rect 42166 615987 42218 616039
rect 42454 615987 42506 616039
rect 42166 613989 42218 614041
rect 42454 613989 42506 614041
rect 42166 613619 42218 613671
rect 42742 613619 42794 613671
rect 42454 613471 42506 613523
rect 59446 613471 59498 613523
rect 649942 613471 649994 613523
rect 679702 613471 679754 613523
rect 654454 613397 654506 613449
rect 669526 613397 669578 613449
rect 42070 612805 42122 612857
rect 42838 612805 42890 612857
rect 42742 607699 42794 607751
rect 51862 607699 51914 607751
rect 42742 606811 42794 606863
rect 53398 606811 53450 606863
rect 671830 603851 671882 603903
rect 675094 603851 675146 603903
rect 672214 603629 672266 603681
rect 674518 603629 674570 603681
rect 675286 603629 675338 603681
rect 673750 602815 673802 602867
rect 674710 602815 674762 602867
rect 675478 602815 675530 602867
rect 673174 602667 673226 602719
rect 675382 602667 675434 602719
rect 663766 602001 663818 602053
rect 675190 602001 675242 602053
rect 672694 601927 672746 601979
rect 675094 601927 675146 601979
rect 51862 601853 51914 601905
rect 59542 601853 59594 601905
rect 672022 599559 672074 599611
rect 675382 599559 675434 599611
rect 671542 599263 671594 599315
rect 675382 599263 675434 599315
rect 654454 599041 654506 599093
rect 669526 599041 669578 599093
rect 672118 598375 672170 598427
rect 675478 598375 675530 598427
rect 672502 597117 672554 597169
rect 675478 597117 675530 597169
rect 675190 596821 675242 596873
rect 675382 596821 675434 596873
rect 42454 589199 42506 589251
rect 45142 589199 45194 589251
rect 670870 587497 670922 587549
rect 676822 587497 676874 587549
rect 53398 587423 53450 587475
rect 59542 587423 59594 587475
rect 663958 586313 664010 586365
rect 674422 586313 674474 586365
rect 40054 585943 40106 585995
rect 42454 585943 42506 585995
rect 666934 585425 666986 585477
rect 674422 585425 674474 585477
rect 43126 585351 43178 585403
rect 43702 585351 43754 585403
rect 671734 584833 671786 584885
rect 674614 584833 674666 584885
rect 42550 584759 42602 584811
rect 43126 584759 43178 584811
rect 655222 584759 655274 584811
rect 674710 584759 674762 584811
rect 42838 584685 42890 584737
rect 50518 584685 50570 584737
rect 41974 584241 42026 584293
rect 43222 584241 43274 584293
rect 41782 584167 41834 584219
rect 42166 584167 42218 584219
rect 42934 584167 42986 584219
rect 41782 583945 41834 583997
rect 672406 583575 672458 583627
rect 674710 583575 674762 583627
rect 675190 582539 675242 582591
rect 676822 582539 676874 582591
rect 42166 582095 42218 582147
rect 42454 582095 42506 582147
rect 42070 581429 42122 581481
rect 42838 581429 42890 581481
rect 42838 581281 42890 581333
rect 43222 581281 43274 581333
rect 42070 580245 42122 580297
rect 43030 580245 43082 580297
rect 42166 578987 42218 579039
rect 43318 578987 43370 579039
rect 672406 578839 672458 578891
rect 672790 578839 672842 578891
rect 42070 578395 42122 578447
rect 42934 578395 42986 578447
rect 42166 577655 42218 577707
rect 43126 577655 43178 577707
rect 43126 577507 43178 577559
rect 43702 577507 43754 577559
rect 671926 575361 671978 575413
rect 674710 575361 674762 575413
rect 671446 574473 671498 574525
rect 674710 574473 674762 574525
rect 42166 574103 42218 574155
rect 42838 574103 42890 574155
rect 672310 573585 672362 573637
rect 674422 573585 674474 573637
rect 42070 573215 42122 573267
rect 43030 573215 43082 573267
rect 654454 573141 654506 573193
rect 661174 573141 661226 573193
rect 672886 572993 672938 573045
rect 674710 572993 674762 573045
rect 42166 572623 42218 572675
rect 42934 572623 42986 572675
rect 671638 571957 671690 572009
rect 674422 571957 674474 572009
rect 672598 571365 672650 571417
rect 674710 571365 674762 571417
rect 42166 570995 42218 571047
rect 43126 570995 43178 571047
rect 42070 570403 42122 570455
rect 42454 570403 42506 570455
rect 42358 570255 42410 570307
rect 59542 570255 59594 570307
rect 42070 569663 42122 569715
rect 42934 569663 42986 569715
rect 650038 567369 650090 567421
rect 679798 567369 679850 567421
rect 34486 564483 34538 564535
rect 53398 564483 53450 564535
rect 654454 564409 654506 564461
rect 666646 564409 666698 564461
rect 672214 564409 672266 564461
rect 674998 564409 675050 564461
rect 672214 564261 672266 564313
rect 672790 564261 672842 564313
rect 42454 563447 42506 563499
rect 50518 563447 50570 563499
rect 673750 561597 673802 561649
rect 675094 561597 675146 561649
rect 674326 559525 674378 559577
rect 675382 559525 675434 559577
rect 53398 558637 53450 558689
rect 59542 558637 59594 558689
rect 673942 558045 673994 558097
rect 675382 558045 675434 558097
rect 660886 555825 660938 555877
rect 675190 555825 675242 555877
rect 674518 555011 674570 555063
rect 675478 555011 675530 555063
rect 675094 554493 675146 554545
rect 675382 554493 675434 554545
rect 674134 553901 674186 553953
rect 675478 553901 675530 553953
rect 674806 553161 674858 553213
rect 675382 553161 675434 553213
rect 674422 551903 674474 551955
rect 675478 551903 675530 551955
rect 675190 551607 675242 551659
rect 675382 551607 675434 551659
rect 654454 550127 654506 550179
rect 663958 550127 664010 550179
rect 675190 550053 675242 550105
rect 675478 550053 675530 550105
rect 674614 548203 674666 548255
rect 675382 548203 675434 548255
rect 42646 546205 42698 546257
rect 45238 546205 45290 546257
rect 42358 545539 42410 545591
rect 42646 545539 42698 545591
rect 42838 544947 42890 544999
rect 42838 544577 42890 544629
rect 40054 544281 40106 544333
rect 42934 544281 42986 544333
rect 50518 543689 50570 543741
rect 59542 543689 59594 543741
rect 43702 541469 43754 541521
rect 53302 541469 53354 541521
rect 655414 541469 655466 541521
rect 674710 541469 674762 541521
rect 672214 541395 672266 541447
rect 673846 541395 673898 541447
rect 661270 541321 661322 541373
rect 674230 541321 674282 541373
rect 674710 541321 674762 541373
rect 675190 541321 675242 541373
rect 41974 541025 42026 541077
rect 43510 541025 43562 541077
rect 41782 540951 41834 541003
rect 42166 540951 42218 541003
rect 43318 540951 43370 541003
rect 41782 540729 41834 540781
rect 664054 540433 664106 540485
rect 674230 540433 674282 540485
rect 42934 540063 42986 540115
rect 43030 539841 43082 539893
rect 42070 538879 42122 538931
rect 43030 538879 43082 538931
rect 654454 538583 654506 538635
rect 661078 538583 661130 538635
rect 674038 538583 674090 538635
rect 675094 538583 675146 538635
rect 42166 538139 42218 538191
rect 43702 538139 43754 538191
rect 42070 537029 42122 537081
rect 42934 537029 42986 537081
rect 42070 535771 42122 535823
rect 42838 535771 42890 535823
rect 42166 535031 42218 535083
rect 42742 535031 42794 535083
rect 42166 534439 42218 534491
rect 43126 534439 43178 534491
rect 43222 534439 43274 534491
rect 43222 534217 43274 534269
rect 42070 533921 42122 533973
rect 43030 533921 43082 533973
rect 43030 533773 43082 533825
rect 43510 533773 43562 533825
rect 42262 532811 42314 532863
rect 42646 532811 42698 532863
rect 672694 532737 672746 532789
rect 673846 532737 673898 532789
rect 671830 532663 671882 532715
rect 673750 532663 673802 532715
rect 42166 531331 42218 531383
rect 43126 531331 43178 531383
rect 42262 530295 42314 530347
rect 42934 530295 42986 530347
rect 42070 530147 42122 530199
rect 42838 530147 42890 530199
rect 672502 529851 672554 529903
rect 673846 529851 673898 529903
rect 671542 529185 671594 529237
rect 673846 529185 673898 529237
rect 42166 527631 42218 527683
rect 43030 527631 43082 527683
rect 42070 527187 42122 527239
rect 42742 527187 42794 527239
rect 42358 527039 42410 527091
rect 59542 527039 59594 527091
rect 654454 527039 654506 527091
rect 669814 527039 669866 527091
rect 672022 526891 672074 526943
rect 673846 526891 673898 526943
rect 672118 526743 672170 526795
rect 673846 526743 673898 526795
rect 42166 526595 42218 526647
rect 42646 526595 42698 526647
rect 650134 521267 650186 521319
rect 679798 521267 679850 521319
rect 674518 518307 674570 518359
rect 674902 518307 674954 518359
rect 654070 517271 654122 517323
rect 663862 517271 663914 517323
rect 50518 512683 50570 512735
rect 59350 512683 59402 512735
rect 673942 508317 673994 508369
rect 674134 508317 674186 508369
rect 674326 508095 674378 508147
rect 674326 507873 674378 507925
rect 674422 507873 674474 507925
rect 674902 507873 674954 507925
rect 654934 504025 654986 504077
rect 666646 504025 666698 504077
rect 53398 498253 53450 498305
rect 57814 498253 57866 498305
rect 666838 497513 666890 497565
rect 674518 497513 674570 497565
rect 669718 496625 669770 496677
rect 674518 496625 674570 496677
rect 655318 495515 655370 495567
rect 674710 495515 674762 495567
rect 53302 483823 53354 483875
rect 59542 483823 59594 483875
rect 654454 480937 654506 480989
rect 666838 480937 666890 480989
rect 650230 478125 650282 478177
rect 679798 478125 679850 478177
rect 654454 470577 654506 470629
rect 660982 470577 661034 470629
rect 50614 469467 50666 469519
rect 59542 469467 59594 469519
rect 656374 457923 656426 457975
rect 663862 457923 663914 457975
rect 45430 455037 45482 455089
rect 59542 455037 59594 455089
rect 654454 446379 654506 446431
rect 669718 446379 669770 446431
rect 45334 440681 45386 440733
rect 57814 440681 57866 440733
rect 42646 436907 42698 436959
rect 50518 436907 50570 436959
rect 42646 436093 42698 436145
rect 53398 436093 53450 436145
rect 654454 434909 654506 434961
rect 664054 434909 664106 434961
rect 53398 426251 53450 426303
rect 59542 426251 59594 426303
rect 654454 423291 654506 423343
rect 669622 423291 669674 423343
rect 42166 419961 42218 420013
rect 42358 419961 42410 420013
rect 42646 418555 42698 418607
rect 44662 418555 44714 418607
rect 37366 416927 37418 416979
rect 42934 416927 42986 416979
rect 40150 416187 40202 416239
rect 43126 416187 43178 416239
rect 40246 414781 40298 414833
rect 42838 414781 42890 414833
rect 37270 414707 37322 414759
rect 43318 414707 43370 414759
rect 41782 413375 41834 413427
rect 41782 413153 41834 413205
rect 53494 411821 53546 411873
rect 59542 411821 59594 411873
rect 42166 411303 42218 411355
rect 42358 411303 42410 411355
rect 42070 410489 42122 410541
rect 47446 410489 47498 410541
rect 42166 409453 42218 409505
rect 42742 409453 42794 409505
rect 42838 409379 42890 409431
rect 43030 409231 43082 409283
rect 42838 409157 42890 409209
rect 669526 409157 669578 409209
rect 674422 409157 674474 409209
rect 655126 409083 655178 409135
rect 674710 409083 674762 409135
rect 43030 409009 43082 409061
rect 43126 409009 43178 409061
rect 43318 409009 43370 409061
rect 654454 408935 654506 408987
rect 669622 408935 669674 408987
rect 661174 408417 661226 408469
rect 674710 408417 674762 408469
rect 42166 408195 42218 408247
rect 42838 408195 42890 408247
rect 42070 407455 42122 407507
rect 42934 407455 42986 407507
rect 42166 406863 42218 406915
rect 43030 406863 43082 406915
rect 42166 403829 42218 403881
rect 43126 403829 43178 403881
rect 42166 403311 42218 403363
rect 42742 403311 42794 403363
rect 654646 397465 654698 397517
rect 661174 397465 661226 397517
rect 42358 393913 42410 393965
rect 50614 393913 50666 393965
rect 42358 393173 42410 393225
rect 45430 393173 45482 393225
rect 42358 392285 42410 392337
rect 53302 392285 53354 392337
rect 650326 391693 650378 391745
rect 679702 391693 679754 391745
rect 654454 385921 654506 385973
rect 669526 385921 669578 385973
rect 674902 384885 674954 384937
rect 675286 384885 675338 384937
rect 674518 384293 674570 384345
rect 675094 384293 675146 384345
rect 674038 383109 674090 383161
rect 675382 383109 675434 383161
rect 45430 383035 45482 383087
rect 59542 383035 59594 383087
rect 674710 378151 674762 378203
rect 675382 378151 675434 378203
rect 674422 377559 674474 377611
rect 675382 377559 675434 377611
rect 654454 377189 654506 377241
rect 666742 377189 666794 377241
rect 674326 376819 674378 376871
rect 675478 376819 675530 376871
rect 673942 375709 673994 375761
rect 675478 375709 675530 375761
rect 42358 375191 42410 375243
rect 47446 375191 47498 375243
rect 37174 371861 37226 371913
rect 43318 371861 43370 371913
rect 37270 371787 37322 371839
rect 43126 371787 43178 371839
rect 37366 371713 37418 371765
rect 42838 371713 42890 371765
rect 40150 371639 40202 371691
rect 42742 371639 42794 371691
rect 40054 371565 40106 371617
rect 42358 371565 42410 371617
rect 41782 370159 41834 370211
rect 41782 369937 41834 369989
rect 50518 368679 50570 368731
rect 59542 368679 59594 368731
rect 42070 368087 42122 368139
rect 43030 368087 43082 368139
rect 43030 367939 43082 367991
rect 43318 367939 43370 367991
rect 42070 367347 42122 367399
rect 50326 367347 50378 367399
rect 42070 366237 42122 366289
rect 42358 366237 42410 366289
rect 42358 366089 42410 366141
rect 43126 366089 43178 366141
rect 42166 364979 42218 365031
rect 42742 364979 42794 365031
rect 661078 364905 661130 364957
rect 674710 364905 674762 364957
rect 42070 364387 42122 364439
rect 42934 364387 42986 364439
rect 663958 363869 664010 363921
rect 674422 363869 674474 363921
rect 42166 363647 42218 363699
rect 42838 363647 42890 363699
rect 654454 363499 654506 363551
rect 660982 363499 661034 363551
rect 669814 363277 669866 363329
rect 674710 363277 674762 363329
rect 42358 360095 42410 360147
rect 43030 360095 43082 360147
rect 47830 354249 47882 354301
rect 59542 354249 59594 354301
rect 42358 350697 42410 350749
rect 53398 350697 53450 350749
rect 42646 349661 42698 349713
rect 53494 349661 53546 349713
rect 42358 349069 42410 349121
rect 45334 349069 45386 349121
rect 650422 345591 650474 345643
rect 679798 345591 679850 345643
rect 674614 340929 674666 340981
rect 675478 340929 675530 340981
rect 53302 339819 53354 339871
rect 59542 339819 59594 339871
rect 654454 339819 654506 339871
rect 666742 339819 666794 339871
rect 674038 339523 674090 339575
rect 675382 339523 675434 339575
rect 674518 336563 674570 336615
rect 675382 336563 675434 336615
rect 674326 332715 674378 332767
rect 675382 332715 675434 332767
rect 674230 332197 674282 332249
rect 675478 332197 675530 332249
rect 42166 331975 42218 332027
rect 47926 331975 47978 332027
rect 674134 331531 674186 331583
rect 675382 331531 675434 331583
rect 39958 331161 40010 331213
rect 41782 331161 41834 331213
rect 37174 330421 37226 330473
rect 40534 330421 40586 330473
rect 654070 329607 654122 329659
rect 663766 329607 663818 329659
rect 40246 328497 40298 328549
rect 43030 328497 43082 328549
rect 40054 328349 40106 328401
rect 43126 328275 43178 328327
rect 43318 328275 43370 328327
rect 43030 328053 43082 328105
rect 40534 327313 40586 327365
rect 42358 327313 42410 327365
rect 41782 327017 41834 327069
rect 41782 326721 41834 326773
rect 53398 325463 53450 325515
rect 59542 325463 59594 325515
rect 42070 324871 42122 324923
rect 42742 324871 42794 324923
rect 42454 324353 42506 324405
rect 43318 324353 43370 324405
rect 42166 324131 42218 324183
rect 53206 324131 53258 324183
rect 42166 323095 42218 323147
rect 42358 323095 42410 323147
rect 42070 321763 42122 321815
rect 43126 321763 43178 321815
rect 42166 321023 42218 321075
rect 43030 321023 43082 321075
rect 42166 320579 42218 320631
rect 42454 320579 42506 320631
rect 655222 319691 655274 319743
rect 674422 319691 674474 319743
rect 666646 318877 666698 318929
rect 674422 318877 674474 318929
rect 666838 318285 666890 318337
rect 674710 318285 674762 318337
rect 45334 311033 45386 311085
rect 59542 311033 59594 311085
rect 42262 307481 42314 307533
rect 45430 307481 45482 307533
rect 42262 306741 42314 306793
rect 50518 306741 50570 306793
rect 42838 305483 42890 305535
rect 58966 305483 59018 305535
rect 650518 299563 650570 299615
rect 679798 299563 679850 299615
rect 674806 299489 674858 299541
rect 676822 299489 676874 299541
rect 674902 299415 674954 299467
rect 676918 299415 676970 299467
rect 675286 299341 675338 299393
rect 677110 299341 677162 299393
rect 45430 296677 45482 296729
rect 59542 296677 59594 296729
rect 674326 295937 674378 295989
rect 675382 295937 675434 295989
rect 674518 295345 674570 295397
rect 675478 295345 675530 295397
rect 673942 294531 673994 294583
rect 675382 294531 675434 294583
rect 674422 291053 674474 291105
rect 675094 291053 675146 291105
rect 42646 289055 42698 289107
rect 48022 289055 48074 289107
rect 41974 288907 42026 288959
rect 42550 288907 42602 288959
rect 674902 288537 674954 288589
rect 675478 288537 675530 288589
rect 39958 287945 40010 287997
rect 41782 287945 41834 287997
rect 674230 287723 674282 287775
rect 675382 287723 675434 287775
rect 674806 287353 674858 287405
rect 675478 287353 675530 287405
rect 37366 286835 37418 286887
rect 42742 286835 42794 286887
rect 674134 286539 674186 286591
rect 675382 286539 675434 286591
rect 40150 285651 40202 285703
rect 43126 285651 43178 285703
rect 40246 285133 40298 285185
rect 42646 285133 42698 285185
rect 41782 283801 41834 283853
rect 42166 283801 42218 283853
rect 43318 283801 43370 283853
rect 41782 283357 41834 283409
rect 654454 282987 654506 283039
rect 660886 282987 660938 283039
rect 45526 282247 45578 282299
rect 59542 282247 59594 282299
rect 42166 281729 42218 281781
rect 42550 281729 42602 281781
rect 42166 281063 42218 281115
rect 47542 281063 47594 281115
rect 42166 279879 42218 279931
rect 42742 279879 42794 279931
rect 42166 278547 42218 278599
rect 42646 278547 42698 278599
rect 42166 277807 42218 277859
rect 43126 277807 43178 277859
rect 43222 277807 43274 277859
rect 43222 277585 43274 277637
rect 42070 277363 42122 277415
rect 42838 277363 42890 277415
rect 303382 276327 303434 276379
rect 435382 276327 435434 276379
rect 117238 276253 117290 276305
rect 397558 276253 397610 276305
rect 120790 276179 120842 276231
rect 398518 276179 398570 276231
rect 73270 276105 73322 276157
rect 386326 276105 386378 276157
rect 113782 276031 113834 276083
rect 396790 276031 396842 276083
rect 303574 275957 303626 276009
rect 439030 275957 439082 276009
rect 303958 275883 304010 275935
rect 442582 275883 442634 275935
rect 304438 275809 304490 275861
rect 446326 275809 446378 275861
rect 305110 275735 305162 275787
rect 449686 275735 449738 275787
rect 305206 275661 305258 275713
rect 453238 275661 453290 275713
rect 421846 275587 421898 275639
rect 649462 275587 649514 275639
rect 306646 275513 306698 275565
rect 464374 275513 464426 275565
rect 307222 275439 307274 275491
rect 467830 275439 467882 275491
rect 307702 275365 307754 275417
rect 471382 275365 471434 275417
rect 307894 275291 307946 275343
rect 475030 275291 475082 275343
rect 308374 275217 308426 275269
rect 478582 275217 478634 275269
rect 308758 275143 308810 275195
rect 481846 275143 481898 275195
rect 309430 275069 309482 275121
rect 485686 275069 485738 275121
rect 64918 274995 64970 275047
rect 181366 274995 181418 275047
rect 309910 274995 309962 275047
rect 489238 274995 489290 275047
rect 573142 274995 573194 275047
rect 649366 274995 649418 275047
rect 310102 274921 310154 274973
rect 492886 274921 492938 274973
rect 669718 274921 669770 274973
rect 674710 274921 674762 274973
rect 310486 274847 310538 274899
rect 496438 274847 496490 274899
rect 311638 274773 311690 274825
rect 503542 274773 503594 274825
rect 310966 274699 311018 274751
rect 499894 274699 499946 274751
rect 42262 274625 42314 274677
rect 42742 274625 42794 274677
rect 312118 274625 312170 274677
rect 507094 274625 507146 274677
rect 312214 274551 312266 274603
rect 510742 274551 510794 274603
rect 312694 274477 312746 274529
rect 514294 274477 514346 274529
rect 313174 274403 313226 274455
rect 517750 274403 517802 274455
rect 313750 274329 313802 274381
rect 521398 274329 521450 274381
rect 314710 274255 314762 274307
rect 528214 274255 528266 274307
rect 314902 274181 314954 274233
rect 532150 274181 532202 274233
rect 42070 274107 42122 274159
rect 43030 274107 43082 274159
rect 315286 274107 315338 274159
rect 535606 274107 535658 274159
rect 315958 274033 316010 274085
rect 539254 274033 539306 274085
rect 663862 274033 663914 274085
rect 674710 274033 674762 274085
rect 316438 273959 316490 274011
rect 542806 273959 542858 274011
rect 316630 273885 316682 273937
rect 546358 273885 546410 273937
rect 358294 273811 358346 273863
rect 429814 273811 429866 273863
rect 42262 273737 42314 273789
rect 43126 273737 43178 273789
rect 302902 273737 302954 273789
rect 432214 273737 432266 273789
rect 262102 273663 262154 273715
rect 337558 273663 337610 273715
rect 358390 273663 358442 273715
rect 433366 273663 433418 273715
rect 306166 273589 306218 273641
rect 460726 273589 460778 273641
rect 239734 273515 239786 273567
rect 370294 273515 370346 273567
rect 375670 273515 375722 273567
rect 488086 273515 488138 273567
rect 240406 273441 240458 273493
rect 377494 273441 377546 273493
rect 380662 273441 380714 273493
rect 550102 273441 550154 273493
rect 241462 273367 241514 273419
rect 384598 273367 384650 273419
rect 242134 273293 242186 273345
rect 391702 273293 391754 273345
rect 664054 273293 664106 273345
rect 674710 273293 674762 273345
rect 243190 273219 243242 273271
rect 398902 273219 398954 273271
rect 243862 273145 243914 273197
rect 406006 273145 406058 273197
rect 244726 273071 244778 273123
rect 413206 273071 413258 273123
rect 245878 272997 245930 273049
rect 419926 272997 419978 273049
rect 246454 272923 246506 272975
rect 427414 272923 427466 272975
rect 247606 272849 247658 272901
rect 434518 272849 434570 272901
rect 229078 272775 229130 272827
rect 284662 272775 284714 272827
rect 322102 272775 322154 272827
rect 230134 272701 230186 272753
rect 291862 272701 291914 272753
rect 322966 272701 323018 272753
rect 327862 272775 327914 272827
rect 582070 272775 582122 272827
rect 230806 272627 230858 272679
rect 298966 272627 299018 272679
rect 323542 272627 323594 272679
rect 589174 272701 589226 272753
rect 231862 272553 231914 272605
rect 306070 272553 306122 272605
rect 324694 272553 324746 272605
rect 596374 272627 596426 272679
rect 64822 272479 64874 272531
rect 72022 272479 72074 272531
rect 261046 272479 261098 272531
rect 327382 272479 327434 272531
rect 232726 272405 232778 272457
rect 313270 272405 313322 272457
rect 325270 272405 325322 272457
rect 603478 272553 603530 272605
rect 327574 272479 327626 272531
rect 545206 272479 545258 272531
rect 233398 272331 233450 272383
rect 320374 272331 320426 272383
rect 326230 272331 326282 272383
rect 610582 272405 610634 272457
rect 64726 272257 64778 272309
rect 66838 272257 66890 272309
rect 234454 272257 234506 272309
rect 327190 272257 327242 272309
rect 617686 272331 617738 272383
rect 624886 272257 624938 272309
rect 266518 272183 266570 272235
rect 591574 272183 591626 272235
rect 267190 272109 267242 272161
rect 595126 272109 595178 272161
rect 228118 272035 228170 272087
rect 277558 272035 277610 272087
rect 302230 272035 302282 272087
rect 428662 272035 428714 272087
rect 238870 271961 238922 272013
rect 363190 271961 363242 272013
rect 364630 271961 364682 272013
rect 393046 271961 393098 272013
rect 227926 271887 227978 271939
rect 274006 271887 274058 271939
rect 301366 271887 301418 271939
rect 387478 271887 387530 271939
rect 387670 271887 387722 271939
rect 421462 271887 421514 271939
rect 237718 271813 237770 271865
rect 356086 271813 356138 271865
rect 374134 271813 374186 271865
rect 387382 271813 387434 271865
rect 393046 271813 393098 271865
rect 426262 271813 426314 271865
rect 237142 271739 237194 271791
rect 348982 271739 349034 271791
rect 356278 271739 356330 271791
rect 415606 271739 415658 271791
rect 227446 271665 227498 271717
rect 270358 271665 270410 271717
rect 300310 271665 300362 271717
rect 410806 271665 410858 271717
rect 299158 271591 299210 271643
rect 403606 271591 403658 271643
rect 235990 271517 236042 271569
rect 341782 271517 341834 271569
rect 362806 271517 362858 271569
rect 383350 271517 383402 271569
rect 387286 271517 387338 271569
rect 394774 271517 394826 271569
rect 327286 271443 327338 271495
rect 588886 271443 588938 271495
rect 235126 271369 235178 271421
rect 334582 271369 334634 271421
rect 378454 271369 378506 271421
rect 407350 271369 407402 271421
rect 298486 271295 298538 271347
rect 396502 271295 396554 271347
rect 237430 271221 237482 271273
rect 331030 271221 331082 271273
rect 376246 271221 376298 271273
rect 459862 271221 459914 271273
rect 294838 271147 294890 271199
rect 367894 271147 367946 271199
rect 377206 271147 377258 271199
rect 387286 271147 387338 271199
rect 387382 271147 387434 271199
rect 472342 271147 472394 271199
rect 296566 271073 296618 271125
rect 382294 271073 382346 271125
rect 295894 270999 295946 271051
rect 375094 270999 375146 271051
rect 379414 270999 379466 271051
rect 394678 270999 394730 271051
rect 394774 270999 394826 271051
rect 502678 270999 502730 271051
rect 297430 270925 297482 270977
rect 389014 270925 389066 270977
rect 247894 270851 247946 270903
rect 327766 270851 327818 270903
rect 328918 270851 328970 270903
rect 562198 270851 562250 270903
rect 320950 270777 321002 270829
rect 327862 270777 327914 270829
rect 327958 270777 328010 270829
rect 570262 270777 570314 270829
rect 216790 270703 216842 270755
rect 228886 270703 228938 270755
rect 230038 270703 230090 270755
rect 333334 270703 333386 270755
rect 382198 270703 382250 270755
rect 124150 270629 124202 270681
rect 220630 270629 220682 270681
rect 220726 270629 220778 270681
rect 327094 270629 327146 270681
rect 329878 270629 329930 270681
rect 345814 270629 345866 270681
rect 351190 270629 351242 270681
rect 372694 270629 372746 270681
rect 374422 270629 374474 270681
rect 387286 270629 387338 270681
rect 387382 270629 387434 270681
rect 390358 270629 390410 270681
rect 394678 270703 394730 270755
rect 403126 270703 403178 270755
rect 626038 270629 626090 270681
rect 105046 270555 105098 270607
rect 139798 270555 139850 270607
rect 160150 270555 160202 270607
rect 101494 270481 101546 270533
rect 139894 270481 139946 270533
rect 98326 270407 98378 270459
rect 139990 270407 140042 270459
rect 94390 270333 94442 270385
rect 140182 270333 140234 270385
rect 89590 270259 89642 270311
rect 140086 270259 140138 270311
rect 176470 270555 176522 270607
rect 178486 270555 178538 270607
rect 180022 270555 180074 270607
rect 181366 270555 181418 270607
rect 172918 270481 172970 270533
rect 175606 270481 175658 270533
rect 174070 270407 174122 270459
rect 195862 270555 195914 270607
rect 206518 270555 206570 270607
rect 217462 270555 217514 270607
rect 187030 270481 187082 270533
rect 216790 270481 216842 270533
rect 216886 270481 216938 270533
rect 220534 270481 220586 270533
rect 182422 270407 182474 270459
rect 195862 270407 195914 270459
rect 196054 270407 196106 270459
rect 337078 270555 337130 270607
rect 357046 270555 357098 270607
rect 397366 270555 397418 270607
rect 397462 270555 397514 270607
rect 400342 270555 400394 270607
rect 403126 270555 403178 270607
rect 604630 270555 604682 270607
rect 228886 270481 228938 270533
rect 405910 270481 405962 270533
rect 407350 270481 407402 270533
rect 597526 270481 597578 270533
rect 236086 270407 236138 270459
rect 337078 270407 337130 270459
rect 357046 270407 357098 270459
rect 387190 270407 387242 270459
rect 387286 270407 387338 270459
rect 436918 270407 436970 270459
rect 459862 270407 459914 270459
rect 579670 270407 579722 270459
rect 168118 270333 168170 270385
rect 195862 270259 195914 270311
rect 195958 270259 196010 270311
rect 213238 270259 213290 270311
rect 213334 270259 213386 270311
rect 220342 270259 220394 270311
rect 405718 270333 405770 270385
rect 508246 270333 508298 270385
rect 601078 270333 601130 270385
rect 237622 270259 237674 270311
rect 337078 270259 337130 270311
rect 357046 270259 357098 270311
rect 380374 270259 380426 270311
rect 380470 270259 380522 270311
rect 402166 270259 402218 270311
rect 402358 270259 402410 270311
rect 554710 270259 554762 270311
rect 562198 270259 562250 270311
rect 646294 270259 646346 270311
rect 84790 270185 84842 270237
rect 140278 270185 140330 270237
rect 152662 270185 152714 270237
rect 394870 270185 394922 270237
rect 400246 270185 400298 270237
rect 568918 270185 568970 270237
rect 588886 270185 588938 270237
rect 632086 270185 632138 270237
rect 80182 270111 80234 270163
rect 140374 270111 140426 270163
rect 161014 270111 161066 270163
rect 403894 270111 403946 270163
rect 408982 270111 409034 270163
rect 422614 270111 422666 270163
rect 521782 270111 521834 270163
rect 622486 270111 622538 270163
rect 75382 270037 75434 270089
rect 139510 270037 139562 270089
rect 153814 270037 153866 270089
rect 68182 269963 68234 270015
rect 139318 269963 139370 270015
rect 142006 269963 142058 270015
rect 380182 269963 380234 270015
rect 135286 269889 135338 269941
rect 155542 269889 155594 269941
rect 166870 269889 166922 269941
rect 182422 269889 182474 269941
rect 182518 269889 182570 269941
rect 195862 269889 195914 269941
rect 195958 269889 196010 269941
rect 209686 269889 209738 269941
rect 209782 269889 209834 269941
rect 219862 269889 219914 269941
rect 219958 269889 220010 269941
rect 236086 269889 236138 269941
rect 237526 269889 237578 269941
rect 337078 269889 337130 269941
rect 337366 269889 337418 269941
rect 356758 269889 356810 269941
rect 357046 269889 357098 269941
rect 380086 269889 380138 269941
rect 127702 269815 127754 269867
rect 387094 269963 387146 270015
rect 387286 269963 387338 270015
rect 403030 269963 403082 270015
rect 403222 270037 403274 270089
rect 408406 270037 408458 270089
rect 405142 269963 405194 270015
rect 406102 269963 406154 270015
rect 411958 270037 412010 270089
rect 446230 270037 446282 270089
rect 576118 270037 576170 270089
rect 409078 269963 409130 270015
rect 583222 269963 583274 270015
rect 382294 269889 382346 269941
rect 408982 269889 409034 269941
rect 409174 269889 409226 269941
rect 593974 269889 594026 269941
rect 380566 269815 380618 269867
rect 388822 269815 388874 269867
rect 391702 269815 391754 269867
rect 590038 269815 590090 269867
rect 114646 269741 114698 269793
rect 383158 269741 383210 269793
rect 383254 269741 383306 269793
rect 407542 269741 407594 269793
rect 407638 269741 407690 269793
rect 608182 269741 608234 269793
rect 74134 269667 74186 269719
rect 367990 269667 368042 269719
rect 380086 269667 380138 269719
rect 382774 269667 382826 269719
rect 382870 269667 382922 269719
rect 633142 269667 633194 269719
rect 90838 269593 90890 269645
rect 388630 269593 388682 269645
rect 388918 269593 388970 269645
rect 611830 269593 611882 269645
rect 87190 269519 87242 269571
rect 81334 269445 81386 269497
rect 385654 269445 385706 269497
rect 386038 269519 386090 269571
rect 618934 269519 618986 269571
rect 388726 269445 388778 269497
rect 388822 269445 388874 269497
rect 394582 269445 394634 269497
rect 394678 269445 394730 269497
rect 629686 269445 629738 269497
rect 78934 269371 78986 269423
rect 382966 269371 383018 269423
rect 69334 269297 69386 269349
rect 376054 269297 376106 269349
rect 380182 269297 380234 269349
rect 383638 269371 383690 269423
rect 383734 269371 383786 269423
rect 383158 269297 383210 269349
rect 71734 269223 71786 269275
rect 385750 269223 385802 269275
rect 385942 269297 385994 269349
rect 407542 269371 407594 269423
rect 636502 269371 636554 269423
rect 391414 269223 391466 269275
rect 391798 269223 391850 269275
rect 394486 269223 394538 269275
rect 394582 269223 394634 269275
rect 640342 269297 640394 269349
rect 108694 269149 108746 269201
rect 139702 269149 139754 269201
rect 155542 269149 155594 269201
rect 182518 269149 182570 269201
rect 182710 269149 182762 269201
rect 405622 269149 405674 269201
rect 643894 269223 643946 269275
rect 112246 269075 112298 269127
rect 139606 269075 139658 269127
rect 181270 269075 181322 269127
rect 380470 269075 380522 269127
rect 382774 269075 382826 269127
rect 388534 269075 388586 269127
rect 388822 269075 388874 269127
rect 115798 269001 115850 269053
rect 139414 269001 139466 269053
rect 185974 269001 186026 269053
rect 405814 269075 405866 269127
rect 407638 269075 407690 269127
rect 472342 269149 472394 269201
rect 561814 269149 561866 269201
rect 570262 269149 570314 269201
rect 639094 269149 639146 269201
rect 452374 269075 452426 269127
rect 488086 269075 488138 269127
rect 572566 269075 572618 269127
rect 119350 268927 119402 268979
rect 140950 268927 141002 268979
rect 184726 268927 184778 268979
rect 387286 268927 387338 268979
rect 387382 268927 387434 268979
rect 400150 268927 400202 268979
rect 406678 268927 406730 268979
rect 502678 269001 502730 269053
rect 586774 269001 586826 269053
rect 448918 268927 448970 268979
rect 478774 268927 478826 268979
rect 558262 268927 558314 268979
rect 135382 268853 135434 268905
rect 259222 268853 259274 268905
rect 283798 268853 283850 268905
rect 133558 268779 133610 268831
rect 140566 268779 140618 268831
rect 175510 268779 175562 268831
rect 187030 268779 187082 268831
rect 195862 268779 195914 268831
rect 218806 268779 218858 268831
rect 219286 268779 219338 268831
rect 122902 268705 122954 268757
rect 140854 268705 140906 268757
rect 213238 268705 213290 268757
rect 219958 268705 220010 268757
rect 226390 268705 226442 268757
rect 324406 268705 324458 268757
rect 131254 268631 131306 268683
rect 135382 268631 135434 268683
rect 212182 268631 212234 268683
rect 313942 268631 313994 268683
rect 331990 268631 332042 268683
rect 337078 268853 337130 268905
rect 357046 268853 357098 268905
rect 371926 268853 371978 268905
rect 543670 268853 543722 268905
rect 550102 268853 550154 268905
rect 615382 268853 615434 268905
rect 349558 268779 349610 268831
rect 358102 268779 358154 268831
rect 371350 268779 371402 268831
rect 536854 268779 536906 268831
rect 337174 268705 337226 268757
rect 339862 268631 339914 268683
rect 350134 268705 350186 268757
rect 365590 268705 365642 268757
rect 370198 268705 370250 268757
rect 529750 268705 529802 268757
rect 356950 268631 357002 268683
rect 373174 268631 373226 268683
rect 522550 268631 522602 268683
rect 217462 268557 217514 268609
rect 219382 268557 219434 268609
rect 247702 268557 247754 268609
rect 252214 268557 252266 268609
rect 269206 268557 269258 268609
rect 331222 268557 331274 268609
rect 337270 268557 337322 268609
rect 356854 268557 356906 268609
rect 368470 268557 368522 268609
rect 515446 268557 515498 268609
rect 223606 268483 223658 268535
rect 238294 268483 238346 268535
rect 240694 268483 240746 268535
rect 267862 268483 267914 268535
rect 272758 268483 272810 268535
rect 334102 268483 334154 268535
rect 367606 268483 367658 268535
rect 508342 268483 508394 268535
rect 126550 268409 126602 268461
rect 140758 268409 140810 268461
rect 218806 268409 218858 268461
rect 237526 268409 237578 268461
rect 279958 268409 280010 268461
rect 334198 268409 334250 268461
rect 336982 268409 337034 268461
rect 346390 268409 346442 268461
rect 366934 268409 366986 268461
rect 501142 268409 501194 268461
rect 130102 268335 130154 268387
rect 140662 268335 140714 268387
rect 224182 268335 224234 268387
rect 245494 268335 245546 268387
rect 264502 268335 264554 268387
rect 282166 268335 282218 268387
rect 286102 268335 286154 268387
rect 296758 268335 296810 268387
rect 298582 268335 298634 268387
rect 338710 268335 338762 268387
rect 365878 268335 365930 268387
rect 494038 268335 494090 268387
rect 209686 268261 209738 268313
rect 237622 268261 237674 268313
rect 271606 268261 271658 268313
rect 282838 268261 282890 268313
rect 259222 268187 259274 268239
rect 279286 268187 279338 268239
rect 294262 268187 294314 268239
rect 339382 268261 339434 268313
rect 365206 268261 365258 268313
rect 486838 268261 486890 268313
rect 301270 268187 301322 268239
rect 339670 268187 339722 268239
rect 364342 268187 364394 268239
rect 479830 268187 479882 268239
rect 287062 268113 287114 268165
rect 298582 268113 298634 268165
rect 308470 268113 308522 268165
rect 343222 268113 343274 268165
rect 363190 268113 363242 268165
rect 472630 268113 472682 268165
rect 287638 268039 287690 268091
rect 307318 268039 307370 268091
rect 315670 268039 315722 268091
rect 341974 268039 342026 268091
rect 362614 268039 362666 268091
rect 465526 268039 465578 268091
rect 322774 267965 322826 268017
rect 344662 267965 344714 268017
rect 361462 267965 361514 268017
rect 458326 267965 458378 268017
rect 222550 267891 222602 267943
rect 231190 267891 231242 267943
rect 319126 267891 319178 267943
rect 341590 267891 341642 267943
rect 360598 267891 360650 267943
rect 450838 267891 450890 267943
rect 66838 267817 66890 267869
rect 137206 267817 137258 267869
rect 140470 267817 140522 267869
rect 147958 267817 148010 267869
rect 149686 267817 149738 267869
rect 151414 267817 151466 267869
rect 152566 267817 152618 267869
rect 158614 267817 158666 267869
rect 161206 267817 161258 267869
rect 162166 267817 162218 267869
rect 164086 267817 164138 267869
rect 165814 267817 165866 267869
rect 166966 267817 167018 267869
rect 191062 267817 191114 267869
rect 192886 267817 192938 267869
rect 222070 267817 222122 267869
rect 227638 267817 227690 267869
rect 258550 267817 258602 267869
rect 275926 267817 275978 267869
rect 278806 267817 278858 267869
rect 283894 267817 283946 267869
rect 285622 267817 285674 267869
rect 293014 267817 293066 267869
rect 324406 267817 324458 267869
rect 330166 267817 330218 267869
rect 344182 267817 344234 267869
rect 347542 267817 347594 267869
rect 359926 267817 359978 267869
rect 444118 267817 444170 267869
rect 72118 267743 72170 267795
rect 139126 267743 139178 267795
rect 140278 267743 140330 267795
rect 181462 267743 181514 267795
rect 191254 267743 191306 267795
rect 250486 267743 250538 267795
rect 250774 267669 250826 267721
rect 258838 267669 258890 267721
rect 259126 267743 259178 267795
rect 447094 267743 447146 267795
rect 455638 267817 455690 267869
rect 447190 267669 447242 267721
rect 455062 267743 455114 267795
rect 511894 267743 511946 267795
rect 463126 267669 463178 267721
rect 210934 267595 210986 267647
rect 275638 267595 275690 267647
rect 317494 267595 317546 267647
rect 321814 267595 321866 267647
rect 321910 267595 321962 267647
rect 524950 267595 525002 267647
rect 251254 267521 251306 267573
rect 251926 267447 251978 267499
rect 258838 267521 258890 267573
rect 447094 267521 447146 267573
rect 447190 267521 447242 267573
rect 459574 267521 459626 267573
rect 252406 267373 252458 267425
rect 466774 267447 466826 267499
rect 470230 267373 470282 267425
rect 473782 267299 473834 267351
rect 207382 267225 207434 267277
rect 258358 267225 258410 267277
rect 258550 267225 258602 267277
rect 275254 267225 275306 267277
rect 289846 267225 289898 267277
rect 325174 267225 325226 267277
rect 325462 267225 325514 267277
rect 549910 267225 549962 267277
rect 225334 267151 225386 267203
rect 247702 267151 247754 267203
rect 252982 267151 253034 267203
rect 215734 267077 215786 267129
rect 253654 267077 253706 267129
rect 253750 267077 253802 267129
rect 258262 267077 258314 267129
rect 191926 267003 191978 267055
rect 217654 267003 217706 267055
rect 222838 267003 222890 267055
rect 253366 267003 253418 267055
rect 254134 267003 254186 267055
rect 258646 267151 258698 267203
rect 477430 267151 477482 267203
rect 258454 267077 258506 267129
rect 484438 267077 484490 267129
rect 189526 266929 189578 266981
rect 223030 266929 223082 266981
rect 254518 266929 254570 266981
rect 480982 267003 481034 267055
rect 203830 266855 203882 266907
rect 252022 266855 252074 266907
rect 204982 266781 205034 266833
rect 256246 266781 256298 266833
rect 487798 266929 487850 266981
rect 256534 266855 256586 266907
rect 274774 266855 274826 266907
rect 276406 266855 276458 266907
rect 294166 266855 294218 266907
rect 318070 266855 318122 266907
rect 321718 266855 321770 266907
rect 321814 266855 321866 266907
rect 553462 266855 553514 266907
rect 491638 266781 491690 266833
rect 200182 266707 200234 266759
rect 274198 266707 274250 266759
rect 288310 266707 288362 266759
rect 314422 266707 314474 266759
rect 318646 266707 318698 266759
rect 321622 266707 321674 266759
rect 321718 266707 321770 266759
rect 557110 266707 557162 266759
rect 201430 266633 201482 266685
rect 253846 266633 253898 266685
rect 254710 266633 254762 266685
rect 495286 266633 495338 266685
rect 196726 266559 196778 266611
rect 273622 266559 273674 266611
rect 289366 266559 289418 266611
rect 321526 266559 321578 266611
rect 321622 266559 321674 266611
rect 560662 266559 560714 266611
rect 197878 266485 197930 266537
rect 255766 266485 255818 266537
rect 193078 266411 193130 266463
rect 250006 266411 250058 266463
rect 250102 266411 250154 266463
rect 138358 266337 138410 266389
rect 254422 266337 254474 266389
rect 255190 266411 255242 266463
rect 498838 266485 498890 266537
rect 548566 266485 548618 266537
rect 573142 266485 573194 266537
rect 266038 266411 266090 266463
rect 299542 266411 299594 266463
rect 259126 266337 259178 266389
rect 288694 266337 288746 266389
rect 317974 266411 318026 266463
rect 318742 266411 318794 266463
rect 564214 266411 564266 266463
rect 314230 266337 314282 266389
rect 319606 266337 319658 266389
rect 319702 266337 319754 266389
rect 571318 266337 571370 266389
rect 194326 266263 194378 266315
rect 329014 266263 329066 266315
rect 372886 266263 372938 266315
rect 551062 266263 551114 266315
rect 208534 266189 208586 266241
rect 250006 266189 250058 266241
rect 257494 266115 257546 266167
rect 257590 266115 257642 266167
rect 272662 266115 272714 266167
rect 272854 266189 272906 266241
rect 445270 266189 445322 266241
rect 273526 266115 273578 266167
rect 274102 266115 274154 266167
rect 441718 266115 441770 266167
rect 254902 266041 254954 266093
rect 256342 266041 256394 266093
rect 256438 266041 256490 266093
rect 394582 266041 394634 266093
rect 394774 266041 394826 266093
rect 394966 266041 395018 266093
rect 249334 265967 249386 266019
rect 388822 265967 388874 266019
rect 218038 265893 218090 265945
rect 276502 265893 276554 265945
rect 300694 265893 300746 265945
rect 414358 265893 414410 265945
rect 249718 265819 249770 265871
rect 256438 265819 256490 265871
rect 267862 265819 267914 265871
rect 334966 265819 335018 265871
rect 356086 265819 356138 265871
rect 406102 265819 406154 265871
rect 221494 265745 221546 265797
rect 276982 265745 277034 265797
rect 294070 265745 294122 265797
rect 360790 265745 360842 265797
rect 362134 265745 362186 265797
rect 397750 265745 397802 265797
rect 225238 265671 225290 265723
rect 277366 265671 277418 265723
rect 293686 265671 293738 265723
rect 357238 265671 357290 265723
rect 373462 265671 373514 265723
rect 402358 265671 402410 265723
rect 214582 265597 214634 265649
rect 275830 265597 275882 265649
rect 275926 265597 275978 265649
rect 337078 265597 337130 265649
rect 355606 265597 355658 265649
rect 403222 265597 403274 265649
rect 228790 265523 228842 265575
rect 232438 265449 232490 265501
rect 272662 265523 272714 265575
rect 279574 265523 279626 265575
rect 293110 265523 293162 265575
rect 353686 265523 353738 265575
rect 354934 265523 354986 265575
rect 404470 265523 404522 265575
rect 243094 265375 243146 265427
rect 257590 265375 257642 265427
rect 277846 265449 277898 265501
rect 292630 265449 292682 265501
rect 350038 265449 350090 265501
rect 367222 265449 367274 265501
rect 394102 265449 394154 265501
rect 278038 265375 278090 265427
rect 292150 265375 292202 265427
rect 346582 265375 346634 265427
rect 354550 265375 354602 265427
rect 401206 265375 401258 265427
rect 235894 265301 235946 265353
rect 278518 265301 278570 265353
rect 292054 265301 292106 265353
rect 342742 265301 342794 265353
rect 357142 265301 357194 265353
rect 382294 265301 382346 265353
rect 382390 265301 382442 265353
rect 391702 265301 391754 265353
rect 239446 265227 239498 265279
rect 279094 265227 279146 265279
rect 291574 265227 291626 265279
rect 339094 265227 339146 265279
rect 358870 265227 358922 265279
rect 374422 265227 374474 265279
rect 374998 265227 375050 265279
rect 400246 265227 400298 265279
rect 246646 265153 246698 265205
rect 280054 265153 280106 265205
rect 290422 265153 290474 265205
rect 318166 265153 318218 265205
rect 141142 265079 141194 265131
rect 151126 265079 151178 265131
rect 181462 265079 181514 265131
rect 191542 265079 191594 265131
rect 250198 265079 250250 265131
rect 280150 265079 280202 265131
rect 291190 265079 291242 265131
rect 335830 265153 335882 265205
rect 367126 265153 367178 265205
rect 390550 265153 390602 265205
rect 318358 265079 318410 265131
rect 332278 265079 332330 265131
rect 369622 265079 369674 265131
rect 373174 265079 373226 265131
rect 377878 265079 377930 265131
rect 380086 265079 380138 265131
rect 380470 265079 380522 265131
rect 388918 265079 388970 265131
rect 254038 265005 254090 265057
rect 280630 265005 280682 265057
rect 290038 265005 290090 265057
rect 328726 265005 328778 265057
rect 87766 264931 87818 264983
rect 106582 264931 106634 264983
rect 126742 264931 126794 264983
rect 141142 264931 141194 264983
rect 151126 264931 151178 264983
rect 168310 264931 168362 264983
rect 168406 264931 168458 264983
rect 66262 264783 66314 264835
rect 168406 264783 168458 264835
rect 168502 264783 168554 264835
rect 181462 264783 181514 264835
rect 202582 264931 202634 264983
rect 218902 264931 218954 264983
rect 253366 264931 253418 264983
rect 332758 264931 332810 264983
rect 333430 264931 333482 264983
rect 334102 264931 334154 264983
rect 338806 264931 338858 264983
rect 350902 265005 350954 265057
rect 346294 264931 346346 264983
rect 348406 264931 348458 264983
rect 351286 264931 351338 264983
rect 365686 265005 365738 265057
rect 379894 265005 379946 265057
rect 381142 265005 381194 265057
rect 386038 265005 386090 265057
rect 369142 264931 369194 264983
rect 372406 264931 372458 264983
rect 547606 264931 547658 264983
rect 191542 264857 191594 264909
rect 216694 264857 216746 264909
rect 223030 264857 223082 264909
rect 415318 264857 415370 264909
rect 216022 264783 216074 264835
rect 227638 264783 227690 264835
rect 249046 264783 249098 264835
rect 250390 264783 250442 264835
rect 438070 264783 438122 264835
rect 106582 264709 106634 264761
rect 126742 264709 126794 264761
rect 188374 264709 188426 264761
rect 414838 264709 414890 264761
rect 178870 264635 178922 264687
rect 412630 264635 412682 264687
rect 177622 264561 177674 264613
rect 412534 264561 412586 264613
rect 67318 264487 67370 264539
rect 87766 264487 87818 264539
rect 171670 264487 171722 264539
rect 410902 264487 410954 264539
rect 170518 264413 170570 264465
rect 410518 264413 410570 264465
rect 164566 264339 164618 264391
rect 409366 264339 409418 264391
rect 42262 264265 42314 264317
rect 53302 264265 53354 264317
rect 163414 264265 163466 264317
rect 408982 264265 409034 264317
rect 156214 264191 156266 264243
rect 407254 264191 407306 264243
rect 157462 264117 157514 264169
rect 407734 264117 407786 264169
rect 150262 264043 150314 264095
rect 406006 264043 406058 264095
rect 149110 263969 149162 264021
rect 405526 263969 405578 264021
rect 405718 263969 405770 264021
rect 410326 263969 410378 264021
rect 145558 263895 145610 263947
rect 404374 263895 404426 263947
rect 405910 263895 405962 263947
rect 412054 263895 412106 263947
rect 146998 263821 147050 263873
rect 405046 263821 405098 263873
rect 405142 263821 405194 263873
rect 406582 263821 406634 263873
rect 132502 263747 132554 263799
rect 401590 263747 401642 263799
rect 403030 263747 403082 263799
rect 414262 263747 414314 263799
rect 107446 263673 107498 263725
rect 395254 263673 395306 263725
rect 395350 263673 395402 263725
rect 396502 263673 396554 263725
rect 398614 263673 398666 263725
rect 403990 263673 404042 263725
rect 405622 263673 405674 263725
rect 413782 263673 413834 263725
rect 91990 263599 92042 263651
rect 391510 263599 391562 263651
rect 394966 263599 395018 263651
rect 408118 263599 408170 263651
rect 42262 263525 42314 263577
rect 53398 263525 53450 263577
rect 76534 263525 76586 263577
rect 387190 263525 387242 263577
rect 388726 263525 388778 263577
rect 390262 263525 390314 263577
rect 390358 263525 390410 263577
rect 394294 263525 394346 263577
rect 394870 263525 394922 263577
rect 406102 263525 406154 263577
rect 195478 263451 195530 263503
rect 218134 263451 218186 263503
rect 223798 263451 223850 263503
rect 241846 263451 241898 263503
rect 256342 263451 256394 263503
rect 336598 263451 336650 263503
rect 353398 263451 353450 263503
rect 367126 263451 367178 263503
rect 371446 263451 371498 263503
rect 540406 263451 540458 263503
rect 191254 263377 191306 263429
rect 198742 263377 198794 263429
rect 224662 263377 224714 263429
rect 227638 263377 227690 263429
rect 253654 263377 253706 263429
rect 331606 263377 331658 263429
rect 334198 263377 334250 263429
rect 339766 263377 339818 263429
rect 353878 263377 353930 263429
rect 367222 263377 367274 263429
rect 370678 263377 370730 263429
rect 533206 263377 533258 263429
rect 199126 263303 199178 263355
rect 218326 263303 218378 263355
rect 255766 263303 255818 263355
rect 329686 263303 329738 263355
rect 331222 263303 331274 263355
rect 338134 263303 338186 263355
rect 340630 263303 340682 263355
rect 346870 263303 346922 263355
rect 349078 263303 349130 263355
rect 354838 263303 354890 263355
rect 355030 263303 355082 263355
rect 365686 263303 365738 263355
rect 369718 263303 369770 263355
rect 526198 263303 526250 263355
rect 252502 263229 252554 263281
rect 258646 263229 258698 263281
rect 286582 263229 286634 263281
rect 300118 263229 300170 263281
rect 327766 263229 327818 263281
rect 335542 263229 335594 263281
rect 357814 263229 357866 263281
rect 364630 263229 364682 263281
rect 369142 263229 369194 263281
rect 518998 263229 519050 263281
rect 254422 263155 254474 263207
rect 402838 263155 402890 263207
rect 406678 263155 406730 263207
rect 414646 263155 414698 263207
rect 253846 263081 253898 263133
rect 330070 263081 330122 263133
rect 330166 263081 330218 263133
rect 332950 263081 333002 263133
rect 339670 263081 339722 263133
rect 342070 263081 342122 263133
rect 349750 263081 349802 263133
rect 362038 263081 362090 263133
rect 367414 263081 367466 263133
rect 504694 263081 504746 263133
rect 223126 263007 223178 263059
rect 234742 263007 234794 263059
rect 257494 263007 257546 263059
rect 330742 263007 330794 263059
rect 331030 263007 331082 263059
rect 334486 263007 334538 263059
rect 338710 263007 338762 263059
rect 340342 263007 340394 263059
rect 354070 263007 354122 263059
rect 362134 263007 362186 263059
rect 366550 263007 366602 263059
rect 497302 263007 497354 263059
rect 261238 262933 261290 262985
rect 326806 262933 326858 262985
rect 326998 262933 327050 262985
rect 345334 262933 345386 262985
rect 351862 262933 351914 262985
rect 355030 262933 355082 262985
rect 365398 262933 365450 262985
rect 490486 262933 490538 262985
rect 248182 262859 248234 262911
rect 274102 262859 274154 262911
rect 285526 262859 285578 262911
rect 289462 262859 289514 262911
rect 290998 262859 291050 262911
rect 341014 262859 341066 262911
rect 352342 262859 352394 262911
rect 362806 262859 362858 262911
rect 364822 262859 364874 262911
rect 483286 262859 483338 262911
rect 248662 262785 248714 262837
rect 272854 262785 272906 262837
rect 294166 262785 294218 262837
rect 339286 262785 339338 262837
rect 339382 262785 339434 262837
rect 341494 262785 341546 262837
rect 341590 262785 341642 262837
rect 344278 262785 344330 262837
rect 363670 262785 363722 262837
rect 476182 262785 476234 262837
rect 257686 262711 257738 262763
rect 281302 262711 281354 262763
rect 282358 262711 282410 262763
rect 284374 262711 284426 262763
rect 297814 262711 297866 262763
rect 341878 262711 341930 262763
rect 341974 262711 342026 262763
rect 344086 262711 344138 262763
rect 362710 262711 362762 262763
rect 468982 262711 469034 262763
rect 42262 262637 42314 262689
rect 47830 262637 47882 262689
rect 260950 262637 261002 262689
rect 275158 262637 275210 262689
rect 283510 262637 283562 262689
rect 287254 262637 287306 262689
rect 303670 262637 303722 262689
rect 304918 262637 304970 262689
rect 342742 262637 342794 262689
rect 362134 262637 362186 262689
rect 461974 262637 462026 262689
rect 268342 262563 268394 262615
rect 282358 262563 282410 262615
rect 285046 262563 285098 262615
rect 285814 262563 285866 262615
rect 299542 262563 299594 262615
rect 337750 262563 337802 262615
rect 361078 262563 361130 262615
rect 454774 262563 454826 262615
rect 287830 262489 287882 262541
rect 310870 262489 310922 262541
rect 312406 262489 312458 262541
rect 343606 262489 343658 262541
rect 367990 262489 368042 262541
rect 455062 262489 455114 262541
rect 281782 262415 281834 262467
rect 313942 262415 313994 262467
rect 331222 262415 331274 262467
rect 360406 262415 360458 262467
rect 447670 262415 447722 262467
rect 317014 262341 317066 262393
rect 325462 262341 325514 262393
rect 327094 262341 327146 262393
rect 399190 262341 399242 262393
rect 400150 262341 400202 262393
rect 409846 262341 409898 262393
rect 351766 262267 351818 262319
rect 375958 262267 376010 262319
rect 376054 262267 376106 262319
rect 384982 262267 385034 262319
rect 385654 262267 385706 262319
rect 388246 262267 388298 262319
rect 388630 262267 388682 262319
rect 390934 262267 390986 262319
rect 391414 262267 391466 262319
rect 396982 262267 397034 262319
rect 397078 262267 397130 262319
rect 401782 262267 401834 262319
rect 402166 262267 402218 262319
rect 413110 262267 413162 262319
rect 144694 262119 144746 262171
rect 146614 262119 146666 262171
rect 221590 262119 221642 262171
rect 223990 262119 224042 262171
rect 247990 262119 248042 262171
rect 250390 262119 250442 262171
rect 256246 262119 256298 262171
rect 330550 262119 330602 262171
rect 251350 262045 251402 262097
rect 336022 262193 336074 262245
rect 359350 262193 359402 262245
rect 244246 261971 244298 262023
rect 335350 262119 335402 262171
rect 352822 262119 352874 262171
rect 357046 262045 357098 262097
rect 362806 262119 362858 262171
rect 384406 262193 384458 262245
rect 385846 262193 385898 262245
rect 386134 262193 386186 262245
rect 390454 262193 390506 262245
rect 390646 262193 390698 262245
rect 396310 262193 396362 262245
rect 382966 262119 383018 262171
rect 388054 262119 388106 262171
rect 389014 262119 389066 262171
rect 394198 262119 394250 262171
rect 394294 262119 394346 262171
rect 400150 262193 400202 262245
rect 400342 262193 400394 262245
rect 411574 262193 411626 262245
rect 396502 262119 396554 262171
rect 403798 262119 403850 262171
rect 403894 262119 403946 262171
rect 408310 262119 408362 262171
rect 440470 262045 440522 262097
rect 382582 261971 382634 262023
rect 382678 261971 382730 262023
rect 394678 261971 394730 262023
rect 262102 261897 262154 261949
rect 263350 261897 263402 261949
rect 324022 261897 324074 261949
rect 346966 261897 347018 261949
rect 362806 261897 362858 261949
rect 419062 261897 419114 261949
rect 243670 261823 243722 261875
rect 402454 261823 402506 261875
rect 244246 261749 244298 261801
rect 409558 261749 409610 261801
rect 245398 261675 245450 261727
rect 416662 261675 416714 261727
rect 245974 261601 246026 261653
rect 423862 261601 423914 261653
rect 246934 261527 246986 261579
rect 431062 261527 431114 261579
rect 521302 261527 521354 261579
rect 548566 261527 548618 261579
rect 239926 261453 239978 261505
rect 373558 261453 373610 261505
rect 374614 261453 374666 261505
rect 565462 261453 565514 261505
rect 320758 261379 320810 261431
rect 578518 261379 578570 261431
rect 229654 261305 229706 261357
rect 288214 261305 288266 261357
rect 321430 261305 321482 261357
rect 585622 261305 585674 261357
rect 230326 261231 230378 261283
rect 295414 261231 295466 261283
rect 231190 261157 231242 261209
rect 302518 261231 302570 261283
rect 308182 261231 308234 261283
rect 318358 261231 318410 261283
rect 322486 261231 322538 261283
rect 592726 261231 592778 261283
rect 298006 261157 298058 261209
rect 316726 261157 316778 261209
rect 323158 261157 323210 261209
rect 599830 261157 599882 261209
rect 232342 261083 232394 261135
rect 309718 261083 309770 261135
rect 318070 261083 318122 261135
rect 338230 261083 338282 261135
rect 346966 261083 347018 261135
rect 607030 261083 607082 261135
rect 225814 261009 225866 261061
rect 255862 261009 255914 261061
rect 260662 261009 260714 261061
rect 541654 261009 541706 261061
rect 225910 260935 225962 260987
rect 259702 260935 259754 260987
rect 261718 260935 261770 260987
rect 552310 260935 552362 260987
rect 232918 260861 232970 260913
rect 298006 260861 298058 260913
rect 305686 260861 305738 260913
rect 318262 260861 318314 260913
rect 325174 260861 325226 260913
rect 614230 260861 614282 260913
rect 234070 260787 234122 260839
rect 323926 260787 323978 260839
rect 325750 260787 325802 260839
rect 620950 260787 621002 260839
rect 226390 260713 226442 260765
rect 262102 260713 262154 260765
rect 262198 260713 262250 260765
rect 555862 260713 555914 260765
rect 234934 260639 234986 260691
rect 318166 260639 318218 260691
rect 318358 260639 318410 260691
rect 328246 260639 328298 260691
rect 328342 260639 328394 260691
rect 642742 260639 642794 260691
rect 240982 260565 241034 260617
rect 381046 260565 381098 260617
rect 381526 260565 381578 260617
rect 521782 260565 521834 260617
rect 239350 260491 239402 260543
rect 366742 260491 366794 260543
rect 378934 260491 378986 260543
rect 508246 260491 508298 260543
rect 228598 260417 228650 260469
rect 280822 260417 280874 260469
rect 301846 260417 301898 260469
rect 425014 260417 425066 260469
rect 238198 260343 238250 260395
rect 359638 260343 359690 260395
rect 373942 260343 373994 260395
rect 478774 260343 478826 260395
rect 226870 260269 226922 260321
rect 266806 260269 266858 260321
rect 301174 260269 301226 260321
rect 417910 260269 417962 260321
rect 237334 260195 237386 260247
rect 352438 260195 352490 260247
rect 376150 260195 376202 260247
rect 446230 260195 446282 260247
rect 236662 260121 236714 260173
rect 345046 260121 345098 260173
rect 376726 260121 376778 260173
rect 409078 260121 409130 260173
rect 299638 260047 299690 260099
rect 407158 260047 407210 260099
rect 235606 259973 235658 260025
rect 318070 259973 318122 260025
rect 318166 259973 318218 260025
rect 331126 259973 331178 260025
rect 378262 259973 378314 260025
rect 409174 259973 409226 260025
rect 233494 259899 233546 259951
rect 72022 259529 72074 259581
rect 77686 259529 77738 259581
rect 298966 259899 299018 259951
rect 400054 259899 400106 259951
rect 308086 259825 308138 259877
rect 308182 259825 308234 259877
rect 328246 259825 328298 259877
rect 334006 259825 334058 259877
rect 379990 259825 380042 259877
rect 405814 259825 405866 259877
rect 298102 259751 298154 259803
rect 392950 259751 393002 259803
rect 394678 259751 394730 259803
rect 395062 259751 395114 259803
rect 296950 259677 297002 259729
rect 385558 259677 385610 259729
rect 296374 259603 296426 259655
rect 378646 259603 378698 259655
rect 295318 259529 295370 259581
rect 371542 259529 371594 259581
rect 294358 259455 294410 259507
rect 364438 259455 364490 259507
rect 308086 259381 308138 259433
rect 318262 259381 318314 259433
rect 457174 259381 457226 259433
rect 242518 259307 242570 259359
rect 395158 259307 395210 259359
rect 241654 259233 241706 259285
rect 388150 259233 388202 259285
rect 146518 259159 146570 259211
rect 146614 259159 146666 259211
rect 639286 256347 639338 256399
rect 679798 256347 679850 256399
rect 675094 253461 675146 253513
rect 678262 253461 678314 253513
rect 72118 253387 72170 253439
rect 77014 253387 77066 253439
rect 674806 251611 674858 251663
rect 676918 251611 676970 251663
rect 674998 251537 675050 251589
rect 676822 251537 676874 251589
rect 673942 250945 673994 250997
rect 675382 250945 675434 250997
rect 198742 250575 198794 250627
rect 207286 250501 207338 250553
rect 674614 250353 674666 250405
rect 675478 250353 675530 250405
rect 674326 247023 674378 247075
rect 675478 247023 675530 247075
rect 139510 246949 139562 247001
rect 141430 246949 141482 247001
rect 674422 246949 674474 247001
rect 675286 246949 675338 247001
rect 257014 246801 257066 246853
rect 327958 246801 328010 246853
rect 262006 246727 262058 246779
rect 331846 246727 331898 246779
rect 252886 246653 252938 246705
rect 328774 246653 328826 246705
rect 258262 246579 258314 246631
rect 332758 246579 332810 246631
rect 65110 246505 65162 246557
rect 204982 246505 205034 246557
rect 257590 246505 257642 246557
rect 334486 246505 334538 246557
rect 47926 246431 47978 246483
rect 204886 246431 204938 246483
rect 256438 246431 256490 246483
rect 336598 246431 336650 246483
rect 48022 246357 48074 246409
rect 204502 246357 204554 246409
rect 255958 246357 256010 246409
rect 338134 246357 338186 246409
rect 47446 246283 47498 246335
rect 207190 246283 207242 246335
rect 255094 246283 255146 246335
rect 339862 246283 339914 246335
rect 44662 246209 44714 246261
rect 204790 246209 204842 246261
rect 254230 246209 254282 246261
rect 341494 246209 341546 246261
rect 277558 246135 277610 246187
rect 364342 246135 364394 246187
rect 139414 246061 139466 246113
rect 141526 246061 141578 246113
rect 276406 246061 276458 246113
rect 362806 246061 362858 246113
rect 674710 246061 674762 246113
rect 675382 246061 675434 246113
rect 253750 245987 253802 246039
rect 343222 245987 343274 246039
rect 273238 245913 273290 245965
rect 360598 245913 360650 245965
rect 251542 245839 251594 245891
rect 348022 245839 348074 245891
rect 139318 245765 139370 245817
rect 143158 245765 143210 245817
rect 252022 245765 252074 245817
rect 346294 245765 346346 245817
rect 250486 245691 250538 245743
rect 349078 245691 349130 245743
rect 249814 245617 249866 245669
rect 350806 245617 350858 245669
rect 248566 245543 248618 245595
rect 354070 245543 354122 245595
rect 249334 245469 249386 245521
rect 352822 245469 352874 245521
rect 263062 245395 263114 245447
rect 372886 245395 372938 245447
rect 80662 245321 80714 245373
rect 100726 245321 100778 245373
rect 247606 245321 247658 245373
rect 355606 245321 355658 245373
rect 262678 245247 262730 245299
rect 373462 245247 373514 245299
rect 246838 245173 246890 245225
rect 357334 245173 357386 245225
rect 246358 245099 246410 245151
rect 358870 245099 358922 245151
rect 158422 245025 158474 245077
rect 168502 245025 168554 245077
rect 261430 245025 261482 245077
rect 376726 245025 376778 245077
rect 260470 244951 260522 245003
rect 378454 244951 378506 245003
rect 420502 244951 420554 245003
rect 440566 244951 440618 245003
rect 204502 244877 204554 244929
rect 205174 244877 205226 244929
rect 214102 244877 214154 244929
rect 259894 244877 259946 244929
rect 379510 244877 379562 244929
rect 42358 244803 42410 244855
rect 214486 244803 214538 244855
rect 259606 244803 259658 244855
rect 380662 244803 380714 244855
rect 268726 244729 268778 244781
rect 318262 244729 318314 244781
rect 217558 244655 217610 244707
rect 257974 244655 258026 244707
rect 267574 244655 267626 244707
rect 218422 244285 218474 244337
rect 256342 244581 256394 244633
rect 236470 244507 236522 244559
rect 268246 244507 268298 244559
rect 278134 244655 278186 244707
rect 318070 244655 318122 244707
rect 278038 244581 278090 244633
rect 336406 244581 336458 244633
rect 270454 244507 270506 244559
rect 318166 244507 318218 244559
rect 325462 244507 325514 244559
rect 326806 244507 326858 244559
rect 338710 244433 338762 244485
rect 261046 244359 261098 244411
rect 335926 244359 335978 244411
rect 398518 244433 398570 244485
rect 250198 244285 250250 244337
rect 258838 244285 258890 244337
rect 277942 244285 277994 244337
rect 337366 244285 337418 244337
rect 210166 244063 210218 244115
rect 287638 244211 287690 244263
rect 294934 244211 294986 244263
rect 306934 244211 306986 244263
rect 307030 244211 307082 244263
rect 325366 244211 325418 244263
rect 325462 244211 325514 244263
rect 348502 244211 348554 244263
rect 352822 244211 352874 244263
rect 254710 244137 254762 244189
rect 356374 244137 356426 244189
rect 251254 244063 251306 244115
rect 355030 244063 355082 244115
rect 77878 243989 77930 244041
rect 149590 243989 149642 244041
rect 219478 243989 219530 244041
rect 254038 243989 254090 244041
rect 256246 243989 256298 244041
rect 357238 243989 357290 244041
rect 77014 243915 77066 243967
rect 152470 243915 152522 243967
rect 248182 243915 248234 243967
rect 353590 243915 353642 243967
rect 44950 243841 45002 243893
rect 204694 243841 204746 243893
rect 220726 243841 220778 243893
rect 250774 243841 250826 243893
rect 252982 243841 253034 243893
rect 355798 243841 355850 243893
rect 45046 243767 45098 243819
rect 204598 243767 204650 243819
rect 40246 243693 40298 243745
rect 41782 243693 41834 243745
rect 45238 243693 45290 243745
rect 206518 243693 206570 243745
rect 246934 243693 246986 243745
rect 348502 243767 348554 243819
rect 360790 243767 360842 243819
rect 397462 243767 397514 243819
rect 44566 243619 44618 243671
rect 204502 243619 204554 243671
rect 41974 243545 42026 243597
rect 42550 243545 42602 243597
rect 47734 243545 47786 243597
rect 212374 243545 212426 243597
rect 245878 243545 245930 243597
rect 351862 243693 351914 243745
rect 360214 243693 360266 243745
rect 395926 243693 395978 243745
rect 254326 243619 254378 243671
rect 258838 243619 258890 243671
rect 354358 243619 354410 243671
rect 362038 243619 362090 243671
rect 401782 243619 401834 243671
rect 350422 243545 350474 243597
rect 362422 243545 362474 243597
rect 402838 243545 402890 243597
rect 45142 243471 45194 243523
rect 212758 243471 212810 243523
rect 240982 243471 241034 243523
rect 349654 243471 349706 243523
rect 363862 243471 363914 243523
rect 405526 243471 405578 243523
rect 44758 243397 44810 243449
rect 211894 243397 211946 243449
rect 239350 243397 239402 243449
rect 349174 243397 349226 243449
rect 361942 243397 361994 243449
rect 401110 243397 401162 243449
rect 44854 243323 44906 243375
rect 212278 243323 212330 243375
rect 242134 243323 242186 243375
rect 254326 243323 254378 243375
rect 243862 243249 243914 243301
rect 351478 243323 351530 243375
rect 364630 243323 364682 243375
rect 407254 243323 407306 243375
rect 264790 243249 264842 243301
rect 313270 243249 313322 243301
rect 316534 243249 316586 243301
rect 381142 243249 381194 243301
rect 265750 243175 265802 243227
rect 311638 243175 311690 243227
rect 315574 243175 315626 243227
rect 348502 243175 348554 243227
rect 368566 243175 368618 243227
rect 378934 243175 378986 243227
rect 266614 243101 266666 243153
rect 310486 243101 310538 243153
rect 326614 243101 326666 243153
rect 374998 243101 375050 243153
rect 268054 243027 268106 243079
rect 294934 243027 294986 243079
rect 268822 242953 268874 243005
rect 305686 243027 305738 243079
rect 295126 242953 295178 243005
rect 302230 242953 302282 243005
rect 265846 242879 265898 242931
rect 278134 242879 278186 242931
rect 282070 242879 282122 242931
rect 312982 243027 313034 243079
rect 326422 243027 326474 243079
rect 326710 243027 326762 243079
rect 377206 243027 377258 243079
rect 326326 242953 326378 243005
rect 326518 242953 326570 243005
rect 372982 242953 373034 243005
rect 262774 242805 262826 242857
rect 278038 242805 278090 242857
rect 283414 242805 283466 242857
rect 263926 242731 263978 242783
rect 277942 242731 277994 242783
rect 293590 242731 293642 242783
rect 296662 242731 296714 242783
rect 270262 242657 270314 242709
rect 295126 242657 295178 242709
rect 298102 242805 298154 242857
rect 316726 242805 316778 242857
rect 298198 242731 298250 242783
rect 325750 242879 325802 242931
rect 330646 242879 330698 242931
rect 361078 242879 361130 242931
rect 317206 242805 317258 242857
rect 323542 242805 323594 242857
rect 331030 242805 331082 242857
rect 362134 242805 362186 242857
rect 318262 242731 318314 242783
rect 339574 242731 339626 242783
rect 348502 242731 348554 242783
rect 368566 242731 368618 242783
rect 674902 242731 674954 242783
rect 675382 242731 675434 242783
rect 324022 242657 324074 242709
rect 330262 242657 330314 242709
rect 360022 242657 360074 242709
rect 282934 242583 282986 242635
rect 275254 242509 275306 242561
rect 309430 242509 309482 242561
rect 316726 242583 316778 242635
rect 317206 242583 317258 242635
rect 318070 242583 318122 242635
rect 337846 242583 337898 242635
rect 324694 242509 324746 242561
rect 330742 242509 330794 242561
rect 361654 242509 361706 242561
rect 139126 242435 139178 242487
rect 140278 242435 140330 242487
rect 269878 242435 269930 242487
rect 302998 242435 303050 242487
rect 293206 242361 293258 242413
rect 140374 242287 140426 242339
rect 141334 242287 141386 242339
rect 268918 242287 268970 242339
rect 304630 242287 304682 242339
rect 326230 242435 326282 242487
rect 318166 242361 318218 242413
rect 340342 242361 340394 242413
rect 674998 242361 675050 242413
rect 675382 242361 675434 242413
rect 313462 242287 313514 242339
rect 326614 242287 326666 242339
rect 283798 242213 283850 242265
rect 298102 242213 298154 242265
rect 314806 242213 314858 242265
rect 326710 242213 326762 242265
rect 37270 242139 37322 242191
rect 42742 242139 42794 242191
rect 40054 242065 40106 242117
rect 42358 242065 42410 242117
rect 37366 241991 37418 242043
rect 43126 241991 43178 242043
rect 140758 241991 140810 242043
rect 141142 241991 141194 242043
rect 40150 241917 40202 241969
rect 43030 241917 43082 241969
rect 44662 241917 44714 241969
rect 206422 241917 206474 241969
rect 206518 241917 206570 241969
rect 207094 241917 207146 241969
rect 213142 241917 213194 241969
rect 244630 241917 244682 241969
rect 43222 241843 43274 241895
rect 43702 241843 43754 241895
rect 140758 241843 140810 241895
rect 152470 241843 152522 241895
rect 41686 241769 41738 241821
rect 43510 241769 43562 241821
rect 140662 241769 140714 241821
rect 221398 241843 221450 241895
rect 234550 241843 234602 241895
rect 240214 241843 240266 241895
rect 259510 241843 259562 241895
rect 271894 241843 271946 241895
rect 286774 241991 286826 242043
rect 293014 242139 293066 242191
rect 325270 242139 325322 242191
rect 287734 242065 287786 242117
rect 298198 242065 298250 242117
rect 320470 242065 320522 242117
rect 339478 242065 339530 242117
rect 292726 241991 292778 242043
rect 324214 241991 324266 242043
rect 286102 241843 286154 241895
rect 289846 241843 289898 241895
rect 289942 241843 289994 241895
rect 295798 241843 295850 241895
rect 296662 241917 296714 241969
rect 307030 241917 307082 241969
rect 330550 241843 330602 241895
rect 331318 241843 331370 241895
rect 338518 241917 338570 241969
rect 383542 241917 383594 241969
rect 338230 241843 338282 241895
rect 352918 241843 352970 241895
rect 368278 241843 368330 241895
rect 223126 241769 223178 241821
rect 233974 241769 234026 241821
rect 239734 241769 239786 241821
rect 216694 241695 216746 241747
rect 228886 241695 228938 241747
rect 241078 241695 241130 241747
rect 245398 241769 245450 241821
rect 273238 241769 273290 241821
rect 275446 241769 275498 241821
rect 291094 241769 291146 241821
rect 291286 241769 291338 241821
rect 298390 241769 298442 241821
rect 328918 241769 328970 241821
rect 338134 241769 338186 241821
rect 338902 241769 338954 241821
rect 353398 241769 353450 241821
rect 261238 241695 261290 241747
rect 271030 241695 271082 241747
rect 286486 241695 286538 241747
rect 289750 241695 289802 241747
rect 296278 241695 296330 241747
rect 318262 241695 318314 241747
rect 334966 241695 335018 241747
rect 337078 241695 337130 241747
rect 345814 241695 345866 241747
rect 226870 241621 226922 241673
rect 232150 241621 232202 241673
rect 227542 241547 227594 241599
rect 244246 241621 244298 241673
rect 281302 241621 281354 241673
rect 289942 241621 289994 241673
rect 290134 241621 290186 241673
rect 236662 241547 236714 241599
rect 248662 241547 248714 241599
rect 271990 241547 272042 241599
rect 288118 241547 288170 241599
rect 228502 241473 228554 241525
rect 238390 241473 238442 241525
rect 238774 241473 238826 241525
rect 225910 241399 225962 241451
rect 232342 241399 232394 241451
rect 225334 241325 225386 241377
rect 232630 241325 232682 241377
rect 217270 241251 217322 241303
rect 229174 241251 229226 241303
rect 236566 241399 236618 241451
rect 237238 241399 237290 241451
rect 247126 241399 247178 241451
rect 235318 241325 235370 241377
rect 245974 241325 246026 241377
rect 247318 241473 247370 241525
rect 262198 241473 262250 241525
rect 264406 241473 264458 241525
rect 275638 241473 275690 241525
rect 283318 241473 283370 241525
rect 289750 241473 289802 241525
rect 290710 241473 290762 241525
rect 297622 241473 297674 241525
rect 273718 241399 273770 241451
rect 286102 241399 286154 241451
rect 286678 241399 286730 241451
rect 296950 241399 297002 241451
rect 262870 241325 262922 241377
rect 271126 241325 271178 241377
rect 286390 241325 286442 241377
rect 220342 241103 220394 241155
rect 236278 241251 236330 241303
rect 244918 241251 244970 241303
rect 272566 241251 272618 241303
rect 286294 241251 286346 241303
rect 239350 241177 239402 241229
rect 247318 241177 247370 241229
rect 273526 241177 273578 241229
rect 286198 241177 286250 241229
rect 289462 241325 289514 241377
rect 289750 241325 289802 241377
rect 300022 241325 300074 241377
rect 286774 241251 286826 241303
rect 298294 241251 298346 241303
rect 229942 241103 229994 241155
rect 240406 241103 240458 241155
rect 240502 241103 240554 241155
rect 264310 241103 264362 241155
rect 275926 241103 275978 241155
rect 287062 241177 287114 241229
rect 291286 241177 291338 241229
rect 291382 241177 291434 241229
rect 226486 241029 226538 241081
rect 239446 241029 239498 241081
rect 247414 241029 247466 241081
rect 267766 241029 267818 241081
rect 277366 241029 277418 241081
rect 286006 241029 286058 241081
rect 286102 241029 286154 241081
rect 294358 241103 294410 241155
rect 294454 241103 294506 241155
rect 297718 241103 297770 241155
rect 286486 241029 286538 241081
rect 300790 241029 300842 241081
rect 223318 240955 223370 241007
rect 235318 240955 235370 241007
rect 42742 240881 42794 240933
rect 43318 240881 43370 240933
rect 224566 240881 224618 240933
rect 243190 240955 243242 241007
rect 243286 240955 243338 241007
rect 264982 240955 265034 241007
rect 272854 240955 272906 241007
rect 285430 240955 285482 241007
rect 285526 240955 285578 241007
rect 290710 240955 290762 241007
rect 290806 240955 290858 241007
rect 298486 240955 298538 241007
rect 223894 240807 223946 240859
rect 236278 240807 236330 240859
rect 222550 240733 222602 240785
rect 237238 240733 237290 240785
rect 221686 240659 221738 240711
rect 249238 240881 249290 240933
rect 271510 240881 271562 240933
rect 281686 240881 281738 240933
rect 283894 240881 283946 240933
rect 296662 240881 296714 240933
rect 318838 241621 318890 241673
rect 335542 241621 335594 241673
rect 338134 241621 338186 241673
rect 354550 241695 354602 241747
rect 334582 241547 334634 241599
rect 348118 241547 348170 241599
rect 348214 241547 348266 241599
rect 358390 241547 358442 241599
rect 378550 241843 378602 241895
rect 385654 241843 385706 241895
rect 387286 241843 387338 241895
rect 372694 241769 372746 241821
rect 386134 241769 386186 241821
rect 377878 241695 377930 241747
rect 387190 241695 387242 241747
rect 387286 241695 387338 241747
rect 397846 241695 397898 241747
rect 373078 241621 373130 241673
rect 384790 241621 384842 241673
rect 384886 241621 384938 241673
rect 398998 241621 399050 241673
rect 389782 241547 389834 241599
rect 674134 241547 674186 241599
rect 675478 241547 675530 241599
rect 317878 241473 317930 241525
rect 333814 241473 333866 241525
rect 338038 241473 338090 241525
rect 355126 241473 355178 241525
rect 370486 241473 370538 241525
rect 384982 241473 385034 241525
rect 385654 241473 385706 241525
rect 388246 241473 388298 241525
rect 328534 241399 328586 241451
rect 357142 241399 357194 241451
rect 329878 241325 329930 241377
rect 359350 241325 359402 241377
rect 362806 241325 362858 241377
rect 385942 241399 385994 241451
rect 386134 241399 386186 241451
rect 399574 241399 399626 241451
rect 372214 241325 372266 241377
rect 383542 241325 383594 241377
rect 383638 241325 383690 241377
rect 389398 241325 389450 241377
rect 301174 241251 301226 241303
rect 316630 241251 316682 241303
rect 327574 241251 327626 241303
rect 338134 241251 338186 241303
rect 338518 241251 338570 241303
rect 346390 241251 346442 241303
rect 381430 241251 381482 241303
rect 392566 241251 392618 241303
rect 328054 241177 328106 241229
rect 338038 241177 338090 241229
rect 338614 241177 338666 241229
rect 344278 241177 344330 241229
rect 301078 241103 301130 241155
rect 315478 241103 315530 241155
rect 332086 241103 332138 241155
rect 302518 241029 302570 241081
rect 315958 241029 316010 241081
rect 317782 241029 317834 241081
rect 332950 241029 333002 241081
rect 319222 240955 319274 241007
rect 332470 240955 332522 241007
rect 333718 240955 333770 241007
rect 322006 240881 322058 240933
rect 335062 240881 335114 240933
rect 41782 240585 41834 240637
rect 221110 240585 221162 240637
rect 250390 240807 250442 240859
rect 276886 240807 276938 240859
rect 237622 240733 237674 240785
rect 266038 240733 266090 240785
rect 238966 240659 239018 240711
rect 266710 240659 266762 240711
rect 225526 240511 225578 240563
rect 228886 240511 228938 240563
rect 228982 240511 229034 240563
rect 237430 240511 237482 240563
rect 226102 240437 226154 240489
rect 229942 240437 229994 240489
rect 230038 240437 230090 240489
rect 237334 240437 237386 240489
rect 41782 240363 41834 240415
rect 224278 240363 224330 240415
rect 227542 240363 227594 240415
rect 222070 240215 222122 240267
rect 234358 240289 234410 240341
rect 228310 240215 228362 240267
rect 235606 240215 235658 240267
rect 226870 240141 226922 240193
rect 228502 240141 228554 240193
rect 228694 240141 228746 240193
rect 234454 240141 234506 240193
rect 227926 240067 227978 240119
rect 231766 240067 231818 240119
rect 226966 239993 227018 240045
rect 228982 239993 229034 240045
rect 229078 239993 229130 240045
rect 230806 239993 230858 240045
rect 218134 239919 218186 239971
rect 225142 239919 225194 239971
rect 227350 239919 227402 239971
rect 230038 239919 230090 239971
rect 230134 239919 230186 239971
rect 230518 239919 230570 239971
rect 229558 239845 229610 239897
rect 232246 239845 232298 239897
rect 229078 239771 229130 239823
rect 233590 239771 233642 239823
rect 220246 239697 220298 239749
rect 252502 240585 252554 240637
rect 276406 240733 276458 240785
rect 278518 240733 278570 240785
rect 285910 240733 285962 240785
rect 280054 240659 280106 240711
rect 285814 240659 285866 240711
rect 287350 240807 287402 240859
rect 315286 240807 315338 240859
rect 324502 240807 324554 240859
rect 334582 240807 334634 240859
rect 334678 240807 334730 240859
rect 287830 240733 287882 240785
rect 290806 240733 290858 240785
rect 290998 240733 291050 240785
rect 321430 240733 321482 240785
rect 288310 240659 288362 240711
rect 289558 240659 289610 240711
rect 237910 240511 237962 240563
rect 243286 240511 243338 240563
rect 244534 240511 244586 240563
rect 273238 240585 273290 240637
rect 284662 240585 284714 240637
rect 286390 240585 286442 240637
rect 299830 240585 299882 240637
rect 273334 240511 273386 240563
rect 281590 240511 281642 240563
rect 281686 240511 281738 240563
rect 285718 240511 285770 240563
rect 289270 240511 289322 240563
rect 295318 240511 295370 240563
rect 300022 240659 300074 240711
rect 318358 240659 318410 240711
rect 315670 240585 315722 240637
rect 327862 240733 327914 240785
rect 328246 240733 328298 240785
rect 338134 240733 338186 240785
rect 326710 240659 326762 240711
rect 338230 240659 338282 240711
rect 323638 240585 323690 240637
rect 337078 240585 337130 240637
rect 338998 241029 339050 241081
rect 363190 241177 363242 241229
rect 373462 241177 373514 241229
rect 384694 241177 384746 241229
rect 384790 241177 384842 241229
rect 400726 241177 400778 241229
rect 374902 241103 374954 241155
rect 403990 241103 404042 241155
rect 359830 241029 359882 241081
rect 384502 241029 384554 241081
rect 363958 240955 364010 241007
rect 375670 240955 375722 241007
rect 406006 241029 406058 241081
rect 384694 240955 384746 241007
rect 401590 240955 401642 241007
rect 364726 240881 364778 240933
rect 374038 240881 374090 240933
rect 402262 240881 402314 240933
rect 367990 240807 368042 240859
rect 384118 240807 384170 240859
rect 414262 240807 414314 240859
rect 370678 240733 370730 240785
rect 375286 240733 375338 240785
rect 405046 240733 405098 240785
rect 338614 240659 338666 240711
rect 366934 240659 366986 240711
rect 372598 240659 372650 240711
rect 384214 240659 384266 240711
rect 384310 240659 384362 240711
rect 414646 240659 414698 240711
rect 369718 240585 369770 240637
rect 376630 240585 376682 240637
rect 407734 240585 407786 240637
rect 317494 240511 317546 240563
rect 319222 240511 319274 240563
rect 327766 240511 327818 240563
rect 327862 240511 327914 240563
rect 332278 240511 332330 240563
rect 332854 240511 332906 240563
rect 365878 240511 365930 240563
rect 374326 240511 374378 240563
rect 403318 240511 403370 240563
rect 674806 240511 674858 240563
rect 675478 240511 675530 240563
rect 238006 240437 238058 240489
rect 240502 240437 240554 240489
rect 276790 240437 276842 240489
rect 280342 240437 280394 240489
rect 280438 240437 280490 240489
rect 295414 240437 295466 240489
rect 324118 240437 324170 240489
rect 334198 240437 334250 240489
rect 334294 240437 334346 240489
rect 368758 240437 368810 240489
rect 376246 240437 376298 240489
rect 406582 240437 406634 240489
rect 549046 240437 549098 240489
rect 650902 240437 650954 240489
rect 279094 240363 279146 240415
rect 294454 240363 294506 240415
rect 321430 240363 321482 240415
rect 327670 240363 327722 240415
rect 327766 240363 327818 240415
rect 336022 240363 336074 240415
rect 338134 240363 338186 240415
rect 356278 240363 356330 240415
rect 370006 240363 370058 240415
rect 386614 240363 386666 240415
rect 275542 240289 275594 240341
rect 240118 240215 240170 240267
rect 260182 240215 260234 240267
rect 277750 240215 277802 240267
rect 285622 240215 285674 240267
rect 278518 240141 278570 240193
rect 284374 240141 284426 240193
rect 279094 240067 279146 240119
rect 283510 240067 283562 240119
rect 272470 239993 272522 240045
rect 273622 239993 273674 240045
rect 278998 239993 279050 240045
rect 280822 239993 280874 240045
rect 273046 239919 273098 239971
rect 276310 239919 276362 239971
rect 279862 239919 279914 239971
rect 280630 239919 280682 239971
rect 268438 239845 268490 239897
rect 274774 239845 274826 239897
rect 279286 239845 279338 239897
rect 282358 239845 282410 239897
rect 286198 240289 286250 240341
rect 288502 240289 288554 240341
rect 288598 240289 288650 240341
rect 294070 240289 294122 240341
rect 302326 240289 302378 240341
rect 326230 240289 326282 240341
rect 302518 240215 302570 240267
rect 324886 240215 324938 240267
rect 329014 240215 329066 240267
rect 329206 240215 329258 240267
rect 329782 240215 329834 240267
rect 333334 240215 333386 240267
rect 338614 240215 338666 240267
rect 342742 240289 342794 240341
rect 343126 240289 343178 240341
rect 381526 240289 381578 240341
rect 393718 240289 393770 240341
rect 342838 240215 342890 240267
rect 381910 240215 381962 240267
rect 394582 240215 394634 240267
rect 285910 240141 285962 240193
rect 288598 240141 288650 240193
rect 288694 240141 288746 240193
rect 298870 240141 298922 240193
rect 298966 240141 299018 240193
rect 302422 240141 302474 240193
rect 325846 240141 325898 240193
rect 286006 240067 286058 240119
rect 286294 239993 286346 240045
rect 291862 239993 291914 240045
rect 292054 240067 292106 240119
rect 300598 240067 300650 240119
rect 300694 240067 300746 240119
rect 304630 240067 304682 240119
rect 324022 240067 324074 240119
rect 331318 240067 331370 240119
rect 293974 239993 294026 240045
rect 295894 239993 295946 240045
rect 302518 239993 302570 240045
rect 303574 239993 303626 240045
rect 305878 239993 305930 240045
rect 310870 239993 310922 240045
rect 313942 239993 313994 240045
rect 323254 239993 323306 240045
rect 338230 240067 338282 240119
rect 338518 240141 338570 240193
rect 366838 240141 366890 240193
rect 377878 240141 377930 240193
rect 380086 240141 380138 240193
rect 390262 240141 390314 240193
rect 331510 239993 331562 240045
rect 338998 239993 339050 240045
rect 344662 240067 344714 240119
rect 368182 240067 368234 240119
rect 378550 240067 378602 240119
rect 378838 240067 378890 240119
rect 387670 240067 387722 240119
rect 388726 240067 388778 240119
rect 396310 240067 396362 240119
rect 342742 239993 342794 240045
rect 382870 239993 382922 240045
rect 386518 239993 386570 240045
rect 386614 239993 386666 240045
rect 393046 239993 393098 240045
rect 285814 239919 285866 239971
rect 294934 239919 294986 239971
rect 296566 239919 296618 239971
rect 302806 239919 302858 239971
rect 302902 239919 302954 239971
rect 305494 239919 305546 239971
rect 309334 239919 309386 239971
rect 309814 239919 309866 239971
rect 310006 239919 310058 239971
rect 311158 239919 311210 239971
rect 311638 239919 311690 239971
rect 327478 239919 327530 239971
rect 290422 239845 290474 239897
rect 290518 239845 290570 239897
rect 292246 239845 292298 239897
rect 292630 239845 292682 239897
rect 300694 239845 300746 239897
rect 301366 239845 301418 239897
rect 305014 239845 305066 239897
rect 321910 239845 321962 239897
rect 330934 239919 330986 239971
rect 331126 239919 331178 239971
rect 332950 239919 333002 239971
rect 334198 239919 334250 239971
rect 347542 239919 347594 239971
rect 382294 239919 382346 239971
rect 385462 239919 385514 239971
rect 327670 239845 327722 239897
rect 341014 239845 341066 239897
rect 382966 239845 383018 239897
rect 388054 239845 388106 239897
rect 279862 239771 279914 239823
rect 281494 239771 281546 239823
rect 281590 239771 281642 239823
rect 289270 239771 289322 239823
rect 289366 239771 289418 239823
rect 299254 239771 299306 239823
rect 299638 239771 299690 239823
rect 304246 239771 304298 239823
rect 311254 239771 311306 239823
rect 314902 239771 314954 239823
rect 322294 239771 322346 239823
rect 329110 239771 329162 239823
rect 329302 239771 329354 239823
rect 348214 239771 348266 239823
rect 371254 239771 371306 239823
rect 388726 239771 388778 239823
rect 222070 239623 222122 239675
rect 236662 239623 236714 239675
rect 236758 239623 236810 239675
rect 247414 239623 247466 239675
rect 224758 239549 224810 239601
rect 242518 239549 242570 239601
rect 243766 239549 243818 239601
rect 277558 239697 277610 239749
rect 278134 239697 278186 239749
rect 284566 239697 284618 239749
rect 284662 239697 284714 239749
rect 290806 239697 290858 239749
rect 290902 239697 290954 239749
rect 300214 239697 300266 239749
rect 321814 239697 321866 239749
rect 276214 239623 276266 239675
rect 285238 239623 285290 239675
rect 277270 239549 277322 239601
rect 287158 239549 287210 239601
rect 223798 239475 223850 239527
rect 233590 239475 233642 239527
rect 246454 239475 246506 239527
rect 276982 239475 277034 239527
rect 281590 239475 281642 239527
rect 282166 239475 282218 239527
rect 296182 239623 296234 239675
rect 297430 239623 297482 239675
rect 302902 239623 302954 239675
rect 305206 239623 305258 239675
rect 306646 239623 306698 239675
rect 310774 239623 310826 239675
rect 313174 239623 313226 239675
rect 321046 239623 321098 239675
rect 328342 239623 328394 239675
rect 330934 239697 330986 239749
rect 343126 239697 343178 239749
rect 374806 239697 374858 239749
rect 386038 239697 386090 239749
rect 341878 239623 341930 239675
rect 370870 239623 370922 239675
rect 383062 239623 383114 239675
rect 288694 239549 288746 239601
rect 222934 239253 222986 239305
rect 280438 239401 280490 239453
rect 291670 239475 291722 239527
rect 291958 239549 292010 239601
rect 297046 239549 297098 239601
rect 301078 239549 301130 239601
rect 320086 239549 320138 239601
rect 338806 239549 338858 239601
rect 380662 239549 380714 239601
rect 390934 239549 390986 239601
rect 637558 239549 637610 239601
rect 650134 239549 650186 239601
rect 298006 239475 298058 239527
rect 303286 239475 303338 239527
rect 310390 239475 310442 239527
rect 312214 239475 312266 239527
rect 369622 239475 369674 239527
rect 392470 239475 392522 239527
rect 638038 239475 638090 239527
rect 650422 239475 650474 239527
rect 288790 239401 288842 239453
rect 290518 239401 290570 239453
rect 290806 239401 290858 239453
rect 295990 239401 296042 239453
rect 325366 239401 325418 239453
rect 245014 239327 245066 239379
rect 273526 239327 273578 239379
rect 274102 239327 274154 239379
rect 285430 239327 285482 239379
rect 290038 239327 290090 239379
rect 299830 239327 299882 239379
rect 304438 239327 304490 239379
rect 306454 239327 306506 239379
rect 326326 239327 326378 239379
rect 368662 239401 368714 239453
rect 390454 239401 390506 239453
rect 637654 239401 637706 239453
rect 650230 239401 650282 239453
rect 229942 239253 229994 239305
rect 231382 239253 231434 239305
rect 275062 239253 275114 239305
rect 292150 239253 292202 239305
rect 292246 239253 292298 239305
rect 301174 239253 301226 239305
rect 319606 239253 319658 239305
rect 336982 239253 337034 239305
rect 349750 239327 349802 239379
rect 369046 239327 369098 239379
rect 391510 239327 391562 239379
rect 494518 239327 494570 239379
rect 497206 239327 497258 239379
rect 638806 239327 638858 239379
rect 649558 239327 649610 239379
rect 352342 239253 352394 239305
rect 370390 239253 370442 239305
rect 394198 239253 394250 239305
rect 639382 239253 639434 239305
rect 649750 239253 649802 239305
rect 140566 239179 140618 239231
rect 216598 239179 216650 239231
rect 233206 239179 233258 239231
rect 277846 239179 277898 239231
rect 281206 239179 281258 239231
rect 282550 239179 282602 239231
rect 287734 239179 287786 239231
rect 288022 239179 288074 239231
rect 293110 239179 293162 239231
rect 294166 239179 294218 239231
rect 301462 239179 301514 239231
rect 322678 239179 322730 239231
rect 328918 239179 328970 239231
rect 329110 239179 329162 239231
rect 343606 239179 343658 239231
rect 371830 239179 371882 239231
rect 396982 239179 397034 239231
rect 505558 239179 505610 239231
rect 674614 239179 674666 239231
rect 675094 239179 675146 239231
rect 228598 239105 228650 239157
rect 231382 239105 231434 239157
rect 237142 239105 237194 239157
rect 238966 239105 239018 239157
rect 274678 239105 274730 239157
rect 287926 239105 287978 239157
rect 288502 239105 288554 239157
rect 301078 239105 301130 239157
rect 319702 239105 319754 239157
rect 337750 239105 337802 239157
rect 381046 239105 381098 239157
rect 391990 239105 392042 239157
rect 510358 239105 510410 239157
rect 674998 239105 675050 239157
rect 144022 239031 144074 239083
rect 174166 239031 174218 239083
rect 208726 239031 208778 239083
rect 215638 239031 215690 239083
rect 222166 239031 222218 239083
rect 227734 239031 227786 239083
rect 236182 239031 236234 239083
rect 236566 239031 236618 239083
rect 238390 239031 238442 239083
rect 277654 239031 277706 239083
rect 286582 239031 286634 239083
rect 294838 239031 294890 239083
rect 302038 239031 302090 239083
rect 327094 239031 327146 239083
rect 338902 239031 338954 239083
rect 379702 239031 379754 239083
rect 388822 239031 388874 239083
rect 420598 239031 420650 239083
rect 421846 239031 421898 239083
rect 541462 239031 541514 239083
rect 549046 239031 549098 239083
rect 639766 239031 639818 239083
rect 649942 239031 649994 239083
rect 140566 238957 140618 239009
rect 264502 238957 264554 239009
rect 314422 238957 314474 239009
rect 325462 238957 325514 239009
rect 396790 238957 396842 239009
rect 140470 238883 140522 238935
rect 141142 238883 141194 238935
rect 235318 238883 235370 238935
rect 270838 238883 270890 238935
rect 271318 238883 271370 238935
rect 340438 238883 340490 238935
rect 384022 238883 384074 238935
rect 384598 238883 384650 238935
rect 266518 238809 266570 238861
rect 338230 238809 338282 238861
rect 235798 238735 235850 238787
rect 269110 238735 269162 238787
rect 256918 238661 256970 238713
rect 277846 238735 277898 238787
rect 278710 238735 278762 238787
rect 339958 238735 340010 238787
rect 276502 238661 276554 238713
rect 336982 238661 337034 238713
rect 247990 238587 248042 238639
rect 42166 238513 42218 238565
rect 42550 238513 42602 238565
rect 217270 238513 217322 238565
rect 259030 238513 259082 238565
rect 261718 238587 261770 238639
rect 336022 238587 336074 238639
rect 264214 238513 264266 238565
rect 264886 238513 264938 238565
rect 337750 238513 337802 238565
rect 237046 238439 237098 238491
rect 257686 238439 257738 238491
rect 259990 238439 260042 238491
rect 335542 238439 335594 238491
rect 219862 238365 219914 238417
rect 253462 238365 253514 238417
rect 255190 238365 255242 238417
rect 356662 238365 356714 238417
rect 218038 238291 218090 238343
rect 257302 238291 257354 238343
rect 263446 238291 263498 238343
rect 276502 238291 276554 238343
rect 277846 238291 277898 238343
rect 357622 238291 357674 238343
rect 218518 238217 218570 238269
rect 255670 238217 255722 238269
rect 220342 238143 220394 238195
rect 251446 238143 251498 238195
rect 253942 238143 253994 238195
rect 355894 238217 355946 238269
rect 252406 238069 252458 238121
rect 355414 238143 355466 238195
rect 264214 238069 264266 238121
rect 353206 238069 353258 238121
rect 249046 237995 249098 238047
rect 353686 237995 353738 238047
rect 42166 237847 42218 237899
rect 50422 237847 50474 237899
rect 243094 237847 243146 237899
rect 350998 237921 351050 237973
rect 257686 237847 257738 237899
rect 347830 237847 347882 237899
rect 361174 237847 361226 237899
rect 399190 237847 399242 237899
rect 241654 237773 241706 237825
rect 350038 237773 350090 237825
rect 361558 237773 361610 237825
rect 400246 237773 400298 237825
rect 244726 237699 244778 237751
rect 351478 237699 351530 237751
rect 363766 237699 363818 237751
rect 404374 237699 404426 237751
rect 140374 237625 140426 237677
rect 140662 237625 140714 237677
rect 239926 237625 239978 237677
rect 349270 237625 349322 237677
rect 363382 237625 363434 237677
rect 403798 237625 403850 237677
rect 233398 237551 233450 237603
rect 346582 237551 346634 237603
rect 364246 237551 364298 237603
rect 406102 237551 406154 237603
rect 277846 237477 277898 237529
rect 312694 237477 312746 237529
rect 316054 237477 316106 237529
rect 380182 237477 380234 237529
rect 266710 237403 266762 237455
rect 309526 237403 309578 237455
rect 316822 237403 316874 237455
rect 381718 237403 381770 237455
rect 140854 237329 140906 237381
rect 141238 237329 141290 237381
rect 266230 237329 266282 237381
rect 310966 237329 311018 237381
rect 315190 237329 315242 237381
rect 377782 237329 377834 237381
rect 267094 237255 267146 237307
rect 308758 237255 308810 237307
rect 313846 237255 313898 237307
rect 375190 237255 375242 237307
rect 140854 237181 140906 237233
rect 141334 237181 141386 237233
rect 267478 237181 267530 237233
rect 307894 237181 307946 237233
rect 317398 237181 317450 237233
rect 382582 237181 382634 237233
rect 269302 237107 269354 237159
rect 303958 237107 304010 237159
rect 313078 237107 313130 237159
rect 374134 237107 374186 237159
rect 269686 237033 269738 237085
rect 278710 237033 278762 237085
rect 286966 237033 287018 237085
rect 302134 237033 302186 237085
rect 314422 237033 314474 237085
rect 376054 237033 376106 237085
rect 235702 236959 235754 237011
rect 269782 236959 269834 237011
rect 274582 236959 274634 237011
rect 305398 236959 305450 237011
rect 312598 236959 312650 237011
rect 372406 236959 372458 237011
rect 265270 236885 265322 236937
rect 277846 236885 277898 236937
rect 270646 236811 270698 236863
rect 301846 236885 301898 236937
rect 302422 236885 302474 236937
rect 303670 236885 303722 236937
rect 312214 236885 312266 236937
rect 371350 236885 371402 236937
rect 284278 236811 284330 236863
rect 322582 236811 322634 236863
rect 284758 236737 284810 236789
rect 320950 236737 321002 236789
rect 42166 236663 42218 236715
rect 43126 236663 43178 236715
rect 284374 236663 284426 236715
rect 321526 236663 321578 236715
rect 285142 236589 285194 236641
rect 319990 236589 320042 236641
rect 286102 236515 286154 236567
rect 318742 236515 318794 236567
rect 43222 236441 43274 236493
rect 43414 236441 43466 236493
rect 291766 236441 291818 236493
rect 323158 236441 323210 236493
rect 43318 236367 43370 236419
rect 43702 236367 43754 236419
rect 286582 236367 286634 236419
rect 317014 236367 317066 236419
rect 290518 236293 290570 236345
rect 319894 236293 319946 236345
rect 144022 236219 144074 236271
rect 165526 236219 165578 236271
rect 286486 236219 286538 236271
rect 317686 236219 317738 236271
rect 144118 236145 144170 236197
rect 168406 236145 168458 236197
rect 290806 236145 290858 236197
rect 320278 236145 320330 236197
rect 273526 236071 273578 236123
rect 361462 236071 361514 236123
rect 257878 235775 257930 235827
rect 333430 235775 333482 235827
rect 257398 235701 257450 235753
rect 335350 235701 335402 235753
rect 248950 235627 249002 235679
rect 329686 235627 329738 235679
rect 256054 235553 256106 235605
rect 337558 235553 337610 235605
rect 255574 235479 255626 235531
rect 339286 235479 339338 235531
rect 42166 235405 42218 235457
rect 43030 235405 43082 235457
rect 254806 235405 254858 235457
rect 340534 235405 340586 235457
rect 253846 235331 253898 235383
rect 342070 235331 342122 235383
rect 253366 235257 253418 235309
rect 344086 235257 344138 235309
rect 675094 235257 675146 235309
rect 679798 235257 679850 235309
rect 252598 235183 252650 235235
rect 345334 235183 345386 235235
rect 674998 235183 675050 235235
rect 679990 235183 680042 235235
rect 251638 235109 251690 235161
rect 346870 235109 346922 235161
rect 257782 235035 257834 235087
rect 358006 235035 358058 235087
rect 251158 234961 251210 235013
rect 348598 234961 348650 235013
rect 258934 234887 258986 234939
rect 358102 234887 358154 234939
rect 42166 234813 42218 234865
rect 42454 234813 42506 234865
rect 250390 234813 250442 234865
rect 350134 234813 350186 234865
rect 210070 234739 210122 234791
rect 383254 234739 383306 234791
rect 42454 234665 42506 234717
rect 43126 234665 43178 234717
rect 249430 234665 249482 234717
rect 351670 234665 351722 234717
rect 264022 234591 264074 234643
rect 370966 234591 371018 234643
rect 248182 234517 248234 234569
rect 354934 234517 354986 234569
rect 263638 234443 263690 234495
rect 371926 234443 371978 234495
rect 247222 234369 247274 234421
rect 356470 234369 356522 234421
rect 246742 234295 246794 234347
rect 357814 234295 357866 234347
rect 245974 234221 246026 234273
rect 359542 234221 359594 234273
rect 42070 234147 42122 234199
rect 42358 234147 42410 234199
rect 262294 234147 262346 234199
rect 374614 234147 374666 234199
rect 261814 234073 261866 234125
rect 375766 234073 375818 234125
rect 260086 233999 260138 234051
rect 379414 233999 379466 234051
rect 260854 233925 260906 233977
rect 377398 233925 377450 233977
rect 243910 233851 243962 233903
rect 363670 233851 363722 233903
rect 258982 233777 259034 233829
rect 381238 233777 381290 233829
rect 207190 233703 207242 233755
rect 213526 233703 213578 233755
rect 220150 233703 220202 233755
rect 258838 233703 258890 233755
rect 382390 233703 382442 233755
rect 210166 233629 210218 233681
rect 212374 233629 212426 233681
rect 358486 233629 358538 233681
rect 210262 233555 210314 233607
rect 212758 233555 212810 233607
rect 216502 233555 216554 233607
rect 414838 233555 414890 233607
rect 144022 233259 144074 233311
rect 171286 233259 171338 233311
rect 204982 233185 205034 233237
rect 206806 233185 206858 233237
rect 645526 233185 645578 233237
rect 649654 233185 649706 233237
rect 204502 233111 204554 233163
rect 206902 233111 206954 233163
rect 645718 233111 645770 233163
rect 649846 233111 649898 233163
rect 204694 233037 204746 233089
rect 206710 233037 206762 233089
rect 645334 233037 645386 233089
rect 650038 233037 650090 233089
rect 645142 232963 645194 233015
rect 650326 232963 650378 233015
rect 645238 232889 645290 232941
rect 650518 232889 650570 232941
rect 204598 232741 204650 232793
rect 206614 232741 206666 232793
rect 144022 230521 144074 230573
rect 151126 230521 151178 230573
rect 144118 230447 144170 230499
rect 162646 230447 162698 230499
rect 141526 230373 141578 230425
rect 201814 230373 201866 230425
rect 139990 230299 140042 230351
rect 141430 230299 141482 230351
rect 201622 230299 201674 230351
rect 172726 230151 172778 230203
rect 178582 230225 178634 230277
rect 178678 230151 178730 230203
rect 201718 230151 201770 230203
rect 139990 230077 140042 230129
rect 141334 230077 141386 230129
rect 143158 230077 143210 230129
rect 146902 230077 146954 230129
rect 166870 230003 166922 230055
rect 172726 230003 172778 230055
rect 139990 229929 140042 229981
rect 661174 229485 661226 229537
rect 674422 229485 674474 229537
rect 669622 228893 669674 228945
rect 674710 228893 674762 228945
rect 141334 227857 141386 227909
rect 669526 227857 669578 227909
rect 674422 227857 674474 227909
rect 140470 227783 140522 227835
rect 140566 227783 140618 227835
rect 140662 227783 140714 227835
rect 140758 227783 140810 227835
rect 144022 227709 144074 227761
rect 188566 227709 188618 227761
rect 144214 227635 144266 227687
rect 194326 227635 194378 227687
rect 139894 227561 139946 227613
rect 140470 227561 140522 227613
rect 140566 227561 140618 227613
rect 140662 227561 140714 227613
rect 140758 227561 140810 227613
rect 144118 227561 144170 227613
rect 197206 227561 197258 227613
rect 141238 227487 141290 227539
rect 201814 227487 201866 227539
rect 140566 227413 140618 227465
rect 197590 227413 197642 227465
rect 140950 227339 141002 227391
rect 201718 227339 201770 227391
rect 140758 227265 140810 227317
rect 201526 227265 201578 227317
rect 140470 227191 140522 227243
rect 201622 227191 201674 227243
rect 144022 225637 144074 225689
rect 156886 225637 156938 225689
rect 144022 224675 144074 224727
rect 179926 224675 179978 224727
rect 140854 224601 140906 224653
rect 201526 224601 201578 224653
rect 140662 224527 140714 224579
rect 201718 224527 201770 224579
rect 141046 224453 141098 224505
rect 201622 224453 201674 224505
rect 146806 224379 146858 224431
rect 201718 224379 201770 224431
rect 149686 224305 149738 224357
rect 201814 224305 201866 224357
rect 152566 224231 152618 224283
rect 209974 224231 210026 224283
rect 209782 223195 209834 223247
rect 210166 223195 210218 223247
rect 144022 221863 144074 221915
rect 177046 221863 177098 221915
rect 144118 221789 144170 221841
rect 202966 221789 203018 221841
rect 146422 221715 146474 221767
rect 146710 221715 146762 221767
rect 155446 221715 155498 221767
rect 198646 221715 198698 221767
rect 161206 221641 161258 221693
rect 201718 221641 201770 221693
rect 164086 221567 164138 221619
rect 209974 221567 210026 221619
rect 166966 221493 167018 221545
rect 201622 221493 201674 221545
rect 169846 221419 169898 221471
rect 201814 221419 201866 221471
rect 42358 221049 42410 221101
rect 45430 221049 45482 221101
rect 42358 220309 42410 220361
rect 45526 220309 45578 220361
rect 42358 219421 42410 219473
rect 45334 219421 45386 219473
rect 144022 218903 144074 218955
rect 174262 218903 174314 218955
rect 140278 218829 140330 218881
rect 197590 218829 197642 218881
rect 175606 218755 175658 218807
rect 209974 218755 210026 218807
rect 178486 218681 178538 218733
rect 201718 218681 201770 218733
rect 181366 218607 181418 218659
rect 198166 218607 198218 218659
rect 184246 218533 184298 218585
rect 210166 218533 210218 218585
rect 144022 216683 144074 216735
rect 154006 216683 154058 216735
rect 140086 215943 140138 215995
rect 201622 215943 201674 215995
rect 139990 215869 140042 215921
rect 210166 215869 210218 215921
rect 140086 215795 140138 215847
rect 201814 215795 201866 215847
rect 140182 215721 140234 215773
rect 201238 215721 201290 215773
rect 187126 215647 187178 215699
rect 201718 215647 201770 215699
rect 192886 215573 192938 215625
rect 209974 215573 210026 215625
rect 144022 213205 144074 213257
rect 168502 213205 168554 213257
rect 144118 213131 144170 213183
rect 171382 213131 171434 213183
rect 140086 213057 140138 213109
rect 201622 213057 201674 213109
rect 139990 212983 140042 213035
rect 140278 212983 140330 213035
rect 201718 212983 201770 213035
rect 209974 212909 210026 212961
rect 144022 210245 144074 210297
rect 148246 210245 148298 210297
rect 645622 210245 645674 210297
rect 646102 210245 646154 210297
rect 679702 210245 679754 210297
rect 674614 210171 674666 210223
rect 676822 210171 676874 210223
rect 209782 208469 209834 208521
rect 210262 208469 210314 208521
rect 144022 207433 144074 207485
rect 162742 207433 162794 207485
rect 144118 207359 144170 207411
rect 165622 207359 165674 207411
rect 146422 207285 146474 207337
rect 146710 207285 146762 207337
rect 674422 205731 674474 205783
rect 675478 205731 675530 205783
rect 675190 205139 675242 205191
rect 675478 205139 675530 205191
rect 675094 204843 675146 204895
rect 674998 204621 675050 204673
rect 42166 204325 42218 204377
rect 44662 204325 44714 204377
rect 146806 201661 146858 201713
rect 185686 201661 185738 201713
rect 144214 201587 144266 201639
rect 200086 201587 200138 201639
rect 40150 201513 40202 201565
rect 42166 201513 42218 201565
rect 674326 201291 674378 201343
rect 675382 201291 675434 201343
rect 37270 200181 37322 200233
rect 43126 200181 43178 200233
rect 146806 198923 146858 198975
rect 159766 198923 159818 198975
rect 37366 198849 37418 198901
rect 43222 198849 43274 198901
rect 40246 198775 40298 198827
rect 43030 198775 43082 198827
rect 146710 198701 146762 198753
rect 191446 198701 191498 198753
rect 674806 197591 674858 197643
rect 675382 197591 675434 197643
rect 42070 197443 42122 197495
rect 42454 197443 42506 197495
rect 41878 197369 41930 197421
rect 41974 197369 42026 197421
rect 42358 197221 42410 197273
rect 41878 197147 41930 197199
rect 674614 196999 674666 197051
rect 675478 196999 675530 197051
rect 674710 196555 674762 196607
rect 675382 196555 675434 196607
rect 146806 195815 146858 195867
rect 182806 195815 182858 195867
rect 42646 195741 42698 195793
rect 43222 195741 43274 195793
rect 42166 195297 42218 195349
rect 42358 195297 42410 195349
rect 42070 194483 42122 194535
rect 47638 194483 47690 194535
rect 42070 193447 42122 193499
rect 43126 193447 43178 193499
rect 146806 193003 146858 193055
rect 148342 193003 148394 193055
rect 42166 192189 42218 192241
rect 43030 192189 43082 192241
rect 42070 191449 42122 191501
rect 42358 191449 42410 191501
rect 42358 191301 42410 191353
rect 42646 191301 42698 191353
rect 146710 190191 146762 190243
rect 148438 190191 148490 190243
rect 146806 190117 146858 190169
rect 200182 190117 200234 190169
rect 42166 187823 42218 187875
rect 42742 187823 42794 187875
rect 146710 187305 146762 187357
rect 148534 187305 148586 187357
rect 146806 187231 146858 187283
rect 194422 187231 194474 187283
rect 42166 187083 42218 187135
rect 42454 187083 42506 187135
rect 42070 186491 42122 186543
rect 42646 186491 42698 186543
rect 144022 184345 144074 184397
rect 151222 184345 151274 184397
rect 655318 184345 655370 184397
rect 674422 184345 674474 184397
rect 660982 183901 661034 183953
rect 674710 183901 674762 183953
rect 666742 182865 666794 182917
rect 674422 182865 674474 182917
rect 144022 181459 144074 181511
rect 185782 181459 185834 181511
rect 144118 178647 144170 178699
rect 148630 178647 148682 178699
rect 144022 178573 144074 178625
rect 191542 178573 191594 178625
rect 144022 175687 144074 175739
rect 188662 175687 188714 175739
rect 144022 172801 144074 172853
rect 182902 172801 182954 172853
rect 144022 170359 144074 170411
rect 159862 170359 159914 170411
rect 209974 169915 210026 169967
rect 210166 169915 210218 169967
rect 209878 169841 209930 169893
rect 209782 169767 209834 169819
rect 209974 169767 210026 169819
rect 209878 169693 209930 169745
rect 647926 167177 647978 167229
rect 674710 167177 674762 167229
rect 144022 167103 144074 167155
rect 156982 167103 157034 167155
rect 144118 167029 144170 167081
rect 148726 167029 148778 167081
rect 646198 164217 646250 164269
rect 674614 164217 674666 164269
rect 144022 164143 144074 164195
rect 148822 164143 148874 164195
rect 645910 164143 645962 164195
rect 674710 164143 674762 164195
rect 675286 164069 675338 164121
rect 677014 164069 677066 164121
rect 674806 163255 674858 163307
rect 676822 163255 676874 163307
rect 144022 161331 144074 161383
rect 148918 161331 148970 161383
rect 144118 161257 144170 161309
rect 197302 161257 197354 161309
rect 674422 160739 674474 160791
rect 675382 160739 675434 160791
rect 675190 159999 675242 160051
rect 675478 159999 675530 160051
rect 674038 159407 674090 159459
rect 675382 159407 675434 159459
rect 144022 158445 144074 158497
rect 149206 158445 149258 158497
rect 144886 157113 144938 157165
rect 146806 157113 146858 157165
rect 674998 157039 675050 157091
rect 675190 157039 675242 157091
rect 144886 156965 144938 157017
rect 146614 156965 146666 157017
rect 674902 156891 674954 156943
rect 675478 156891 675530 156943
rect 144022 155559 144074 155611
rect 149302 155559 149354 155611
rect 144022 152747 144074 152799
rect 177142 152747 177194 152799
rect 144118 152673 144170 152725
rect 180022 152673 180074 152725
rect 674326 152599 674378 152651
rect 675382 152599 675434 152651
rect 674806 152155 674858 152207
rect 675478 152155 675530 152207
rect 674518 151415 674570 151467
rect 675382 151415 675434 151467
rect 144118 149861 144170 149913
rect 149398 149861 149450 149913
rect 144022 149787 144074 149839
rect 174358 149787 174410 149839
rect 209782 149787 209834 149839
rect 209974 149787 210026 149839
rect 144022 149639 144074 149691
rect 144310 149639 144362 149691
rect 144310 149491 144362 149543
rect 144502 149491 144554 149543
rect 209974 148233 210026 148285
rect 210166 148233 210218 148285
rect 144022 146975 144074 147027
rect 149494 146975 149546 147027
rect 144214 146901 144266 146953
rect 171478 146901 171530 146953
rect 210070 146975 210122 147027
rect 210262 146827 210314 146879
rect 209974 146753 210026 146805
rect 210070 146679 210122 146731
rect 144694 144311 144746 144363
rect 144886 144311 144938 144363
rect 144214 144015 144266 144067
rect 154102 144015 154154 144067
rect 144694 141351 144746 141403
rect 144406 141203 144458 141255
rect 149590 141203 149642 141255
rect 144214 141129 144266 141181
rect 168598 141129 168650 141181
rect 146518 141055 146570 141107
rect 144214 140981 144266 141033
rect 147190 140981 147242 141033
rect 146038 140463 146090 140515
rect 146710 140463 146762 140515
rect 144214 138539 144266 138591
rect 655222 138539 655274 138591
rect 674710 138539 674762 138591
rect 655126 138391 655178 138443
rect 674422 138391 674474 138443
rect 144214 138317 144266 138369
rect 149686 138317 149738 138369
rect 144406 138243 144458 138295
rect 165718 138243 165770 138295
rect 144406 138095 144458 138147
rect 144886 136911 144938 136963
rect 144502 136763 144554 136815
rect 144886 136763 144938 136815
rect 146518 136615 146570 136667
rect 144406 136245 144458 136297
rect 144694 136245 144746 136297
rect 144598 136171 144650 136223
rect 144598 135949 144650 136001
rect 655414 135579 655466 135631
rect 674614 135579 674666 135631
rect 144502 135431 144554 135483
rect 147094 135431 147146 135483
rect 646486 135357 646538 135409
rect 674710 135357 674762 135409
rect 143926 134099 143978 134151
rect 144406 134099 144458 134151
rect 146710 134099 146762 134151
rect 146998 134099 147050 134151
rect 144502 132693 144554 132745
rect 162934 132693 162986 132745
rect 144406 132545 144458 132597
rect 208822 132545 208874 132597
rect 144214 132471 144266 132523
rect 208918 132471 208970 132523
rect 143926 132397 143978 132449
rect 144502 132397 144554 132449
rect 144214 130103 144266 130155
rect 151318 130103 151370 130155
rect 144214 129585 144266 129637
rect 209014 129585 209066 129637
rect 144214 129437 144266 129489
rect 144694 129437 144746 129489
rect 146518 129363 146570 129415
rect 144694 129289 144746 129341
rect 146902 126995 146954 127047
rect 148150 126995 148202 127047
rect 209974 126995 210026 127047
rect 146902 126773 146954 126825
rect 148054 126773 148106 126825
rect 146518 126699 146570 126751
rect 200278 126699 200330 126751
rect 209974 126699 210026 126751
rect 210166 126699 210218 126751
rect 210262 126699 210314 126751
rect 146902 126625 146954 126677
rect 147190 126625 147242 126677
rect 144790 125293 144842 125345
rect 146614 125293 146666 125345
rect 144598 124479 144650 124531
rect 146038 124479 146090 124531
rect 144598 123961 144650 124013
rect 194518 123961 194570 124013
rect 144790 123887 144842 123939
rect 197398 123887 197450 123939
rect 647830 121223 647882 121275
rect 674710 121223 674762 121275
rect 144598 121149 144650 121201
rect 203062 121149 203114 121201
rect 647926 121149 647978 121201
rect 674806 121149 674858 121201
rect 647830 121075 647882 121127
rect 674614 121075 674666 121127
rect 144790 121001 144842 121053
rect 209110 121001 209162 121053
rect 674806 119965 674858 120017
rect 675190 119965 675242 120017
rect 674134 118929 674186 118981
rect 674422 118929 674474 118981
rect 144598 118559 144650 118611
rect 191638 118559 191690 118611
rect 144598 118263 144650 118315
rect 185878 118263 185930 118315
rect 144790 118115 144842 118167
rect 209206 118115 209258 118167
rect 674614 118041 674666 118093
rect 676822 118041 676874 118093
rect 144790 117967 144842 118019
rect 146614 117967 146666 118019
rect 674422 117967 674474 118019
rect 676918 117967 676970 118019
rect 146230 116635 146282 116687
rect 146614 116635 146666 116687
rect 146230 115599 146282 115651
rect 146902 115377 146954 115429
rect 146710 115303 146762 115355
rect 209302 115303 209354 115355
rect 144598 115229 144650 115281
rect 209398 115229 209450 115281
rect 146902 114859 146954 114911
rect 146518 114267 146570 114319
rect 146998 114267 147050 114319
rect 146518 114119 146570 114171
rect 674134 114119 674186 114171
rect 675382 114119 675434 114171
rect 674038 113601 674090 113653
rect 675190 113601 675242 113653
rect 674230 113305 674282 113357
rect 675094 113305 675146 113357
rect 144790 113231 144842 113283
rect 146902 113231 146954 113283
rect 647926 112861 647978 112913
rect 665206 112861 665258 112913
rect 144598 112491 144650 112543
rect 188758 112491 188810 112543
rect 144790 112417 144842 112469
rect 203158 112417 203210 112469
rect 144598 112343 144650 112395
rect 209494 112343 209546 112395
rect 674326 111159 674378 111211
rect 675382 111159 675434 111211
rect 146518 111085 146570 111137
rect 146230 110937 146282 110989
rect 146518 110937 146570 110989
rect 146230 110789 146282 110841
rect 144790 109531 144842 109583
rect 162838 109531 162890 109583
rect 144598 109457 144650 109509
rect 182998 109457 183050 109509
rect 144790 109383 144842 109435
rect 146038 109383 146090 109435
rect 144598 107459 144650 107511
rect 160150 107459 160202 107511
rect 674518 107311 674570 107363
rect 675382 107311 675434 107363
rect 674614 106941 674666 106993
rect 675478 106941 675530 106993
rect 143926 106719 143978 106771
rect 144790 106719 144842 106771
rect 146230 106645 146282 106697
rect 144790 106571 144842 106623
rect 146038 106571 146090 106623
rect 193942 106571 193994 106623
rect 144022 106497 144074 106549
rect 146230 106497 146282 106549
rect 143926 106349 143978 106401
rect 144310 106349 144362 106401
rect 673942 106127 673994 106179
rect 675382 106127 675434 106179
rect 144118 105979 144170 106031
rect 146038 105979 146090 106031
rect 674422 105165 674474 105217
rect 675382 105165 675434 105217
rect 144022 104351 144074 104403
rect 159958 104351 160010 104403
rect 144022 104203 144074 104255
rect 157078 104203 157130 104255
rect 144118 103685 144170 103737
rect 209590 103685 209642 103737
rect 146614 103611 146666 103663
rect 201718 103611 201770 103663
rect 144790 103537 144842 103589
rect 199990 103537 200042 103589
rect 146518 103463 146570 103515
rect 210166 103463 210218 103515
rect 146710 103389 146762 103441
rect 146998 103389 147050 103441
rect 144022 100873 144074 100925
rect 149014 100873 149066 100925
rect 144118 100799 144170 100851
rect 209686 100799 209738 100851
rect 201814 100725 201866 100777
rect 144310 100651 144362 100703
rect 146902 100651 146954 100703
rect 201622 100651 201674 100703
rect 151126 100577 151178 100629
rect 201718 100577 201770 100629
rect 159766 100503 159818 100555
rect 210166 100503 210218 100555
rect 185686 100429 185738 100481
rect 201718 100429 201770 100481
rect 144022 98283 144074 98335
rect 160054 98283 160106 98335
rect 144022 97987 144074 98039
rect 177238 97987 177290 98039
rect 144118 97913 144170 97965
rect 180118 97913 180170 97965
rect 156886 97765 156938 97817
rect 210166 97765 210218 97817
rect 168502 97691 168554 97743
rect 201814 97691 201866 97743
rect 171382 97617 171434 97669
rect 201622 97617 201674 97669
rect 174262 97543 174314 97595
rect 201718 97543 201770 97595
rect 154006 97469 154058 97521
rect 210166 97469 210218 97521
rect 663190 96433 663242 96485
rect 665206 96433 665258 96485
rect 144406 95397 144458 95449
rect 146614 95397 146666 95449
rect 146518 95101 146570 95153
rect 171574 95101 171626 95153
rect 144022 95027 144074 95079
rect 174454 95027 174506 95079
rect 162742 94879 162794 94931
rect 201718 94879 201770 94931
rect 165622 94805 165674 94857
rect 210166 94805 210218 94857
rect 144598 94657 144650 94709
rect 201622 94657 201674 94709
rect 193942 94065 193994 94117
rect 209590 94065 209642 94117
rect 646486 92659 646538 92711
rect 659830 92659 659882 92711
rect 647542 92585 647594 92637
rect 661750 92585 661802 92637
rect 647350 92511 647402 92563
rect 660694 92511 660746 92563
rect 646102 92437 646154 92489
rect 663094 92437 663146 92489
rect 647830 92289 647882 92341
rect 662518 92289 662570 92341
rect 144118 92215 144170 92267
rect 154006 92215 154058 92267
rect 647254 92215 647306 92267
rect 661174 92215 661226 92267
rect 144022 92141 144074 92193
rect 168502 92141 168554 92193
rect 646582 92141 646634 92193
rect 658870 92141 658922 92193
rect 146230 92067 146282 92119
rect 201718 92067 201770 92119
rect 146038 91993 146090 92045
rect 197686 91993 197738 92045
rect 151222 91919 151274 91971
rect 201622 91919 201674 91971
rect 185782 91845 185834 91897
rect 201814 91845 201866 91897
rect 144118 91179 144170 91231
rect 144310 91179 144362 91231
rect 144022 89403 144074 89455
rect 151126 89403 151178 89455
rect 144118 89329 144170 89381
rect 163126 89329 163178 89381
rect 146230 89255 146282 89307
rect 165814 89255 165866 89307
rect 144118 89181 144170 89233
rect 144790 89181 144842 89233
rect 156982 89181 157034 89233
rect 201814 89181 201866 89233
rect 159862 89107 159914 89159
rect 201622 89107 201674 89159
rect 182902 89033 182954 89085
rect 201526 89033 201578 89085
rect 188662 88959 188714 89011
rect 198742 88959 198794 89011
rect 191542 88885 191594 88937
rect 201718 88885 201770 88937
rect 646294 87553 646346 87605
rect 650998 87553 651050 87605
rect 652342 87331 652394 87383
rect 659350 87331 659402 87383
rect 658006 87257 658058 87309
rect 657046 87109 657098 87161
rect 647926 87035 647978 87087
rect 663286 87035 663338 87087
rect 646390 86739 646442 86791
rect 651094 86739 651146 86791
rect 144022 86443 144074 86495
rect 162742 86443 162794 86495
rect 144598 86369 144650 86421
rect 144886 86369 144938 86421
rect 154102 86369 154154 86421
rect 201910 86369 201962 86421
rect 171478 86295 171530 86347
rect 201526 86295 201578 86347
rect 174358 86221 174410 86273
rect 201814 86221 201866 86273
rect 177142 86147 177194 86199
rect 201622 86147 201674 86199
rect 180022 86073 180074 86125
rect 201718 86073 201770 86125
rect 144022 84963 144074 85015
rect 201718 84963 201770 85015
rect 646486 84889 646538 84941
rect 650902 84889 650954 84941
rect 145942 83631 145994 83683
rect 146230 83631 146282 83683
rect 151318 83483 151370 83535
rect 194614 83483 194666 83535
rect 162934 83409 162986 83461
rect 201622 83409 201674 83461
rect 165718 83335 165770 83387
rect 201718 83335 201770 83387
rect 168598 83261 168650 83313
rect 201046 83261 201098 83313
rect 646294 83113 646346 83165
rect 657046 83113 657098 83165
rect 144022 82077 144074 82129
rect 197782 82077 197834 82129
rect 646102 81855 646154 81907
rect 663286 81855 663338 81907
rect 646006 81781 646058 81833
rect 663382 81781 663434 81833
rect 647638 81633 647690 81685
rect 661078 81633 661130 81685
rect 647926 81411 647978 81463
rect 657526 81411 657578 81463
rect 144022 80745 144074 80797
rect 163030 80745 163082 80797
rect 144118 80671 144170 80723
rect 144694 80671 144746 80723
rect 659446 80671 659498 80723
rect 659542 80671 659594 80723
rect 185878 80597 185930 80649
rect 201718 80597 201770 80649
rect 191638 80523 191690 80575
rect 200374 80523 200426 80575
rect 646870 80227 646922 80279
rect 656950 80227 657002 80279
rect 647926 79339 647978 79391
rect 660694 79339 660746 79391
rect 640726 79191 640778 79243
rect 663190 79191 663242 79243
rect 646870 78895 646922 78947
rect 658870 78895 658922 78947
rect 646870 78303 646922 78355
rect 651190 78303 651242 78355
rect 646486 78229 646538 78281
rect 662518 78229 662570 78281
rect 144022 77859 144074 77911
rect 165622 77859 165674 77911
rect 144118 77785 144170 77837
rect 185686 77785 185738 77837
rect 149014 77711 149066 77763
rect 201526 77711 201578 77763
rect 647926 77711 647978 77763
rect 662902 77711 662954 77763
rect 157078 77637 157130 77689
rect 201814 77637 201866 77689
rect 646678 77637 646730 77689
rect 658294 77637 658346 77689
rect 160150 77563 160202 77615
rect 195574 77563 195626 77615
rect 646294 77563 646346 77615
rect 650902 77563 650954 77615
rect 182998 77489 183050 77541
rect 201622 77489 201674 77541
rect 647830 77489 647882 77541
rect 650998 77489 651050 77541
rect 185686 77415 185738 77467
rect 201718 77415 201770 77467
rect 647446 77415 647498 77467
rect 659446 77415 659498 77467
rect 188758 77341 188810 77393
rect 210262 77341 210314 77393
rect 144118 76527 144170 76579
rect 144598 76527 144650 76579
rect 144406 76453 144458 76505
rect 144214 76305 144266 76357
rect 144406 76305 144458 76357
rect 144598 76305 144650 76357
rect 145174 76305 145226 76357
rect 144790 76231 144842 76283
rect 146038 76231 146090 76283
rect 145174 76157 145226 76209
rect 647926 76083 647978 76135
rect 661750 76083 661802 76135
rect 646486 75639 646538 75691
rect 656854 75639 656906 75691
rect 144118 74973 144170 75025
rect 160150 74973 160202 75025
rect 144022 74899 144074 74951
rect 155542 74899 155594 74951
rect 144118 74825 144170 74877
rect 208726 74825 208778 74877
rect 154006 74751 154058 74803
rect 201718 74751 201770 74803
rect 171574 74677 171626 74729
rect 200950 74677 201002 74729
rect 174454 74603 174506 74655
rect 198358 74603 198410 74655
rect 177238 74529 177290 74581
rect 201046 74529 201098 74581
rect 180118 74455 180170 74507
rect 210262 74455 210314 74507
rect 144790 72679 144842 72731
rect 145366 72679 145418 72731
rect 144118 72605 144170 72657
rect 144310 72605 144362 72657
rect 145366 72531 145418 72583
rect 146806 72531 146858 72583
rect 646294 72531 646346 72583
rect 663286 72531 663338 72583
rect 144310 72457 144362 72509
rect 146230 72457 146282 72509
rect 646102 72383 646154 72435
rect 663478 72383 663530 72435
rect 146230 72309 146282 72361
rect 146518 72309 146570 72361
rect 145174 72161 145226 72213
rect 146518 72161 146570 72213
rect 647158 72161 647210 72213
rect 660118 72161 660170 72213
rect 144022 72013 144074 72065
rect 154102 72013 154154 72065
rect 146902 71939 146954 71991
rect 200470 71939 200522 71991
rect 208630 71939 208682 71991
rect 209206 71939 209258 71991
rect 151126 71865 151178 71917
rect 201814 71865 201866 71917
rect 163126 71791 163178 71843
rect 201622 71791 201674 71843
rect 165814 71717 165866 71769
rect 209974 71717 210026 71769
rect 168502 71643 168554 71695
rect 201718 71643 201770 71695
rect 144022 70237 144074 70289
rect 149782 70237 149834 70289
rect 145174 69497 145226 69549
rect 145558 69497 145610 69549
rect 144214 69349 144266 69401
rect 145558 69349 145610 69401
rect 144022 69127 144074 69179
rect 201526 69053 201578 69105
rect 149782 68979 149834 69031
rect 201814 68979 201866 69031
rect 154102 68905 154154 68957
rect 201622 68905 201674 68957
rect 155542 68831 155594 68883
rect 201718 68831 201770 68883
rect 160150 68757 160202 68809
rect 194710 68757 194762 68809
rect 144022 66981 144074 67033
rect 152662 66981 152714 67033
rect 144214 66537 144266 66589
rect 158326 66537 158378 66589
rect 144886 66315 144938 66367
rect 145558 66315 145610 66367
rect 144022 66241 144074 66293
rect 144214 66167 144266 66219
rect 144694 66167 144746 66219
rect 200182 66167 200234 66219
rect 152662 66093 152714 66145
rect 201718 66093 201770 66145
rect 145558 66019 145610 66071
rect 145846 66019 145898 66071
rect 158326 66019 158378 66071
rect 201622 66019 201674 66071
rect 146038 65575 146090 65627
rect 146230 65575 146282 65627
rect 146230 64835 146282 64887
rect 201718 64835 201770 64887
rect 144022 64761 144074 64813
rect 193750 64761 193802 64813
rect 146902 63355 146954 63407
rect 201718 63355 201770 63407
rect 208726 63059 208778 63111
rect 209590 63059 209642 63111
rect 209686 62837 209738 62889
rect 210166 62837 210218 62889
rect 144022 62171 144074 62223
rect 151414 62171 151466 62223
rect 208246 61949 208298 62001
rect 208918 61949 208970 62001
rect 208534 61875 208586 61927
rect 209014 61875 209066 61927
rect 208150 61801 208202 61853
rect 208822 61801 208874 61853
rect 147958 60765 148010 60817
rect 148246 60765 148298 60817
rect 169942 60765 169994 60817
rect 201718 60765 201770 60817
rect 167062 60691 167114 60743
rect 194134 60691 194186 60743
rect 164182 60617 164234 60669
rect 209974 60617 210026 60669
rect 152470 60543 152522 60595
rect 201622 60543 201674 60595
rect 148438 60469 148490 60521
rect 199318 60469 199370 60521
rect 146902 60395 146954 60447
rect 201718 60395 201770 60447
rect 151414 60321 151466 60373
rect 209974 60321 210026 60373
rect 146518 60247 146570 60299
rect 169942 60247 169994 60299
rect 208630 59137 208682 59189
rect 209014 59137 209066 59189
rect 144022 58989 144074 59041
rect 201622 58989 201674 59041
rect 144118 58619 144170 58671
rect 144214 58397 144266 58449
rect 144022 57509 144074 57561
rect 167062 57509 167114 57561
rect 144118 57435 144170 57487
rect 164182 57435 164234 57487
rect 144022 54623 144074 54675
rect 152470 54623 152522 54675
rect 210070 54327 210122 54379
rect 213814 54327 213866 54379
rect 214198 54327 214250 54379
rect 216022 54327 216074 54379
rect 209782 54253 209834 54305
rect 216406 54253 216458 54305
rect 206614 54179 206666 54231
rect 218230 54179 218282 54231
rect 144022 54105 144074 54157
rect 148438 54105 148490 54157
rect 206518 54105 206570 54157
rect 220438 54105 220490 54157
rect 209494 54031 209546 54083
rect 218230 54031 218282 54083
rect 206998 53957 207050 54009
rect 218422 53957 218474 54009
rect 206902 53883 206954 53935
rect 216214 53883 216266 53935
rect 210646 53809 210698 53861
rect 206422 53735 206474 53787
rect 209398 53661 209450 53713
rect 210262 53587 210314 53639
rect 210358 53513 210410 53565
rect 217798 53513 217850 53565
rect 219430 53587 219482 53639
rect 221446 53587 221498 53639
rect 231766 53587 231818 53639
rect 246742 53661 246794 53713
rect 282262 53735 282314 53787
rect 282070 53661 282122 53713
rect 345622 53661 345674 53713
rect 241846 53513 241898 53565
rect 241942 53513 241994 53565
rect 380182 53513 380234 53565
rect 209590 53439 209642 53491
rect 217270 53439 217322 53491
rect 218422 53439 218474 53491
rect 219574 53439 219626 53491
rect 220630 53439 220682 53491
rect 289174 53439 289226 53491
rect 417622 53439 417674 53491
rect 440566 53439 440618 53491
rect 208726 53365 208778 53417
rect 217558 53365 217610 53417
rect 206710 53291 206762 53343
rect 217366 53291 217418 53343
rect 206806 53217 206858 53269
rect 215542 53217 215594 53269
rect 210166 53143 210218 53195
rect 262102 53365 262154 53417
rect 262198 53365 262250 53417
rect 463702 53365 463754 53417
rect 246742 53291 246794 53343
rect 209974 53069 210026 53121
rect 221782 53069 221834 53121
rect 262390 53217 262442 53269
rect 282358 53217 282410 53269
rect 283606 53217 283658 53269
rect 316918 53291 316970 53343
rect 383158 53291 383210 53343
rect 383254 53291 383306 53343
rect 423286 53291 423338 53343
rect 463606 53291 463658 53343
rect 498742 53291 498794 53343
rect 293782 53217 293834 53269
rect 293686 53143 293738 53195
rect 296566 53143 296618 53195
rect 296758 53143 296810 53195
rect 328534 53143 328586 53195
rect 273622 53069 273674 53121
rect 313846 53069 313898 53121
rect 316726 53069 316778 53121
rect 328630 53069 328682 53121
rect 354262 53143 354314 53195
rect 417622 53217 417674 53269
rect 440566 53217 440618 53269
rect 509878 53217 509930 53269
rect 525910 53217 525962 53269
rect 509686 53143 509738 53195
rect 374326 53069 374378 53121
rect 443542 53069 443594 53121
rect 463606 53069 463658 53121
rect 211798 52995 211850 53047
rect 261910 52995 261962 53047
rect 207094 52921 207146 52973
rect 219286 52921 219338 52973
rect 221782 52921 221834 52973
rect 231766 52921 231818 52973
rect 282358 52921 282410 52973
rect 293686 52921 293738 52973
rect 293782 52921 293834 52973
rect 313846 52921 313898 52973
rect 210070 52847 210122 52899
rect 218806 52847 218858 52899
rect 273622 52847 273674 52899
rect 283606 52847 283658 52899
rect 165622 52551 165674 52603
rect 216118 52551 216170 52603
rect 162838 52403 162890 52455
rect 217942 52403 217994 52455
rect 212278 52181 212330 52233
rect 220438 52181 220490 52233
rect 160054 52107 160106 52159
rect 215734 52107 215786 52159
rect 163030 52033 163082 52085
rect 220918 52033 220970 52085
rect 159958 51959 160010 52011
rect 216886 51959 216938 52011
rect 223606 51959 223658 52011
rect 241174 51959 241226 52011
rect 162742 51885 162794 51937
rect 227542 51885 227594 51937
rect 625750 51885 625802 51937
rect 639670 51885 639722 51937
rect 209878 51811 209930 51863
rect 214486 51811 214538 51863
rect 220438 51811 220490 51863
rect 645526 51811 645578 51863
rect 208342 51737 208394 51789
rect 213334 51737 213386 51789
rect 219478 51737 219530 51789
rect 645718 51737 645770 51789
rect 208438 51663 208490 51715
rect 214102 51663 214154 51715
rect 145750 51589 145802 51641
rect 223606 51589 223658 51641
rect 211126 51515 211178 51567
rect 348406 51589 348458 51641
rect 348502 51589 348554 51641
rect 362902 51663 362954 51715
rect 383062 51515 383114 51567
rect 403222 51663 403274 51715
rect 423382 51515 423434 51567
rect 434902 51663 434954 51715
rect 509686 51663 509738 51715
rect 520246 51663 520298 51715
rect 459286 51589 459338 51641
rect 489622 51589 489674 51641
rect 520246 51515 520298 51567
rect 550006 51589 550058 51641
rect 550102 51589 550154 51641
rect 558838 51663 558890 51715
rect 558838 51515 558890 51567
rect 601942 51663 601994 51715
rect 622006 51589 622058 51641
rect 625750 51589 625802 51641
rect 211510 51441 211562 51493
rect 219478 51441 219530 51493
rect 144982 51367 145034 51419
rect 233782 51367 233834 51419
rect 145462 51293 145514 51345
rect 235990 51293 236042 51345
rect 145654 51219 145706 51271
rect 235030 51219 235082 51271
rect 146134 51145 146186 51197
rect 231958 51145 232010 51197
rect 146422 51071 146474 51123
rect 231190 51071 231242 51123
rect 146326 50997 146378 51049
rect 231574 50997 231626 51049
rect 146806 50923 146858 50975
rect 230518 50923 230570 50975
rect 498742 50923 498794 50975
rect 504022 50923 504074 50975
rect 145078 50849 145130 50901
rect 228982 50849 229034 50901
rect 289174 50849 289226 50901
rect 302422 50849 302474 50901
rect 159382 50775 159434 50827
rect 243862 50775 243914 50827
rect 145270 50701 145322 50753
rect 228406 50701 228458 50753
rect 146710 50627 146762 50679
rect 229750 50627 229802 50679
rect 145366 50553 145418 50605
rect 229366 50553 229418 50605
rect 144118 50479 144170 50531
rect 144886 50405 144938 50457
rect 145942 50331 145994 50383
rect 224950 50405 225002 50457
rect 146038 50257 146090 50309
rect 210838 50257 210890 50309
rect 226102 50331 226154 50383
rect 227158 50257 227210 50309
rect 145846 50183 145898 50235
rect 225718 50183 225770 50235
rect 144214 50109 144266 50161
rect 223126 50109 223178 50161
rect 144406 50035 144458 50087
rect 223510 50035 223562 50087
rect 144502 49961 144554 50013
rect 224182 49961 224234 50013
rect 145174 49887 145226 49939
rect 235606 49887 235658 49939
rect 145558 49813 145610 49865
rect 234646 49813 234698 49865
rect 144310 49739 144362 49791
rect 232438 49739 232490 49791
rect 210838 49665 210890 49717
rect 226774 49665 226826 49717
rect 144598 49591 144650 49643
rect 234550 49591 234602 49643
rect 144790 49517 144842 49569
rect 236758 49517 236810 49569
rect 218614 49073 218666 49125
rect 208630 48925 208682 48977
rect 345622 48999 345674 49051
rect 353590 48999 353642 49051
rect 463702 48999 463754 49051
rect 471382 48999 471434 49051
rect 625078 48999 625130 49051
rect 640726 48999 640778 49051
rect 645622 48925 645674 48977
rect 209302 48777 209354 48829
rect 219094 48777 219146 48829
rect 209014 48629 209066 48681
rect 219766 48629 219818 48681
rect 224086 48851 224138 48903
rect 645334 48851 645386 48903
rect 222934 48777 222986 48829
rect 645142 48777 645194 48829
rect 222166 48703 222218 48755
rect 645238 48703 645290 48755
rect 226390 48629 226442 48681
rect 504022 48629 504074 48681
rect 512566 48629 512618 48681
rect 203062 48555 203114 48607
rect 208726 48555 208778 48607
rect 208822 48555 208874 48607
rect 220534 48555 220586 48607
rect 191446 48481 191498 48533
rect 240790 48481 240842 48533
rect 182806 48407 182858 48459
rect 199222 48407 199274 48459
rect 200086 48407 200138 48459
rect 241270 48407 241322 48459
rect 148822 48333 148874 48385
rect 227926 48333 227978 48385
rect 149302 48259 149354 48311
rect 230134 48259 230186 48311
rect 380182 48259 380234 48311
rect 394582 48259 394634 48311
rect 149398 48185 149450 48237
rect 208630 48185 208682 48237
rect 208726 48185 208778 48237
rect 220150 48185 220202 48237
rect 149494 48111 149546 48163
rect 208438 48111 208490 48163
rect 208534 48111 208586 48163
rect 221974 48111 222026 48163
rect 149590 48037 149642 48089
rect 208054 48037 208106 48089
rect 208246 48037 208298 48089
rect 222358 48037 222410 48089
rect 149686 47963 149738 48015
rect 208150 47963 208202 48015
rect 222742 47963 222794 48015
rect 223894 47889 223946 47941
rect 199222 47815 199274 47867
rect 240406 47815 240458 47867
rect 148150 47667 148202 47719
rect 221686 47741 221738 47793
rect 148054 47593 148106 47645
rect 221302 47667 221354 47719
rect 177046 47593 177098 47645
rect 238582 47593 238634 47645
rect 208054 47519 208106 47571
rect 224566 47519 224618 47571
rect 208438 47445 208490 47497
rect 225334 47445 225386 47497
rect 149206 47371 149258 47423
rect 233398 47371 233450 47423
rect 197206 46853 197258 46905
rect 239062 46853 239114 46905
rect 148918 46779 148970 46831
rect 234166 46779 234218 46831
rect 148630 46705 148682 46757
rect 230614 46705 230666 46757
rect 148342 46631 148394 46683
rect 232822 46631 232874 46683
rect 148534 46557 148586 46609
rect 232342 46557 232394 46609
rect 148726 46483 148778 46535
rect 228022 46483 228074 46535
rect 179926 46409 179978 46461
rect 238966 46409 239018 46461
rect 148246 46335 148298 46387
rect 236854 46335 236906 46387
rect 147958 46113 148010 46165
rect 236374 46113 236426 46165
rect 212854 44781 212906 44833
rect 408886 44781 408938 44833
rect 213910 44707 213962 44759
rect 457750 44707 457802 44759
rect 141814 44633 141866 44685
rect 155542 44633 155594 44685
rect 214678 44633 214730 44685
rect 509782 44633 509834 44685
rect 509782 43227 509834 43279
rect 394582 43153 394634 43205
rect 408982 43153 409034 43205
rect 521590 43153 521642 43205
rect 212470 42339 212522 42391
rect 310102 42339 310154 42391
rect 207286 42117 207338 42169
rect 405238 42117 405290 42169
rect 512566 42117 512618 42169
rect 520342 42117 520394 42169
rect 213526 42043 213578 42095
rect 460054 42043 460106 42095
rect 514870 41747 514922 41799
rect 214294 41673 214346 41725
<< metal2 >>
rect 439222 1005797 439274 1005803
rect 439222 1005739 439274 1005745
rect 466582 1005797 466634 1005803
rect 466582 1005739 466634 1005745
rect 371830 1005723 371882 1005729
rect 371830 1005665 371882 1005671
rect 92374 1005575 92426 1005581
rect 92374 1005517 92426 1005523
rect 92386 1005304 92414 1005517
rect 108598 1005501 108650 1005507
rect 108596 1005466 108598 1005475
rect 357910 1005501 357962 1005507
rect 108650 1005466 108652 1005475
rect 93622 1005427 93674 1005433
rect 108596 1005401 108652 1005410
rect 114164 1005466 114220 1005475
rect 308756 1005466 308812 1005475
rect 114164 1005401 114166 1005410
rect 93622 1005369 93674 1005375
rect 114218 1005401 114220 1005410
rect 298102 1005427 298154 1005433
rect 114166 1005369 114218 1005375
rect 308756 1005401 308758 1005410
rect 298102 1005369 298154 1005375
rect 308810 1005401 308812 1005410
rect 321044 1005466 321100 1005475
rect 321428 1005466 321484 1005475
rect 321100 1005424 321428 1005452
rect 321044 1005401 321100 1005410
rect 321428 1005401 321484 1005410
rect 325460 1005466 325516 1005475
rect 325460 1005401 325516 1005410
rect 357908 1005466 357910 1005475
rect 365014 1005501 365066 1005507
rect 357962 1005466 357964 1005475
rect 357908 1005401 357964 1005410
rect 364148 1005466 364204 1005475
rect 364148 1005401 364150 1005410
rect 308758 1005369 308810 1005375
rect 92290 1005276 92414 1005304
rect 81044 995846 81100 995855
rect 80784 995804 81044 995832
rect 92290 995832 92318 1005276
rect 93046 999655 93098 999661
rect 93046 999597 93098 999603
rect 82032 995813 82334 995832
rect 87552 995813 87902 995832
rect 82032 995807 82346 995813
rect 82032 995804 82294 995807
rect 81044 995781 81100 995790
rect 87552 995807 87914 995813
rect 87552 995804 87862 995807
rect 82294 995749 82346 995755
rect 87862 995749 87914 995755
rect 92098 995804 92318 995832
rect 91510 995733 91562 995739
rect 85940 995698 85996 995707
rect 85728 995656 85940 995684
rect 91248 995681 91510 995684
rect 91248 995675 91562 995681
rect 91248 995656 91550 995675
rect 85940 995633 85996 995642
rect 77088 995508 77342 995536
rect 69142 995215 69194 995221
rect 69142 995157 69194 995163
rect 61844 993922 61900 993931
rect 61844 993857 61900 993866
rect 45046 985521 45098 985527
rect 45046 985463 45098 985469
rect 44950 985151 45002 985157
rect 44950 985093 45002 985099
rect 44854 985077 44906 985083
rect 44854 985019 44906 985025
rect 42934 985003 42986 985009
rect 42934 984945 42986 984951
rect 42082 968771 42110 969252
rect 42068 968762 42124 968771
rect 42068 968697 42124 968706
rect 41794 967143 41822 967402
rect 42946 967323 42974 984945
rect 44758 983745 44810 983751
rect 44758 983687 44810 983693
rect 44566 983671 44618 983677
rect 44566 983613 44618 983619
rect 42166 967317 42218 967323
rect 42166 967259 42218 967265
rect 42934 967317 42986 967323
rect 42934 967259 42986 967265
rect 41780 967134 41836 967143
rect 41780 967069 41836 967078
rect 42178 966736 42206 967259
rect 41794 965071 41822 965552
rect 41780 965062 41836 965071
rect 41780 964997 41836 965006
rect 42178 964035 42206 964368
rect 42164 964026 42220 964035
rect 42164 963961 42220 963970
rect 41794 963443 41822 963702
rect 41780 963434 41836 963443
rect 41780 963369 41836 963378
rect 42178 962851 42206 963081
rect 42164 962842 42220 962851
rect 42164 962777 42220 962786
rect 42548 962546 42604 962555
rect 41890 962111 41918 962518
rect 42548 962481 42604 962490
rect 41876 962102 41932 962111
rect 41876 962037 41932 962046
rect 42356 962102 42412 962111
rect 42356 962037 42412 962046
rect 42070 961397 42122 961403
rect 42070 961339 42122 961345
rect 42082 961260 42110 961339
rect 42370 960737 42398 962037
rect 42562 961403 42590 962481
rect 42550 961397 42602 961403
rect 42550 961339 42602 961345
rect 42166 960731 42218 960737
rect 42166 960673 42218 960679
rect 42358 960731 42410 960737
rect 42358 960673 42410 960679
rect 42178 960594 42206 960673
rect 41794 959743 41822 960045
rect 41780 959734 41836 959743
rect 41780 959669 41836 959678
rect 41794 959151 41822 959410
rect 41780 959142 41836 959151
rect 41780 959077 41836 959086
rect 41986 958411 42014 958744
rect 41972 958402 42028 958411
rect 41972 958337 42028 958346
rect 41794 957819 41822 958226
rect 41780 957810 41836 957819
rect 41780 957745 41836 957754
rect 41794 956191 41822 956376
rect 41780 956182 41836 956191
rect 41780 956117 41836 956126
rect 42082 955335 42110 955710
rect 42070 955329 42122 955335
rect 42070 955271 42122 955277
rect 42178 954669 42206 955077
rect 42166 954663 42218 954669
rect 42166 954605 42218 954611
rect 42164 949374 42220 949383
rect 42164 949309 42220 949318
rect 42178 947713 42206 949309
rect 42370 948601 42398 960673
rect 42562 953231 42590 961339
rect 43126 956217 43178 956223
rect 43126 956159 43178 956165
rect 42934 955329 42986 955335
rect 42934 955271 42986 955277
rect 42838 954663 42890 954669
rect 42838 954605 42890 954611
rect 42548 953222 42604 953231
rect 42548 953157 42604 953166
rect 42358 948595 42410 948601
rect 42358 948537 42410 948543
rect 42646 948595 42698 948601
rect 42646 948537 42698 948543
rect 42356 948486 42412 948495
rect 42356 948421 42412 948430
rect 42370 947787 42398 948421
rect 42358 947781 42410 947787
rect 42358 947723 42410 947729
rect 42166 947707 42218 947713
rect 42166 947649 42218 947655
rect 42658 947607 42686 948537
rect 42644 947598 42700 947607
rect 42644 947533 42700 947542
rect 40340 946562 40396 946571
rect 40340 946497 40396 946506
rect 40052 945082 40108 945091
rect 40052 945017 40108 945026
rect 40066 820179 40094 945017
rect 40354 820771 40382 946497
rect 42850 942279 42878 954605
rect 42836 942270 42892 942279
rect 42836 942205 42892 942214
rect 42946 939171 42974 955271
rect 43138 947903 43166 956159
rect 43124 947894 43180 947903
rect 43124 947829 43180 947838
rect 43028 947006 43084 947015
rect 43028 946941 43084 946950
rect 42932 939162 42988 939171
rect 42932 939097 42988 939106
rect 43042 933103 43070 946941
rect 44578 944795 44606 983613
rect 44770 945683 44798 983687
rect 44756 945674 44812 945683
rect 44756 945609 44812 945618
rect 44564 944786 44620 944795
rect 44564 944721 44620 944730
rect 43028 933094 43084 933103
rect 43028 933029 43084 933038
rect 42356 932650 42412 932659
rect 42356 932585 42412 932594
rect 42370 931031 42398 932585
rect 42356 931022 42412 931031
rect 42356 930957 42358 930966
rect 42410 930957 42412 930966
rect 44566 930983 44618 930989
rect 42358 930925 42410 930931
rect 44566 930925 44618 930931
rect 43124 907194 43180 907203
rect 43124 907129 43180 907138
rect 43138 887223 43166 907129
rect 43124 887214 43180 887223
rect 43124 887149 43180 887158
rect 42358 823905 42410 823911
rect 42356 823870 42358 823879
rect 42410 823870 42412 823879
rect 42356 823805 42412 823814
rect 42452 822686 42508 822695
rect 42452 822621 42508 822630
rect 42358 822277 42410 822283
rect 42356 822242 42358 822251
rect 42410 822242 42412 822251
rect 42356 822177 42412 822186
rect 42466 821913 42494 822621
rect 42454 821907 42506 821913
rect 42454 821849 42506 821855
rect 43220 821206 43276 821215
rect 43220 821141 43276 821150
rect 40340 820762 40396 820771
rect 40340 820697 40396 820706
rect 40052 820170 40108 820179
rect 40052 820105 40108 820114
rect 37460 819134 37516 819143
rect 37460 819069 37516 819078
rect 37474 817788 37502 819069
rect 41684 817950 41740 817959
rect 41684 817885 41740 817894
rect 37282 817760 37502 817788
rect 37282 802123 37310 817760
rect 40148 816766 40204 816775
rect 40148 816701 40204 816710
rect 37364 812770 37420 812779
rect 37364 812705 37420 812714
rect 37378 802271 37406 812705
rect 40162 803487 40190 816701
rect 40244 815878 40300 815887
rect 40244 815813 40300 815822
rect 40150 803481 40202 803487
rect 40150 803423 40202 803429
rect 37364 802262 37420 802271
rect 37364 802197 37420 802206
rect 37268 802114 37324 802123
rect 37268 802049 37324 802058
rect 40258 801975 40286 815813
rect 41588 815286 41644 815295
rect 41588 815221 41644 815230
rect 40244 801966 40300 801975
rect 40244 801901 40300 801910
rect 41602 800527 41630 815221
rect 41698 800601 41726 817885
rect 41972 814398 42028 814407
rect 41972 814333 42028 814342
rect 41876 813658 41932 813667
rect 41876 813593 41932 813602
rect 41780 809662 41836 809671
rect 41780 809597 41836 809606
rect 41686 800595 41738 800601
rect 41686 800537 41738 800543
rect 41590 800521 41642 800527
rect 41590 800463 41642 800469
rect 41794 800347 41822 809597
rect 41780 800338 41836 800347
rect 41780 800273 41836 800282
rect 41890 800231 41918 813593
rect 41986 802451 42014 814333
rect 42356 812326 42412 812335
rect 42356 812261 42412 812270
rect 42068 811142 42124 811151
rect 42068 811077 42124 811086
rect 41974 802445 42026 802451
rect 41974 802387 42026 802393
rect 42082 800347 42110 811077
rect 42164 808330 42220 808339
rect 42164 808265 42220 808274
rect 42068 800338 42124 800347
rect 42068 800273 42124 800282
rect 41878 800225 41930 800231
rect 41878 800167 41930 800173
rect 42178 800176 42206 808265
rect 42260 805222 42316 805231
rect 42260 805157 42262 805166
rect 42314 805157 42316 805166
rect 42262 805125 42314 805131
rect 42370 804449 42398 812261
rect 43124 810402 43180 810411
rect 43124 810337 43180 810346
rect 43028 809366 43084 809375
rect 43028 809301 43084 809310
rect 42452 807590 42508 807599
rect 42452 807525 42508 807534
rect 42358 804443 42410 804449
rect 42358 804385 42410 804391
rect 42466 804153 42494 807525
rect 42934 804443 42986 804449
rect 42934 804385 42986 804391
rect 42454 804147 42506 804153
rect 42454 804089 42506 804095
rect 42742 804147 42794 804153
rect 42742 804089 42794 804095
rect 42452 803594 42508 803603
rect 42508 803552 42590 803580
rect 42452 803529 42508 803538
rect 42454 803481 42506 803487
rect 42454 803423 42506 803429
rect 42178 800148 42302 800176
rect 42274 800051 42302 800148
rect 42260 800042 42316 800051
rect 42260 799977 42316 799986
rect 41878 799781 41930 799787
rect 41878 799723 41930 799729
rect 41890 799422 41918 799723
rect 42466 798085 42494 803423
rect 42166 798079 42218 798085
rect 42166 798021 42218 798027
rect 42454 798079 42506 798085
rect 42454 798021 42506 798027
rect 42178 797605 42206 798021
rect 42452 797970 42508 797979
rect 42452 797905 42508 797914
rect 42070 797339 42122 797345
rect 42070 797281 42122 797287
rect 42082 796980 42110 797281
rect 42166 796303 42218 796309
rect 42166 796245 42218 796251
rect 42178 795765 42206 796245
rect 42166 795045 42218 795051
rect 42166 794987 42218 794993
rect 42178 794569 42206 794987
rect 41780 794270 41836 794279
rect 41780 794205 41836 794214
rect 41794 793946 41822 794205
rect 42466 793867 42494 797905
rect 42166 793861 42218 793867
rect 42166 793803 42218 793809
rect 42454 793861 42506 793867
rect 42454 793803 42506 793809
rect 42178 793280 42206 793803
rect 42166 793195 42218 793201
rect 42166 793137 42218 793143
rect 42178 792729 42206 793137
rect 42262 792159 42314 792165
rect 42262 792101 42314 792107
rect 42166 792011 42218 792017
rect 42166 791953 42218 791959
rect 42178 791444 42206 791953
rect 41808 791430 42206 791444
rect 41794 791416 42192 791430
rect 41794 791319 41822 791416
rect 41780 791310 41836 791319
rect 41780 791245 41836 791254
rect 42164 791014 42220 791023
rect 42164 790949 42220 790958
rect 42178 790797 42206 790949
rect 42274 790260 42302 792101
rect 42454 792011 42506 792017
rect 42562 791999 42590 803552
rect 42754 795051 42782 804089
rect 42838 802445 42890 802451
rect 42838 802387 42890 802393
rect 42742 795045 42794 795051
rect 42742 794987 42794 794993
rect 42740 794862 42796 794871
rect 42740 794797 42796 794806
rect 42754 792979 42782 794797
rect 42850 793201 42878 802387
rect 42838 793195 42890 793201
rect 42838 793137 42890 793143
rect 42838 793047 42890 793053
rect 42838 792989 42890 792995
rect 42742 792973 42794 792979
rect 42742 792915 42794 792921
rect 42506 791971 42590 791999
rect 42454 791953 42506 791959
rect 42452 791902 42508 791911
rect 42452 791837 42508 791846
rect 42192 790232 42302 790260
rect 42262 790161 42314 790167
rect 42262 790103 42314 790109
rect 42166 789939 42218 789945
rect 42166 789881 42218 789887
rect 42178 789580 42206 789881
rect 42166 789495 42218 789501
rect 42166 789437 42218 789443
rect 42178 788957 42206 789437
rect 42274 788410 42302 790103
rect 42192 788382 42302 788410
rect 42166 787053 42218 787059
rect 42166 786995 42218 787001
rect 42178 786546 42206 786995
rect 42166 786461 42218 786467
rect 42166 786403 42218 786409
rect 42178 785921 42206 786403
rect 42466 785801 42494 791837
rect 42740 791754 42796 791763
rect 42740 791689 42796 791698
rect 42754 786467 42782 791689
rect 42850 790167 42878 792989
rect 42838 790161 42890 790167
rect 42838 790103 42890 790109
rect 42946 789501 42974 804385
rect 43042 801637 43070 809301
rect 43030 801631 43082 801637
rect 43030 801573 43082 801579
rect 43030 801483 43082 801489
rect 43030 801425 43082 801431
rect 43042 797345 43070 801425
rect 43030 797339 43082 797345
rect 43030 797281 43082 797287
rect 43030 797191 43082 797197
rect 43030 797133 43082 797139
rect 43042 793127 43070 797133
rect 43138 796309 43166 810337
rect 43126 796303 43178 796309
rect 43126 796245 43178 796251
rect 43126 796155 43178 796161
rect 43126 796097 43178 796103
rect 43030 793121 43082 793127
rect 43030 793063 43082 793069
rect 43030 792973 43082 792979
rect 43030 792915 43082 792921
rect 43042 789945 43070 792915
rect 43138 792165 43166 796097
rect 43126 792159 43178 792165
rect 43126 792101 43178 792107
rect 43126 792011 43178 792017
rect 43126 791953 43178 791959
rect 43030 789939 43082 789945
rect 43030 789881 43082 789887
rect 42934 789495 42986 789501
rect 42934 789437 42986 789443
rect 43138 787059 43166 791953
rect 43126 787053 43178 787059
rect 43126 786995 43178 787001
rect 42742 786461 42794 786467
rect 42742 786403 42794 786409
rect 42070 785795 42122 785801
rect 42070 785737 42122 785743
rect 42454 785795 42506 785801
rect 42454 785737 42506 785743
rect 42082 785288 42110 785737
rect 42740 780506 42796 780515
rect 42740 780441 42742 780450
rect 42794 780441 42796 780450
rect 42742 780409 42794 780415
rect 42454 779949 42506 779955
rect 42452 779914 42454 779923
rect 42506 779914 42508 779923
rect 42452 779849 42508 779858
rect 42742 778913 42794 778919
rect 42740 778878 42742 778887
rect 42794 778878 42796 778887
rect 42740 778813 42796 778822
rect 43234 777259 43262 821141
rect 43414 801631 43466 801637
rect 43414 801573 43466 801579
rect 43318 800521 43370 800527
rect 43318 800463 43370 800469
rect 43330 797197 43358 800463
rect 43318 797191 43370 797197
rect 43318 797133 43370 797139
rect 43426 796161 43454 801573
rect 43510 800595 43562 800601
rect 43510 800537 43562 800543
rect 43414 796155 43466 796161
rect 43414 796097 43466 796103
rect 43522 792017 43550 800537
rect 43510 792011 43562 792017
rect 43510 791953 43562 791959
rect 43316 777990 43372 777999
rect 43316 777925 43372 777934
rect 43220 777250 43276 777259
rect 43220 777185 43276 777194
rect 42836 774882 42892 774891
rect 42836 774817 42892 774826
rect 38996 773550 39052 773559
rect 38996 773485 39052 773494
rect 38804 772662 38860 772671
rect 38804 772597 38860 772606
rect 37364 769554 37420 769563
rect 37364 769489 37420 769498
rect 37378 758611 37406 769489
rect 38818 760239 38846 772597
rect 39010 760345 39038 773485
rect 42452 771182 42508 771191
rect 42452 771117 42508 771126
rect 41780 770442 41836 770451
rect 41780 770377 41836 770386
rect 38998 760339 39050 760345
rect 38998 760281 39050 760287
rect 38804 760230 38860 760239
rect 38804 760165 38860 760174
rect 37364 758602 37420 758611
rect 37364 758537 37420 758546
rect 41794 757015 41822 770377
rect 41876 769110 41932 769119
rect 41876 769045 41932 769054
rect 41890 757015 41918 769045
rect 41972 767926 42028 767935
rect 41972 767861 42028 767870
rect 41986 757163 42014 767861
rect 42068 765262 42124 765271
rect 42068 765197 42124 765206
rect 41974 757157 42026 757163
rect 41974 757099 42026 757105
rect 42082 757089 42110 765197
rect 42466 757311 42494 771117
rect 42740 763782 42796 763791
rect 42740 763717 42796 763726
rect 42754 762311 42782 763717
rect 42740 762302 42796 762311
rect 42740 762237 42742 762246
rect 42794 762237 42796 762246
rect 42742 762205 42794 762211
rect 42742 760339 42794 760345
rect 42742 760281 42794 760287
rect 42454 757305 42506 757311
rect 42454 757247 42506 757253
rect 42070 757083 42122 757089
rect 42070 757025 42122 757031
rect 41782 757009 41834 757015
rect 41782 756951 41834 756957
rect 41878 757009 41930 757015
rect 41878 756951 41930 756957
rect 41782 756787 41834 756793
rect 41782 756729 41834 756735
rect 41794 756245 41822 756729
rect 42754 754943 42782 760281
rect 42070 754937 42122 754943
rect 42070 754879 42122 754885
rect 42742 754937 42794 754943
rect 42742 754879 42794 754885
rect 42082 754430 42110 754879
rect 42454 754345 42506 754351
rect 42454 754287 42506 754293
rect 42166 754123 42218 754129
rect 42166 754065 42218 754071
rect 42178 753764 42206 754065
rect 42070 753087 42122 753093
rect 42070 753029 42122 753035
rect 42082 752580 42110 753029
rect 41780 751794 41836 751803
rect 41780 751729 41836 751738
rect 41794 751396 41822 751729
rect 42070 751237 42122 751243
rect 42070 751179 42122 751185
rect 42082 750730 42110 751179
rect 42166 750423 42218 750429
rect 42166 750365 42218 750371
rect 42178 750064 42206 750365
rect 42070 749979 42122 749985
rect 42070 749921 42122 749927
rect 42082 749546 42110 749921
rect 42262 748943 42314 748949
rect 42262 748885 42314 748891
rect 41780 748686 41836 748695
rect 41780 748621 41836 748630
rect 41794 748214 41822 748621
rect 41986 747363 42014 747622
rect 42164 747502 42220 747511
rect 42164 747437 42220 747446
rect 41972 747354 42028 747363
rect 41972 747289 42028 747298
rect 42178 747030 42206 747437
rect 42274 746415 42302 748885
rect 42192 746387 42302 746415
rect 42070 746131 42122 746137
rect 42070 746073 42122 746079
rect 42082 745772 42110 746073
rect 42466 745693 42494 754287
rect 42850 751951 42878 774817
rect 42932 772514 42988 772523
rect 42932 772449 42988 772458
rect 42946 754351 42974 772449
rect 43124 767778 43180 767787
rect 43124 767713 43180 767722
rect 43028 767038 43084 767047
rect 43028 766973 43084 766982
rect 43042 758144 43070 766973
rect 43138 759383 43166 767713
rect 43126 759377 43178 759383
rect 43126 759319 43178 759325
rect 43042 758116 43262 758144
rect 43030 757823 43082 757829
rect 43030 757765 43082 757771
rect 42934 754345 42986 754351
rect 42934 754287 42986 754293
rect 43042 754129 43070 757765
rect 43030 754123 43082 754129
rect 43030 754065 43082 754071
rect 43234 752372 43262 758116
rect 43138 752344 43262 752372
rect 42836 751942 42892 751951
rect 43138 751909 43166 752344
rect 43222 752273 43274 752279
rect 43222 752215 43274 752221
rect 42836 751877 42892 751886
rect 43126 751903 43178 751909
rect 43126 751845 43178 751851
rect 42934 751829 42986 751835
rect 43234 751780 43262 752215
rect 42934 751771 42986 751777
rect 42836 751646 42892 751655
rect 42836 751581 42892 751590
rect 42742 751015 42794 751021
rect 42742 750957 42794 750963
rect 42754 748949 42782 750957
rect 42742 748943 42794 748949
rect 42742 748885 42794 748891
rect 42740 746910 42796 746919
rect 42740 746845 42796 746854
rect 42166 745687 42218 745693
rect 42166 745629 42218 745635
rect 42454 745687 42506 745693
rect 42454 745629 42506 745635
rect 42178 745180 42206 745629
rect 42166 743837 42218 743843
rect 42166 743779 42218 743785
rect 42178 743365 42206 743779
rect 42070 743097 42122 743103
rect 42070 743039 42122 743045
rect 42082 742738 42110 743039
rect 42754 742659 42782 746845
rect 42850 743843 42878 751581
rect 42946 751243 42974 751771
rect 43042 751752 43262 751780
rect 42934 751237 42986 751243
rect 42934 751179 42986 751185
rect 43042 749985 43070 751752
rect 43126 751681 43178 751687
rect 43126 751623 43178 751629
rect 43138 750429 43166 751623
rect 43126 750423 43178 750429
rect 43126 750365 43178 750371
rect 43126 750275 43178 750281
rect 43126 750217 43178 750223
rect 43030 749979 43082 749985
rect 43030 749921 43082 749927
rect 42932 747206 42988 747215
rect 42932 747141 42988 747150
rect 42838 743837 42890 743843
rect 42838 743779 42890 743785
rect 42946 743103 42974 747141
rect 43138 746137 43166 750217
rect 43126 746131 43178 746137
rect 43126 746073 43178 746079
rect 42934 743097 42986 743103
rect 42934 743039 42986 743045
rect 42166 742653 42218 742659
rect 42166 742595 42218 742601
rect 42742 742653 42794 742659
rect 42742 742595 42794 742601
rect 42178 742072 42206 742595
rect 42644 737290 42700 737299
rect 42644 737225 42646 737234
rect 42698 737225 42700 737234
rect 42646 737193 42698 737199
rect 42358 736733 42410 736739
rect 42356 736698 42358 736707
rect 42410 736698 42412 736707
rect 42356 736633 42412 736642
rect 42068 735958 42124 735967
rect 42068 735893 42124 735902
rect 40148 730334 40204 730343
rect 40148 730269 40204 730278
rect 37364 726338 37420 726347
rect 37364 726273 37420 726282
rect 37378 717023 37406 726273
rect 37364 717014 37420 717023
rect 37364 716949 37420 716958
rect 40162 715945 40190 730269
rect 40244 729594 40300 729603
rect 40244 729529 40300 729538
rect 40258 716727 40286 729529
rect 41684 728854 41740 728863
rect 41684 728789 41740 728798
rect 41588 727226 41644 727235
rect 41588 727161 41644 727170
rect 40244 716718 40300 716727
rect 40244 716653 40300 716662
rect 40150 715939 40202 715945
rect 40150 715881 40202 715887
rect 41602 714095 41630 727161
rect 41698 714095 41726 728789
rect 41972 727966 42028 727975
rect 41972 727901 42028 727910
rect 41780 725894 41836 725903
rect 41780 725829 41836 725838
rect 41590 714089 41642 714095
rect 41590 714031 41642 714037
rect 41686 714089 41738 714095
rect 41686 714031 41738 714037
rect 41794 714021 41822 725829
rect 41986 716135 42014 727901
rect 42082 725903 42110 735893
rect 42356 735514 42412 735523
rect 42356 735449 42358 735458
rect 42410 735449 42412 735458
rect 42358 735417 42410 735423
rect 43220 734922 43276 734931
rect 43220 734857 43276 734866
rect 42932 731666 42988 731675
rect 42932 731601 42988 731610
rect 42068 725894 42124 725903
rect 42068 725829 42124 725838
rect 42068 724710 42124 724719
rect 42068 724645 42124 724654
rect 41972 716126 42028 716135
rect 41972 716061 42028 716070
rect 41878 715939 41930 715945
rect 41878 715881 41930 715887
rect 41782 714015 41834 714021
rect 41782 713957 41834 713963
rect 41890 713915 41918 715881
rect 42082 713915 42110 724645
rect 42164 724118 42220 724127
rect 42164 724053 42220 724062
rect 42178 722180 42206 724053
rect 42178 722152 42398 722180
rect 41876 713906 41932 713915
rect 41876 713841 41932 713850
rect 42068 713906 42124 713915
rect 42068 713841 42124 713850
rect 41782 713571 41834 713577
rect 41782 713513 41834 713519
rect 41794 713064 41822 713513
rect 41876 711686 41932 711695
rect 41876 711621 41932 711630
rect 41890 711214 41918 711621
rect 42166 710833 42218 710839
rect 42166 710775 42218 710781
rect 42178 710548 42206 710775
rect 42370 709951 42398 722152
rect 42946 711801 42974 731601
rect 43028 722194 43084 722203
rect 43028 722129 43084 722138
rect 42934 711795 42986 711801
rect 42934 711737 42986 711743
rect 42836 710798 42892 710807
rect 42836 710733 42892 710742
rect 42166 709945 42218 709951
rect 42166 709887 42218 709893
rect 42358 709945 42410 709951
rect 42358 709887 42410 709893
rect 42178 709364 42206 709887
rect 41780 708578 41836 708587
rect 41780 708513 41836 708522
rect 41794 708180 41822 708513
rect 42550 707947 42602 707953
rect 42550 707889 42602 707895
rect 42164 707838 42220 707847
rect 42164 707773 42220 707782
rect 42178 707514 42206 707773
rect 42166 707429 42218 707435
rect 42166 707371 42218 707377
rect 42178 706881 42206 707371
rect 41780 706802 41836 706811
rect 41780 706737 41836 706746
rect 41794 706330 41822 706737
rect 42164 706210 42220 706219
rect 42164 706145 42220 706154
rect 42178 705881 42206 706145
rect 42166 705875 42218 705881
rect 42166 705817 42218 705823
rect 42262 705653 42314 705659
rect 42262 705595 42314 705601
rect 41794 704739 41822 705041
rect 41780 704730 41836 704739
rect 41780 704665 41836 704674
rect 41794 704147 41822 704406
rect 41780 704138 41836 704147
rect 41780 704073 41836 704082
rect 42274 703859 42302 705595
rect 42192 703831 42302 703859
rect 42260 703694 42316 703703
rect 42260 703629 42316 703638
rect 42070 703581 42122 703587
rect 42070 703523 42122 703529
rect 42082 703222 42110 703523
rect 42166 702915 42218 702921
rect 42166 702857 42218 702863
rect 42178 702556 42206 702857
rect 42166 702323 42218 702329
rect 42166 702265 42218 702271
rect 42178 702005 42206 702265
rect 42274 700891 42302 703629
rect 42562 702329 42590 707889
rect 42850 703661 42878 710733
rect 43042 707435 43070 722129
rect 43234 711283 43262 734857
rect 43330 734043 43358 777925
rect 43414 759377 43466 759383
rect 43414 759319 43466 759325
rect 43426 753093 43454 759319
rect 43606 757305 43658 757311
rect 43606 757247 43658 757253
rect 43510 757083 43562 757089
rect 43510 757025 43562 757031
rect 43414 753087 43466 753093
rect 43414 753029 43466 753035
rect 43522 752076 43550 757025
rect 43618 752279 43646 757247
rect 43798 757157 43850 757163
rect 43798 757099 43850 757105
rect 43702 756935 43754 756941
rect 43702 756877 43754 756883
rect 43606 752273 43658 752279
rect 43606 752215 43658 752221
rect 43426 752048 43550 752076
rect 43426 751687 43454 752048
rect 43714 751928 43742 756877
rect 43522 751900 43742 751928
rect 43414 751681 43466 751687
rect 43414 751623 43466 751629
rect 43522 750281 43550 751900
rect 43810 751780 43838 757099
rect 43618 751752 43838 751780
rect 43618 751021 43646 751752
rect 43606 751015 43658 751021
rect 43606 750957 43658 750963
rect 43510 750275 43562 750281
rect 43510 750217 43562 750223
rect 43316 734034 43372 734043
rect 43316 733969 43372 733978
rect 43316 720566 43372 720575
rect 43316 720501 43372 720510
rect 43330 719095 43358 720501
rect 43316 719086 43372 719095
rect 43316 719021 43372 719030
rect 43330 717277 43358 719021
rect 43318 717271 43370 717277
rect 43318 717213 43370 717219
rect 43510 714089 43562 714095
rect 43510 714031 43562 714037
rect 43522 711524 43550 714031
rect 43606 714015 43658 714021
rect 43606 713957 43658 713963
rect 43426 711496 43550 711524
rect 43222 711277 43274 711283
rect 43222 711219 43274 711225
rect 43426 707953 43454 711496
rect 43510 711425 43562 711431
rect 43510 711367 43562 711373
rect 43414 707947 43466 707953
rect 43414 707889 43466 707895
rect 43030 707429 43082 707435
rect 43030 707371 43082 707377
rect 43030 707281 43082 707287
rect 43030 707223 43082 707229
rect 42934 706467 42986 706473
rect 42934 706409 42986 706415
rect 42838 703655 42890 703661
rect 42838 703597 42890 703603
rect 42836 703546 42892 703555
rect 42836 703481 42892 703490
rect 42550 702323 42602 702329
rect 42550 702265 42602 702271
rect 42260 700882 42316 700891
rect 42260 700817 42316 700826
rect 42070 700621 42122 700627
rect 42070 700563 42122 700569
rect 42260 700586 42316 700595
rect 42082 700188 42110 700563
rect 42260 700521 42316 700530
rect 42166 700103 42218 700109
rect 42166 700045 42218 700051
rect 42178 699522 42206 700045
rect 42274 699388 42302 700521
rect 42850 700109 42878 703481
rect 42946 700627 42974 706409
rect 43042 702921 43070 707223
rect 43522 706473 43550 711367
rect 43618 707287 43646 713957
rect 43702 711277 43754 711283
rect 43702 711219 43754 711225
rect 43606 707281 43658 707287
rect 43606 707223 43658 707229
rect 43510 706467 43562 706473
rect 43510 706409 43562 706415
rect 43030 702915 43082 702921
rect 43030 702857 43082 702863
rect 43714 701312 43742 711219
rect 43234 701284 43742 701312
rect 42934 700621 42986 700627
rect 42934 700563 42986 700569
rect 42838 700103 42890 700109
rect 42838 700045 42890 700051
rect 42358 699881 42410 699887
rect 42358 699823 42410 699829
rect 42178 699360 42302 699388
rect 42178 698856 42206 699360
rect 42370 693491 42398 699823
rect 42644 694074 42700 694083
rect 42644 694009 42646 694018
rect 42698 694009 42700 694018
rect 42646 693977 42698 693983
rect 42356 693482 42412 693491
rect 42356 693417 42412 693426
rect 41396 692742 41452 692751
rect 41396 692677 41452 692686
rect 40244 687118 40300 687127
rect 40244 687053 40300 687062
rect 40258 672433 40286 687053
rect 41300 680014 41356 680023
rect 41300 679949 41356 679958
rect 40246 672427 40298 672433
rect 40246 672369 40298 672375
rect 41314 670953 41342 679949
rect 41410 670995 41438 692677
rect 42646 692481 42698 692487
rect 42644 692446 42646 692455
rect 42698 692446 42700 692455
rect 42644 692381 42700 692390
rect 43234 690827 43262 701284
rect 43508 691706 43564 691715
rect 43508 691641 43564 691650
rect 43220 690818 43276 690827
rect 43220 690753 43276 690762
rect 41876 688302 41932 688311
rect 41876 688237 41932 688246
rect 41780 684010 41836 684019
rect 41780 683945 41836 683954
rect 41396 670986 41452 670995
rect 41302 670947 41354 670953
rect 41396 670921 41452 670930
rect 41302 670889 41354 670895
rect 41794 670657 41822 683945
rect 41890 674579 41918 688237
rect 42740 686082 42796 686091
rect 42740 686017 42796 686026
rect 42068 684898 42124 684907
rect 42068 684833 42124 684842
rect 41972 679570 42028 679579
rect 41972 679505 42028 679514
rect 41878 674573 41930 674579
rect 41878 674515 41930 674521
rect 41878 672427 41930 672433
rect 41878 672369 41930 672375
rect 41890 670657 41918 672369
rect 41986 670731 42014 679505
rect 42082 671989 42110 684833
rect 42164 682678 42220 682687
rect 42164 682613 42220 682622
rect 42070 671983 42122 671989
rect 42070 671925 42122 671931
rect 41974 670725 42026 670731
rect 42178 670699 42206 682613
rect 42260 681494 42316 681503
rect 42260 681429 42316 681438
rect 42274 670805 42302 681429
rect 42356 677202 42412 677211
rect 42356 677137 42412 677146
rect 42370 675731 42398 677137
rect 42754 676355 42782 686017
rect 43124 678238 43180 678247
rect 43124 678173 43180 678182
rect 42742 676349 42794 676355
rect 42742 676291 42794 676297
rect 42646 676053 42698 676059
rect 42646 675995 42698 676001
rect 42356 675722 42412 675731
rect 42356 675657 42358 675666
rect 42410 675657 42412 675666
rect 42358 675625 42410 675631
rect 42454 671983 42506 671989
rect 42454 671925 42506 671931
rect 42262 670799 42314 670805
rect 42262 670741 42314 670747
rect 41974 670667 42026 670673
rect 42164 670690 42220 670699
rect 41782 670651 41834 670657
rect 41782 670593 41834 670599
rect 41878 670651 41930 670657
rect 42164 670625 42220 670634
rect 41878 670593 41930 670599
rect 41782 670355 41834 670361
rect 41782 670297 41834 670303
rect 41794 669848 41822 670297
rect 42466 669367 42494 671925
rect 42658 670995 42686 675995
rect 43138 674672 43166 678173
rect 43042 674644 43166 674672
rect 42644 670986 42700 670995
rect 42644 670921 42700 670930
rect 42934 670947 42986 670953
rect 42934 670889 42986 670895
rect 42946 670676 42974 670889
rect 43042 670824 43070 674644
rect 43126 674573 43178 674579
rect 43126 674515 43178 674521
rect 43138 670972 43166 674515
rect 43318 673833 43370 673839
rect 43318 673775 43370 673781
rect 43138 670953 43262 670972
rect 43138 670947 43274 670953
rect 43138 670944 43222 670947
rect 43222 670889 43274 670895
rect 43042 670796 43262 670824
rect 43126 670725 43178 670731
rect 42946 670648 43070 670676
rect 43126 670667 43178 670673
rect 42934 670577 42986 670583
rect 42934 670519 42986 670525
rect 42452 669358 42508 669367
rect 42452 669293 42508 669302
rect 42548 668914 42604 668923
rect 42604 668872 42686 668900
rect 42548 668849 42604 668858
rect 42548 668766 42604 668775
rect 42548 668701 42604 668710
rect 42166 668579 42218 668585
rect 42166 668521 42218 668527
rect 42178 667998 42206 668521
rect 42166 667913 42218 667919
rect 42166 667855 42218 667861
rect 42178 667361 42206 667855
rect 41780 666694 41836 666703
rect 41780 666629 41836 666638
rect 41794 666148 41822 666629
rect 42166 665397 42218 665403
rect 42166 665339 42218 665345
rect 42178 664964 42206 665339
rect 42166 664879 42218 664885
rect 42166 664821 42218 664827
rect 42178 664298 42206 664821
rect 42562 663997 42590 668701
rect 42070 663991 42122 663997
rect 42070 663933 42122 663939
rect 42550 663991 42602 663997
rect 42550 663933 42602 663939
rect 42082 663706 42110 663933
rect 42658 663424 42686 668872
rect 42946 668585 42974 670519
rect 42934 668579 42986 668585
rect 42934 668521 42986 668527
rect 42934 668431 42986 668437
rect 42934 668373 42986 668379
rect 42836 666546 42892 666555
rect 42836 666481 42892 666490
rect 42562 663405 42686 663424
rect 42166 663399 42218 663405
rect 42166 663341 42218 663347
rect 42550 663399 42686 663405
rect 42602 663396 42686 663399
rect 42550 663341 42602 663347
rect 42178 663114 42206 663341
rect 42262 662437 42314 662443
rect 42262 662379 42314 662385
rect 42178 661523 42206 661856
rect 42164 661514 42220 661523
rect 42164 661449 42220 661458
rect 41890 660783 41918 661190
rect 42070 661105 42122 661111
rect 42070 661047 42122 661053
rect 41876 660774 41932 660783
rect 41876 660709 41932 660718
rect 42082 660672 42110 661047
rect 42274 660020 42302 662379
rect 42192 659992 42302 660020
rect 42850 659927 42878 666481
rect 42946 665403 42974 668373
rect 42934 665397 42986 665403
rect 42934 665339 42986 665345
rect 42934 665249 42986 665255
rect 42934 665191 42986 665197
rect 42946 662443 42974 665191
rect 43042 664885 43070 670648
rect 43030 664879 43082 664885
rect 43030 664821 43082 664827
rect 43028 664770 43084 664779
rect 43028 664705 43084 664714
rect 42934 662437 42986 662443
rect 42934 662379 42986 662385
rect 42934 662289 42986 662295
rect 42934 662231 42986 662237
rect 42166 659921 42218 659927
rect 42166 659863 42218 659869
rect 42838 659921 42890 659927
rect 42838 659863 42890 659869
rect 42178 659340 42206 659863
rect 42070 659107 42122 659113
rect 42070 659049 42122 659055
rect 42082 658822 42110 659049
rect 42178 656893 42206 656972
rect 42946 656893 42974 662231
rect 43042 659113 43070 664705
rect 43138 661111 43166 670667
rect 43234 668437 43262 670796
rect 43222 668431 43274 668437
rect 43222 668373 43274 668379
rect 43330 667919 43358 673775
rect 43414 670799 43466 670805
rect 43414 670741 43466 670747
rect 43318 667913 43370 667919
rect 43318 667855 43370 667861
rect 43426 665255 43454 670741
rect 43414 665249 43466 665255
rect 43414 665191 43466 665197
rect 43126 661105 43178 661111
rect 43126 661047 43178 661053
rect 43030 659107 43082 659113
rect 43030 659049 43082 659055
rect 42166 656887 42218 656893
rect 42166 656829 42218 656835
rect 42934 656887 42986 656893
rect 42934 656829 42986 656835
rect 41780 656778 41836 656787
rect 41780 656713 41836 656722
rect 42838 656739 42890 656745
rect 41794 656306 41822 656713
rect 42838 656681 42890 656687
rect 41780 656186 41836 656195
rect 41780 656121 41836 656130
rect 41794 655677 41822 656121
rect 42850 650867 42878 656681
rect 42836 650858 42892 650867
rect 42836 650793 42892 650802
rect 42452 649822 42508 649831
rect 42452 649757 42454 649766
rect 42506 649757 42508 649766
rect 42454 649725 42506 649731
rect 42454 649561 42506 649567
rect 42452 649526 42454 649535
rect 42506 649526 42508 649535
rect 42452 649461 42508 649470
rect 43220 648490 43276 648499
rect 43220 648425 43276 648434
rect 43124 645382 43180 645391
rect 43124 645317 43180 645326
rect 40052 643902 40108 643911
rect 40052 643837 40108 643846
rect 40066 627885 40094 643837
rect 41876 642422 41932 642431
rect 41876 642357 41932 642366
rect 41780 640794 41836 640803
rect 41780 640729 41836 640738
rect 41492 638426 41548 638435
rect 41492 638361 41548 638370
rect 40054 627879 40106 627885
rect 40054 627821 40106 627827
rect 41506 627737 41534 638361
rect 41494 627731 41546 627737
rect 41494 627673 41546 627679
rect 41794 627441 41822 640729
rect 41890 627483 41918 642357
rect 42164 641682 42220 641691
rect 42164 641617 42220 641626
rect 41972 639462 42028 639471
rect 41972 639397 42028 639406
rect 41876 627474 41932 627483
rect 41782 627435 41834 627441
rect 41986 627441 42014 639397
rect 42068 636798 42124 636807
rect 42068 636733 42124 636742
rect 42082 627441 42110 636733
rect 42178 627483 42206 641617
rect 43028 636650 43084 636659
rect 43028 636585 43084 636594
rect 42644 635762 42700 635771
rect 42644 635697 42700 635706
rect 42452 632506 42508 632515
rect 42452 632441 42454 632450
rect 42506 632441 42508 632450
rect 42454 632409 42506 632415
rect 42454 627953 42506 627959
rect 42454 627895 42506 627901
rect 42164 627474 42220 627483
rect 41876 627409 41932 627418
rect 41974 627435 42026 627441
rect 41782 627377 41834 627383
rect 41974 627377 42026 627383
rect 42070 627435 42122 627441
rect 42164 627409 42220 627418
rect 42070 627377 42122 627383
rect 41782 627213 41834 627219
rect 41782 627155 41834 627161
rect 41794 626632 41822 627155
rect 42166 625363 42218 625369
rect 42166 625305 42218 625311
rect 42178 624782 42206 625305
rect 42466 624703 42494 627895
rect 42658 627663 42686 635697
rect 42932 635022 42988 635031
rect 42932 634957 42988 634966
rect 42946 628052 42974 634957
rect 43042 628200 43070 636585
rect 43138 632177 43166 645317
rect 43126 632171 43178 632177
rect 43126 632113 43178 632119
rect 43042 628172 43166 628200
rect 42946 628024 43070 628052
rect 42934 627879 42986 627885
rect 42934 627821 42986 627827
rect 42646 627657 42698 627663
rect 42646 627599 42698 627605
rect 42946 625369 42974 627821
rect 43042 627589 43070 628024
rect 43138 627927 43166 628172
rect 43124 627918 43180 627927
rect 43124 627853 43180 627862
rect 43126 627731 43178 627737
rect 43126 627673 43178 627679
rect 43030 627583 43082 627589
rect 43030 627525 43082 627531
rect 43030 627435 43082 627441
rect 43030 627377 43082 627383
rect 42934 625363 42986 625369
rect 42934 625305 42986 625311
rect 42934 625215 42986 625221
rect 42934 625157 42986 625163
rect 42166 624697 42218 624703
rect 42166 624639 42218 624645
rect 42454 624697 42506 624703
rect 42454 624639 42506 624645
rect 42178 624161 42206 624639
rect 42452 623922 42508 623931
rect 42370 623880 42452 623908
rect 42164 623478 42220 623487
rect 42164 623413 42220 623422
rect 42178 622965 42206 623413
rect 42166 622255 42218 622261
rect 42166 622197 42218 622203
rect 42178 621748 42206 622197
rect 42166 621663 42218 621669
rect 42166 621605 42218 621611
rect 42178 621125 42206 621605
rect 42070 620923 42122 620929
rect 42070 620865 42122 620871
rect 42082 620490 42110 620865
rect 42068 620222 42124 620231
rect 42068 620157 42124 620166
rect 42082 619929 42110 620157
rect 42370 618654 42398 623880
rect 42452 623857 42508 623866
rect 42454 623809 42506 623815
rect 42454 623751 42506 623757
rect 42466 623501 42494 623751
rect 42466 623473 42590 623501
rect 42452 623330 42508 623339
rect 42452 623265 42508 623274
rect 42000 618640 42398 618654
rect 41986 618626 42398 618640
rect 41986 618455 42014 618626
rect 41972 618446 42028 618455
rect 41972 618381 42028 618390
rect 41794 617863 41822 617974
rect 41780 617854 41836 617863
rect 41780 617789 41836 617798
rect 42070 617667 42122 617673
rect 42070 617609 42122 617615
rect 42082 617456 42110 617609
rect 42166 617371 42218 617377
rect 42166 617313 42218 617319
rect 42178 616790 42206 617313
rect 42166 616705 42218 616711
rect 42166 616647 42218 616653
rect 42178 616157 42206 616647
rect 42466 616045 42494 623265
rect 42166 616039 42218 616045
rect 42166 615981 42218 615987
rect 42454 616039 42506 616045
rect 42454 615981 42506 615987
rect 42178 615606 42206 615981
rect 42562 614140 42590 623473
rect 42946 620929 42974 625157
rect 43042 621669 43070 627377
rect 43030 621663 43082 621669
rect 43030 621605 43082 621611
rect 43030 621515 43082 621521
rect 43030 621457 43082 621463
rect 42934 620923 42986 620929
rect 42934 620865 42986 620871
rect 42932 620814 42988 620823
rect 42932 620749 42988 620758
rect 42740 618298 42796 618307
rect 42740 618233 42796 618242
rect 42466 614112 42590 614140
rect 42466 614047 42494 614112
rect 42166 614041 42218 614047
rect 42166 613983 42218 613989
rect 42454 614041 42506 614047
rect 42454 613983 42506 613989
rect 42178 613756 42206 613983
rect 42754 613677 42782 618233
rect 42836 618150 42892 618159
rect 42836 618085 42892 618094
rect 42166 613671 42218 613677
rect 42166 613613 42218 613619
rect 42742 613671 42794 613677
rect 42742 613613 42794 613619
rect 42178 613121 42206 613613
rect 42454 613523 42506 613529
rect 42454 613465 42506 613471
rect 42070 612857 42122 612863
rect 42070 612799 42122 612805
rect 42082 612498 42110 612799
rect 42466 606319 42494 613465
rect 42850 612863 42878 618085
rect 42946 617673 42974 620749
rect 42934 617667 42986 617673
rect 42934 617609 42986 617615
rect 43042 616711 43070 621457
rect 43138 617377 43166 627673
rect 43126 617371 43178 617377
rect 43126 617313 43178 617319
rect 43030 616705 43082 616711
rect 43030 616647 43082 616653
rect 42838 612857 42890 612863
rect 42838 612799 42890 612805
rect 42742 607751 42794 607757
rect 42740 607716 42742 607725
rect 42794 607716 42796 607725
rect 42740 607651 42796 607660
rect 42740 606902 42796 606911
rect 42740 606837 42742 606846
rect 42794 606837 42796 606846
rect 42742 606805 42794 606811
rect 42452 606310 42508 606319
rect 42452 606245 42508 606254
rect 43234 604691 43262 648425
rect 43522 647611 43550 691641
rect 43606 670947 43658 670953
rect 43606 670889 43658 670895
rect 43618 662295 43646 670889
rect 43606 662289 43658 662295
rect 43606 662231 43658 662237
rect 43508 647602 43564 647611
rect 43508 647537 43564 647546
rect 43796 647010 43852 647019
rect 43796 646945 43852 646954
rect 43604 646122 43660 646131
rect 43604 646057 43660 646066
rect 43318 627657 43370 627663
rect 43318 627599 43370 627605
rect 43330 625221 43358 627599
rect 43414 627583 43466 627589
rect 43414 627525 43466 627531
rect 43318 625215 43370 625221
rect 43318 625157 43370 625163
rect 43426 622261 43454 627525
rect 43510 627361 43562 627367
rect 43510 627303 43562 627309
rect 43414 622255 43466 622261
rect 43414 622197 43466 622203
rect 43522 621521 43550 627303
rect 43510 621515 43562 621521
rect 43510 621457 43562 621463
rect 43508 605274 43564 605283
rect 43508 605209 43564 605218
rect 43220 604682 43276 604691
rect 43220 604617 43276 604626
rect 43412 603794 43468 603803
rect 43412 603729 43468 603738
rect 43124 602166 43180 602175
rect 43124 602101 43180 602110
rect 40052 600686 40108 600695
rect 40052 600621 40108 600630
rect 40066 586001 40094 600621
rect 43028 599650 43084 599659
rect 43028 599585 43084 599594
rect 41876 598466 41932 598475
rect 41876 598401 41932 598410
rect 41780 597578 41836 597587
rect 41780 597513 41836 597522
rect 40054 585995 40106 586001
rect 40054 585937 40106 585943
rect 41794 584225 41822 597513
rect 41890 584267 41918 598401
rect 42068 596246 42124 596255
rect 42068 596181 42124 596190
rect 41972 595210 42028 595219
rect 41972 595145 42028 595154
rect 41986 584299 42014 595145
rect 41974 584293 42026 584299
rect 41876 584258 41932 584267
rect 41782 584219 41834 584225
rect 42082 584267 42110 596181
rect 42836 594914 42892 594923
rect 42836 594849 42892 594858
rect 42164 593730 42220 593739
rect 42164 593665 42220 593674
rect 41974 584235 42026 584241
rect 42068 584258 42124 584267
rect 41876 584193 41932 584202
rect 42178 584225 42206 593665
rect 42548 593582 42604 593591
rect 42604 593540 42686 593568
rect 42548 593517 42604 593526
rect 42548 592398 42604 592407
rect 42548 592333 42604 592342
rect 42452 590622 42508 590631
rect 42452 590557 42508 590566
rect 42466 589299 42494 590557
rect 42452 589290 42508 589299
rect 42452 589225 42454 589234
rect 42506 589225 42508 589234
rect 42454 589193 42506 589199
rect 42454 585995 42506 586001
rect 42454 585937 42506 585943
rect 42466 584563 42494 585937
rect 42562 584817 42590 592333
rect 42550 584811 42602 584817
rect 42550 584753 42602 584759
rect 42548 584702 42604 584711
rect 42658 584688 42686 593540
rect 42850 585132 42878 594849
rect 42932 591806 42988 591815
rect 42932 591741 42988 591750
rect 42946 585280 42974 591741
rect 43042 585451 43070 599585
rect 43028 585442 43084 585451
rect 43138 585409 43166 602101
rect 43028 585377 43084 585386
rect 43126 585403 43178 585409
rect 43126 585345 43178 585351
rect 42946 585252 43166 585280
rect 42850 585104 43070 585132
rect 42604 584660 42686 584688
rect 42838 584737 42890 584743
rect 42838 584679 42890 584685
rect 42548 584637 42604 584646
rect 42452 584554 42508 584563
rect 42452 584489 42508 584498
rect 42452 584258 42508 584267
rect 42068 584193 42124 584202
rect 42166 584219 42218 584225
rect 41782 584161 41834 584167
rect 42452 584193 42508 584202
rect 42166 584161 42218 584167
rect 41782 583997 41834 584003
rect 41782 583939 41834 583945
rect 41794 583445 41822 583939
rect 42466 582153 42494 584193
rect 42166 582147 42218 582153
rect 42166 582089 42218 582095
rect 42454 582147 42506 582153
rect 42454 582089 42506 582095
rect 42178 581605 42206 582089
rect 42850 581487 42878 584679
rect 42934 584219 42986 584225
rect 42934 584161 42986 584167
rect 42070 581481 42122 581487
rect 42070 581423 42122 581429
rect 42838 581481 42890 581487
rect 42838 581423 42890 581429
rect 42082 580974 42110 581423
rect 42838 581333 42890 581339
rect 42838 581275 42890 581281
rect 42070 580297 42122 580303
rect 42070 580239 42122 580245
rect 42082 579790 42110 580239
rect 42166 579039 42218 579045
rect 42166 578981 42218 578987
rect 42178 578569 42206 578981
rect 42070 578447 42122 578453
rect 42070 578389 42122 578395
rect 42082 577940 42110 578389
rect 42166 577707 42218 577713
rect 42166 577649 42218 577655
rect 42178 577274 42206 577649
rect 41780 577154 41836 577163
rect 41780 577089 41836 577098
rect 41794 576756 41822 577089
rect 42260 575970 42316 575979
rect 42260 575905 42316 575914
rect 41986 575239 42014 575424
rect 41972 575230 42028 575239
rect 41972 575165 42028 575174
rect 41794 574647 41822 574797
rect 41780 574638 41836 574647
rect 41780 574573 41836 574582
rect 42274 574254 42302 575905
rect 42192 574226 42302 574254
rect 42850 574161 42878 581275
rect 42946 578453 42974 584161
rect 43042 580303 43070 585104
rect 43138 584984 43166 585252
rect 43138 584956 43358 584984
rect 43126 584811 43178 584817
rect 43126 584753 43178 584759
rect 43030 580297 43082 580303
rect 43030 580239 43082 580245
rect 43028 580114 43084 580123
rect 43028 580049 43084 580058
rect 42934 578447 42986 578453
rect 42934 578389 42986 578395
rect 42932 578338 42988 578347
rect 42932 578273 42988 578282
rect 42166 574155 42218 574161
rect 42166 574097 42218 574103
rect 42838 574155 42890 574161
rect 42838 574097 42890 574103
rect 42178 573574 42206 574097
rect 42452 574046 42508 574055
rect 42452 573981 42508 573990
rect 42070 573267 42122 573273
rect 42070 573209 42122 573215
rect 42082 572982 42110 573209
rect 42166 572675 42218 572681
rect 42166 572617 42218 572623
rect 42178 572390 42206 572617
rect 42166 571047 42218 571053
rect 42166 570989 42218 570995
rect 42178 570540 42206 570989
rect 42466 570461 42494 573981
rect 42836 573898 42892 573907
rect 42836 573833 42892 573842
rect 42850 572552 42878 573833
rect 42946 572681 42974 578273
rect 43042 573273 43070 580049
rect 43138 577713 43166 584753
rect 43222 584293 43274 584299
rect 43222 584235 43274 584241
rect 43234 581339 43262 584235
rect 43222 581333 43274 581339
rect 43222 581275 43274 581281
rect 43330 579045 43358 584956
rect 43318 579039 43370 579045
rect 43318 578981 43370 578987
rect 43126 577707 43178 577713
rect 43126 577649 43178 577655
rect 43126 577559 43178 577565
rect 43126 577501 43178 577507
rect 43030 573267 43082 573273
rect 43030 573209 43082 573215
rect 42934 572675 42986 572681
rect 42934 572617 42986 572623
rect 42850 572524 42974 572552
rect 42070 570455 42122 570461
rect 42070 570397 42122 570403
rect 42454 570455 42506 570461
rect 42454 570397 42506 570403
rect 42082 569948 42110 570397
rect 42358 570307 42410 570313
rect 42358 570249 42410 570255
rect 42070 569715 42122 569721
rect 42070 569657 42122 569663
rect 42082 569282 42110 569657
rect 34484 564722 34540 564731
rect 34484 564657 34540 564666
rect 34498 564541 34526 564657
rect 34486 564535 34538 564541
rect 34486 564477 34538 564483
rect 42370 563103 42398 570249
rect 42946 569721 42974 572524
rect 43138 571053 43166 577501
rect 43126 571047 43178 571053
rect 43126 570989 43178 570995
rect 42934 569715 42986 569721
rect 42934 569657 42986 569663
rect 42452 563538 42508 563547
rect 42452 563473 42454 563482
rect 42506 563473 42508 563482
rect 42454 563441 42506 563447
rect 42356 563094 42412 563103
rect 42356 563029 42412 563038
rect 43220 562058 43276 562067
rect 43220 561993 43276 562002
rect 41972 558654 42028 558663
rect 41972 558589 42028 558598
rect 40052 557470 40108 557479
rect 40052 557405 40108 557414
rect 37364 553622 37420 553631
rect 37364 553557 37420 553566
rect 37378 542975 37406 553557
rect 40066 544339 40094 557405
rect 40148 556730 40204 556739
rect 40148 556665 40204 556674
rect 40054 544333 40106 544339
rect 40162 544307 40190 556665
rect 41876 555990 41932 555999
rect 41876 555925 41932 555934
rect 41684 555250 41740 555259
rect 41684 555185 41740 555194
rect 40054 544275 40106 544281
rect 40148 544298 40204 544307
rect 40148 544233 40204 544242
rect 37364 542966 37420 542975
rect 37364 542901 37420 542910
rect 41698 541347 41726 555185
rect 41780 554362 41836 554371
rect 41780 554297 41836 554306
rect 41684 541338 41740 541347
rect 41684 541273 41740 541282
rect 41794 541009 41822 554297
rect 41890 541199 41918 555925
rect 41876 541190 41932 541199
rect 41876 541125 41932 541134
rect 41986 541083 42014 558589
rect 42068 553030 42124 553039
rect 42068 552965 42124 552974
rect 41974 541077 42026 541083
rect 42082 541051 42110 552965
rect 42356 551994 42412 552003
rect 42356 551929 42412 551938
rect 42164 550070 42220 550079
rect 42164 550005 42220 550014
rect 41974 541019 42026 541025
rect 42068 541042 42124 541051
rect 41782 541003 41834 541009
rect 42178 541009 42206 550005
rect 42370 545597 42398 551929
rect 43028 551698 43084 551707
rect 43028 551633 43084 551642
rect 42932 551106 42988 551115
rect 42932 551041 42988 551050
rect 42836 548590 42892 548599
rect 42836 548525 42892 548534
rect 42644 546296 42700 546305
rect 42644 546231 42646 546240
rect 42698 546231 42700 546240
rect 42646 546199 42698 546205
rect 42358 545591 42410 545597
rect 42358 545533 42410 545539
rect 42646 545591 42698 545597
rect 42646 545533 42698 545539
rect 42068 540977 42124 540986
rect 42166 541003 42218 541009
rect 41782 540945 41834 540951
rect 42166 540945 42218 540951
rect 41782 540781 41834 540787
rect 41782 540723 41834 540729
rect 41794 540245 41822 540723
rect 42070 538931 42122 538937
rect 42070 538873 42122 538879
rect 42082 538424 42110 538873
rect 42166 538191 42218 538197
rect 42166 538133 42218 538139
rect 42178 537758 42206 538133
rect 42070 537081 42122 537087
rect 42070 537023 42122 537029
rect 42082 536574 42110 537023
rect 42070 535823 42122 535829
rect 42070 535765 42122 535771
rect 42082 535390 42110 535765
rect 42166 535083 42218 535089
rect 42166 535025 42218 535031
rect 42178 534724 42206 535025
rect 42166 534491 42218 534497
rect 42166 534433 42218 534439
rect 42178 534058 42206 534433
rect 42070 533973 42122 533979
rect 42070 533915 42122 533921
rect 42082 533540 42110 533915
rect 42658 532869 42686 545533
rect 42850 545005 42878 548525
rect 42838 544999 42890 545005
rect 42838 544941 42890 544947
rect 42946 544876 42974 551041
rect 42754 544848 42974 544876
rect 42754 535089 42782 544848
rect 42838 544629 42890 544635
rect 42838 544571 42890 544577
rect 42850 535829 42878 544571
rect 42934 544333 42986 544339
rect 42934 544275 42986 544281
rect 42946 540121 42974 544275
rect 42934 540115 42986 540121
rect 42934 540057 42986 540063
rect 43042 539992 43070 551633
rect 43124 549330 43180 549339
rect 43124 549265 43180 549274
rect 42946 539964 43070 539992
rect 42946 537087 42974 539964
rect 43030 539893 43082 539899
rect 43030 539835 43082 539841
rect 43042 538937 43070 539835
rect 43030 538931 43082 538937
rect 43030 538873 43082 538879
rect 43028 538822 43084 538831
rect 43028 538757 43084 538766
rect 42934 537081 42986 537087
rect 42934 537023 42986 537029
rect 42932 536898 42988 536907
rect 42932 536833 42988 536842
rect 42838 535823 42890 535829
rect 42838 535765 42890 535771
rect 42836 535714 42892 535723
rect 42836 535649 42892 535658
rect 42742 535083 42794 535089
rect 42742 535025 42794 535031
rect 42262 532863 42314 532869
rect 42262 532805 42314 532811
rect 42646 532863 42698 532869
rect 42646 532805 42698 532811
rect 41890 532023 41918 532241
rect 41876 532014 41932 532023
rect 41876 531949 41932 531958
rect 41794 531283 41822 531616
rect 42166 531383 42218 531389
rect 42166 531325 42218 531331
rect 41780 531274 41836 531283
rect 41780 531209 41836 531218
rect 42178 531024 42206 531325
rect 42274 530415 42302 532805
rect 42740 532606 42796 532615
rect 42740 532541 42796 532550
rect 42644 532310 42700 532319
rect 42644 532245 42700 532254
rect 42192 530387 42302 530415
rect 42262 530347 42314 530353
rect 42262 530289 42314 530295
rect 42070 530199 42122 530205
rect 42070 530141 42122 530147
rect 42082 529766 42110 530141
rect 42274 529219 42302 530289
rect 42192 529191 42302 529219
rect 42166 527683 42218 527689
rect 42166 527625 42218 527631
rect 42178 527365 42206 527625
rect 42070 527239 42122 527245
rect 42070 527181 42122 527187
rect 42082 526732 42110 527181
rect 42358 527091 42410 527097
rect 42358 527033 42410 527039
rect 42166 526647 42218 526653
rect 42166 526589 42218 526595
rect 42178 526066 42206 526589
rect 42370 435527 42398 527033
rect 42658 526653 42686 532245
rect 42754 527245 42782 532541
rect 42850 530205 42878 535649
rect 42946 530353 42974 536833
rect 43042 533979 43070 538757
rect 43138 534497 43166 549265
rect 43234 534497 43262 561993
rect 43426 560587 43454 603729
rect 43522 561623 43550 605209
rect 43618 602915 43646 646057
rect 43702 632171 43754 632177
rect 43702 632113 43754 632119
rect 43714 623815 43742 632113
rect 43702 623809 43754 623815
rect 43702 623751 43754 623757
rect 43810 603803 43838 646945
rect 43796 603794 43852 603803
rect 43796 603729 43852 603738
rect 43604 602906 43660 602915
rect 43604 602841 43660 602850
rect 43508 561614 43564 561623
rect 43508 561549 43564 561558
rect 43412 560578 43468 560587
rect 43412 560513 43468 560522
rect 43318 541003 43370 541009
rect 43318 540945 43370 540951
rect 43126 534491 43178 534497
rect 43126 534433 43178 534439
rect 43222 534491 43274 534497
rect 43222 534433 43274 534439
rect 43330 534368 43358 540945
rect 43138 534340 43358 534368
rect 43030 533973 43082 533979
rect 43030 533915 43082 533921
rect 43030 533825 43082 533831
rect 43030 533767 43082 533773
rect 42934 530347 42986 530353
rect 42934 530289 42986 530295
rect 42838 530199 42890 530205
rect 42838 530141 42890 530147
rect 43042 527689 43070 533767
rect 43138 531389 43166 534340
rect 43222 534269 43274 534275
rect 43222 534211 43274 534217
rect 43126 531383 43178 531389
rect 43126 531325 43178 531331
rect 43030 527683 43082 527689
rect 43030 527625 43082 527631
rect 42742 527239 42794 527245
rect 42742 527181 42794 527187
rect 42646 526647 42698 526653
rect 42646 526589 42698 526595
rect 42646 436959 42698 436965
rect 42644 436924 42646 436933
rect 42698 436924 42700 436933
rect 42644 436859 42700 436868
rect 42646 436145 42698 436151
rect 42644 436110 42646 436119
rect 42698 436110 42700 436119
rect 42644 436045 42700 436054
rect 42356 435518 42412 435527
rect 42356 435453 42412 435462
rect 43234 433603 43262 534211
rect 43220 433594 43276 433603
rect 43220 433529 43276 433538
rect 43426 433011 43454 560513
rect 43618 559847 43646 602841
rect 43702 585403 43754 585409
rect 43702 585345 43754 585351
rect 43714 577565 43742 585345
rect 43702 577559 43754 577565
rect 43702 577501 43754 577507
rect 43604 559838 43660 559847
rect 43604 559773 43660 559782
rect 43510 541077 43562 541083
rect 43510 541019 43562 541025
rect 43522 533831 43550 541019
rect 43510 533825 43562 533831
rect 43510 533767 43562 533773
rect 43508 434482 43564 434491
rect 43508 434417 43564 434426
rect 43412 433002 43468 433011
rect 43412 432937 43468 432946
rect 42164 429894 42220 429903
rect 42164 429829 42220 429838
rect 41780 426786 41836 426795
rect 41780 426721 41836 426730
rect 37364 424418 37420 424427
rect 37364 424353 37420 424362
rect 37268 422050 37324 422059
rect 37268 421985 37324 421994
rect 37282 414765 37310 421985
rect 37378 416985 37406 424353
rect 40148 423234 40204 423243
rect 40148 423169 40204 423178
rect 37366 416979 37418 416985
rect 37366 416921 37418 416927
rect 40162 416245 40190 423169
rect 40244 420570 40300 420579
rect 40244 420505 40300 420514
rect 40150 416239 40202 416245
rect 40150 416181 40202 416187
rect 40258 414839 40286 420505
rect 40246 414833 40298 414839
rect 40246 414775 40298 414781
rect 37270 414759 37322 414765
rect 37270 414701 37322 414707
rect 41794 413433 41822 426721
rect 42178 420019 42206 429829
rect 43522 429140 43550 434417
rect 43618 432123 43646 559773
rect 43702 541521 43754 541527
rect 43702 541463 43754 541469
rect 43714 538197 43742 541463
rect 43702 538191 43754 538197
rect 43702 538133 43754 538139
rect 43604 432114 43660 432123
rect 43604 432049 43660 432058
rect 43234 429112 43550 429140
rect 42740 424122 42796 424131
rect 42740 424057 42796 424066
rect 42644 420126 42700 420135
rect 42644 420061 42700 420070
rect 42166 420013 42218 420019
rect 42166 419955 42218 419961
rect 42358 420013 42410 420019
rect 42358 419955 42410 419961
rect 41782 413427 41834 413433
rect 41782 413369 41834 413375
rect 41782 413205 41834 413211
rect 41782 413147 41834 413153
rect 41794 412624 41822 413147
rect 42370 411361 42398 419955
rect 42658 418655 42686 420061
rect 42644 418646 42700 418655
rect 42644 418581 42646 418590
rect 42698 418581 42700 418590
rect 42646 418549 42698 418555
rect 42166 411355 42218 411361
rect 42166 411297 42218 411303
rect 42358 411355 42410 411361
rect 42358 411297 42410 411303
rect 42178 410805 42206 411297
rect 42070 410541 42122 410547
rect 42070 410483 42122 410489
rect 42082 410182 42110 410483
rect 42754 409511 42782 424057
rect 43028 421310 43084 421319
rect 43028 421245 43084 421254
rect 42934 416979 42986 416985
rect 42934 416921 42986 416927
rect 42838 414833 42890 414839
rect 42838 414775 42890 414781
rect 42166 409505 42218 409511
rect 42166 409447 42218 409453
rect 42742 409505 42794 409511
rect 42742 409447 42794 409453
rect 42178 408965 42206 409447
rect 42850 409437 42878 414775
rect 42838 409431 42890 409437
rect 42838 409373 42890 409379
rect 42946 409308 42974 416921
rect 42754 409280 42974 409308
rect 43042 409289 43070 421245
rect 43126 416239 43178 416245
rect 43126 416181 43178 416187
rect 43030 409283 43082 409289
rect 42166 408247 42218 408253
rect 42166 408189 42218 408195
rect 42178 407769 42206 408189
rect 42070 407507 42122 407513
rect 42070 407449 42122 407455
rect 42082 407148 42110 407449
rect 42166 406915 42218 406921
rect 42166 406857 42218 406863
rect 42178 406482 42206 406857
rect 41780 406066 41836 406075
rect 41780 406001 41836 406010
rect 41794 405929 41822 406001
rect 41972 404882 42028 404891
rect 41972 404817 42028 404826
rect 41986 404646 42014 404817
rect 41986 404632 42302 404646
rect 42000 404618 42302 404632
rect 41794 403855 41822 403997
rect 42166 403881 42218 403887
rect 41780 403846 41836 403855
rect 42166 403823 42218 403829
rect 41780 403781 41836 403790
rect 42178 403448 42206 403823
rect 42166 403363 42218 403369
rect 42166 403305 42218 403311
rect 42178 402782 42206 403305
rect 42164 402662 42220 402671
rect 42164 402597 42220 402606
rect 42178 402157 42206 402597
rect 41780 401922 41836 401931
rect 41780 401857 41836 401866
rect 41794 401598 41822 401857
rect 41780 400146 41836 400155
rect 41780 400081 41836 400090
rect 41794 399748 41822 400081
rect 42274 400007 42302 404618
rect 42754 403369 42782 409280
rect 43030 409225 43082 409231
rect 42838 409209 42890 409215
rect 43138 409160 43166 416181
rect 42838 409151 42890 409157
rect 42850 408253 42878 409151
rect 42946 409132 43166 409160
rect 42838 408247 42890 408253
rect 42838 408189 42890 408195
rect 42946 407513 42974 409132
rect 43030 409061 43082 409067
rect 43030 409003 43082 409009
rect 43126 409061 43178 409067
rect 43126 409003 43178 409009
rect 42934 407507 42986 407513
rect 42934 407449 42986 407455
rect 43042 406921 43070 409003
rect 43030 406915 43082 406921
rect 43030 406857 43082 406863
rect 43138 403887 43166 409003
rect 43126 403881 43178 403887
rect 43126 403823 43178 403829
rect 42742 403363 42794 403369
rect 42742 403305 42794 403311
rect 42260 399998 42316 400007
rect 42260 399933 42316 399942
rect 41780 399554 41836 399563
rect 41780 399489 41836 399498
rect 41794 399121 41822 399489
rect 41780 398814 41836 398823
rect 41780 398749 41836 398758
rect 41794 398490 41822 398749
rect 42358 393965 42410 393971
rect 42356 393930 42358 393939
rect 42410 393930 42412 393939
rect 42356 393865 42412 393874
rect 42358 393225 42410 393231
rect 42356 393190 42358 393199
rect 42410 393190 42412 393199
rect 42356 393125 42412 393134
rect 42358 392337 42410 392343
rect 42356 392302 42358 392311
rect 42410 392302 42412 392311
rect 42356 392237 42412 392246
rect 43234 391400 43262 429112
rect 43318 414759 43370 414765
rect 43318 414701 43370 414707
rect 43330 409067 43358 414701
rect 43318 409061 43370 409067
rect 43318 409003 43370 409009
rect 43138 391372 43262 391400
rect 43138 390979 43166 391372
rect 43220 391266 43276 391275
rect 43220 391201 43276 391210
rect 43124 390970 43180 390979
rect 43124 390905 43180 390914
rect 43028 387270 43084 387279
rect 43028 387205 43084 387214
rect 35924 384458 35980 384467
rect 35924 384393 35980 384402
rect 35938 371591 35966 384393
rect 41780 383570 41836 383579
rect 41780 383505 41836 383514
rect 37172 381202 37228 381211
rect 37172 381137 37228 381146
rect 37186 371919 37214 381137
rect 40052 380462 40108 380471
rect 40052 380397 40108 380406
rect 37268 378834 37324 378843
rect 37268 378769 37324 378778
rect 37174 371913 37226 371919
rect 37174 371855 37226 371861
rect 37282 371845 37310 378769
rect 37364 378094 37420 378103
rect 37364 378029 37420 378038
rect 37270 371839 37322 371845
rect 37270 371781 37322 371787
rect 37378 371771 37406 378029
rect 37366 371765 37418 371771
rect 37366 371707 37418 371713
rect 40066 371623 40094 380397
rect 40148 377502 40204 377511
rect 40148 377437 40204 377446
rect 40162 371697 40190 377437
rect 40150 371691 40202 371697
rect 40150 371633 40202 371639
rect 40054 371617 40106 371623
rect 35924 371582 35980 371591
rect 40054 371559 40106 371565
rect 35924 371517 35980 371526
rect 41794 370217 41822 383505
rect 42932 380314 42988 380323
rect 42932 380249 42988 380258
rect 42356 376762 42412 376771
rect 42356 376697 42412 376706
rect 42370 375291 42398 376697
rect 42356 375282 42412 375291
rect 42356 375217 42358 375226
rect 42410 375217 42412 375226
rect 42358 375185 42410 375191
rect 42838 371765 42890 371771
rect 42838 371707 42890 371713
rect 42742 371691 42794 371697
rect 42742 371633 42794 371639
rect 42358 371617 42410 371623
rect 42358 371559 42410 371565
rect 41782 370211 41834 370217
rect 41782 370153 41834 370159
rect 41782 369989 41834 369995
rect 41782 369931 41834 369937
rect 41794 369445 41822 369931
rect 42070 368139 42122 368145
rect 42070 368081 42122 368087
rect 42082 367632 42110 368081
rect 42070 367399 42122 367405
rect 42070 367341 42122 367347
rect 42082 366966 42110 367341
rect 42370 366295 42398 371559
rect 42070 366289 42122 366295
rect 42070 366231 42122 366237
rect 42358 366289 42410 366295
rect 42358 366231 42410 366237
rect 42082 365782 42110 366231
rect 42358 366141 42410 366147
rect 42358 366083 42410 366089
rect 42166 365031 42218 365037
rect 42166 364973 42218 364979
rect 42178 364569 42206 364973
rect 42070 364439 42122 364445
rect 42070 364381 42122 364387
rect 42082 363932 42110 364381
rect 42166 363699 42218 363705
rect 42166 363641 42218 363647
rect 42178 363266 42206 363641
rect 42068 362850 42124 362859
rect 42068 362785 42124 362794
rect 42082 362748 42110 362785
rect 41876 361962 41932 361971
rect 41876 361897 41932 361906
rect 41890 361416 41918 361897
rect 41780 361370 41836 361379
rect 41780 361305 41836 361314
rect 41794 360824 41822 361305
rect 42370 360246 42398 366083
rect 42754 365037 42782 371633
rect 42742 365031 42794 365037
rect 42742 364973 42794 364979
rect 42850 363705 42878 371707
rect 42946 364445 42974 380249
rect 43042 368145 43070 387205
rect 43126 371839 43178 371845
rect 43126 371781 43178 371787
rect 43030 368139 43082 368145
rect 43030 368081 43082 368087
rect 43030 367991 43082 367997
rect 43030 367933 43082 367939
rect 42934 364439 42986 364445
rect 42934 364381 42986 364387
rect 42838 363699 42890 363705
rect 42838 363641 42890 363647
rect 42192 360218 42398 360246
rect 43042 360153 43070 367933
rect 43138 366147 43166 371781
rect 43126 366141 43178 366147
rect 43126 366083 43178 366089
rect 42358 360147 42410 360153
rect 42358 360089 42410 360095
rect 43030 360147 43082 360153
rect 43030 360089 43082 360095
rect 42370 359615 42398 360089
rect 42192 359587 42398 359615
rect 41780 359446 41836 359455
rect 41780 359381 41836 359390
rect 41794 358974 41822 359381
rect 41780 358706 41836 358715
rect 41780 358641 41836 358650
rect 41794 358382 41822 358641
rect 41876 356930 41932 356939
rect 41876 356865 41932 356874
rect 41890 356565 41918 356865
rect 41780 356486 41836 356495
rect 41780 356421 41836 356430
rect 41794 355940 41822 356421
rect 41780 355598 41836 355607
rect 41780 355533 41836 355542
rect 41794 355274 41822 355533
rect 42358 350749 42410 350755
rect 42356 350714 42358 350723
rect 42410 350714 42412 350723
rect 42356 350649 42412 350658
rect 42646 349713 42698 349719
rect 42644 349678 42646 349687
rect 42698 349678 42700 349687
rect 42644 349613 42700 349622
rect 42358 349121 42410 349127
rect 42356 349086 42358 349095
rect 42410 349086 42412 349095
rect 42356 349021 42412 349030
rect 43234 347763 43262 391201
rect 43318 371913 43370 371919
rect 43318 371855 43370 371861
rect 43330 367997 43358 371855
rect 43318 367991 43370 367997
rect 43318 367933 43370 367939
rect 43220 347754 43276 347763
rect 43220 347689 43276 347698
rect 43220 347606 43276 347615
rect 43220 347541 43276 347550
rect 42740 344128 42796 344137
rect 42740 344063 42796 344072
rect 39956 340354 40012 340363
rect 39956 340289 40012 340298
rect 37172 337394 37228 337403
rect 37172 337329 37228 337338
rect 37186 330479 37214 337329
rect 39970 331219 39998 340289
rect 42356 337986 42412 337995
rect 42356 337921 42412 337930
rect 40052 337246 40108 337255
rect 40052 337181 40108 337190
rect 39958 331213 40010 331219
rect 39958 331155 40010 331161
rect 37174 330473 37226 330479
rect 37174 330415 37226 330421
rect 40066 328407 40094 337181
rect 40244 334138 40300 334147
rect 40244 334073 40300 334082
rect 40258 328555 40286 334073
rect 42164 333546 42220 333555
rect 42164 333481 42220 333490
rect 42178 332075 42206 333481
rect 42164 332066 42220 332075
rect 42164 332001 42166 332010
rect 42218 332001 42220 332010
rect 42166 331969 42218 331975
rect 41782 331213 41834 331219
rect 41782 331155 41834 331161
rect 40534 330473 40586 330479
rect 40534 330415 40586 330421
rect 40246 328549 40298 328555
rect 40246 328491 40298 328497
rect 40054 328401 40106 328407
rect 40054 328343 40106 328349
rect 40546 327371 40574 330415
rect 40534 327365 40586 327371
rect 40534 327307 40586 327313
rect 41794 327075 41822 331155
rect 42370 327487 42398 337921
rect 42356 327478 42412 327487
rect 42356 327413 42412 327422
rect 42358 327365 42410 327371
rect 42358 327307 42410 327313
rect 41782 327069 41834 327075
rect 41782 327011 41834 327017
rect 41782 326773 41834 326779
rect 41782 326715 41834 326721
rect 41794 326266 41822 326715
rect 42070 324923 42122 324929
rect 42070 324865 42122 324871
rect 42082 324416 42110 324865
rect 42166 324183 42218 324189
rect 42166 324125 42218 324131
rect 42178 323750 42206 324125
rect 42370 323153 42398 327307
rect 42754 324929 42782 344063
rect 43124 335470 43180 335479
rect 43124 335405 43180 335414
rect 43030 328549 43082 328555
rect 43030 328491 43082 328497
rect 43042 328204 43070 328491
rect 43138 328333 43166 335405
rect 43126 328327 43178 328333
rect 43126 328269 43178 328275
rect 43042 328176 43166 328204
rect 43030 328105 43082 328111
rect 43030 328047 43082 328053
rect 42742 324923 42794 324929
rect 42742 324865 42794 324871
rect 42454 324405 42506 324411
rect 42454 324347 42506 324353
rect 42166 323147 42218 323153
rect 42166 323089 42218 323095
rect 42358 323147 42410 323153
rect 42358 323089 42410 323095
rect 42178 322566 42206 323089
rect 42356 323038 42412 323047
rect 42356 322973 42412 322982
rect 42070 321815 42122 321821
rect 42070 321757 42122 321763
rect 42082 321382 42110 321757
rect 42166 321075 42218 321081
rect 42166 321017 42218 321023
rect 42178 320716 42206 321017
rect 42166 320631 42218 320637
rect 42166 320573 42218 320579
rect 42178 320081 42206 320573
rect 41780 319782 41836 319791
rect 41780 319717 41836 319726
rect 41794 319532 41822 319717
rect 41876 318746 41932 318755
rect 41876 318681 41932 318690
rect 41890 318241 41918 318681
rect 41780 318006 41836 318015
rect 41780 317941 41836 317950
rect 41794 317608 41822 317941
rect 42164 317414 42220 317423
rect 42164 317349 42220 317358
rect 42178 317045 42206 317349
rect 42370 317104 42398 322973
rect 42466 320637 42494 324347
rect 43042 321081 43070 328047
rect 43138 321821 43166 328176
rect 43126 321815 43178 321821
rect 43126 321757 43178 321763
rect 43030 321075 43082 321081
rect 43030 321017 43082 321023
rect 42454 320631 42506 320637
rect 42454 320573 42506 320579
rect 42274 317076 42398 317104
rect 42178 316364 42206 316424
rect 42274 316364 42302 317076
rect 42178 316336 42302 316364
rect 41780 316230 41836 316239
rect 41780 316165 41836 316174
rect 41794 315758 41822 316165
rect 41780 315490 41836 315499
rect 41780 315425 41836 315434
rect 41794 315205 41822 315425
rect 41780 313714 41836 313723
rect 41780 313649 41836 313658
rect 41794 313390 41822 313649
rect 41780 313270 41836 313279
rect 41780 313205 41836 313214
rect 41794 312724 41822 313205
rect 41780 312382 41836 312391
rect 41780 312317 41836 312326
rect 41794 312058 41822 312317
rect 42262 307533 42314 307539
rect 42260 307498 42262 307507
rect 42314 307498 42316 307507
rect 42260 307433 42316 307442
rect 42262 306793 42314 306799
rect 42260 306758 42262 306767
rect 42314 306758 42316 306767
rect 42260 306693 42316 306702
rect 42836 305722 42892 305731
rect 42836 305657 42892 305666
rect 42850 305541 42878 305657
rect 42838 305535 42890 305541
rect 42838 305477 42890 305483
rect 43234 304103 43262 347541
rect 43318 328327 43370 328333
rect 43318 328269 43370 328275
rect 43330 324411 43358 328269
rect 43318 324405 43370 324411
rect 43318 324347 43370 324353
rect 43220 304094 43276 304103
rect 43220 304029 43276 304038
rect 43220 303946 43276 303955
rect 43220 303881 43276 303890
rect 41972 300394 42028 300403
rect 41972 300329 42028 300338
rect 39956 297286 40012 297295
rect 39956 297221 40012 297230
rect 37364 294030 37420 294039
rect 37364 293965 37420 293974
rect 37378 286893 37406 293965
rect 39970 288003 39998 297221
rect 40148 294030 40204 294039
rect 40148 293965 40204 293974
rect 39958 287997 40010 288003
rect 39958 287939 40010 287945
rect 37366 286887 37418 286893
rect 37366 286829 37418 286835
rect 40162 285709 40190 293965
rect 40244 290922 40300 290931
rect 40244 290857 40300 290866
rect 40150 285703 40202 285709
rect 40150 285645 40202 285651
rect 40258 285191 40286 290857
rect 41986 288965 42014 300329
rect 42164 294770 42220 294779
rect 42164 294705 42220 294714
rect 41974 288959 42026 288965
rect 41974 288901 42026 288907
rect 41782 287997 41834 288003
rect 41782 287939 41834 287945
rect 40246 285185 40298 285191
rect 40246 285127 40298 285133
rect 41794 283859 41822 287939
rect 42178 283859 42206 294705
rect 42260 292698 42316 292707
rect 42260 292633 42316 292642
rect 41782 283853 41834 283859
rect 41782 283795 41834 283801
rect 42166 283853 42218 283859
rect 42166 283795 42218 283801
rect 42274 283679 42302 292633
rect 42836 292254 42892 292263
rect 42836 292189 42892 292198
rect 42548 290330 42604 290339
rect 42548 290265 42604 290274
rect 42562 289132 42590 290265
rect 42644 289146 42700 289155
rect 42562 289104 42644 289132
rect 42644 289081 42646 289090
rect 42698 289081 42700 289090
rect 42646 289049 42698 289055
rect 42550 288959 42602 288965
rect 42550 288901 42602 288907
rect 42260 283670 42316 283679
rect 42260 283605 42316 283614
rect 41782 283409 41834 283415
rect 41782 283351 41834 283357
rect 41794 283050 41822 283351
rect 42562 281787 42590 288901
rect 42742 286887 42794 286893
rect 42742 286829 42794 286835
rect 42646 285185 42698 285191
rect 42646 285127 42698 285133
rect 42166 281781 42218 281787
rect 42166 281723 42218 281729
rect 42550 281781 42602 281787
rect 42550 281723 42602 281729
rect 42178 281200 42206 281723
rect 42548 281598 42604 281607
rect 42548 281533 42604 281542
rect 42166 281115 42218 281121
rect 42166 281057 42218 281063
rect 42178 280534 42206 281057
rect 42166 279931 42218 279937
rect 42166 279873 42218 279879
rect 42178 279350 42206 279873
rect 42166 278599 42218 278605
rect 42166 278541 42218 278547
rect 42178 278166 42206 278541
rect 42562 278476 42590 281533
rect 42658 278605 42686 285127
rect 42754 279937 42782 286829
rect 42742 279931 42794 279937
rect 42742 279873 42794 279879
rect 42646 278599 42698 278605
rect 42646 278541 42698 278547
rect 42562 278448 42782 278476
rect 42166 277859 42218 277865
rect 42166 277801 42218 277807
rect 42178 277500 42206 277801
rect 42070 277415 42122 277421
rect 42070 277357 42122 277363
rect 42082 276908 42110 277357
rect 41780 276566 41836 276575
rect 41780 276501 41836 276510
rect 41794 276316 41822 276501
rect 41972 275234 42028 275243
rect 41972 275169 42028 275178
rect 41986 275072 42014 275169
rect 41986 275058 42192 275072
rect 42000 275044 42206 275058
rect 42178 274776 42206 275044
rect 42178 274748 42398 274776
rect 42262 274677 42314 274683
rect 41780 274642 41836 274651
rect 42262 274619 42314 274625
rect 41780 274577 41836 274586
rect 41794 274406 41822 274577
rect 41794 274392 42096 274406
rect 41808 274378 42110 274392
rect 42082 274165 42110 274378
rect 42070 274159 42122 274165
rect 42070 274101 42122 274107
rect 42274 273859 42302 274619
rect 42192 273831 42302 273859
rect 42262 273789 42314 273795
rect 42262 273731 42314 273737
rect 42274 273222 42302 273731
rect 42192 273194 42302 273222
rect 41780 272866 41836 272875
rect 41780 272801 41836 272810
rect 41794 272542 41822 272801
rect 41780 272422 41836 272431
rect 41780 272357 41836 272366
rect 41794 272024 41822 272357
rect 41780 270646 41836 270655
rect 41780 270581 41836 270590
rect 41794 270174 41822 270581
rect 42260 270498 42316 270507
rect 42370 270484 42398 274748
rect 42754 274683 42782 278448
rect 42850 277421 42878 292189
rect 43126 285703 43178 285709
rect 43126 285645 43178 285651
rect 43138 277865 43166 285645
rect 43234 277865 43262 303881
rect 43318 283853 43370 283859
rect 43318 283795 43370 283801
rect 43126 277859 43178 277865
rect 43126 277801 43178 277807
rect 43222 277859 43274 277865
rect 43222 277801 43274 277807
rect 43330 277736 43358 283795
rect 43138 277708 43358 277736
rect 42838 277415 42890 277421
rect 42838 277357 42890 277363
rect 42742 274677 42794 274683
rect 42742 274619 42794 274625
rect 43030 274159 43082 274165
rect 43030 274101 43082 274107
rect 43042 273592 43070 274101
rect 43138 273795 43166 277708
rect 43222 277637 43274 277643
rect 43222 277579 43274 277585
rect 43126 273789 43178 273795
rect 43126 273731 43178 273737
rect 43042 273564 43166 273592
rect 42316 270456 42398 270484
rect 42260 270433 42316 270442
rect 41780 270054 41836 270063
rect 41780 269989 41836 269998
rect 41794 269508 41822 269989
rect 41780 269166 41836 269175
rect 41780 269101 41836 269110
rect 41794 268877 41822 269101
rect 42262 264317 42314 264323
rect 42260 264282 42262 264291
rect 42314 264282 42316 264291
rect 42260 264217 42316 264226
rect 42262 263577 42314 263583
rect 42260 263542 42262 263551
rect 42314 263542 42316 263551
rect 42260 263477 42316 263486
rect 42262 262689 42314 262695
rect 42260 262654 42262 262663
rect 42314 262654 42316 262663
rect 42260 262589 42316 262598
rect 41780 259546 41836 259555
rect 41780 259481 41836 259490
rect 40244 254070 40300 254079
rect 40244 254005 40300 254014
rect 37364 250814 37420 250823
rect 37364 250749 37420 250758
rect 40052 250814 40108 250823
rect 40052 250749 40108 250758
rect 37268 249186 37324 249195
rect 37268 249121 37324 249130
rect 37282 242197 37310 249121
rect 37270 242191 37322 242197
rect 37270 242133 37322 242139
rect 37378 242049 37406 250749
rect 40066 242123 40094 250749
rect 40148 248002 40204 248011
rect 40148 247937 40204 247946
rect 40054 242117 40106 242123
rect 40054 242059 40106 242065
rect 37366 242043 37418 242049
rect 37366 241985 37418 241991
rect 40162 241975 40190 247937
rect 40258 243751 40286 254005
rect 41794 243844 41822 259481
rect 43028 259398 43084 259407
rect 43028 259333 43084 259342
rect 41972 257178 42028 257187
rect 41972 257113 42028 257122
rect 41698 243816 41822 243844
rect 40246 243745 40298 243751
rect 40246 243687 40298 243693
rect 40150 241969 40202 241975
rect 40150 241911 40202 241917
rect 41698 241827 41726 243816
rect 41782 243745 41834 243751
rect 41782 243687 41834 243693
rect 41686 241821 41738 241827
rect 41686 241763 41738 241769
rect 41794 240643 41822 243687
rect 41986 243603 42014 257113
rect 42068 251554 42124 251563
rect 42068 251489 42124 251498
rect 41974 243597 42026 243603
rect 41974 243539 42026 243545
rect 42082 240759 42110 251489
rect 42260 248446 42316 248455
rect 42260 248381 42316 248390
rect 42068 240750 42124 240759
rect 42068 240685 42124 240694
rect 41782 240637 41834 240643
rect 41782 240579 41834 240585
rect 42274 240588 42302 248381
rect 42356 245486 42412 245495
rect 42356 245421 42412 245430
rect 42370 244861 42398 245421
rect 42358 244855 42410 244861
rect 42358 244797 42410 244803
rect 42550 243597 42602 243603
rect 42550 243539 42602 243545
rect 42358 242117 42410 242123
rect 42358 242059 42410 242065
rect 42370 240759 42398 242059
rect 42356 240750 42412 240759
rect 42356 240685 42412 240694
rect 42274 240560 42398 240588
rect 41782 240415 41834 240421
rect 41782 240357 41834 240363
rect 41794 239834 41822 240357
rect 42166 238565 42218 238571
rect 42166 238507 42218 238513
rect 42178 237984 42206 238507
rect 42166 237899 42218 237905
rect 42166 237841 42218 237847
rect 42178 237361 42206 237841
rect 42166 236715 42218 236721
rect 42166 236657 42218 236663
rect 42178 236165 42206 236657
rect 42166 235457 42218 235463
rect 42166 235399 42218 235405
rect 42178 234950 42206 235399
rect 42166 234865 42218 234871
rect 42166 234807 42218 234813
rect 42178 234325 42206 234807
rect 42370 234205 42398 240560
rect 42562 238571 42590 243539
rect 43042 242216 43070 259333
rect 43138 245347 43166 273564
rect 43234 260887 43262 277579
rect 43412 261618 43468 261627
rect 43412 261553 43468 261562
rect 43220 260878 43276 260887
rect 43220 260813 43276 260822
rect 43124 245338 43180 245347
rect 43124 245273 43180 245282
rect 43138 243423 43166 245273
rect 43124 243414 43180 243423
rect 43124 243349 43180 243358
rect 42742 242191 42794 242197
rect 43042 242188 43262 242216
rect 42742 242133 42794 242139
rect 42754 240939 42782 242133
rect 43126 242043 43178 242049
rect 43126 241985 43178 241991
rect 43030 241969 43082 241975
rect 43030 241911 43082 241917
rect 42742 240933 42794 240939
rect 42742 240875 42794 240881
rect 42550 238565 42602 238571
rect 42550 238507 42602 238513
rect 42452 237938 42508 237947
rect 42452 237873 42508 237882
rect 42466 234871 42494 237873
rect 43042 235463 43070 241911
rect 43138 236721 43166 241985
rect 43234 241901 43262 242188
rect 43222 241895 43274 241901
rect 43222 241837 43274 241843
rect 43318 240933 43370 240939
rect 43318 240875 43370 240881
rect 43126 236715 43178 236721
rect 43126 236657 43178 236663
rect 43330 236592 43358 240875
rect 43138 236564 43358 236592
rect 43030 235457 43082 235463
rect 43030 235399 43082 235405
rect 42454 234865 42506 234871
rect 42454 234807 42506 234813
rect 43138 234723 43166 236564
rect 43426 236499 43454 261553
rect 44578 243677 44606 930925
rect 44758 805183 44810 805189
rect 44758 805125 44810 805131
rect 44662 418607 44714 418613
rect 44662 418549 44714 418555
rect 44674 246267 44702 418549
rect 44662 246261 44714 246267
rect 44662 246203 44714 246209
rect 44566 243671 44618 243677
rect 44566 243613 44618 243619
rect 44770 243455 44798 805125
rect 44866 801489 44894 985019
rect 44854 801483 44906 801489
rect 44854 801425 44906 801431
rect 44854 762263 44906 762269
rect 44854 762205 44906 762211
rect 44758 243449 44810 243455
rect 44758 243391 44810 243397
rect 44866 243381 44894 762205
rect 44962 757829 44990 985093
rect 44950 757823 45002 757829
rect 44950 757765 45002 757771
rect 44950 717271 45002 717277
rect 44950 717213 45002 717219
rect 44962 243899 44990 717213
rect 45058 673839 45086 985463
rect 50518 985447 50570 985453
rect 50518 985389 50570 985395
rect 47830 985373 47882 985379
rect 47830 985315 47882 985321
rect 45142 985225 45194 985231
rect 45142 985167 45194 985173
rect 45154 710839 45182 985167
rect 47446 983819 47498 983825
rect 47446 983761 47498 983767
rect 47458 946275 47486 983761
rect 47542 947781 47594 947787
rect 47542 947723 47594 947729
rect 47444 946266 47500 946275
rect 47444 946201 47500 946210
rect 47554 930249 47582 947723
rect 47542 930243 47594 930249
rect 47542 930185 47594 930191
rect 47446 913001 47498 913007
rect 47446 912943 47498 912949
rect 45142 710833 45194 710839
rect 45142 710775 45194 710781
rect 45046 673833 45098 673839
rect 45046 673775 45098 673781
rect 45046 632467 45098 632473
rect 45046 632409 45098 632415
rect 44950 243893 45002 243899
rect 44950 243835 45002 243841
rect 45058 243825 45086 632409
rect 45142 589251 45194 589257
rect 45142 589193 45194 589199
rect 45046 243819 45098 243825
rect 45046 243761 45098 243767
rect 45154 243529 45182 589193
rect 45238 546257 45290 546263
rect 45238 546199 45290 546205
rect 45250 243751 45278 546199
rect 45430 455089 45482 455095
rect 45430 455031 45482 455037
rect 45334 440733 45386 440739
rect 45334 440675 45386 440681
rect 45346 349127 45374 440675
rect 45442 393231 45470 455031
rect 47458 410547 47486 912943
rect 47542 815099 47594 815105
rect 47542 815041 47594 815047
rect 47554 779955 47582 815041
rect 47542 779949 47594 779955
rect 47542 779891 47594 779897
rect 47542 743097 47594 743103
rect 47542 743039 47594 743045
rect 47446 410541 47498 410547
rect 47446 410483 47498 410489
rect 45430 393225 45482 393231
rect 45430 393167 45482 393173
rect 45430 383087 45482 383093
rect 45430 383029 45482 383035
rect 45334 349121 45386 349127
rect 45334 349063 45386 349069
rect 45334 311085 45386 311091
rect 45334 311027 45386 311033
rect 45238 243745 45290 243751
rect 45238 243687 45290 243693
rect 45142 243523 45194 243529
rect 45142 243465 45194 243471
rect 44854 243375 44906 243381
rect 44854 243317 44906 243323
rect 44662 241969 44714 241975
rect 44662 241911 44714 241917
rect 43702 241895 43754 241901
rect 43702 241837 43754 241843
rect 43510 241821 43562 241827
rect 43510 241763 43562 241769
rect 43222 236493 43274 236499
rect 43222 236435 43274 236441
rect 43414 236493 43466 236499
rect 43414 236435 43466 236441
rect 42454 234717 42506 234723
rect 42454 234659 42506 234665
rect 43126 234717 43178 234723
rect 43126 234659 43178 234665
rect 42070 234199 42122 234205
rect 42070 234141 42122 234147
rect 42358 234199 42410 234205
rect 42358 234141 42410 234147
rect 42082 233692 42110 234141
rect 41780 233350 41836 233359
rect 41780 233285 41836 233294
rect 41794 233129 41822 233285
rect 41890 231731 41918 231842
rect 41876 231722 41932 231731
rect 41876 231657 41932 231666
rect 41794 231139 41822 231176
rect 41780 231130 41836 231139
rect 41780 231065 41836 231074
rect 42466 230672 42494 234659
rect 42192 230644 42494 230672
rect 42068 230538 42124 230547
rect 42068 230473 42124 230482
rect 42082 229992 42110 230473
rect 41780 229650 41836 229659
rect 41780 229585 41836 229594
rect 41794 229357 41822 229585
rect 41780 229058 41836 229067
rect 41780 228993 41836 229002
rect 41794 228808 41822 228993
rect 41780 227282 41836 227291
rect 41780 227217 41836 227226
rect 41794 226958 41822 227217
rect 41780 226838 41836 226847
rect 41780 226773 41836 226782
rect 41794 226321 41822 226773
rect 41780 225950 41836 225959
rect 41780 225885 41836 225894
rect 41794 225700 41822 225885
rect 42358 221101 42410 221107
rect 42356 221066 42358 221075
rect 42410 221066 42412 221075
rect 42356 221001 42412 221010
rect 42358 220361 42410 220367
rect 42356 220326 42358 220335
rect 42410 220326 42412 220335
rect 42356 220261 42412 220270
rect 42358 219473 42410 219479
rect 42356 219438 42358 219447
rect 42410 219438 42412 219447
rect 42356 219373 42412 219382
rect 43234 217671 43262 236435
rect 43318 236419 43370 236425
rect 43318 236361 43370 236367
rect 43220 217662 43276 217671
rect 43220 217597 43276 217606
rect 43330 216191 43358 236361
rect 43522 216931 43550 241763
rect 43714 236425 43742 241837
rect 43702 236419 43754 236425
rect 43702 236361 43754 236367
rect 43508 216922 43564 216931
rect 43508 216857 43564 216866
rect 43316 216182 43372 216191
rect 43316 216117 43372 216126
rect 41972 213962 42028 213971
rect 41972 213897 42028 213906
rect 41876 210854 41932 210863
rect 41876 210789 41932 210798
rect 37268 207746 37324 207755
rect 37268 207681 37324 207690
rect 37282 200239 37310 207681
rect 40148 207154 40204 207163
rect 40148 207089 40204 207098
rect 37364 206118 37420 206127
rect 37364 206053 37420 206062
rect 37270 200233 37322 200239
rect 37270 200175 37322 200181
rect 37378 198907 37406 206053
rect 40162 201571 40190 207089
rect 40244 204638 40300 204647
rect 40244 204573 40300 204582
rect 40150 201565 40202 201571
rect 40150 201507 40202 201513
rect 37366 198901 37418 198907
rect 37366 198843 37418 198849
rect 40258 198833 40286 204573
rect 40246 198827 40298 198833
rect 40246 198769 40298 198775
rect 41890 197427 41918 210789
rect 41986 197427 42014 213897
rect 43124 209818 43180 209827
rect 43124 209753 43180 209762
rect 42068 208338 42124 208347
rect 42068 208273 42124 208282
rect 42082 197501 42110 208273
rect 42356 205526 42412 205535
rect 42356 205461 42412 205470
rect 42166 204377 42218 204383
rect 42164 204342 42166 204351
rect 42218 204342 42220 204351
rect 42164 204277 42220 204286
rect 42178 203019 42206 204277
rect 42164 203010 42220 203019
rect 42164 202945 42220 202954
rect 42166 201565 42218 201571
rect 42166 201507 42218 201513
rect 42178 197691 42206 201507
rect 42164 197682 42220 197691
rect 42164 197617 42220 197626
rect 42070 197495 42122 197501
rect 42070 197437 42122 197443
rect 41878 197421 41930 197427
rect 41878 197363 41930 197369
rect 41974 197421 42026 197427
rect 42370 197395 42398 205461
rect 43138 200332 43166 209753
rect 44674 204383 44702 241911
rect 45346 219479 45374 311027
rect 45442 307539 45470 383029
rect 47446 375243 47498 375249
rect 47446 375185 47498 375191
rect 45430 307533 45482 307539
rect 45430 307475 45482 307481
rect 45430 296729 45482 296735
rect 45430 296671 45482 296677
rect 45442 221107 45470 296671
rect 45526 282299 45578 282305
rect 45526 282241 45578 282247
rect 45430 221101 45482 221107
rect 45430 221043 45482 221049
rect 45538 220367 45566 282241
rect 47458 246341 47486 375185
rect 47554 281121 47582 743039
rect 47734 675683 47786 675689
rect 47734 675625 47786 675631
rect 47638 627879 47690 627885
rect 47638 627821 47690 627827
rect 47542 281115 47594 281121
rect 47542 281057 47594 281063
rect 47446 246335 47498 246341
rect 47446 246277 47498 246283
rect 45526 220361 45578 220367
rect 45526 220303 45578 220309
rect 45334 219473 45386 219479
rect 45334 219415 45386 219421
rect 44662 204377 44714 204383
rect 44662 204319 44714 204325
rect 42946 200304 43166 200332
rect 42454 197495 42506 197501
rect 42454 197437 42506 197443
rect 41974 197363 42026 197369
rect 42356 197386 42412 197395
rect 42356 197321 42412 197330
rect 42358 197273 42410 197279
rect 42358 197215 42410 197221
rect 41878 197199 41930 197205
rect 41878 197141 41930 197147
rect 41890 196618 41918 197141
rect 42370 195355 42398 197215
rect 42166 195349 42218 195355
rect 42166 195291 42218 195297
rect 42358 195349 42410 195355
rect 42358 195291 42410 195297
rect 42178 194805 42206 195291
rect 42356 195166 42412 195175
rect 42356 195101 42412 195110
rect 42070 194535 42122 194541
rect 42070 194477 42122 194483
rect 42082 194176 42110 194477
rect 42070 193499 42122 193505
rect 42070 193441 42122 193447
rect 42082 192992 42110 193441
rect 42166 192241 42218 192247
rect 42166 192183 42218 192189
rect 42178 191769 42206 192183
rect 42370 191507 42398 195101
rect 42070 191501 42122 191507
rect 42070 191443 42122 191449
rect 42358 191501 42410 191507
rect 42358 191443 42410 191449
rect 42082 191142 42110 191443
rect 42358 191353 42410 191359
rect 42358 191295 42410 191301
rect 42068 191022 42124 191031
rect 42068 190957 42124 190966
rect 42082 190476 42110 190957
rect 41780 190134 41836 190143
rect 41780 190069 41836 190078
rect 41794 189929 41822 190069
rect 41876 189098 41932 189107
rect 41876 189033 41932 189042
rect 41890 188626 41918 189033
rect 42370 188492 42398 191295
rect 42274 188464 42398 188492
rect 41780 188358 41836 188367
rect 41780 188293 41836 188302
rect 41794 188011 41822 188293
rect 41794 187997 42192 188011
rect 41808 187983 42206 187997
rect 42178 187881 42206 187983
rect 42166 187875 42218 187881
rect 42166 187817 42218 187823
rect 42274 187456 42302 188464
rect 42192 187428 42302 187456
rect 42466 187141 42494 197437
rect 42646 195793 42698 195799
rect 42646 195735 42698 195741
rect 42658 191359 42686 195735
rect 42646 191353 42698 191359
rect 42646 191295 42698 191301
rect 42946 188196 42974 200304
rect 43126 200233 43178 200239
rect 43126 200175 43178 200181
rect 43030 198827 43082 198833
rect 43030 198769 43082 198775
rect 43042 192247 43070 198769
rect 43138 193505 43166 200175
rect 43222 198901 43274 198907
rect 43222 198843 43274 198849
rect 43234 195799 43262 198843
rect 43222 195793 43274 195799
rect 43222 195735 43274 195741
rect 47650 194541 47678 627821
rect 47746 243603 47774 675625
rect 47842 627959 47870 985315
rect 50326 947707 50378 947713
rect 50326 947649 50378 947655
rect 50338 944605 50366 947649
rect 50326 944599 50378 944605
rect 50326 944541 50378 944547
rect 50422 884215 50474 884221
rect 50422 884157 50474 884163
rect 50326 858315 50378 858321
rect 50326 858257 50378 858263
rect 47830 627953 47882 627959
rect 47830 627895 47882 627901
rect 50338 367405 50366 858257
rect 50434 823911 50462 884157
rect 50422 823905 50474 823911
rect 50422 823847 50474 823853
rect 50422 757527 50474 757533
rect 50422 757469 50474 757475
rect 50434 736739 50462 757469
rect 50422 736733 50474 736739
rect 50422 736675 50474 736681
rect 50422 728667 50474 728673
rect 50422 728609 50474 728615
rect 50434 692487 50462 728609
rect 50422 692481 50474 692487
rect 50422 692423 50474 692429
rect 50422 685525 50474 685531
rect 50422 685467 50474 685473
rect 50326 367399 50378 367405
rect 50326 367341 50378 367347
rect 47830 354301 47882 354307
rect 47830 354243 47882 354249
rect 47842 262695 47870 354243
rect 47926 332027 47978 332033
rect 47926 331969 47978 331975
rect 47830 262689 47882 262695
rect 47830 262631 47882 262637
rect 47938 246489 47966 331969
rect 48022 289107 48074 289113
rect 48022 289049 48074 289055
rect 47926 246483 47978 246489
rect 47926 246425 47978 246431
rect 48034 246415 48062 289049
rect 48022 246409 48074 246415
rect 48022 246351 48074 246357
rect 47734 243597 47786 243603
rect 47734 243539 47786 243545
rect 50434 237905 50462 685467
rect 50530 584743 50558 985389
rect 59540 973202 59596 973211
rect 59540 973137 59596 973146
rect 59554 970653 59582 973137
rect 53302 970647 53354 970653
rect 53302 970589 53354 970595
rect 59542 970647 59594 970653
rect 59542 970589 59594 970595
rect 53206 901531 53258 901537
rect 53206 901473 53258 901479
rect 50614 829529 50666 829535
rect 50614 829471 50666 829477
rect 50626 780473 50654 829471
rect 53218 822283 53246 901473
rect 53206 822277 53258 822283
rect 53206 822219 53258 822225
rect 53206 800669 53258 800675
rect 53206 800611 53258 800617
rect 50614 780467 50666 780473
rect 50614 780409 50666 780415
rect 51862 649783 51914 649789
rect 51862 649725 51914 649731
rect 51874 644535 51902 649725
rect 51862 644529 51914 644535
rect 51862 644471 51914 644477
rect 51862 607751 51914 607757
rect 51862 607693 51914 607699
rect 51874 601911 51902 607693
rect 51862 601905 51914 601911
rect 51862 601847 51914 601853
rect 50518 584737 50570 584743
rect 50518 584679 50570 584685
rect 50518 563499 50570 563505
rect 50518 563441 50570 563447
rect 50530 543747 50558 563441
rect 50518 543741 50570 543747
rect 50518 543683 50570 543689
rect 50518 512735 50570 512741
rect 50518 512677 50570 512683
rect 50530 436965 50558 512677
rect 50614 469519 50666 469525
rect 50614 469461 50666 469467
rect 50518 436959 50570 436965
rect 50518 436901 50570 436907
rect 50626 393971 50654 469461
rect 50614 393965 50666 393971
rect 50614 393907 50666 393913
rect 50518 368731 50570 368737
rect 50518 368673 50570 368679
rect 50530 306799 50558 368673
rect 53218 324189 53246 800611
rect 53314 541527 53342 970589
rect 61858 962111 61886 993857
rect 62036 992146 62092 992155
rect 62036 992081 62092 992090
rect 62050 962555 62078 992081
rect 69154 987895 69182 995157
rect 77314 993667 77342 995508
rect 77698 993815 77726 995522
rect 77686 993809 77738 993815
rect 78370 993783 78398 995522
rect 77686 993751 77738 993757
rect 78356 993774 78412 993783
rect 80194 993741 80222 995522
rect 81408 995517 81662 995536
rect 81408 995511 81674 995517
rect 81408 995508 81622 995511
rect 81622 995453 81674 995459
rect 82594 995115 82622 995522
rect 83232 995508 83486 995536
rect 82580 995106 82636 995115
rect 82580 995041 82636 995050
rect 82594 993931 82622 995041
rect 82580 993922 82636 993931
rect 82580 993857 82636 993866
rect 78356 993709 78412 993718
rect 80182 993735 80234 993741
rect 80182 993677 80234 993683
rect 77302 993661 77354 993667
rect 83458 993635 83486 995508
rect 84514 994671 84542 995522
rect 85104 995508 85406 995536
rect 86352 995508 86462 995536
rect 88752 995508 89054 995536
rect 89424 995508 89822 995536
rect 85378 995411 85406 995508
rect 85364 995402 85420 995411
rect 85364 995337 85420 995346
rect 86434 995263 86462 995508
rect 86420 995254 86476 995263
rect 86420 995189 86476 995198
rect 89026 995073 89054 995508
rect 89794 995443 89822 995508
rect 92098 995443 92126 995804
rect 89782 995437 89834 995443
rect 89782 995379 89834 995385
rect 92086 995437 92138 995443
rect 92086 995379 92138 995385
rect 89014 995067 89066 995073
rect 89014 995009 89066 995015
rect 84500 994662 84556 994671
rect 84500 994597 84556 994606
rect 93058 993635 93086 999597
rect 77302 993603 77354 993609
rect 83444 993626 83500 993635
rect 83444 993561 83500 993570
rect 93044 993626 93100 993635
rect 93044 993561 93100 993570
rect 83458 992155 83486 993561
rect 83444 992146 83500 992155
rect 83444 992081 83500 992090
rect 69142 987889 69194 987895
rect 69142 987831 69194 987837
rect 64918 987815 64970 987821
rect 64918 987757 64970 987763
rect 64726 980859 64778 980865
rect 64726 980801 64778 980807
rect 62036 962546 62092 962555
rect 62036 962481 62092 962490
rect 61844 962102 61900 962111
rect 61844 962037 61900 962046
rect 59540 958846 59596 958855
rect 59540 958781 59596 958790
rect 59554 956223 59582 958781
rect 59542 956217 59594 956223
rect 59542 956159 59594 956165
rect 59540 944638 59596 944647
rect 59540 944573 59542 944582
rect 59594 944573 59596 944582
rect 59542 944541 59594 944547
rect 59542 930243 59594 930249
rect 59542 930185 59594 930191
rect 59554 930143 59582 930185
rect 59540 930134 59596 930143
rect 59540 930069 59596 930078
rect 59540 915778 59596 915787
rect 59540 915713 59596 915722
rect 59554 913007 59582 915713
rect 59542 913001 59594 913007
rect 59542 912943 59594 912949
rect 58196 901570 58252 901579
rect 58196 901505 58198 901514
rect 58250 901505 58252 901514
rect 58198 901473 58250 901479
rect 59540 887066 59596 887075
rect 59540 887001 59596 887010
rect 59554 884221 59582 887001
rect 59542 884215 59594 884221
rect 59542 884157 59594 884163
rect 58964 872562 59020 872571
rect 58964 872497 59020 872506
rect 53398 843885 53450 843891
rect 53398 843827 53450 843833
rect 53410 778919 53438 843827
rect 58978 821913 59006 872497
rect 59540 858354 59596 858363
rect 59540 858289 59542 858298
rect 59594 858289 59596 858298
rect 59542 858257 59594 858263
rect 59540 843998 59596 844007
rect 59540 843933 59596 843942
rect 59554 843891 59582 843933
rect 59542 843885 59594 843891
rect 59542 843827 59594 843833
rect 59540 829642 59596 829651
rect 59540 829577 59596 829586
rect 59554 829535 59582 829577
rect 59542 829529 59594 829535
rect 59542 829471 59594 829477
rect 58966 821907 59018 821913
rect 58966 821849 59018 821855
rect 59540 815286 59596 815295
rect 59540 815221 59596 815230
rect 59554 815105 59582 815221
rect 59542 815099 59594 815105
rect 59542 815041 59594 815047
rect 59540 800782 59596 800791
rect 59540 800717 59596 800726
rect 59554 800675 59582 800717
rect 59542 800669 59594 800675
rect 59542 800611 59594 800617
rect 58964 786574 59020 786583
rect 58964 786509 59020 786518
rect 53398 778913 53450 778919
rect 53398 778855 53450 778861
rect 53398 771883 53450 771889
rect 53398 771825 53450 771831
rect 53410 737257 53438 771825
rect 53398 737251 53450 737257
rect 53398 737193 53450 737199
rect 58978 735481 59006 786509
rect 59540 772070 59596 772079
rect 59540 772005 59596 772014
rect 59554 771889 59582 772005
rect 59542 771883 59594 771889
rect 59542 771825 59594 771831
rect 59540 757714 59596 757723
rect 59540 757649 59596 757658
rect 59554 757533 59582 757649
rect 59542 757527 59594 757533
rect 59542 757469 59594 757475
rect 59540 743358 59596 743367
rect 59540 743293 59596 743302
rect 59554 743103 59582 743293
rect 59542 743097 59594 743103
rect 59542 743039 59594 743045
rect 58966 735475 59018 735481
rect 58966 735417 59018 735423
rect 58388 729002 58444 729011
rect 58388 728937 58444 728946
rect 58402 728673 58430 728937
rect 58390 728667 58442 728673
rect 58390 728609 58442 728615
rect 58388 714646 58444 714655
rect 58388 714581 58444 714590
rect 58402 714317 58430 714581
rect 53398 714311 53450 714317
rect 53398 714253 53450 714259
rect 58390 714311 58442 714317
rect 58390 714253 58442 714259
rect 53410 694041 53438 714253
rect 57812 700290 57868 700299
rect 57812 700225 57868 700234
rect 57826 699887 57854 700225
rect 57814 699881 57866 699887
rect 57814 699823 57866 699829
rect 53398 694035 53450 694041
rect 53398 693977 53450 693983
rect 59540 685934 59596 685943
rect 59540 685869 59596 685878
rect 59554 685531 59582 685869
rect 59542 685525 59594 685531
rect 59542 685467 59594 685473
rect 59444 671578 59500 671587
rect 59444 671513 59500 671522
rect 59458 671101 59486 671513
rect 53398 671095 53450 671101
rect 53398 671037 53450 671043
rect 59446 671095 59498 671101
rect 59446 671037 59498 671043
rect 53410 649567 53438 671037
rect 59540 657222 59596 657231
rect 59540 657157 59596 657166
rect 59554 656745 59582 657157
rect 59542 656739 59594 656745
rect 59542 656681 59594 656687
rect 53398 649561 53450 649567
rect 53398 649503 53450 649509
rect 59254 644529 59306 644535
rect 59254 644471 59306 644477
rect 59266 642875 59294 644471
rect 59252 642866 59308 642875
rect 59252 642801 59308 642810
rect 58004 628510 58060 628519
rect 58004 628445 58060 628454
rect 58018 627885 58046 628445
rect 58006 627879 58058 627885
rect 58006 627821 58058 627827
rect 59444 614006 59500 614015
rect 59444 613941 59500 613950
rect 59458 613529 59486 613941
rect 59446 613523 59498 613529
rect 59446 613465 59498 613471
rect 53398 606863 53450 606869
rect 53398 606805 53450 606811
rect 53410 587481 53438 606805
rect 59542 601905 59594 601911
rect 59542 601847 59594 601853
rect 59554 599807 59582 601847
rect 59540 599798 59596 599807
rect 59540 599733 59596 599742
rect 53398 587475 53450 587481
rect 53398 587417 53450 587423
rect 59542 587475 59594 587481
rect 59542 587417 59594 587423
rect 59554 585451 59582 587417
rect 59540 585442 59596 585451
rect 59540 585377 59596 585386
rect 59540 570938 59596 570947
rect 59540 570873 59596 570882
rect 59554 570313 59582 570873
rect 59542 570307 59594 570313
rect 59542 570249 59594 570255
rect 53398 564535 53450 564541
rect 53398 564477 53450 564483
rect 53410 558695 53438 564477
rect 53398 558689 53450 558695
rect 53398 558631 53450 558637
rect 59542 558689 59594 558695
rect 59542 558631 59594 558637
rect 59554 556739 59582 558631
rect 59540 556730 59596 556739
rect 59540 556665 59596 556674
rect 59542 543741 59594 543747
rect 59542 543683 59594 543689
rect 59554 542383 59582 543683
rect 59540 542374 59596 542383
rect 59540 542309 59596 542318
rect 53302 541521 53354 541527
rect 53302 541463 53354 541469
rect 59540 527870 59596 527879
rect 59540 527805 59596 527814
rect 59554 527097 59582 527805
rect 59542 527091 59594 527097
rect 59542 527033 59594 527039
rect 59348 513514 59404 513523
rect 59348 513449 59404 513458
rect 59362 512741 59390 513449
rect 59350 512735 59402 512741
rect 59350 512677 59402 512683
rect 57812 499158 57868 499167
rect 57812 499093 57868 499102
rect 57826 498311 57854 499093
rect 53398 498305 53450 498311
rect 53398 498247 53450 498253
rect 57814 498305 57866 498311
rect 57814 498247 57866 498253
rect 53302 483875 53354 483881
rect 53302 483817 53354 483823
rect 53314 392343 53342 483817
rect 53410 436151 53438 498247
rect 59540 484802 59596 484811
rect 59540 484737 59596 484746
rect 59554 483881 59582 484737
rect 59542 483875 59594 483881
rect 59542 483817 59594 483823
rect 59540 470446 59596 470455
rect 59540 470381 59596 470390
rect 59554 469525 59582 470381
rect 59542 469519 59594 469525
rect 59542 469461 59594 469467
rect 59540 456090 59596 456099
rect 59540 456025 59596 456034
rect 59554 455095 59582 456025
rect 59542 455089 59594 455095
rect 59542 455031 59594 455037
rect 57812 441586 57868 441595
rect 57812 441521 57868 441530
rect 57826 440739 57854 441521
rect 57814 440733 57866 440739
rect 57814 440675 57866 440681
rect 53398 436145 53450 436151
rect 53398 436087 53450 436093
rect 59540 427378 59596 427387
rect 59540 427313 59596 427322
rect 59554 426309 59582 427313
rect 53398 426303 53450 426309
rect 53398 426245 53450 426251
rect 59542 426303 59594 426309
rect 59542 426245 59594 426251
rect 53302 392337 53354 392343
rect 53302 392279 53354 392285
rect 53410 350755 53438 426245
rect 59540 412874 59596 412883
rect 59540 412809 59596 412818
rect 59554 411879 59582 412809
rect 53494 411873 53546 411879
rect 53494 411815 53546 411821
rect 59542 411873 59594 411879
rect 59542 411815 59594 411821
rect 53398 350749 53450 350755
rect 53398 350691 53450 350697
rect 53506 349719 53534 411815
rect 58964 398666 59020 398675
rect 58964 398601 59020 398610
rect 53494 349713 53546 349719
rect 53494 349655 53546 349661
rect 53302 339871 53354 339877
rect 53302 339813 53354 339819
rect 53206 324183 53258 324189
rect 53206 324125 53258 324131
rect 50518 306793 50570 306799
rect 50518 306735 50570 306741
rect 53314 264323 53342 339813
rect 53398 325515 53450 325521
rect 53398 325457 53450 325463
rect 53302 264317 53354 264323
rect 53302 264259 53354 264265
rect 53410 263583 53438 325457
rect 58978 305541 59006 398601
rect 59540 384162 59596 384171
rect 59540 384097 59596 384106
rect 59554 383093 59582 384097
rect 59542 383087 59594 383093
rect 59542 383029 59594 383035
rect 59540 369806 59596 369815
rect 59540 369741 59596 369750
rect 59554 368737 59582 369741
rect 59542 368731 59594 368737
rect 59542 368673 59594 368679
rect 59540 355598 59596 355607
rect 59540 355533 59596 355542
rect 59554 354307 59582 355533
rect 59542 354301 59594 354307
rect 59542 354243 59594 354249
rect 59540 341094 59596 341103
rect 59540 341029 59596 341038
rect 59554 339877 59582 341029
rect 59542 339871 59594 339877
rect 59542 339813 59594 339819
rect 59540 326738 59596 326747
rect 59540 326673 59596 326682
rect 59554 325521 59582 326673
rect 59542 325515 59594 325521
rect 59542 325457 59594 325463
rect 59540 312382 59596 312391
rect 59540 312317 59596 312326
rect 59554 311091 59582 312317
rect 59542 311085 59594 311091
rect 59542 311027 59594 311033
rect 58966 305535 59018 305541
rect 58966 305477 59018 305483
rect 59540 298026 59596 298035
rect 59540 297961 59596 297970
rect 59554 296735 59582 297961
rect 59542 296729 59594 296735
rect 59542 296671 59594 296677
rect 59540 283670 59596 283679
rect 59540 283605 59596 283614
rect 59554 282305 59582 283605
rect 59542 282299 59594 282305
rect 59542 282241 59594 282247
rect 64738 272315 64766 980801
rect 64822 980711 64874 980717
rect 64822 980653 64874 980659
rect 64834 272537 64862 980653
rect 64930 275053 64958 987757
rect 93634 986415 93662 1005369
rect 217268 1005318 217324 1005327
rect 217268 1005253 217270 1005262
rect 217322 1005253 217324 1005262
rect 218900 1005318 218956 1005327
rect 218900 1005253 218902 1005262
rect 217270 1005221 217322 1005227
rect 218954 1005253 218956 1005262
rect 223124 1005318 223180 1005327
rect 223124 1005253 223180 1005262
rect 218902 1005221 218954 1005227
rect 93718 1005205 93770 1005211
rect 115222 1005205 115274 1005211
rect 93718 1005147 93770 1005153
rect 115220 1005170 115222 1005179
rect 115274 1005170 115276 1005179
rect 73462 986409 73514 986415
rect 73462 986351 73514 986357
rect 93622 986409 93674 986415
rect 93622 986351 93674 986357
rect 65014 983893 65066 983899
rect 65014 983835 65066 983841
rect 64918 275047 64970 275053
rect 64918 274989 64970 274995
rect 64822 272531 64874 272537
rect 64822 272473 64874 272479
rect 64726 272309 64778 272315
rect 64726 272251 64778 272257
rect 53398 263577 53450 263583
rect 53398 263519 53450 263525
rect 65026 246235 65054 983835
rect 65110 983597 65162 983603
rect 65110 983539 65162 983545
rect 65122 246563 65150 983539
rect 65206 983523 65258 983529
rect 65206 983465 65258 983471
rect 65110 246557 65162 246563
rect 65110 246499 65162 246505
rect 65218 246383 65246 983465
rect 73474 981462 73502 986351
rect 93730 985897 93758 1005147
rect 115220 1005105 115276 1005114
rect 221876 1005170 221932 1005179
rect 221876 1005105 221932 1005114
rect 144022 1002541 144074 1002547
rect 150358 1002541 150410 1002547
rect 144022 1002483 144074 1002489
rect 150356 1002506 150358 1002515
rect 150410 1002506 150412 1002515
rect 143926 1002393 143978 1002399
rect 143926 1002335 143978 1002341
rect 143734 1002319 143786 1002325
rect 143734 1002261 143786 1002267
rect 127414 999655 127466 999661
rect 127414 999597 127466 999603
rect 115318 996177 115370 996183
rect 115318 996119 115370 996125
rect 126742 996177 126794 996183
rect 126742 996119 126794 996125
rect 115222 996103 115274 996109
rect 115222 996045 115274 996051
rect 100628 995994 100684 996003
rect 100628 995929 100630 995938
rect 100682 995929 100684 995938
rect 107252 995994 107308 996003
rect 107252 995929 107308 995938
rect 100630 995897 100682 995903
rect 94678 995881 94730 995887
rect 99958 995881 100010 995887
rect 94678 995823 94730 995829
rect 94868 995846 94924 995855
rect 94690 995411 94718 995823
rect 94868 995781 94924 995790
rect 99956 995846 99958 995855
rect 100010 995846 100012 995855
rect 99956 995781 100012 995790
rect 102164 995846 102220 995855
rect 102164 995781 102166 995790
rect 94882 995411 94910 995781
rect 102218 995781 102220 995790
rect 105332 995846 105388 995855
rect 105332 995781 105388 995790
rect 106486 995807 106538 995813
rect 102166 995749 102218 995755
rect 105346 995739 105374 995781
rect 106486 995749 106538 995755
rect 105334 995733 105386 995739
rect 94964 995698 95020 995707
rect 94964 995633 95020 995642
rect 98996 995698 99052 995707
rect 105334 995675 105386 995681
rect 98996 995633 99052 995642
rect 94676 995402 94732 995411
rect 94676 995337 94732 995346
rect 94868 995402 94924 995411
rect 94868 995337 94924 995346
rect 89590 985891 89642 985897
rect 89590 985833 89642 985839
rect 93718 985891 93770 985897
rect 93718 985833 93770 985839
rect 80578 985592 80798 985620
rect 80578 985305 80606 985592
rect 80770 985527 80798 985592
rect 80758 985521 80810 985527
rect 80758 985463 80810 985469
rect 80566 985299 80618 985305
rect 80566 985241 80618 985247
rect 89602 981462 89630 985833
rect 94978 983899 95006 995633
rect 99010 995263 99038 995633
rect 102164 995550 102220 995559
rect 102164 995485 102166 995494
rect 102218 995485 102220 995494
rect 102166 995453 102218 995459
rect 98996 995254 99052 995263
rect 98996 995189 99052 995198
rect 100724 995254 100780 995263
rect 100724 995189 100780 995198
rect 100738 993815 100766 995189
rect 100726 993809 100778 993815
rect 100726 993751 100778 993757
rect 100822 985521 100874 985527
rect 100820 985486 100822 985495
rect 100874 985486 100876 985495
rect 100820 985421 100876 985430
rect 94966 983893 95018 983899
rect 94966 983835 95018 983841
rect 106498 981624 106526 995749
rect 106580 995254 106636 995263
rect 106580 995189 106636 995198
rect 106594 994671 106622 995189
rect 106580 994662 106636 994671
rect 106580 994597 106636 994606
rect 107266 993741 107294 995929
rect 113494 995881 113546 995887
rect 113300 995846 113356 995855
rect 113300 995781 113302 995790
rect 113354 995781 113356 995790
rect 113492 995846 113494 995855
rect 113546 995846 113548 995855
rect 113492 995781 113548 995790
rect 113302 995749 113354 995755
rect 115234 995559 115262 996045
rect 115220 995550 115276 995559
rect 115220 995485 115276 995494
rect 108212 995254 108268 995263
rect 108212 995189 108268 995198
rect 108404 995254 108460 995263
rect 108404 995189 108460 995198
rect 107254 993735 107306 993741
rect 107254 993677 107306 993683
rect 108226 993667 108254 995189
rect 108418 993783 108446 995189
rect 108404 993774 108460 993783
rect 108404 993709 108460 993718
rect 108214 993661 108266 993667
rect 108214 993603 108266 993609
rect 115234 983751 115262 995485
rect 115330 995411 115358 996119
rect 120982 996029 121034 996035
rect 120982 995971 121034 995977
rect 118102 995807 118154 995813
rect 118102 995749 118154 995755
rect 115316 995402 115372 995411
rect 115316 995337 115372 995346
rect 115222 983745 115274 983751
rect 115222 983687 115274 983693
rect 115330 983677 115358 995337
rect 118114 983825 118142 995749
rect 120994 995707 121022 995971
rect 120980 995698 121036 995707
rect 120980 995633 121036 995642
rect 126754 995443 126782 996119
rect 127426 995739 127454 999597
rect 143746 999532 143774 1002261
rect 143830 1000839 143882 1000845
rect 143830 1000781 143882 1000787
rect 143650 999504 143774 999532
rect 131732 995846 131788 995855
rect 131616 995804 131732 995832
rect 132144 995813 132446 995832
rect 133440 995813 133694 995832
rect 142656 995813 143006 995832
rect 132144 995807 132458 995813
rect 132144 995804 132406 995807
rect 131732 995781 131788 995790
rect 133440 995807 133706 995813
rect 133440 995804 133654 995807
rect 132406 995749 132458 995755
rect 142656 995807 143018 995813
rect 142656 995804 142966 995807
rect 133654 995749 133706 995755
rect 142966 995749 143018 995755
rect 127414 995733 127466 995739
rect 127414 995675 127466 995681
rect 134326 995733 134378 995739
rect 141046 995733 141098 995739
rect 136724 995698 136780 995707
rect 134378 995681 134640 995684
rect 134326 995675 134640 995681
rect 134338 995670 134640 995675
rect 134338 995656 134654 995670
rect 136464 995656 136724 995684
rect 126742 995437 126794 995443
rect 126742 995379 126794 995385
rect 128482 993741 128510 995522
rect 129120 995508 129374 995536
rect 129346 993815 129374 995508
rect 129334 993809 129386 993815
rect 129334 993751 129386 993757
rect 128470 993735 128522 993741
rect 128470 993677 128522 993683
rect 129730 993667 129758 995522
rect 132816 995508 133118 995536
rect 134016 995508 134270 995536
rect 133090 995411 133118 995508
rect 133076 995402 133132 995411
rect 133076 995337 133132 995346
rect 134242 995115 134270 995508
rect 134228 995106 134284 995115
rect 134228 995041 134284 995050
rect 134626 994819 134654 995656
rect 138960 995665 139358 995684
rect 140784 995681 141046 995684
rect 140784 995675 141098 995681
rect 138960 995659 139370 995665
rect 138960 995656 139318 995659
rect 136724 995633 136780 995642
rect 140784 995656 141086 995675
rect 139318 995601 139370 995607
rect 137974 995585 138026 995591
rect 137396 995550 137452 995559
rect 135936 995508 136190 995536
rect 137136 995508 137396 995536
rect 134612 994810 134668 994819
rect 134612 994745 134668 994754
rect 136162 994079 136190 995508
rect 137760 995533 137974 995536
rect 137760 995527 138026 995533
rect 137760 995508 138014 995527
rect 140160 995508 140414 995536
rect 137396 995485 137452 995494
rect 136148 994070 136204 994079
rect 136148 994005 136204 994014
rect 140386 993783 140414 995508
rect 143650 995115 143678 999504
rect 143734 999433 143786 999439
rect 143734 999375 143786 999381
rect 143746 995813 143774 999375
rect 143734 995807 143786 995813
rect 143734 995749 143786 995755
rect 143842 995739 143870 1000781
rect 143830 995733 143882 995739
rect 143830 995675 143882 995681
rect 143938 995665 143966 1002335
rect 143926 995659 143978 995665
rect 143926 995601 143978 995607
rect 144034 995591 144062 1002483
rect 150356 1002441 150412 1002450
rect 153622 1002393 153674 1002399
rect 153620 1002358 153622 1002367
rect 153674 1002358 153676 1002367
rect 153620 1002293 153676 1002302
rect 178486 1002319 178538 1002325
rect 178486 1002261 178538 1002267
rect 160244 1000878 160300 1000887
rect 160244 1000813 160246 1000822
rect 160298 1000813 160300 1000822
rect 160246 1000781 160298 1000787
rect 144214 999581 144266 999587
rect 158614 999581 158666 999587
rect 144214 999523 144266 999529
rect 155156 999546 155212 999555
rect 144118 999507 144170 999513
rect 144118 999449 144170 999455
rect 144130 995961 144158 999449
rect 144118 995955 144170 995961
rect 144118 995897 144170 995903
rect 144226 995855 144254 999523
rect 155156 999481 155158 999490
rect 155210 999481 155212 999490
rect 158612 999546 158614 999555
rect 158666 999546 158668 999555
rect 158612 999481 158668 999490
rect 155158 999449 155210 999455
rect 156886 999433 156938 999439
rect 156884 999398 156886 999407
rect 156938 999398 156940 999407
rect 156884 999333 156940 999342
rect 144310 996325 144362 996331
rect 162262 996325 162314 996331
rect 144310 996267 144362 996273
rect 162260 996290 162262 996299
rect 162314 996290 162316 996299
rect 144212 995846 144268 995855
rect 144212 995781 144268 995790
rect 144022 995585 144074 995591
rect 144022 995527 144074 995533
rect 144322 995443 144350 996267
rect 162260 996225 162316 996234
rect 163124 996142 163180 996151
rect 163124 996077 163126 996086
rect 163178 996077 163180 996086
rect 177046 996103 177098 996109
rect 163126 996045 163178 996051
rect 177046 996045 177098 996051
rect 164566 996029 164618 996035
rect 145268 995994 145324 996003
rect 145268 995929 145324 995938
rect 149108 995994 149164 996003
rect 149492 995994 149548 996003
rect 149164 995952 149492 995980
rect 149108 995929 149164 995938
rect 149492 995929 149548 995938
rect 152084 995994 152140 996003
rect 152084 995929 152086 995938
rect 144310 995437 144362 995443
rect 144310 995379 144362 995385
rect 143636 995106 143692 995115
rect 143636 995041 143692 995050
rect 141238 994549 141290 994555
rect 141236 994514 141238 994523
rect 141290 994514 141292 994523
rect 141236 994449 141292 994458
rect 140372 993774 140428 993783
rect 140372 993709 140428 993718
rect 129718 993661 129770 993667
rect 129718 993603 129770 993609
rect 138262 986409 138314 986415
rect 138262 986351 138314 986357
rect 120886 985521 120938 985527
rect 120884 985486 120886 985495
rect 120938 985486 120940 985495
rect 120884 985421 120940 985430
rect 122038 985447 122090 985453
rect 122038 985389 122090 985395
rect 118102 983819 118154 983825
rect 118102 983761 118154 983767
rect 115318 983671 115370 983677
rect 115318 983613 115370 983619
rect 106402 981596 106526 981624
rect 106402 981476 106430 981596
rect 105840 981448 106430 981476
rect 122050 981462 122078 985389
rect 138274 981462 138302 986351
rect 145282 983603 145310 995929
rect 152138 995929 152140 995938
rect 164180 995994 164236 996003
rect 164180 995929 164182 995938
rect 152086 995897 152138 995903
rect 164234 995929 164236 995938
rect 164564 995994 164566 996003
rect 164618 995994 164620 996003
rect 164564 995929 164620 995938
rect 164182 995897 164234 995903
rect 177058 995887 177086 996045
rect 177046 995881 177098 995887
rect 165620 995846 165676 995855
rect 164086 995807 164138 995813
rect 165620 995781 165622 995790
rect 164086 995749 164138 995755
rect 165674 995781 165676 995790
rect 166292 995846 166348 995855
rect 177046 995823 177098 995829
rect 178498 995813 178526 1002261
rect 208436 1000878 208492 1000887
rect 195094 1000839 195146 1000845
rect 208436 1000813 208438 1000822
rect 195094 1000781 195146 1000787
rect 208490 1000813 208492 1000822
rect 208438 1000781 208490 1000787
rect 185108 995846 185164 995855
rect 166292 995781 166348 995790
rect 178486 995807 178538 995813
rect 165622 995749 165674 995755
rect 163990 995733 164042 995739
rect 163990 995675 164042 995681
rect 152564 995254 152620 995263
rect 152564 995189 152620 995198
rect 156692 995254 156748 995263
rect 156692 995189 156748 995198
rect 159572 995254 159628 995263
rect 159572 995189 159628 995198
rect 161204 995254 161260 995263
rect 161204 995189 161260 995198
rect 146996 994662 147052 994671
rect 146996 994597 147052 994606
rect 147010 994555 147038 994597
rect 146998 994549 147050 994555
rect 146998 994491 147050 994497
rect 152578 993815 152606 995189
rect 156706 994079 156734 995189
rect 158420 994662 158476 994671
rect 158420 994597 158422 994606
rect 158474 994597 158476 994606
rect 158422 994565 158474 994571
rect 156692 994070 156748 994079
rect 156692 994005 156748 994014
rect 152566 993809 152618 993815
rect 152566 993751 152618 993757
rect 159586 993741 159614 995189
rect 159574 993735 159626 993741
rect 159574 993677 159626 993683
rect 161218 993667 161246 995189
rect 161206 993661 161258 993667
rect 161206 993603 161258 993609
rect 164002 986045 164030 995675
rect 164098 986415 164126 995749
rect 166306 995739 166334 995781
rect 184848 995804 185108 995832
rect 188084 995846 188140 995855
rect 185218 995818 185424 995832
rect 185218 995813 185438 995818
rect 185108 995781 185164 995790
rect 185206 995807 185438 995813
rect 178486 995749 178538 995755
rect 185258 995804 185438 995807
rect 187872 995804 188084 995832
rect 185206 995749 185258 995755
rect 166294 995733 166346 995739
rect 166294 995675 166346 995681
rect 170228 995698 170284 995707
rect 184176 995665 184382 995684
rect 184176 995659 184394 995665
rect 184176 995656 184342 995659
rect 170228 995633 170284 995642
rect 164086 986409 164138 986415
rect 164086 986351 164138 986357
rect 154486 986039 154538 986045
rect 154486 985981 154538 985987
rect 163990 986039 164042 986045
rect 163990 985981 164042 985987
rect 146806 985521 146858 985527
rect 146858 985469 147038 985472
rect 146806 985463 147038 985469
rect 146818 985453 147038 985463
rect 146818 985447 147050 985453
rect 146818 985444 146998 985447
rect 146998 985389 147050 985395
rect 145270 983597 145322 983603
rect 145270 983539 145322 983545
rect 154498 981462 154526 985981
rect 170242 981476 170270 995633
rect 184342 995601 184394 995607
rect 178484 994662 178540 994671
rect 178484 994597 178486 994606
rect 178538 994597 178540 994606
rect 178486 994565 178538 994571
rect 179842 993741 179870 995522
rect 180514 993963 180542 995522
rect 181152 995508 181406 995536
rect 180502 993957 180554 993963
rect 180502 993899 180554 993905
rect 181378 993815 181406 995508
rect 183010 993889 183038 995522
rect 183552 995508 183806 995536
rect 183778 995411 183806 995508
rect 183764 995402 183820 995411
rect 183764 995337 183820 995346
rect 182998 993883 183050 993889
rect 182998 993825 183050 993831
rect 181366 993809 181418 993815
rect 181366 993751 181418 993757
rect 179830 993735 179882 993741
rect 179830 993677 179882 993683
rect 185410 993667 185438 995804
rect 190368 995813 190622 995832
rect 190368 995807 190634 995813
rect 190368 995804 190582 995807
rect 188084 995781 188140 995790
rect 190582 995749 190634 995755
rect 195106 995739 195134 1000781
rect 201622 996695 201674 996701
rect 201622 996637 201674 996643
rect 195766 996547 195818 996553
rect 195766 996489 195818 996495
rect 194422 995733 194474 995739
rect 194064 995681 194422 995684
rect 194064 995675 194474 995681
rect 195094 995733 195146 995739
rect 195094 995675 195146 995681
rect 195380 995698 195436 995707
rect 194064 995656 194462 995675
rect 195778 995665 195806 996489
rect 198550 996177 198602 996183
rect 198550 996119 198602 996125
rect 198562 996003 198590 996119
rect 198646 996029 198698 996035
rect 198548 995994 198604 996003
rect 198646 995971 198698 995977
rect 198548 995929 198604 995938
rect 198658 995855 198686 995971
rect 198644 995846 198700 995855
rect 198644 995781 198700 995790
rect 198646 995733 198698 995739
rect 198646 995675 198698 995681
rect 195380 995633 195436 995642
rect 195766 995659 195818 995665
rect 189428 995550 189484 995559
rect 185794 995508 186048 995536
rect 185794 994671 185822 995508
rect 185780 994662 185836 994671
rect 185780 994597 185836 994606
rect 185794 994079 185822 994597
rect 187330 994227 187358 995522
rect 188544 995508 188894 995536
rect 189168 995508 189428 995536
rect 188866 995411 188894 995508
rect 189428 995485 189484 995494
rect 188852 995402 188908 995411
rect 188852 995337 188908 995346
rect 187316 994218 187372 994227
rect 187316 994153 187372 994162
rect 185780 994070 185836 994079
rect 185780 994005 185836 994014
rect 191554 993931 191582 995522
rect 192192 995508 192446 995536
rect 192418 995263 192446 995508
rect 192404 995254 192460 995263
rect 192404 995189 192460 995198
rect 191540 993922 191596 993931
rect 191540 993857 191596 993866
rect 185398 993661 185450 993667
rect 185398 993603 185450 993609
rect 186934 985373 186986 985379
rect 186934 985315 186986 985321
rect 170242 981448 170736 981476
rect 186946 981462 186974 985315
rect 195394 983529 195422 995633
rect 195766 995601 195818 995607
rect 198658 994967 198686 995675
rect 201634 995263 201662 996637
rect 205652 996586 205708 996595
rect 205652 996521 205654 996530
rect 205706 996521 205708 996530
rect 211700 996586 211756 996595
rect 211700 996521 211702 996530
rect 205654 996489 205706 996495
rect 211754 996521 211756 996530
rect 211702 996489 211754 996495
rect 203638 996177 203690 996183
rect 203636 996142 203638 996151
rect 214102 996177 214154 996183
rect 203690 996142 203692 996151
rect 203636 996077 203692 996086
rect 213332 996142 213388 996151
rect 214102 996119 214154 996125
rect 213332 996077 213334 996086
rect 213386 996077 213388 996086
rect 213334 996045 213386 996051
rect 202966 996029 203018 996035
rect 202964 995994 202966 996003
rect 213046 996029 213098 996035
rect 203018 995994 203020 996003
rect 202964 995929 203020 995938
rect 206612 995994 206668 996003
rect 213046 995971 213098 995977
rect 206612 995929 206668 995938
rect 201812 995846 201868 995855
rect 201812 995781 201868 995790
rect 204980 995846 205036 995855
rect 204980 995781 204982 995790
rect 201718 995659 201770 995665
rect 201718 995601 201770 995607
rect 201620 995254 201676 995263
rect 201620 995189 201676 995198
rect 198644 994958 198700 994967
rect 198644 994893 198700 994902
rect 201730 993963 201758 995601
rect 201826 995559 201854 995781
rect 205034 995781 205036 995790
rect 204982 995749 205034 995755
rect 206626 995739 206654 995929
rect 206614 995733 206666 995739
rect 206614 995675 206666 995681
rect 206996 995698 207052 995707
rect 206996 995633 206998 995642
rect 207050 995633 207052 995642
rect 206998 995601 207050 995607
rect 201812 995550 201868 995559
rect 201812 995485 201868 995494
rect 212660 995550 212716 995559
rect 212660 995485 212716 995494
rect 207380 995254 207436 995263
rect 207380 995189 207436 995198
rect 211028 995254 211084 995263
rect 211028 995189 211084 995198
rect 207284 995106 207340 995115
rect 207284 995041 207340 995050
rect 201718 993957 201770 993963
rect 201718 993899 201770 993905
rect 207298 993889 207326 995041
rect 207394 994227 207422 995189
rect 207380 994218 207436 994227
rect 207380 994153 207436 994162
rect 207286 993883 207338 993889
rect 207286 993825 207338 993831
rect 211042 993741 211070 995189
rect 212674 993815 212702 995485
rect 212662 993809 212714 993815
rect 212662 993751 212714 993757
rect 211030 993735 211082 993741
rect 211030 993677 211082 993683
rect 213058 986341 213086 995971
rect 214114 995887 214142 996119
rect 216886 996029 216938 996035
rect 215636 995994 215692 996003
rect 215636 995929 215638 995938
rect 215690 995929 215692 995938
rect 216884 995994 216886 996003
rect 216938 995994 216940 996003
rect 216884 995929 216940 995938
rect 218902 995955 218954 995961
rect 215638 995897 215690 995903
rect 218902 995897 218954 995903
rect 214102 995881 214154 995887
rect 214100 995846 214102 995855
rect 214154 995846 214156 995855
rect 214100 995781 214156 995790
rect 218914 995707 218942 995897
rect 218900 995698 218956 995707
rect 218900 995633 218956 995642
rect 221890 987229 221918 1005105
rect 223138 987821 223166 1005253
rect 246836 1005170 246892 1005179
rect 246836 1005105 246892 1005114
rect 246550 1002467 246602 1002473
rect 246550 1002409 246602 1002415
rect 246562 999532 246590 1002409
rect 246742 1002319 246794 1002325
rect 246742 1002261 246794 1002267
rect 246466 999504 246590 999532
rect 246646 999581 246698 999587
rect 246646 999523 246698 999529
rect 246466 995855 246494 999504
rect 246550 999433 246602 999439
rect 246550 999375 246602 999381
rect 239540 995846 239596 995855
rect 239280 995804 239540 995832
rect 246452 995846 246508 995855
rect 240576 995813 240926 995832
rect 245424 995813 245726 995832
rect 240576 995807 240938 995813
rect 240576 995804 240886 995807
rect 239540 995781 239596 995790
rect 245424 995807 245738 995813
rect 245424 995804 245686 995807
rect 240886 995749 240938 995755
rect 246562 995813 246590 999375
rect 246452 995781 246508 995790
rect 246550 995807 246602 995813
rect 245686 995749 245738 995755
rect 246550 995749 246602 995755
rect 246658 995739 246686 999523
rect 246754 995887 246782 1002261
rect 246742 995881 246794 995887
rect 246742 995823 246794 995829
rect 243190 995733 243242 995739
rect 241844 995698 241900 995707
rect 241776 995656 241844 995684
rect 242976 995681 243190 995684
rect 242976 995675 243242 995681
rect 246646 995733 246698 995739
rect 246646 995675 246698 995681
rect 242976 995656 243230 995675
rect 241844 995633 241900 995642
rect 240212 995550 240268 995559
rect 231264 995508 231518 995536
rect 231936 995508 232190 995536
rect 231490 994227 231518 995508
rect 231476 994218 231532 994227
rect 231476 994153 231532 994162
rect 232162 993889 232190 995508
rect 232150 993883 232202 993889
rect 232150 993825 232202 993831
rect 232546 993741 232574 995522
rect 234370 993815 234398 995522
rect 234946 993963 234974 995522
rect 235584 995508 235838 995536
rect 236256 995517 236510 995536
rect 236256 995511 236522 995517
rect 236256 995508 236470 995511
rect 235810 995443 235838 995508
rect 236470 995453 236522 995459
rect 235798 995437 235850 995443
rect 235798 995379 235850 995385
rect 234934 993957 234986 993963
rect 234934 993899 234986 993905
rect 234358 993809 234410 993815
rect 234358 993751 234410 993757
rect 232534 993735 232586 993741
rect 232534 993677 232586 993683
rect 236770 993667 236798 995522
rect 237442 995115 237470 995522
rect 237428 995106 237484 995115
rect 237428 995041 237484 995050
rect 237442 994079 237470 995041
rect 238690 994671 238718 995522
rect 239952 995508 240212 995536
rect 246850 995536 246878 1005105
rect 254036 1002506 254092 1002515
rect 254036 1002441 254038 1002450
rect 254090 1002441 254092 1002450
rect 254038 1002409 254090 1002415
rect 253172 1002358 253228 1002367
rect 253172 1002293 253174 1002302
rect 253226 1002293 253228 1002302
rect 253174 1002261 253226 1002267
rect 298114 999661 298142 1005369
rect 298390 1005353 298442 1005359
rect 309622 1005353 309674 1005359
rect 298390 1005295 298442 1005301
rect 307988 1005318 308044 1005327
rect 298294 1005279 298346 1005285
rect 298294 1005221 298346 1005227
rect 298102 999655 298154 999661
rect 262114 999615 262238 999643
rect 262114 999587 262142 999615
rect 262102 999581 262154 999587
rect 262102 999523 262154 999529
rect 250486 999507 250538 999513
rect 250486 999449 250538 999455
rect 240212 995485 240268 995494
rect 243586 995263 243614 995522
rect 246466 995508 246878 995536
rect 243572 995254 243628 995263
rect 243572 995189 243628 995198
rect 238676 994662 238732 994671
rect 238676 994597 238732 994606
rect 237428 994070 237484 994079
rect 237428 994005 237484 994014
rect 236758 993661 236810 993667
rect 236758 993603 236810 993609
rect 246466 990929 246494 995508
rect 247606 995437 247658 995443
rect 247604 995402 247606 995411
rect 247658 995402 247660 995411
rect 247604 995337 247660 995346
rect 250498 995263 250526 999449
rect 259606 999433 259658 999439
rect 259604 999398 259606 999407
rect 259658 999398 259660 999407
rect 259604 999333 259660 999342
rect 259124 995994 259180 996003
rect 259124 995929 259180 995938
rect 261428 995994 261484 996003
rect 261428 995929 261484 995938
rect 261812 995994 261868 996003
rect 261812 995929 261868 995938
rect 259138 995887 259166 995929
rect 253366 995881 253418 995887
rect 259126 995881 259178 995887
rect 253366 995823 253418 995829
rect 254804 995846 254860 995855
rect 250484 995254 250540 995263
rect 250676 995254 250732 995263
rect 250484 995189 250540 995198
rect 250594 995212 250676 995240
rect 250594 995092 250622 995212
rect 250676 995189 250732 995198
rect 250498 995064 250622 995092
rect 250498 993963 250526 995064
rect 250486 993957 250538 993963
rect 250486 993899 250538 993905
rect 253378 993889 253406 995823
rect 254804 995781 254860 995790
rect 255956 995846 256012 995855
rect 259126 995823 259178 995829
rect 260468 995846 260524 995855
rect 255956 995781 256012 995790
rect 260468 995781 260524 995790
rect 254818 995517 254846 995781
rect 255970 995559 255998 995781
rect 255956 995550 256012 995559
rect 254806 995511 254858 995517
rect 255956 995485 256012 995494
rect 254806 995453 254858 995459
rect 260482 994671 260510 995781
rect 260468 994662 260524 994671
rect 260468 994597 260524 994606
rect 253366 993883 253418 993889
rect 253366 993825 253418 993831
rect 261442 993815 261470 995929
rect 261826 994227 261854 995929
rect 262210 995147 262238 999615
rect 298102 999597 298154 999603
rect 263060 999546 263116 999555
rect 263060 999481 263062 999490
rect 263114 999481 263116 999490
rect 298102 999507 298154 999513
rect 263062 999449 263114 999455
rect 298102 999449 298154 999455
rect 266806 996177 266858 996183
rect 265940 996142 265996 996151
rect 265940 996077 265942 996086
rect 265994 996077 265996 996086
rect 266804 996142 266806 996151
rect 266858 996142 266860 996151
rect 266804 996077 266860 996086
rect 265942 996045 265994 996051
rect 265078 996029 265130 996035
rect 265076 995994 265078 996003
rect 265130 995994 265132 996003
rect 265076 995929 265132 995938
rect 266996 995994 267052 996003
rect 266996 995929 266998 995938
rect 267050 995929 267052 995938
rect 266998 995897 267050 995903
rect 268628 995846 268684 995855
rect 268628 995781 268684 995790
rect 273620 995846 273676 995855
rect 292436 995846 292492 995855
rect 283536 995813 283742 995832
rect 283536 995807 283754 995813
rect 283536 995804 283702 995807
rect 273620 995781 273676 995790
rect 264020 995402 264076 995411
rect 264020 995337 264076 995346
rect 262198 995141 262250 995147
rect 262198 995083 262250 995089
rect 261812 994218 261868 994227
rect 261812 994153 261868 994162
rect 261430 993809 261482 993815
rect 261430 993751 261482 993757
rect 264034 993741 264062 995337
rect 264022 993735 264074 993741
rect 264022 993677 264074 993683
rect 241942 990923 241994 990929
rect 241942 990865 241994 990871
rect 246454 990923 246506 990929
rect 246454 990865 246506 990871
rect 241954 987895 241982 990865
rect 241942 987889 241994 987895
rect 241942 987831 241994 987837
rect 223126 987815 223178 987821
rect 223126 987757 223178 987763
rect 235606 987815 235658 987821
rect 235606 987757 235658 987763
rect 236278 987815 236330 987821
rect 236278 987757 236330 987763
rect 219478 987223 219530 987229
rect 219478 987165 219530 987171
rect 221878 987223 221930 987229
rect 221878 987165 221930 987171
rect 203158 986335 203210 986341
rect 203158 986277 203210 986283
rect 213046 986335 213098 986341
rect 213046 986277 213098 986283
rect 201526 985521 201578 985527
rect 201622 985521 201674 985527
rect 201578 985469 201622 985472
rect 201526 985463 201674 985469
rect 201538 985444 201662 985463
rect 195382 983523 195434 983529
rect 195382 983465 195434 983471
rect 203170 981462 203198 986277
rect 218914 985592 219038 985620
rect 218914 985527 218942 985592
rect 218902 985521 218954 985527
rect 218902 985463 218954 985469
rect 219010 985379 219038 985592
rect 218998 985373 219050 985379
rect 218998 985315 219050 985321
rect 217366 983523 217418 983529
rect 217366 983465 217418 983471
rect 130390 981081 130442 981087
rect 106498 981013 106622 981032
rect 130390 981023 130442 981029
rect 161300 981046 161356 981055
rect 106486 981007 106634 981013
rect 106538 981004 106582 981007
rect 106486 980949 106538 980955
rect 106582 980949 106634 980955
rect 130402 980939 130430 981023
rect 161300 980981 161302 980990
rect 161354 980981 161356 980990
rect 171284 981046 171340 981055
rect 171284 980981 171340 980990
rect 161302 980949 161354 980955
rect 130390 980933 130442 980939
rect 130390 980875 130442 980881
rect 171298 980865 171326 980981
rect 178486 980933 178538 980939
rect 178486 980875 178538 980881
rect 146902 980859 146954 980865
rect 146902 980801 146954 980807
rect 171286 980859 171338 980865
rect 171286 980801 171338 980807
rect 106486 980785 106538 980791
rect 106582 980785 106634 980791
rect 106538 980733 106582 980736
rect 106486 980727 106634 980733
rect 146806 980785 146858 980791
rect 146914 980736 146942 980801
rect 178498 980791 178526 980875
rect 217378 980791 217406 983465
rect 219490 981462 219518 987165
rect 235618 981462 235646 987757
rect 236290 983529 236318 987757
rect 239158 985447 239210 985453
rect 239158 985389 239210 985395
rect 251830 985447 251882 985453
rect 251830 985389 251882 985395
rect 239060 985338 239116 985347
rect 239170 985305 239198 985389
rect 239540 985338 239596 985347
rect 239060 985273 239116 985282
rect 239158 985299 239210 985305
rect 239074 985231 239102 985273
rect 239540 985273 239596 985282
rect 239158 985241 239210 985247
rect 239554 985231 239582 985273
rect 239062 985225 239114 985231
rect 239542 985225 239594 985231
rect 239062 985167 239114 985173
rect 239156 985190 239212 985199
rect 239542 985167 239594 985173
rect 239732 985190 239788 985199
rect 239156 985125 239158 985134
rect 239210 985125 239212 985134
rect 239732 985125 239734 985134
rect 239158 985093 239210 985099
rect 239786 985125 239788 985134
rect 239734 985093 239786 985099
rect 239062 985077 239114 985083
rect 239446 985077 239498 985083
rect 239114 985025 239446 985028
rect 239062 985019 239498 985025
rect 239074 985000 239486 985019
rect 236278 983523 236330 983529
rect 236278 983465 236330 983471
rect 251842 981462 251870 985389
rect 268642 981476 268670 995781
rect 273634 986193 273662 995781
rect 292176 995804 292436 995832
rect 293588 995846 293644 995855
rect 293376 995804 293588 995832
rect 292436 995781 292492 995790
rect 297072 995813 297374 995832
rect 298114 995813 298142 999449
rect 298198 996547 298250 996553
rect 298198 996489 298250 996495
rect 297072 995807 297386 995813
rect 297072 995804 297334 995807
rect 293588 995781 293644 995790
rect 283702 995749 283754 995755
rect 297334 995749 297386 995755
rect 298102 995807 298154 995813
rect 298102 995749 298154 995755
rect 298210 995739 298238 996489
rect 298306 995855 298334 1005221
rect 298292 995846 298348 995855
rect 298292 995781 298348 995790
rect 294838 995733 294890 995739
rect 273716 995698 273772 995707
rect 291092 995698 291148 995707
rect 286560 995665 286814 995684
rect 286560 995659 286826 995665
rect 286560 995656 286774 995659
rect 273716 995633 273772 995642
rect 273730 986415 273758 995633
rect 290880 995656 291092 995684
rect 294576 995681 294838 995684
rect 294576 995675 294890 995681
rect 298198 995733 298250 995739
rect 298198 995675 298250 995681
rect 294576 995656 294878 995675
rect 298402 995665 298430 1005295
rect 307988 1005253 307990 1005262
rect 308042 1005253 308044 1005262
rect 309620 1005318 309622 1005327
rect 309674 1005318 309676 1005327
rect 309620 1005253 309676 1005262
rect 318644 1005318 318700 1005327
rect 318644 1005253 318646 1005262
rect 307990 1005221 308042 1005227
rect 318698 1005253 318700 1005262
rect 318646 1005221 318698 1005227
rect 325474 1005211 325502 1005401
rect 364202 1005401 364204 1005410
rect 365012 1005466 365014 1005475
rect 365066 1005466 365068 1005475
rect 365012 1005401 365068 1005410
rect 371062 1005427 371114 1005433
rect 364150 1005369 364202 1005375
rect 371062 1005369 371114 1005375
rect 366742 1005353 366794 1005359
rect 365780 1005318 365836 1005327
rect 331126 1005279 331178 1005285
rect 365780 1005253 365782 1005262
rect 331126 1005221 331178 1005227
rect 365834 1005253 365836 1005262
rect 366740 1005318 366742 1005327
rect 366794 1005318 366796 1005327
rect 366740 1005253 366796 1005262
rect 365782 1005221 365834 1005227
rect 299926 1005205 299978 1005211
rect 315190 1005205 315242 1005211
rect 299926 1005147 299978 1005153
rect 315188 1005170 315190 1005179
rect 325462 1005205 325514 1005211
rect 315242 1005170 315244 1005179
rect 299638 1002541 299690 1002547
rect 299638 1002483 299690 1002489
rect 299542 1002467 299594 1002473
rect 299542 1002409 299594 1002415
rect 298580 1002358 298636 1002367
rect 298580 1002293 298636 1002302
rect 298486 999655 298538 999661
rect 298486 999597 298538 999603
rect 298390 995659 298442 995665
rect 291092 995633 291148 995642
rect 286774 995601 286826 995607
rect 298390 995601 298442 995607
rect 298498 995591 298526 999597
rect 287542 995585 287594 995591
rect 282850 993667 282878 995522
rect 284160 995508 284414 995536
rect 287184 995533 287542 995536
rect 298486 995585 298538 995591
rect 291764 995550 291820 995559
rect 287184 995527 287594 995533
rect 284386 995443 284414 995508
rect 284374 995437 284426 995443
rect 284374 995379 284426 995385
rect 286018 994227 286046 995522
rect 287184 995508 287582 995527
rect 287856 995517 287966 995536
rect 287856 995511 287978 995517
rect 287856 995508 287926 995511
rect 288384 995508 288446 995536
rect 287926 995453 287978 995459
rect 286004 994218 286060 994227
rect 286004 994153 286060 994162
rect 279286 993661 279338 993667
rect 279284 993626 279286 993635
rect 282838 993661 282890 993667
rect 279338 993626 279340 993635
rect 288418 993635 288446 995508
rect 288802 995508 289056 995536
rect 288802 995115 288830 995508
rect 288788 995106 288844 995115
rect 288788 995041 288844 995050
rect 288802 994079 288830 995041
rect 290338 994523 290366 995522
rect 291504 995508 291764 995536
rect 295200 995508 295454 995536
rect 298486 995527 298538 995533
rect 291764 995485 291820 995494
rect 290324 994514 290380 994523
rect 290324 994449 290380 994458
rect 295426 994375 295454 995508
rect 295412 994366 295468 994375
rect 295412 994301 295468 994310
rect 288788 994070 288844 994079
rect 288788 994005 288844 994014
rect 282838 993603 282890 993609
rect 288404 993626 288460 993635
rect 279284 993561 279340 993570
rect 288404 993561 288460 993570
rect 288418 992155 288446 993561
rect 288404 992146 288460 992155
rect 288404 992081 288460 992090
rect 298594 991669 298622 1002293
rect 299446 999433 299498 999439
rect 299446 999375 299498 999381
rect 299458 995887 299486 999375
rect 299446 995881 299498 995887
rect 299446 995823 299498 995829
rect 299554 995707 299582 1002409
rect 299540 995698 299596 995707
rect 299540 995633 299596 995642
rect 299650 995559 299678 1002483
rect 299830 1002393 299882 1002399
rect 299830 1002335 299882 1002341
rect 299734 1002319 299786 1002325
rect 299734 1002261 299786 1002267
rect 299746 996003 299774 1002261
rect 299732 995994 299788 996003
rect 299732 995929 299788 995938
rect 299636 995550 299692 995559
rect 299842 995517 299870 1002335
rect 299636 995485 299692 995494
rect 299830 995511 299882 995517
rect 299830 995453 299882 995459
rect 299938 995443 299966 1005147
rect 325462 1005147 325514 1005153
rect 315188 1005105 315244 1005114
rect 307606 1002541 307658 1002547
rect 305588 1002506 305644 1002515
rect 305588 1002441 305590 1002450
rect 305642 1002441 305644 1002450
rect 307604 1002506 307606 1002515
rect 307658 1002506 307660 1002515
rect 307604 1002441 307660 1002450
rect 305590 1002409 305642 1002415
rect 306550 1002393 306602 1002399
rect 304724 1002358 304780 1002367
rect 304724 1002293 304726 1002302
rect 304778 1002293 304780 1002302
rect 306548 1002358 306550 1002367
rect 306602 1002358 306604 1002367
rect 306548 1002293 306604 1002302
rect 304726 1002261 304778 1002267
rect 311156 999546 311212 999555
rect 311156 999481 311158 999490
rect 311210 999481 311212 999490
rect 311158 999449 311210 999455
rect 310294 999433 310346 999439
rect 310292 999398 310294 999407
rect 310346 999398 310348 999407
rect 310292 999333 310348 999342
rect 320950 997953 321002 997959
rect 320950 997895 321002 997901
rect 320182 996473 320234 996479
rect 320182 996415 320234 996421
rect 318646 996177 318698 996183
rect 317108 996142 317164 996151
rect 317108 996077 317110 996086
rect 317162 996077 317164 996086
rect 318644 996142 318646 996151
rect 318698 996142 318700 996151
rect 318644 996077 318700 996086
rect 317110 996045 317162 996051
rect 320194 996035 320222 996415
rect 320962 996109 320990 997895
rect 331138 997885 331166 1005221
rect 371074 1005211 371102 1005369
rect 371842 1005211 371870 1005665
rect 383638 1005649 383690 1005655
rect 439234 1005600 439262 1005739
rect 440662 1005723 440714 1005729
rect 440662 1005665 440714 1005671
rect 446422 1005723 446474 1005729
rect 446422 1005665 446474 1005671
rect 383638 1005591 383690 1005597
rect 380566 1005501 380618 1005507
rect 380566 1005443 380618 1005449
rect 380470 1005427 380522 1005433
rect 380470 1005369 380522 1005375
rect 380374 1005353 380426 1005359
rect 380374 1005295 380426 1005301
rect 380278 1005279 380330 1005285
rect 380278 1005221 380330 1005227
rect 331222 1005205 331274 1005211
rect 363478 1005205 363530 1005211
rect 331222 1005147 331274 1005153
rect 363476 1005170 363478 1005179
rect 371062 1005205 371114 1005211
rect 363530 1005170 363532 1005179
rect 331126 997879 331178 997885
rect 331126 997821 331178 997827
rect 320950 996103 321002 996109
rect 320950 996045 321002 996051
rect 316342 996029 316394 996035
rect 313844 995994 313900 996003
rect 313844 995929 313900 995938
rect 316340 995994 316342 996003
rect 320182 996029 320234 996035
rect 316394 995994 316396 996003
rect 320182 995971 320234 995977
rect 326804 995994 326860 996003
rect 316340 995929 316396 995938
rect 326804 995929 326860 995938
rect 310292 995698 310348 995707
rect 310292 995633 310348 995642
rect 299926 995437 299978 995443
rect 299926 995379 299978 995385
rect 310306 994523 310334 995633
rect 311060 995254 311116 995263
rect 311060 995189 311116 995198
rect 310292 994514 310348 994523
rect 310292 994449 310348 994458
rect 311074 994227 311102 995189
rect 311060 994218 311116 994227
rect 311060 994153 311116 994162
rect 313858 993667 313886 995929
rect 323924 995698 323980 995707
rect 323924 995633 323980 995642
rect 313846 993661 313898 993667
rect 313846 993603 313898 993609
rect 285142 991663 285194 991669
rect 285142 991605 285194 991611
rect 298582 991663 298634 991669
rect 298582 991605 298634 991611
rect 273718 986409 273770 986415
rect 273718 986351 273770 986357
rect 273622 986187 273674 986193
rect 273622 986129 273674 986135
rect 284278 986187 284330 986193
rect 284278 986129 284330 986135
rect 279382 985373 279434 985379
rect 279382 985315 279434 985321
rect 279394 982345 279422 985315
rect 273622 982339 273674 982345
rect 273622 982281 273674 982287
rect 279382 982339 279434 982345
rect 279382 982281 279434 982287
rect 268176 981448 268670 981476
rect 247618 980865 247742 980884
rect 238966 980859 239018 980865
rect 238966 980801 239018 980807
rect 247606 980859 247754 980865
rect 247658 980856 247702 980859
rect 247606 980801 247658 980807
rect 247702 980801 247754 980807
rect 146858 980733 146942 980736
rect 146806 980727 146942 980733
rect 178486 980785 178538 980791
rect 178486 980727 178538 980733
rect 217366 980785 217418 980791
rect 217366 980727 217418 980733
rect 217558 980785 217610 980791
rect 217654 980785 217706 980791
rect 217610 980745 217654 980773
rect 217558 980727 217610 980733
rect 218902 980785 218954 980791
rect 217654 980727 217706 980733
rect 218900 980750 218902 980759
rect 238978 980759 239006 980801
rect 273634 980791 273662 982281
rect 284290 981462 284318 986129
rect 285154 985379 285182 991605
rect 323938 986415 323966 995633
rect 326818 986489 326846 995929
rect 331234 992187 331262 1005147
rect 371062 1005147 371114 1005153
rect 371830 1005205 371882 1005211
rect 371830 1005147 371882 1005153
rect 380182 1005205 380234 1005211
rect 380182 1005147 380234 1005153
rect 363476 1005105 363532 1005114
rect 359926 1004021 359978 1004027
rect 359924 1003986 359926 1003995
rect 380086 1004021 380138 1004027
rect 359978 1003986 359980 1003995
rect 380086 1003963 380138 1003969
rect 359924 1003921 359980 1003930
rect 359062 1003873 359114 1003879
rect 358388 1003838 358444 1003847
rect 358388 1003773 358390 1003782
rect 358442 1003773 358444 1003782
rect 359060 1003838 359062 1003847
rect 377494 1003873 377546 1003879
rect 359114 1003838 359116 1003847
rect 377494 1003815 377546 1003821
rect 359060 1003773 359116 1003782
rect 377398 1003799 377450 1003805
rect 358390 1003741 358442 1003747
rect 377398 1003741 377450 1003747
rect 360694 1003725 360746 1003731
rect 360692 1003690 360694 1003699
rect 377302 1003725 377354 1003731
rect 360746 1003690 360748 1003699
rect 377302 1003667 377354 1003673
rect 360692 1003625 360748 1003634
rect 361556 1000878 361612 1000887
rect 361556 1000813 361558 1000822
rect 361610 1000813 361612 1000822
rect 361558 1000781 361610 1000787
rect 377314 999661 377342 1003667
rect 377302 999655 377354 999661
rect 377302 999597 377354 999603
rect 356278 998101 356330 998107
rect 356276 998066 356278 998075
rect 368758 998101 368810 998107
rect 356330 998066 356332 998075
rect 356276 998001 356332 998010
rect 357044 998066 357100 998075
rect 368758 998043 368810 998049
rect 357044 998001 357046 998010
rect 357098 998001 357100 998010
rect 368662 998027 368714 998033
rect 357046 997969 357098 997975
rect 368662 997969 368714 997975
rect 367894 997953 367946 997959
rect 367892 997918 367894 997927
rect 367946 997918 367948 997927
rect 367892 997853 367948 997862
rect 367126 996473 367178 996479
rect 367126 996415 367178 996421
rect 367138 996035 367166 996415
rect 367126 996029 367178 996035
rect 362324 995994 362380 996003
rect 362324 995929 362380 995938
rect 367124 995994 367126 996003
rect 367178 995994 367180 996003
rect 367124 995929 367180 995938
rect 343892 995698 343948 995707
rect 343892 995633 343948 995642
rect 343906 995221 343934 995633
rect 343894 995215 343946 995221
rect 343894 995157 343946 995163
rect 362338 993667 362366 995929
rect 368674 993889 368702 997969
rect 368662 993883 368714 993889
rect 368662 993825 368714 993831
rect 368770 993741 368798 998043
rect 369044 997918 369100 997927
rect 369044 997853 369046 997862
rect 369098 997853 369100 997862
rect 369046 997821 369098 997827
rect 377410 996923 377438 1003741
rect 377398 996917 377450 996923
rect 377398 996859 377450 996865
rect 377506 996627 377534 1003815
rect 377494 996621 377546 996627
rect 377494 996563 377546 996569
rect 380098 996572 380126 1003963
rect 380194 999587 380222 1005147
rect 380182 999581 380234 999587
rect 380182 999523 380234 999529
rect 374518 996547 374570 996553
rect 380098 996544 380222 996572
rect 374518 996489 374570 996495
rect 371542 996177 371594 996183
rect 371542 996119 371594 996125
rect 370580 995994 370636 996003
rect 370580 995929 370582 995938
rect 370634 995929 370636 995938
rect 370582 995897 370634 995903
rect 371348 995846 371404 995855
rect 371348 995781 371350 995790
rect 371402 995781 371404 995790
rect 371350 995749 371402 995755
rect 371554 995707 371582 996119
rect 374422 995807 374474 995813
rect 374422 995749 374474 995755
rect 371540 995698 371596 995707
rect 371540 995633 371596 995642
rect 368758 993735 368810 993741
rect 368758 993677 368810 993683
rect 362326 993661 362378 993667
rect 362326 993603 362378 993609
rect 331222 992181 331274 992187
rect 331222 992123 331274 992129
rect 332566 992181 332618 992187
rect 332566 992123 332618 992129
rect 326806 986483 326858 986489
rect 326806 986425 326858 986431
rect 300502 986409 300554 986415
rect 300502 986351 300554 986357
rect 323926 986409 323978 986415
rect 323926 986351 323978 986357
rect 285142 985373 285194 985379
rect 285142 985315 285194 985321
rect 300514 981462 300542 986351
rect 316726 985225 316778 985231
rect 316726 985167 316778 985173
rect 316738 981462 316766 985167
rect 332578 981476 332606 992123
rect 374434 986563 374462 995749
rect 374530 995221 374558 996489
rect 377300 995994 377356 996003
rect 374614 995955 374666 995961
rect 377300 995929 377356 995938
rect 374614 995897 374666 995903
rect 374518 995215 374570 995221
rect 374518 995157 374570 995163
rect 374422 986557 374474 986563
rect 374422 986499 374474 986505
rect 349174 986483 349226 986489
rect 349174 986425 349226 986431
rect 332578 981448 332976 981476
rect 349186 981462 349214 986425
rect 374626 986415 374654 995897
rect 377314 986489 377342 995929
rect 380194 995855 380222 996544
rect 380180 995846 380236 995855
rect 380180 995781 380236 995790
rect 380290 995707 380318 1005221
rect 380386 999513 380414 1005295
rect 380482 999957 380510 1005369
rect 380470 999951 380522 999957
rect 380470 999893 380522 999899
rect 380374 999507 380426 999513
rect 380374 999449 380426 999455
rect 380578 999439 380606 1005443
rect 383446 1000839 383498 1000845
rect 383446 1000781 383498 1000787
rect 383254 999951 383306 999957
rect 383254 999893 383306 999899
rect 383158 999655 383210 999661
rect 383158 999597 383210 999603
rect 382966 999507 383018 999513
rect 382966 999449 383018 999455
rect 380566 999433 380618 999439
rect 380566 999375 380618 999381
rect 381718 997953 381770 997959
rect 381718 997895 381770 997901
rect 381730 996109 381758 997895
rect 382870 996917 382922 996923
rect 382870 996859 382922 996865
rect 382774 996621 382826 996627
rect 382774 996563 382826 996569
rect 381718 996103 381770 996109
rect 381718 996045 381770 996051
rect 380276 995698 380332 995707
rect 380276 995633 380332 995642
rect 382786 994999 382814 996563
rect 382882 995443 382910 996859
rect 382978 995887 383006 999449
rect 382966 995881 383018 995887
rect 382966 995823 383018 995829
rect 383170 995517 383198 999597
rect 383266 995591 383294 999893
rect 383350 999581 383402 999587
rect 383350 999523 383402 999529
rect 383362 995961 383390 999523
rect 383350 995955 383402 995961
rect 383350 995897 383402 995903
rect 383458 995665 383486 1000781
rect 383542 999433 383594 999439
rect 383542 999375 383594 999381
rect 383554 995739 383582 999375
rect 383650 995813 383678 1005591
rect 439138 1005572 439262 1005600
rect 430774 1005501 430826 1005507
rect 430870 1005501 430922 1005507
rect 430774 1005443 430826 1005449
rect 430868 1005466 430870 1005475
rect 430922 1005466 430924 1005475
rect 439138 1005452 439166 1005572
rect 424534 1005353 424586 1005359
rect 424532 1005318 424534 1005327
rect 430786 1005327 430814 1005443
rect 430868 1005401 430924 1005410
rect 439042 1005424 439166 1005452
rect 439222 1005427 439274 1005433
rect 424586 1005318 424588 1005327
rect 424532 1005253 424588 1005262
rect 425300 1005318 425356 1005327
rect 425300 1005253 425302 1005262
rect 425354 1005253 425356 1005262
rect 430772 1005318 430828 1005327
rect 439042 1005285 439070 1005424
rect 439222 1005369 439274 1005375
rect 439414 1005427 439466 1005433
rect 439414 1005369 439466 1005375
rect 430772 1005253 430828 1005262
rect 439030 1005279 439082 1005285
rect 425302 1005221 425354 1005227
rect 439030 1005221 439082 1005227
rect 439234 1005211 439262 1005369
rect 426070 1005205 426122 1005211
rect 426068 1005170 426070 1005179
rect 437590 1005205 437642 1005211
rect 426122 1005170 426124 1005179
rect 426068 1005105 426124 1005114
rect 433172 1005170 433228 1005179
rect 433172 1005105 433174 1005114
rect 433226 1005105 433228 1005114
rect 435572 1005170 435628 1005179
rect 437878 1005205 437930 1005211
rect 437642 1005153 437878 1005156
rect 437590 1005147 437930 1005153
rect 439222 1005205 439274 1005211
rect 439222 1005147 439274 1005153
rect 437602 1005128 437918 1005147
rect 435572 1005105 435628 1005114
rect 433174 1005073 433226 1005079
rect 435586 1005063 435614 1005105
rect 435574 1005057 435626 1005063
rect 435574 1004999 435626 1005005
rect 423380 1003986 423436 1003995
rect 423380 1003921 423382 1003930
rect 423434 1003921 423436 1003930
rect 423382 1003889 423434 1003895
rect 426454 1003873 426506 1003879
rect 426452 1003838 426454 1003847
rect 426506 1003838 426508 1003847
rect 422518 1003799 422570 1003805
rect 426452 1003773 426508 1003782
rect 422518 1003741 422570 1003747
rect 399958 999433 400010 999439
rect 399958 999375 400010 999381
rect 388820 995846 388876 995855
rect 384418 995813 384672 995832
rect 383638 995807 383690 995813
rect 383638 995749 383690 995755
rect 384406 995807 384672 995813
rect 384458 995804 384672 995807
rect 385968 995813 386078 995832
rect 385968 995807 386090 995813
rect 385968 995804 386038 995807
rect 384406 995749 384458 995755
rect 388876 995804 388992 995832
rect 389410 995813 389664 995832
rect 389398 995807 389664 995813
rect 388820 995781 388876 995790
rect 386038 995749 386090 995755
rect 389450 995804 389664 995807
rect 396336 995813 396638 995832
rect 399970 995813 399998 999375
rect 422530 995855 422558 1003741
rect 428086 1003725 428138 1003731
rect 428084 1003690 428086 1003699
rect 428138 1003690 428140 1003699
rect 428084 1003625 428140 1003634
rect 434132 1001174 434188 1001183
rect 434132 1001109 434134 1001118
rect 434186 1001109 434188 1001118
rect 434134 1001077 434186 1001083
rect 432500 1001026 432556 1001035
rect 432500 1000961 432502 1000970
rect 432554 1000961 432556 1000970
rect 432502 1000929 432554 1000935
rect 428950 1000913 429002 1000919
rect 427316 1000878 427372 1000887
rect 427316 1000813 427318 1000822
rect 427370 1000813 427372 1000822
rect 428948 1000878 428950 1000887
rect 429002 1000878 429004 1000887
rect 428948 1000813 429004 1000822
rect 427318 1000781 427370 1000787
rect 436340 996290 436396 996299
rect 436340 996225 436396 996234
rect 436354 996183 436382 996225
rect 436342 996177 436394 996183
rect 436438 996177 436490 996183
rect 436342 996119 436394 996125
rect 436436 996142 436438 996151
rect 436490 996142 436492 996151
rect 436436 996077 436492 996086
rect 439426 996035 439454 1005369
rect 440674 1005063 440702 1005665
rect 446434 1005507 446462 1005665
rect 466486 1005575 466538 1005581
rect 466486 1005517 466538 1005523
rect 446326 1005501 446378 1005507
rect 446326 1005443 446378 1005449
rect 446422 1005501 446474 1005507
rect 446422 1005443 446474 1005449
rect 440662 1005057 440714 1005063
rect 440662 1004999 440714 1005005
rect 440674 996109 440702 1004999
rect 446338 1002325 446366 1005443
rect 460822 1005353 460874 1005359
rect 460822 1005295 460874 1005301
rect 453334 1003947 453386 1003953
rect 453334 1003889 453386 1003895
rect 446326 1002319 446378 1002325
rect 446326 1002261 446378 1002267
rect 453346 1000475 453374 1003889
rect 453334 1000469 453386 1000475
rect 453334 1000411 453386 1000417
rect 460834 1000401 460862 1005295
rect 463702 1003873 463754 1003879
rect 463702 1003815 463754 1003821
rect 461014 1003799 461066 1003805
rect 461014 1003741 461066 1003747
rect 460918 1002245 460970 1002251
rect 460918 1002187 460970 1002193
rect 460822 1000395 460874 1000401
rect 460822 1000337 460874 1000343
rect 460822 999359 460874 999365
rect 460822 999301 460874 999307
rect 440662 996103 440714 996109
rect 440662 996045 440714 996051
rect 434134 996029 434186 996035
rect 429716 995994 429772 996003
rect 429716 995929 429772 995938
rect 434132 995994 434134 996003
rect 439414 996029 439466 996035
rect 434186 995994 434188 996003
rect 439414 995971 439466 995977
rect 445076 995994 445132 996003
rect 434132 995929 434188 995938
rect 445076 995929 445132 995938
rect 422516 995846 422572 995855
rect 396336 995807 396650 995813
rect 396336 995804 396598 995807
rect 389398 995749 389450 995755
rect 396598 995749 396650 995755
rect 399958 995807 400010 995813
rect 422516 995781 422572 995790
rect 399958 995749 400010 995755
rect 383542 995733 383594 995739
rect 387478 995733 387530 995739
rect 383542 995675 383594 995681
rect 384994 995665 385296 995684
rect 396692 995698 396748 995707
rect 387530 995681 387792 995684
rect 387478 995675 387792 995681
rect 383446 995659 383498 995665
rect 383446 995601 383498 995607
rect 384982 995659 385296 995665
rect 385034 995656 385296 995659
rect 387490 995656 387792 995675
rect 396748 995656 397008 995684
rect 396692 995633 396748 995642
rect 384982 995601 385034 995607
rect 383254 995585 383306 995591
rect 391702 995585 391754 995591
rect 383254 995527 383306 995533
rect 388066 995517 388368 995536
rect 391754 995533 392112 995536
rect 391702 995527 392112 995533
rect 383158 995511 383210 995517
rect 383158 995453 383210 995459
rect 388054 995511 388368 995517
rect 388106 995508 388368 995511
rect 388054 995453 388106 995459
rect 382870 995437 382922 995443
rect 382870 995379 382922 995385
rect 382774 994993 382826 994999
rect 382774 994935 382826 994941
rect 390178 993635 390206 995522
rect 390850 994079 390878 995522
rect 391714 995508 392112 995527
rect 390836 994070 390892 994079
rect 390836 994005 390892 994014
rect 392674 993889 392702 995522
rect 393058 995508 393312 995536
rect 393730 995508 393984 995536
rect 393058 995443 393086 995508
rect 393046 995437 393098 995443
rect 393046 995379 393098 995385
rect 392662 993883 392714 993889
rect 392662 993825 392714 993831
rect 393730 993741 393758 995508
rect 395170 994999 395198 995522
rect 395158 994993 395210 994999
rect 395158 994935 395210 994941
rect 393718 993735 393770 993741
rect 393718 993677 393770 993683
rect 398818 993667 398846 995522
rect 429730 993667 429758 995929
rect 438740 995846 438796 995855
rect 438740 995781 438742 995790
rect 438794 995781 438796 995790
rect 444886 995807 444938 995813
rect 438742 995749 438794 995755
rect 444886 995749 444938 995755
rect 440660 995698 440716 995707
rect 440660 995633 440716 995642
rect 398806 993661 398858 993667
rect 390164 993626 390220 993635
rect 398806 993603 398858 993609
rect 429718 993661 429770 993667
rect 429718 993603 429770 993609
rect 390164 993561 390220 993570
rect 390178 992155 390206 993561
rect 390164 992146 390220 992155
rect 390164 992081 390220 992090
rect 397846 986557 397898 986563
rect 397846 986499 397898 986505
rect 377302 986483 377354 986489
rect 377302 986425 377354 986431
rect 365398 986409 365450 986415
rect 365398 986351 365450 986357
rect 374614 986409 374666 986415
rect 374614 986351 374666 986357
rect 365410 981462 365438 986351
rect 381622 985151 381674 985157
rect 381622 985093 381674 985099
rect 381634 981462 381662 985093
rect 397858 981462 397886 986499
rect 414070 986483 414122 986489
rect 414070 986425 414122 986431
rect 414082 981462 414110 986425
rect 440674 986415 440702 995633
rect 430294 986409 430346 986415
rect 430294 986351 430346 986357
rect 440662 986409 440714 986415
rect 440662 986351 440714 986357
rect 430306 981462 430334 986351
rect 444898 985157 444926 995749
rect 445090 986489 445118 995929
rect 460834 995443 460862 999301
rect 460930 996997 460958 1002187
rect 461026 999291 461054 1003741
rect 463714 1001067 463742 1003815
rect 463702 1001061 463754 1001067
rect 463702 1001003 463754 1001009
rect 463702 1000469 463754 1000475
rect 463702 1000411 463754 1000417
rect 461014 999285 461066 999291
rect 461014 999227 461066 999233
rect 460918 996991 460970 996997
rect 460918 996933 460970 996939
rect 460822 995437 460874 995443
rect 460822 995379 460874 995385
rect 463714 994999 463742 1000411
rect 466498 995411 466526 1005517
rect 466594 1002251 466622 1005739
rect 471862 1005501 471914 1005507
rect 471862 1005443 471914 1005449
rect 501140 1005466 501196 1005475
rect 470902 1005427 470954 1005433
rect 470902 1005369 470954 1005375
rect 466582 1002245 466634 1002251
rect 466582 1002187 466634 1002193
rect 470914 996035 470942 1005369
rect 471478 1005279 471530 1005285
rect 471478 1005221 471530 1005227
rect 470902 996029 470954 996035
rect 470902 995971 470954 995977
rect 471490 995559 471518 1005221
rect 471670 1005205 471722 1005211
rect 471670 1005147 471722 1005153
rect 471574 999285 471626 999291
rect 471574 999227 471626 999233
rect 471476 995550 471532 995559
rect 471476 995485 471532 995494
rect 466484 995402 466540 995411
rect 471586 995369 471614 999227
rect 466484 995337 466540 995346
rect 471574 995363 471626 995369
rect 471574 995305 471626 995311
rect 463702 994993 463754 994999
rect 463702 994935 463754 994941
rect 471682 994925 471710 1005147
rect 471766 1001061 471818 1001067
rect 471766 1001003 471818 1001009
rect 471778 995517 471806 1001003
rect 471874 995961 471902 1005443
rect 501140 1005401 501142 1005410
rect 501194 1005401 501196 1005410
rect 518326 1005427 518378 1005433
rect 501142 1005369 501194 1005375
rect 518326 1005369 518378 1005375
rect 504596 1005318 504652 1005327
rect 504596 1005253 504598 1005262
rect 504650 1005253 504652 1005262
rect 504598 1005221 504650 1005227
rect 518338 1005211 518366 1005369
rect 554518 1005353 554570 1005359
rect 554516 1005318 554518 1005327
rect 572854 1005353 572906 1005359
rect 554570 1005318 554572 1005327
rect 521398 1005279 521450 1005285
rect 554516 1005253 554572 1005262
rect 555764 1005318 555820 1005327
rect 572854 1005295 572906 1005301
rect 555764 1005253 555766 1005262
rect 521398 1005221 521450 1005227
rect 555818 1005253 555820 1005262
rect 555766 1005221 555818 1005227
rect 500758 1005205 500810 1005211
rect 500756 1005170 500758 1005179
rect 512566 1005205 512618 1005211
rect 500810 1005170 500812 1005179
rect 512566 1005147 512618 1005153
rect 518326 1005205 518378 1005211
rect 518326 1005147 518378 1005153
rect 500756 1005105 500812 1005114
rect 499990 1003799 500042 1003805
rect 499990 1003741 500042 1003747
rect 472054 1003725 472106 1003731
rect 472054 1003667 472106 1003673
rect 471958 1002245 472010 1002251
rect 471958 1002187 472010 1002193
rect 471970 996003 471998 1002187
rect 471956 995994 472012 996003
rect 471862 995955 471914 995961
rect 471956 995929 472012 995938
rect 471862 995897 471914 995903
rect 472066 995707 472094 1003667
rect 489526 1002319 489578 1002325
rect 489526 1002261 489578 1002267
rect 472642 1001141 472766 1001160
rect 472630 1001135 472766 1001141
rect 472682 1001132 472766 1001135
rect 472630 1001077 472682 1001083
rect 472630 1000987 472682 1000993
rect 472630 1000929 472682 1000935
rect 472534 1000913 472586 1000919
rect 472534 1000855 472586 1000861
rect 472342 1000839 472394 1000845
rect 472342 1000781 472394 1000787
rect 472150 1000395 472202 1000401
rect 472150 1000337 472202 1000343
rect 472052 995698 472108 995707
rect 472052 995633 472108 995642
rect 471766 995511 471818 995517
rect 471766 995453 471818 995459
rect 472162 995295 472190 1000337
rect 472246 996991 472298 996997
rect 472246 996933 472298 996939
rect 472258 995855 472286 996933
rect 472244 995846 472300 995855
rect 472244 995781 472300 995790
rect 472354 995665 472382 1000781
rect 472546 995739 472574 1000855
rect 472642 995813 472670 1000929
rect 472630 995807 472682 995813
rect 472630 995749 472682 995755
rect 472534 995733 472586 995739
rect 472534 995675 472586 995681
rect 472342 995659 472394 995665
rect 472342 995601 472394 995607
rect 472738 995591 472766 1001132
rect 488852 999546 488908 999555
rect 488852 999481 488908 999490
rect 480980 995846 481036 995855
rect 473314 995813 473664 995832
rect 473302 995807 473664 995813
rect 473354 995804 473664 995807
rect 485684 995846 485740 995855
rect 481036 995804 481104 995832
rect 480980 995781 481036 995790
rect 485740 995804 486000 995832
rect 485684 995781 485740 995790
rect 473302 995749 473354 995755
rect 474070 995733 474122 995739
rect 488866 995707 488894 999481
rect 477044 995698 477100 995707
rect 474122 995681 474336 995684
rect 474070 995675 474336 995681
rect 474082 995656 474336 995675
rect 479924 995698 479980 995707
rect 477100 995656 477360 995684
rect 477730 995665 477984 995684
rect 479856 995670 479924 995684
rect 477718 995659 477984 995665
rect 477044 995633 477100 995642
rect 477770 995656 477984 995659
rect 479446 995659 479498 995665
rect 477718 995601 477770 995607
rect 479446 995601 479498 995607
rect 479842 995656 479924 995670
rect 472726 995585 472778 995591
rect 472726 995527 472778 995533
rect 474646 995585 474698 995591
rect 474698 995533 474960 995536
rect 474646 995527 474960 995533
rect 474658 995508 474960 995527
rect 476482 995508 476784 995536
rect 476482 995411 476510 995508
rect 476468 995402 476524 995411
rect 476468 995337 476524 995346
rect 478642 995295 478670 995522
rect 472150 995289 472202 995295
rect 472150 995231 472202 995237
rect 478630 995289 478682 995295
rect 478630 995231 478682 995237
rect 471670 994919 471722 994925
rect 471670 994861 471722 994867
rect 469460 993626 469516 993635
rect 479170 993593 479198 995522
rect 479458 995369 479486 995601
rect 479446 995363 479498 995369
rect 479446 995305 479498 995311
rect 479842 994079 479870 995656
rect 479924 995633 479980 995642
rect 488852 995698 488908 995707
rect 488852 995633 488908 995642
rect 482036 995550 482092 995559
rect 481666 994925 481694 995522
rect 482092 995508 482352 995536
rect 482722 995508 482976 995536
rect 483874 995517 484176 995536
rect 483862 995511 484176 995517
rect 482036 995485 482092 995494
rect 482722 994999 482750 995508
rect 483914 995508 484176 995511
rect 485376 995508 485630 995536
rect 483862 995453 483914 995459
rect 482710 994993 482762 994999
rect 482710 994935 482762 994941
rect 481654 994919 481706 994925
rect 481654 994861 481706 994867
rect 485602 994079 485630 995508
rect 479828 994070 479884 994079
rect 479828 994005 479884 994014
rect 485588 994070 485644 994079
rect 485588 994005 485644 994014
rect 487810 993667 487838 995522
rect 487798 993661 487850 993667
rect 487798 993603 487850 993609
rect 489538 993593 489566 1002261
rect 497590 999581 497642 999587
rect 497588 999546 497590 999555
rect 497642 999546 497644 999555
rect 497588 999481 497644 999490
rect 500002 995855 500030 1003741
rect 503446 1002541 503498 1002547
rect 502772 1002506 502828 1002515
rect 502772 1002441 502774 1002450
rect 502826 1002441 502828 1002450
rect 503444 1002506 503446 1002515
rect 503498 1002506 503500 1002515
rect 503444 1002441 503500 1002450
rect 502774 1002409 502826 1002415
rect 505078 1002393 505130 1002399
rect 505076 1002358 505078 1002367
rect 505130 1002358 505132 1002367
rect 505076 1002293 505132 1002302
rect 511028 1001322 511084 1001331
rect 511028 1001257 511030 1001266
rect 511082 1001257 511084 1001266
rect 511030 1001225 511082 1001231
rect 509398 1001061 509450 1001067
rect 509396 1001026 509398 1001035
rect 509450 1001026 509452 1001035
rect 509396 1000961 509452 1000970
rect 507766 1000765 507818 1000771
rect 507764 1000730 507766 1000739
rect 507818 1000730 507820 1000739
rect 507764 1000665 507820 1000674
rect 506324 999546 506380 999555
rect 506324 999481 506326 999490
rect 506378 999481 506380 999490
rect 506326 999449 506378 999455
rect 502388 999398 502444 999407
rect 512578 999384 512606 1005147
rect 515542 1003799 515594 1003805
rect 515542 1003741 515594 1003747
rect 515446 1002541 515498 1002547
rect 515446 1002483 515498 1002489
rect 513526 1002467 513578 1002473
rect 513526 1002409 513578 1002415
rect 513538 1001659 513566 1002409
rect 513526 1001653 513578 1001659
rect 513526 1001595 513578 1001601
rect 515458 1001585 515486 1002483
rect 515446 1001579 515498 1001585
rect 515446 1001521 515498 1001527
rect 512578 999356 512798 999384
rect 502388 999333 502390 999342
rect 502442 999333 502444 999342
rect 502390 999301 502442 999307
rect 510262 996621 510314 996627
rect 508628 996586 508684 996595
rect 508628 996521 508630 996530
rect 508682 996521 508684 996530
rect 510260 996586 510262 996595
rect 510314 996586 510316 996595
rect 510260 996521 510316 996530
rect 508630 996489 508682 996495
rect 511126 996251 511178 996257
rect 511126 996193 511178 996199
rect 511138 996003 511166 996193
rect 511124 995994 511180 996003
rect 511124 995929 511126 995938
rect 511178 995929 511180 995938
rect 511126 995897 511178 995903
rect 511894 995881 511946 995887
rect 499988 995846 500044 995855
rect 499988 995781 500044 995790
rect 511892 995846 511894 995855
rect 511946 995846 511948 995855
rect 511892 995781 511948 995790
rect 506612 995254 506668 995263
rect 506612 995189 506668 995198
rect 506626 993741 506654 995189
rect 512770 993815 512798 999356
rect 515554 999291 515582 1003741
rect 519190 1002319 519242 1002325
rect 519190 1002261 519242 1002267
rect 518326 1001653 518378 1001659
rect 518326 1001595 518378 1001601
rect 516886 1001579 516938 1001585
rect 516886 1001521 516938 1001527
rect 516692 1001322 516748 1001331
rect 516692 1001257 516694 1001266
rect 516746 1001257 516748 1001266
rect 516694 1001225 516746 1001231
rect 516694 1001061 516746 1001067
rect 516692 1001026 516694 1001035
rect 516746 1001026 516748 1001035
rect 516692 1000961 516748 1000970
rect 516694 1000765 516746 1000771
rect 516692 1000730 516694 1000739
rect 516746 1000730 516748 1000739
rect 516692 1000665 516748 1000674
rect 516692 999842 516748 999851
rect 516692 999777 516748 999786
rect 516706 999587 516734 999777
rect 516694 999581 516746 999587
rect 516694 999523 516746 999529
rect 516788 999546 516844 999555
rect 516788 999481 516790 999490
rect 516842 999481 516844 999490
rect 516790 999449 516842 999455
rect 516692 999398 516748 999407
rect 516898 999365 516926 1001521
rect 516692 999333 516694 999342
rect 516746 999333 516748 999342
rect 516886 999359 516938 999365
rect 516694 999301 516746 999307
rect 516886 999301 516938 999307
rect 515542 999285 515594 999291
rect 515542 999227 515594 999233
rect 518338 999236 518366 1001595
rect 518338 999208 518558 999236
rect 513430 996177 513482 996183
rect 513428 996142 513430 996151
rect 513482 996142 513484 996151
rect 513428 996077 513484 996086
rect 513430 996029 513482 996035
rect 513428 995994 513430 996003
rect 513482 995994 513484 996003
rect 513428 995929 513484 995938
rect 518420 995698 518476 995707
rect 518420 995633 518476 995642
rect 512758 993809 512810 993815
rect 512758 993751 512810 993757
rect 506614 993735 506666 993741
rect 506614 993677 506666 993683
rect 469460 993561 469462 993570
rect 469514 993561 469516 993570
rect 479158 993587 479210 993593
rect 469462 993529 469514 993535
rect 479158 993529 479210 993535
rect 489526 993587 489578 993593
rect 489526 993529 489578 993535
rect 518434 987821 518462 995633
rect 518530 995369 518558 999208
rect 518612 995550 518668 995559
rect 518612 995485 518668 995494
rect 518518 995363 518570 995369
rect 518518 995305 518570 995311
rect 518422 987815 518474 987821
rect 518422 987757 518474 987763
rect 445078 986483 445130 986489
rect 445078 986425 445130 986431
rect 478966 986483 479018 986489
rect 478966 986425 479018 986431
rect 444886 985151 444938 985157
rect 444886 985093 444938 985099
rect 462742 985151 462794 985157
rect 462742 985093 462794 985099
rect 446518 985077 446570 985083
rect 446518 985019 446570 985025
rect 446530 981462 446558 985019
rect 462754 981462 462782 985093
rect 478978 981462 479006 986425
rect 518626 986415 518654 995485
rect 519202 994925 519230 1002261
rect 521410 999703 521438 1005221
rect 521590 1005205 521642 1005211
rect 553750 1005205 553802 1005211
rect 521590 1005147 521642 1005153
rect 553748 1005170 553750 1005179
rect 553802 1005170 553804 1005179
rect 521494 1002393 521546 1002399
rect 521494 1002335 521546 1002341
rect 521396 999694 521452 999703
rect 521396 999629 521452 999638
rect 521506 999555 521534 1002335
rect 521602 999999 521630 1005147
rect 553748 1005105 553804 1005114
rect 552598 1003873 552650 1003879
rect 552596 1003838 552598 1003847
rect 572662 1003873 572714 1003879
rect 552650 1003838 552652 1003847
rect 552596 1003773 552652 1003782
rect 556532 1003838 556588 1003847
rect 572662 1003815 572714 1003821
rect 556532 1003773 556534 1003782
rect 556586 1003773 556588 1003782
rect 556534 1003741 556586 1003747
rect 551734 1003725 551786 1003731
rect 551732 1003690 551734 1003699
rect 551786 1003690 551788 1003699
rect 551732 1003625 551788 1003634
rect 559222 1002689 559274 1002695
rect 559220 1002654 559222 1002663
rect 566326 1002689 566378 1002695
rect 559274 1002654 559276 1002663
rect 559220 1002589 559276 1002598
rect 559988 1002654 560044 1002663
rect 566326 1002631 566378 1002637
rect 559988 1002589 559990 1002598
rect 560042 1002589 560044 1002598
rect 566134 1002615 566186 1002621
rect 559990 1002557 560042 1002563
rect 566134 1002557 566186 1002563
rect 562198 1002541 562250 1002547
rect 562196 1002506 562198 1002515
rect 562250 1002506 562252 1002515
rect 562196 1002441 562252 1002450
rect 564596 1002506 564652 1002515
rect 564596 1002441 564598 1002450
rect 564650 1002441 564652 1002450
rect 564598 1002409 564650 1002415
rect 560470 1002393 560522 1002399
rect 544244 1002358 544300 1002367
rect 544244 1002293 544300 1002302
rect 560468 1002358 560470 1002367
rect 564790 1002393 564842 1002399
rect 560522 1002358 560524 1002367
rect 560468 1002293 560524 1002302
rect 561524 1002358 561580 1002367
rect 564790 1002335 564842 1002341
rect 561524 1002293 561526 1002302
rect 523604 1001322 523660 1001331
rect 523604 1001257 523660 1001266
rect 523508 1000730 523564 1000739
rect 523508 1000665 523564 1000674
rect 521588 999990 521644 999999
rect 521588 999925 521644 999934
rect 523316 999842 523372 999851
rect 523316 999777 523372 999786
rect 521492 999546 521548 999555
rect 521492 999481 521548 999490
rect 521108 999398 521164 999407
rect 520918 999359 520970 999365
rect 521108 999333 521164 999342
rect 520918 999301 520970 999307
rect 520930 995559 520958 999301
rect 521014 996621 521066 996627
rect 521014 996563 521066 996569
rect 520916 995550 520972 995559
rect 520916 995485 520972 995494
rect 521026 995295 521054 996563
rect 521122 995961 521150 999333
rect 521206 996547 521258 996553
rect 521206 996489 521258 996495
rect 521110 995955 521162 995961
rect 521110 995897 521162 995903
rect 521218 995855 521246 996489
rect 521300 995994 521356 996003
rect 521300 995929 521356 995938
rect 521204 995846 521260 995855
rect 521204 995781 521260 995790
rect 521014 995289 521066 995295
rect 521014 995231 521066 995237
rect 519190 994919 519242 994925
rect 519190 994861 519242 994867
rect 521314 986489 521342 995929
rect 523330 995411 523358 999777
rect 523414 999285 523466 999291
rect 523414 999227 523466 999233
rect 523316 995402 523372 995411
rect 523316 995337 523372 995346
rect 523426 994999 523454 999227
rect 523522 996003 523550 1000665
rect 523508 995994 523564 996003
rect 523508 995929 523564 995938
rect 523618 995707 523646 1001257
rect 523700 1001026 523756 1001035
rect 523700 1000961 523756 1000970
rect 523604 995698 523660 995707
rect 523604 995633 523660 995642
rect 523714 995591 523742 1000961
rect 523892 999990 523948 999999
rect 523892 999925 523948 999934
rect 523796 999398 523852 999407
rect 523796 999333 523852 999342
rect 523810 995665 523838 999333
rect 523906 995887 523934 999925
rect 523988 999694 524044 999703
rect 523988 999629 524044 999638
rect 523894 995881 523946 995887
rect 523894 995823 523946 995829
rect 524002 995739 524030 999629
rect 524084 999546 524140 999555
rect 524084 999481 524140 999490
rect 524098 995813 524126 999481
rect 540310 999433 540362 999439
rect 540310 999375 540362 999381
rect 527924 995846 527980 995855
rect 524086 995807 524138 995813
rect 532244 995846 532300 995855
rect 527980 995804 528192 995832
rect 528418 995813 528768 995832
rect 529858 995813 530064 995832
rect 528406 995807 528768 995813
rect 527924 995781 527980 995790
rect 524086 995749 524138 995755
rect 528458 995804 528768 995807
rect 529846 995807 530064 995813
rect 528406 995749 528458 995755
rect 529898 995804 530064 995807
rect 532300 995804 532512 995832
rect 536784 995813 537182 995832
rect 540322 995813 540350 999375
rect 536784 995807 537194 995813
rect 536784 995804 537142 995807
rect 532244 995781 532300 995790
rect 529846 995749 529898 995755
rect 537142 995749 537194 995755
rect 540310 995807 540362 995813
rect 540310 995749 540362 995755
rect 523990 995733 524042 995739
rect 528982 995733 529034 995739
rect 526100 995698 526156 995707
rect 523990 995675 524042 995681
rect 525442 995665 525744 995684
rect 523798 995659 523850 995665
rect 523798 995601 523850 995607
rect 525430 995659 525744 995665
rect 525482 995656 525744 995659
rect 526156 995656 526368 995684
rect 532822 995733 532874 995739
rect 529034 995681 529392 995684
rect 528982 995675 529392 995681
rect 532874 995681 533088 995684
rect 532822 995675 533088 995681
rect 528994 995656 529392 995675
rect 532834 995656 533088 995675
rect 526100 995633 526156 995642
rect 525430 995601 525482 995607
rect 523702 995585 523754 995591
rect 523702 995527 523754 995533
rect 524758 995585 524810 995591
rect 535316 995550 535372 995559
rect 524810 995533 525072 995536
rect 524758 995527 525072 995533
rect 524770 995508 525072 995527
rect 530338 995508 530592 995536
rect 530914 995522 531216 995536
rect 530914 995508 531230 995522
rect 523414 994993 523466 994999
rect 523414 994935 523466 994941
rect 530338 994925 530366 995508
rect 530914 995411 530942 995508
rect 530900 995402 530956 995411
rect 530900 995337 530956 995346
rect 530326 994919 530378 994925
rect 530326 994861 530378 994867
rect 530338 993667 530366 994861
rect 531202 994227 531230 995508
rect 533698 995369 533726 995522
rect 533686 995363 533738 995369
rect 533686 995305 533738 995311
rect 531188 994218 531244 994227
rect 531188 994153 531244 994162
rect 534370 993815 534398 995522
rect 535372 995508 535584 995536
rect 535316 995485 535372 995494
rect 537394 995295 537422 995522
rect 538978 995508 539232 995536
rect 537382 995289 537434 995295
rect 537382 995231 537434 995237
rect 537526 995289 537578 995295
rect 537526 995231 537578 995237
rect 537538 994999 537566 995231
rect 537526 994993 537578 994999
rect 537526 994935 537578 994941
rect 534358 993809 534410 993815
rect 534358 993751 534410 993757
rect 538978 993741 539006 995508
rect 538966 993735 539018 993741
rect 538966 993677 539018 993683
rect 530326 993661 530378 993667
rect 530326 993603 530378 993609
rect 527638 987815 527690 987821
rect 527638 987757 527690 987763
rect 521302 986483 521354 986489
rect 521302 986425 521354 986431
rect 495190 986409 495242 986415
rect 495190 986351 495242 986357
rect 518614 986409 518666 986415
rect 518614 986351 518666 986357
rect 495202 981462 495230 986351
rect 511414 985003 511466 985009
rect 511414 984945 511466 984951
rect 511426 981462 511454 984945
rect 527650 981462 527678 987757
rect 543766 986483 543818 986489
rect 543766 986425 543818 986431
rect 543778 981462 543806 986425
rect 544258 983529 544286 1002293
rect 561578 1002293 561580 1002302
rect 564694 1002319 564746 1002325
rect 561526 1002261 561578 1002267
rect 564694 1002261 564746 1002267
rect 564706 999513 564734 1002261
rect 564694 999507 564746 999513
rect 564694 999449 564746 999455
rect 561526 999433 561578 999439
rect 561526 999375 561578 999381
rect 555284 998066 555340 998075
rect 555284 998001 555286 998010
rect 555338 998001 555340 998010
rect 555286 997969 555338 997975
rect 561538 997959 561566 999375
rect 561526 997953 561578 997959
rect 557300 997918 557356 997927
rect 561526 997895 561578 997901
rect 557300 997853 557302 997862
rect 557354 997853 557356 997862
rect 557302 997821 557354 997827
rect 564802 997589 564830 1002335
rect 566146 1001511 566174 1002557
rect 566134 1001505 566186 1001511
rect 566134 1001447 566186 1001453
rect 566338 999439 566366 1002631
rect 567574 1002541 567626 1002547
rect 567574 1002483 567626 1002489
rect 566326 999433 566378 999439
rect 566326 999375 566378 999381
rect 564790 997583 564842 997589
rect 564790 997525 564842 997531
rect 562774 996177 562826 996183
rect 562774 996119 562826 996125
rect 562786 995707 562814 996119
rect 563542 996103 563594 996109
rect 563542 996045 563594 996051
rect 563554 995707 563582 996045
rect 564790 996029 564842 996035
rect 564788 995994 564790 996003
rect 564842 995994 564844 996003
rect 564788 995929 564844 995938
rect 562772 995698 562828 995707
rect 562772 995633 562828 995642
rect 563540 995698 563596 995707
rect 563540 995633 563542 995642
rect 562786 995591 562814 995633
rect 563594 995633 563596 995642
rect 567382 995659 567434 995665
rect 563542 995601 563594 995607
rect 567382 995601 567434 995607
rect 562774 995585 562826 995591
rect 562774 995527 562826 995533
rect 557972 995402 558028 995411
rect 557972 995337 558028 995346
rect 557986 993741 558014 995337
rect 557974 993735 558026 993741
rect 557974 993677 558026 993683
rect 560086 986409 560138 986415
rect 560086 986351 560138 986357
rect 544246 983523 544298 983529
rect 544246 983465 544298 983471
rect 560098 981462 560126 986351
rect 567394 983603 567422 995601
rect 567478 995585 567530 995591
rect 567478 995527 567530 995533
rect 567490 983677 567518 995527
rect 567586 994523 567614 1002483
rect 568726 1002467 568778 1002473
rect 568726 1002409 568778 1002415
rect 567766 1001505 567818 1001511
rect 567766 1001447 567818 1001453
rect 567778 997737 567806 1001447
rect 567766 997731 567818 997737
rect 567766 997673 567818 997679
rect 567572 994514 567628 994523
rect 567572 994449 567628 994458
rect 568738 983751 568766 1002409
rect 570454 999359 570506 999365
rect 570454 999301 570506 999307
rect 570646 999359 570698 999365
rect 570646 999301 570698 999307
rect 570356 995698 570412 995707
rect 570356 995633 570412 995642
rect 570262 995067 570314 995073
rect 570262 995009 570314 995015
rect 570274 987821 570302 995009
rect 570262 987815 570314 987821
rect 570262 987757 570314 987763
rect 570370 986563 570398 995633
rect 570466 994375 570494 999301
rect 570548 995550 570604 995559
rect 570548 995485 570604 995494
rect 570452 994366 570508 994375
rect 570452 994301 570508 994310
rect 570358 986557 570410 986563
rect 570358 986499 570410 986505
rect 570562 986415 570590 995485
rect 570658 993963 570686 999301
rect 570742 998027 570794 998033
rect 570742 997969 570794 997975
rect 570646 993957 570698 993963
rect 570646 993899 570698 993905
rect 570754 993815 570782 997969
rect 572674 993889 572702 1003815
rect 572758 1003725 572810 1003731
rect 572758 1003667 572810 1003673
rect 572770 994037 572798 1003667
rect 572866 1001363 572894 1005295
rect 573046 1005279 573098 1005285
rect 573046 1005221 573098 1005227
rect 572950 1005205 573002 1005211
rect 572950 1005147 573002 1005153
rect 572962 1001881 572990 1005147
rect 573058 1002251 573086 1005221
rect 574006 1003799 574058 1003805
rect 574006 1003741 574058 1003747
rect 573046 1002245 573098 1002251
rect 573046 1002187 573098 1002193
rect 573910 1002245 573962 1002251
rect 573910 1002187 573962 1002193
rect 572950 1001875 573002 1001881
rect 572950 1001817 573002 1001823
rect 573238 1001875 573290 1001881
rect 573238 1001817 573290 1001823
rect 572854 1001357 572906 1001363
rect 572854 1001299 572906 1001305
rect 573140 995846 573196 995855
rect 573140 995781 573196 995790
rect 572758 994031 572810 994037
rect 572758 993973 572810 993979
rect 572662 993883 572714 993889
rect 572662 993825 572714 993831
rect 570742 993809 570794 993815
rect 570742 993751 570794 993757
rect 573154 986489 573182 995781
rect 573250 994671 573278 1001817
rect 573922 997663 573950 1002187
rect 574018 997811 574046 1003741
rect 574486 1001357 574538 1001363
rect 574486 1001299 574538 1001305
rect 574006 997805 574058 997811
rect 574006 997747 574058 997753
rect 573910 997657 573962 997663
rect 573910 997599 573962 997605
rect 573236 994662 573292 994671
rect 573236 994597 573292 994606
rect 574498 994185 574526 1001299
rect 610582 999729 610634 999735
rect 610582 999671 610634 999677
rect 625750 999729 625802 999735
rect 625750 999671 625802 999677
rect 604726 999581 604778 999587
rect 604726 999523 604778 999529
rect 593302 999507 593354 999513
rect 593302 999449 593354 999455
rect 590518 999433 590570 999439
rect 590518 999375 590570 999381
rect 590530 997811 590558 999375
rect 593314 997885 593342 999449
rect 593302 997879 593354 997885
rect 593302 997821 593354 997827
rect 590518 997805 590570 997811
rect 590518 997747 590570 997753
rect 604738 997737 604766 999523
rect 604726 997731 604778 997737
rect 604726 997673 604778 997679
rect 610594 997589 610622 999671
rect 613462 999655 613514 999661
rect 613462 999597 613514 999603
rect 625462 999655 625514 999661
rect 625462 999597 625514 999603
rect 613474 997663 613502 999597
rect 616342 997953 616394 997959
rect 616342 997895 616394 997901
rect 613462 997657 613514 997663
rect 613462 997599 613514 997605
rect 610582 997583 610634 997589
rect 610582 997525 610634 997531
rect 616354 995073 616382 997895
rect 625474 995961 625502 999597
rect 625558 999581 625610 999587
rect 625558 999523 625610 999529
rect 625462 995955 625514 995961
rect 625462 995897 625514 995903
rect 625570 995665 625598 999523
rect 625654 999433 625706 999439
rect 625654 999375 625706 999381
rect 625666 995887 625694 999375
rect 625654 995881 625706 995887
rect 625654 995823 625706 995829
rect 625762 995739 625790 999671
rect 625846 999507 625898 999513
rect 625846 999449 625898 999455
rect 625858 995813 625886 999449
rect 627106 995813 627504 995832
rect 630178 995813 630576 995832
rect 630946 995813 631200 995832
rect 625846 995807 625898 995813
rect 625846 995749 625898 995755
rect 627094 995807 627504 995813
rect 627146 995804 627504 995807
rect 630166 995807 630576 995813
rect 627094 995749 627146 995755
rect 630218 995804 630576 995807
rect 630934 995807 631200 995813
rect 630166 995749 630218 995755
rect 630986 995804 631200 995807
rect 630934 995749 630986 995755
rect 625750 995733 625802 995739
rect 625750 995675 625802 995681
rect 626518 995733 626570 995739
rect 626570 995681 626880 995684
rect 626518 995675 626880 995681
rect 625558 995659 625610 995665
rect 626530 995656 626880 995675
rect 629602 995665 630000 995684
rect 629590 995659 630000 995665
rect 625558 995601 625610 995607
rect 629642 995656 630000 995659
rect 629590 995601 629642 995607
rect 616342 995067 616394 995073
rect 616342 995009 616394 995015
rect 628162 994523 628190 995522
rect 629206 995511 629258 995517
rect 629206 995453 629258 995459
rect 628148 994514 628204 994523
rect 628148 994449 628204 994458
rect 574486 994179 574538 994185
rect 574486 994121 574538 994127
rect 604724 994070 604780 994079
rect 604724 994005 604780 994014
rect 604738 988265 604766 994005
rect 622004 993774 622060 993783
rect 622004 993709 622060 993718
rect 604726 988259 604778 988265
rect 604726 988201 604778 988207
rect 618550 988259 618602 988265
rect 618550 988201 618602 988207
rect 576310 987815 576362 987821
rect 576310 987757 576362 987763
rect 573142 986483 573194 986489
rect 573142 986425 573194 986431
rect 570550 986409 570602 986415
rect 570550 986351 570602 986357
rect 568726 983745 568778 983751
rect 568726 983687 568778 983693
rect 567478 983671 567530 983677
rect 567478 983613 567530 983619
rect 567382 983597 567434 983603
rect 567382 983539 567434 983545
rect 576322 981462 576350 987757
rect 592438 986557 592490 986563
rect 592438 986499 592490 986505
rect 592450 981462 592478 986499
rect 608758 986483 608810 986489
rect 608758 986425 608810 986431
rect 608770 981462 608798 986425
rect 618562 983825 618590 988201
rect 622018 986489 622046 993709
rect 629218 990929 629246 995453
rect 630742 995437 630794 995443
rect 630742 995379 630794 995385
rect 629206 990923 629258 990929
rect 629206 990865 629258 990871
rect 630754 986563 630782 995379
rect 631810 994671 631838 995522
rect 631796 994662 631852 994671
rect 631796 994597 631852 994606
rect 631028 994218 631084 994227
rect 631028 994153 631084 994162
rect 630838 993661 630890 993667
rect 630838 993603 630890 993609
rect 630742 986557 630794 986563
rect 630742 986499 630794 986505
rect 622006 986483 622058 986489
rect 622006 986425 622058 986431
rect 624982 986409 625034 986415
rect 624982 986351 625034 986357
rect 630742 986409 630794 986415
rect 630742 986351 630794 986357
rect 618550 983819 618602 983825
rect 618550 983761 618602 983767
rect 624994 981462 625022 986351
rect 273622 980785 273674 980791
rect 218954 980750 218956 980759
rect 106498 980708 106622 980727
rect 146818 980708 146942 980727
rect 218900 980685 218956 980694
rect 238964 980750 239020 980759
rect 273622 980727 273674 980733
rect 630754 980736 630782 986351
rect 630850 980865 630878 993603
rect 631042 986415 631070 994153
rect 632386 993667 632414 995522
rect 632770 995508 633024 995536
rect 632770 994227 632798 995508
rect 634306 994375 634334 995522
rect 634292 994366 634348 994375
rect 634292 994301 634348 994310
rect 632756 994218 632812 994227
rect 632756 994153 632812 994162
rect 634882 993889 634910 995522
rect 635266 995508 635520 995536
rect 635266 994185 635294 995508
rect 635254 994179 635306 994185
rect 635254 994121 635306 994127
rect 636130 994037 636158 995522
rect 636118 994031 636170 994037
rect 636118 993973 636170 993979
rect 634870 993883 634922 993889
rect 634870 993825 634922 993831
rect 637378 993815 637406 995522
rect 638544 995508 638942 995536
rect 637366 993809 637418 993815
rect 637366 993751 637418 993757
rect 638914 993667 638942 995508
rect 639202 993963 639230 995522
rect 640342 995067 640394 995073
rect 640342 995009 640394 995015
rect 639190 993957 639242 993963
rect 639190 993899 639242 993905
rect 632374 993661 632426 993667
rect 632374 993603 632426 993609
rect 638902 993661 638954 993667
rect 638902 993603 638954 993609
rect 640354 989523 640382 995009
rect 641026 993741 641054 995522
rect 645142 995289 645194 995295
rect 645142 995231 645194 995237
rect 641014 993735 641066 993741
rect 641014 993677 641066 993683
rect 643606 993661 643658 993667
rect 643606 993603 643658 993609
rect 642166 990923 642218 990929
rect 642166 990865 642218 990871
rect 642178 990652 642206 990865
rect 642178 990624 642302 990652
rect 640342 989517 640394 989523
rect 640342 989459 640394 989465
rect 639382 986557 639434 986563
rect 639382 986499 639434 986505
rect 631030 986409 631082 986415
rect 631030 986351 631082 986357
rect 639394 981383 639422 986499
rect 641110 986483 641162 986489
rect 641110 986425 641162 986431
rect 641122 981462 641150 986425
rect 642274 985009 642302 990624
rect 642262 985003 642314 985009
rect 642262 984945 642314 984951
rect 643618 981827 643646 993603
rect 645154 987821 645182 995231
rect 649942 995215 649994 995221
rect 649942 995157 649994 995163
rect 645238 995141 645290 995147
rect 645238 995083 645290 995089
rect 645250 988561 645278 995083
rect 649556 993922 649612 993931
rect 649556 993857 649612 993866
rect 645238 988555 645290 988561
rect 645238 988497 645290 988503
rect 645142 987815 645194 987821
rect 645142 987757 645194 987763
rect 649366 987815 649418 987821
rect 649366 987757 649418 987763
rect 643606 981821 643658 981827
rect 643606 981763 643658 981769
rect 639382 981377 639434 981383
rect 639382 981319 639434 981325
rect 630838 980859 630890 980865
rect 630838 980801 630890 980807
rect 630934 980785 630986 980791
rect 630754 980733 630934 980736
rect 630754 980727 630986 980733
rect 630754 980708 630974 980727
rect 238964 980685 239020 980694
rect 435394 276385 435696 276404
rect 303382 276379 303434 276385
rect 303382 276321 303434 276327
rect 435382 276379 435696 276385
rect 435434 276376 435696 276379
rect 435382 276321 435434 276327
rect 117238 276305 117290 276311
rect 116976 276253 117238 276256
rect 116976 276247 117290 276253
rect 116976 276228 117278 276247
rect 120528 276237 120830 276256
rect 120528 276231 120842 276237
rect 120528 276228 120790 276231
rect 120790 276173 120842 276179
rect 73270 276157 73322 276163
rect 73008 276105 73270 276108
rect 73008 276099 73322 276105
rect 73008 276080 73310 276099
rect 113520 276089 113822 276108
rect 113520 276083 113834 276089
rect 113520 276080 113782 276083
rect 113782 276025 113834 276031
rect 67056 275784 67358 275812
rect 82608 275784 82910 275812
rect 98064 275784 98366 275812
rect 128976 275784 129278 275812
rect 144432 275784 144734 275812
rect 155088 275784 155486 275812
rect 159888 275784 160190 275812
rect 175344 275784 175550 275812
rect 190800 275784 191102 275812
rect 206256 275784 206558 275812
rect 65904 275636 66302 275664
rect 66274 264841 66302 275636
rect 66838 272309 66890 272315
rect 66838 272251 66890 272257
rect 66850 267875 66878 272251
rect 66838 267869 66890 267875
rect 66838 267811 66890 267817
rect 66262 264835 66314 264841
rect 66262 264777 66314 264783
rect 67330 264545 67358 275784
rect 68194 270021 68222 275650
rect 68182 270015 68234 270021
rect 68182 269957 68234 269963
rect 69346 269355 69374 275650
rect 69334 269349 69386 269355
rect 69334 269291 69386 269297
rect 67318 264539 67370 264545
rect 67318 264481 67370 264487
rect 70594 262811 70622 275650
rect 71746 269281 71774 275650
rect 72022 272531 72074 272537
rect 72022 272473 72074 272479
rect 71734 269275 71786 269281
rect 71734 269217 71786 269223
rect 70580 262802 70636 262811
rect 70580 262737 70636 262746
rect 72034 259587 72062 272473
rect 74146 269725 74174 275650
rect 75394 270095 75422 275650
rect 75382 270089 75434 270095
rect 75382 270031 75434 270037
rect 74134 269719 74186 269725
rect 74134 269661 74186 269667
rect 72118 267795 72170 267801
rect 72118 267737 72170 267743
rect 72022 259581 72074 259587
rect 72022 259523 72074 259529
rect 72130 253445 72158 267737
rect 76546 263583 76574 275650
rect 77794 269323 77822 275650
rect 78946 269429 78974 275650
rect 80194 270169 80222 275650
rect 80182 270163 80234 270169
rect 80182 270105 80234 270111
rect 81346 269503 81374 275650
rect 81334 269497 81386 269503
rect 81334 269439 81386 269445
rect 78934 269423 78986 269429
rect 78934 269365 78986 269371
rect 77780 269314 77836 269323
rect 77780 269249 77836 269258
rect 82882 263847 82910 275784
rect 83650 264143 83678 275650
rect 84802 270243 84830 275650
rect 84790 270237 84842 270243
rect 84790 270179 84842 270185
rect 83636 264134 83692 264143
rect 83636 264069 83692 264078
rect 86050 263995 86078 275650
rect 87202 269577 87230 275650
rect 87190 269571 87242 269577
rect 87190 269513 87242 269519
rect 88450 269471 88478 275650
rect 89602 270317 89630 275650
rect 89590 270311 89642 270317
rect 89590 270253 89642 270259
rect 90850 269651 90878 275650
rect 90838 269645 90890 269651
rect 90838 269587 90890 269593
rect 88436 269462 88492 269471
rect 88436 269397 88492 269406
rect 87766 264983 87818 264989
rect 87766 264925 87818 264931
rect 87778 264545 87806 264925
rect 87766 264539 87818 264545
rect 87766 264481 87818 264487
rect 86036 263986 86092 263995
rect 86036 263921 86092 263930
rect 82868 263838 82924 263847
rect 82868 263773 82924 263782
rect 92002 263657 92030 275650
rect 93250 264291 93278 275650
rect 94402 270391 94430 275650
rect 94390 270385 94442 270391
rect 94390 270327 94442 270333
rect 95650 269767 95678 275650
rect 95636 269758 95692 269767
rect 95636 269693 95692 269702
rect 96802 269619 96830 275650
rect 98338 270465 98366 275784
rect 98326 270459 98378 270465
rect 98326 270401 98378 270407
rect 96788 269610 96844 269619
rect 96788 269545 96844 269554
rect 99202 264587 99230 275650
rect 99188 264578 99244 264587
rect 99188 264513 99244 264522
rect 100258 264439 100286 275650
rect 101506 270539 101534 275650
rect 101494 270533 101546 270539
rect 101494 270475 101546 270481
rect 102658 270063 102686 275650
rect 102644 270054 102700 270063
rect 102644 269989 102700 269998
rect 103906 269915 103934 275650
rect 105058 270613 105086 275650
rect 105046 270607 105098 270613
rect 105046 270549 105098 270555
rect 103892 269906 103948 269915
rect 103892 269841 103948 269850
rect 106306 264735 106334 275650
rect 106582 264983 106634 264989
rect 106582 264925 106634 264931
rect 106594 264767 106622 264925
rect 106582 264761 106634 264767
rect 106292 264726 106348 264735
rect 106582 264703 106634 264709
rect 106292 264661 106348 264670
rect 100244 264430 100300 264439
rect 100244 264365 100300 264374
rect 93236 264282 93292 264291
rect 93236 264217 93292 264226
rect 107458 263731 107486 275650
rect 108706 269207 108734 275650
rect 109858 270211 109886 275650
rect 111106 270359 111134 275650
rect 111092 270350 111148 270359
rect 111092 270285 111148 270294
rect 109844 270202 109900 270211
rect 109844 270137 109900 270146
rect 108694 269201 108746 269207
rect 108694 269143 108746 269149
rect 112258 269133 112286 275650
rect 114658 269799 114686 275650
rect 114646 269793 114698 269799
rect 114646 269735 114698 269741
rect 112246 269127 112298 269133
rect 112246 269069 112298 269075
rect 115810 269059 115838 275650
rect 115798 269053 115850 269059
rect 115798 268995 115850 269001
rect 118114 264883 118142 275650
rect 119362 268985 119390 275650
rect 121762 270507 121790 275650
rect 121748 270498 121804 270507
rect 121748 270433 121804 270442
rect 119350 268979 119402 268985
rect 119350 268921 119402 268927
rect 122914 268763 122942 275650
rect 124162 270687 124190 275650
rect 124150 270681 124202 270687
rect 124150 270623 124202 270629
rect 122902 268757 122954 268763
rect 122902 268699 122954 268705
rect 118100 264874 118156 264883
rect 118100 264809 118156 264818
rect 107446 263725 107498 263731
rect 107446 263667 107498 263673
rect 91990 263651 92042 263657
rect 91990 263593 92042 263599
rect 76534 263577 76586 263583
rect 76534 263519 76586 263525
rect 125314 263403 125342 275650
rect 126562 268467 126590 275650
rect 127714 269873 127742 275650
rect 129250 270655 129278 275784
rect 129236 270646 129292 270655
rect 129236 270581 129292 270590
rect 127702 269867 127754 269873
rect 127702 269809 127754 269815
rect 126550 268461 126602 268467
rect 126550 268403 126602 268409
rect 130114 268393 130142 275650
rect 131266 268689 131294 275650
rect 131254 268683 131306 268689
rect 131254 268625 131306 268631
rect 130102 268387 130154 268393
rect 130102 268329 130154 268335
rect 126742 264983 126794 264989
rect 126742 264925 126794 264931
rect 126754 264767 126782 264925
rect 126742 264761 126794 264767
rect 126742 264703 126794 264709
rect 132514 263805 132542 275650
rect 133570 268837 133598 275650
rect 134832 275636 135326 275664
rect 135298 269947 135326 275636
rect 135286 269941 135338 269947
rect 135286 269883 135338 269889
rect 135970 269175 135998 275650
rect 135956 269166 136012 269175
rect 135956 269101 136012 269110
rect 135382 268905 135434 268911
rect 135382 268847 135434 268853
rect 133558 268831 133610 268837
rect 133558 268773 133610 268779
rect 135394 268689 135422 268847
rect 135382 268683 135434 268689
rect 135382 268625 135434 268631
rect 137218 267875 137246 275650
rect 137206 267869 137258 267875
rect 137206 267811 137258 267817
rect 138370 266395 138398 275650
rect 139234 275636 139632 275664
rect 140784 275636 141086 275664
rect 139126 267795 139178 267801
rect 139126 267737 139178 267743
rect 138358 266389 138410 266395
rect 138358 266331 138410 266337
rect 132502 263799 132554 263805
rect 132502 263741 132554 263747
rect 125300 263394 125356 263403
rect 125300 263329 125356 263338
rect 77686 259581 77738 259587
rect 77686 259523 77738 259529
rect 77698 256128 77726 259523
rect 77698 256100 77918 256128
rect 72118 253439 72170 253445
rect 72118 253381 72170 253387
rect 77014 253439 77066 253445
rect 77014 253381 77066 253387
rect 65204 246374 65260 246383
rect 65204 246309 65260 246318
rect 65012 246226 65068 246235
rect 65012 246161 65068 246170
rect 77026 243973 77054 253381
rect 77890 244047 77918 256100
rect 80662 245373 80714 245379
rect 80660 245338 80662 245347
rect 100726 245373 100778 245379
rect 80714 245338 80716 245347
rect 100726 245315 100778 245321
rect 80660 245273 80716 245282
rect 100738 245199 100766 245315
rect 100724 245190 100780 245199
rect 100724 245125 100780 245134
rect 126548 245190 126604 245199
rect 126740 245190 126796 245199
rect 126604 245148 126740 245176
rect 126548 245125 126604 245134
rect 126740 245125 126796 245134
rect 77878 244041 77930 244047
rect 77878 243983 77930 243989
rect 77014 243967 77066 243973
rect 77014 243909 77066 243915
rect 139138 242493 139166 267737
rect 139234 263255 139262 275636
rect 139798 270607 139850 270613
rect 139798 270549 139850 270555
rect 139510 270089 139562 270095
rect 139510 270031 139562 270037
rect 139318 270015 139370 270021
rect 139318 269957 139370 269963
rect 139220 263246 139276 263255
rect 139220 263181 139276 263190
rect 139330 245823 139358 269957
rect 139414 269053 139466 269059
rect 139414 268995 139466 269001
rect 139426 246119 139454 268995
rect 139522 247007 139550 270031
rect 139702 269201 139754 269207
rect 139702 269143 139754 269149
rect 139606 269127 139658 269133
rect 139606 269069 139658 269075
rect 139510 247001 139562 247007
rect 139510 246943 139562 246949
rect 139414 246113 139466 246119
rect 139414 246055 139466 246061
rect 139318 245817 139370 245823
rect 139318 245759 139370 245765
rect 139126 242487 139178 242493
rect 139126 242429 139178 242435
rect 50422 237899 50474 237905
rect 50422 237841 50474 237847
rect 139618 237628 139646 269069
rect 139426 237600 139646 237628
rect 139426 229340 139454 237600
rect 139426 229312 139550 229340
rect 139522 212912 139550 229312
rect 139714 215132 139742 269143
rect 139810 229932 139838 270549
rect 139894 270533 139946 270539
rect 139894 270475 139946 270481
rect 139906 230117 139934 270475
rect 139990 270459 140042 270465
rect 139990 270401 140042 270407
rect 140002 230357 140030 270401
rect 140182 270385 140234 270391
rect 140182 270327 140234 270333
rect 140086 270311 140138 270317
rect 140086 270253 140138 270259
rect 139990 230351 140042 230357
rect 139990 230293 140042 230299
rect 139990 230129 140042 230135
rect 139906 230089 139990 230117
rect 139990 230071 140042 230077
rect 139990 229981 140042 229987
rect 139810 229904 139934 229932
rect 139990 229923 140042 229929
rect 139906 229636 139934 229904
rect 139810 229608 139934 229636
rect 139810 215724 139838 229608
rect 139894 227613 139946 227619
rect 139894 227555 139946 227561
rect 139906 215798 139934 227555
rect 140002 215927 140030 229923
rect 140098 216001 140126 270253
rect 140086 215995 140138 216001
rect 140086 215937 140138 215943
rect 139990 215921 140042 215927
rect 139990 215863 140042 215869
rect 140086 215847 140138 215853
rect 139906 215795 140086 215798
rect 139906 215789 140138 215795
rect 139906 215770 140126 215789
rect 140194 215779 140222 270327
rect 140278 270237 140330 270243
rect 140278 270179 140330 270185
rect 140290 267801 140318 270179
rect 140374 270163 140426 270169
rect 140374 270105 140426 270111
rect 140278 267795 140330 267801
rect 140278 267737 140330 267743
rect 140278 242487 140330 242493
rect 140278 242429 140330 242435
rect 140290 218887 140318 242429
rect 140386 242345 140414 270105
rect 140950 268979 141002 268985
rect 140950 268921 141002 268927
rect 140566 268831 140618 268837
rect 140566 268773 140618 268779
rect 140470 267869 140522 267875
rect 140470 267811 140522 267817
rect 140374 242339 140426 242345
rect 140374 242281 140426 242287
rect 140482 242216 140510 267811
rect 140386 242188 140510 242216
rect 140386 237683 140414 242188
rect 140578 242068 140606 268773
rect 140854 268757 140906 268763
rect 140854 268699 140906 268705
rect 140758 268461 140810 268467
rect 140758 268403 140810 268409
rect 140662 268387 140714 268393
rect 140662 268329 140714 268335
rect 140482 242040 140606 242068
rect 140482 239108 140510 242040
rect 140674 241920 140702 268329
rect 140770 242049 140798 268403
rect 140758 242043 140810 242049
rect 140758 241985 140810 241991
rect 140578 241892 140702 241920
rect 140758 241895 140810 241901
rect 140578 239237 140606 241892
rect 140758 241837 140810 241843
rect 140662 241821 140714 241827
rect 140662 241763 140714 241769
rect 140674 239279 140702 241763
rect 140660 239270 140716 239279
rect 140566 239231 140618 239237
rect 140660 239205 140716 239214
rect 140566 239173 140618 239179
rect 140770 239131 140798 241837
rect 140756 239122 140812 239131
rect 140482 239080 140702 239108
rect 140566 239009 140618 239015
rect 140566 238951 140618 238957
rect 140674 238960 140702 239080
rect 140756 239057 140812 239066
rect 140470 238935 140522 238941
rect 140470 238877 140522 238883
rect 140374 237677 140426 237683
rect 140374 237619 140426 237625
rect 140482 227841 140510 238877
rect 140578 227841 140606 238951
rect 140674 238932 140798 238960
rect 140662 237677 140714 237683
rect 140662 237619 140714 237625
rect 140674 227841 140702 237619
rect 140770 227841 140798 238932
rect 140866 237387 140894 268699
rect 140854 237381 140906 237387
rect 140854 237323 140906 237329
rect 140854 237233 140906 237239
rect 140854 237175 140906 237181
rect 140470 227835 140522 227841
rect 140470 227777 140522 227783
rect 140566 227835 140618 227841
rect 140566 227777 140618 227783
rect 140662 227835 140714 227841
rect 140662 227777 140714 227783
rect 140758 227835 140810 227841
rect 140758 227777 140810 227783
rect 140470 227613 140522 227619
rect 140470 227555 140522 227561
rect 140566 227613 140618 227619
rect 140566 227555 140618 227561
rect 140662 227613 140714 227619
rect 140662 227555 140714 227561
rect 140758 227613 140810 227619
rect 140758 227555 140810 227561
rect 140482 227249 140510 227555
rect 140578 227471 140606 227555
rect 140566 227465 140618 227471
rect 140566 227407 140618 227413
rect 140470 227243 140522 227249
rect 140470 227185 140522 227191
rect 140674 224585 140702 227555
rect 140770 227323 140798 227555
rect 140758 227317 140810 227323
rect 140758 227259 140810 227265
rect 140866 224659 140894 237175
rect 140962 227397 140990 268921
rect 141058 229821 141086 275636
rect 142018 270021 142046 275650
rect 142006 270015 142058 270021
rect 142006 269957 142058 269963
rect 143170 268879 143198 275650
rect 143156 268870 143212 268879
rect 143156 268805 143212 268814
rect 141142 265131 141194 265137
rect 141142 265073 141194 265079
rect 141154 264989 141182 265073
rect 141142 264983 141194 264989
rect 141142 264925 141194 264931
rect 144706 262177 144734 275784
rect 145570 263953 145598 275650
rect 146736 275636 147038 275664
rect 145558 263947 145610 263953
rect 145558 263889 145610 263895
rect 147010 263879 147038 275636
rect 147970 267875 147998 275650
rect 147958 267869 148010 267875
rect 147958 267811 148010 267817
rect 149122 264027 149150 275650
rect 149686 267869 149738 267875
rect 149686 267811 149738 267817
rect 149110 264021 149162 264027
rect 149110 263963 149162 263969
rect 146998 263873 147050 263879
rect 146998 263815 147050 263821
rect 144694 262171 144746 262177
rect 144694 262113 144746 262119
rect 146614 262171 146666 262177
rect 146614 262113 146666 262119
rect 146626 259217 146654 262113
rect 146518 259211 146570 259217
rect 146518 259153 146570 259159
rect 146614 259211 146666 259217
rect 146614 259153 146666 259159
rect 141430 247001 141482 247007
rect 141430 246943 141482 246949
rect 141334 242339 141386 242345
rect 141334 242281 141386 242287
rect 141142 242043 141194 242049
rect 141142 241985 141194 241991
rect 141154 238941 141182 241985
rect 141142 238935 141194 238941
rect 141142 238877 141194 238883
rect 141238 237381 141290 237387
rect 141238 237323 141290 237329
rect 141058 229793 141182 229821
rect 141154 227416 141182 229793
rect 141250 227545 141278 237323
rect 141346 237239 141374 242281
rect 141334 237233 141386 237239
rect 141334 237175 141386 237181
rect 141442 230357 141470 246943
rect 141526 246113 141578 246119
rect 141526 246055 141578 246061
rect 141538 230431 141566 246055
rect 143158 245817 143210 245823
rect 143158 245759 143210 245765
rect 141526 230425 141578 230431
rect 141526 230367 141578 230373
rect 141430 230351 141482 230357
rect 141430 230293 141482 230299
rect 143170 230135 143198 245759
rect 146036 240602 146092 240611
rect 146036 240537 146092 240546
rect 144020 239862 144076 239871
rect 144020 239797 144076 239806
rect 144034 239089 144062 239797
rect 144022 239083 144074 239089
rect 144022 239025 144074 239031
rect 144116 238678 144172 238687
rect 144116 238613 144172 238622
rect 144020 236310 144076 236319
rect 144020 236245 144022 236254
rect 144074 236245 144076 236254
rect 144022 236213 144074 236219
rect 144130 236203 144158 238613
rect 144118 236197 144170 236203
rect 144118 236139 144170 236145
rect 144020 233646 144076 233655
rect 144020 233581 144076 233590
rect 144034 233317 144062 233581
rect 144022 233311 144074 233317
rect 144022 233253 144074 233259
rect 144116 232166 144172 232175
rect 144116 232101 144172 232110
rect 144020 231426 144076 231435
rect 144020 231361 144076 231370
rect 144034 230579 144062 231361
rect 144022 230573 144074 230579
rect 144022 230515 144074 230521
rect 144130 230505 144158 232101
rect 144118 230499 144170 230505
rect 144118 230441 144170 230447
rect 144212 230242 144268 230251
rect 144212 230177 144268 230186
rect 141334 230129 141386 230135
rect 141334 230071 141386 230077
rect 143158 230129 143210 230135
rect 143158 230071 143210 230077
rect 141346 227915 141374 230071
rect 144020 228466 144076 228475
rect 144020 228401 144076 228410
rect 141334 227909 141386 227915
rect 141334 227851 141386 227857
rect 144034 227767 144062 228401
rect 144022 227761 144074 227767
rect 144022 227703 144074 227709
rect 144116 227726 144172 227735
rect 144226 227693 144254 230177
rect 144116 227661 144172 227670
rect 144214 227687 144266 227693
rect 144130 227619 144158 227661
rect 144214 227629 144266 227635
rect 144118 227613 144170 227619
rect 144118 227555 144170 227561
rect 141238 227539 141290 227545
rect 141238 227481 141290 227487
rect 140950 227391 141002 227397
rect 140950 227333 141002 227339
rect 141058 227388 141182 227416
rect 140854 224653 140906 224659
rect 140854 224595 140906 224601
rect 140662 224579 140714 224585
rect 140662 224521 140714 224527
rect 141058 224511 141086 227388
rect 144020 226690 144076 226699
rect 144020 226625 144076 226634
rect 144034 225695 144062 226625
rect 144022 225689 144074 225695
rect 144022 225631 144074 225637
rect 144020 225062 144076 225071
rect 144020 224997 144076 225006
rect 144034 224733 144062 224997
rect 144022 224727 144074 224733
rect 144022 224669 144074 224675
rect 141046 224505 141098 224511
rect 141046 224447 141098 224453
rect 144116 223730 144172 223739
rect 144116 223665 144172 223674
rect 144020 222990 144076 222999
rect 144020 222925 144076 222934
rect 144034 221921 144062 222925
rect 144022 221915 144074 221921
rect 144022 221857 144074 221863
rect 144130 221847 144158 223665
rect 144118 221841 144170 221847
rect 144118 221783 144170 221789
rect 144020 220178 144076 220187
rect 144020 220113 144076 220122
rect 144034 218961 144062 220113
rect 144022 218955 144074 218961
rect 144022 218897 144074 218903
rect 140278 218881 140330 218887
rect 140278 218823 140330 218829
rect 144020 218254 144076 218263
rect 144020 218189 144076 218198
rect 144034 216741 144062 218189
rect 144022 216735 144074 216741
rect 144022 216677 144074 216683
rect 140182 215773 140234 215779
rect 139810 215696 140126 215724
rect 140182 215715 140234 215721
rect 140098 215576 140126 215696
rect 140098 215548 140318 215576
rect 139714 215104 140030 215132
rect 140002 213041 140030 215104
rect 140086 213109 140138 213115
rect 140086 213051 140138 213057
rect 139990 213035 140042 213041
rect 139990 212977 140042 212983
rect 140098 212912 140126 213051
rect 140290 213041 140318 215548
rect 144116 215294 144172 215303
rect 144116 215229 144172 215238
rect 144020 213370 144076 213379
rect 144020 213305 144076 213314
rect 144034 213263 144062 213305
rect 144022 213257 144074 213263
rect 144022 213199 144074 213205
rect 144130 213189 144158 215229
rect 145364 214554 145420 214563
rect 145364 214489 145420 214498
rect 144118 213183 144170 213189
rect 144118 213125 144170 213131
rect 140278 213035 140330 213041
rect 140278 212977 140330 212983
rect 139522 212884 140126 212912
rect 144020 211742 144076 211751
rect 144020 211677 144076 211686
rect 144034 210303 144062 211677
rect 144022 210297 144074 210303
rect 144022 210239 144074 210245
rect 144116 209818 144172 209827
rect 144116 209753 144172 209762
rect 144022 207485 144074 207491
rect 144020 207450 144022 207459
rect 144074 207450 144076 207459
rect 144130 207417 144158 209753
rect 144020 207385 144076 207394
rect 144118 207411 144170 207417
rect 144118 207353 144170 207359
rect 144212 203306 144268 203315
rect 144212 203241 144268 203250
rect 144226 201645 144254 203241
rect 144214 201639 144266 201645
rect 144214 201581 144266 201587
rect 144788 196646 144844 196655
rect 144788 196581 144844 196590
rect 144596 194870 144652 194879
rect 144596 194805 144652 194814
rect 47638 194535 47690 194541
rect 47638 194477 47690 194483
rect 43126 193499 43178 193505
rect 43126 193441 43178 193447
rect 43030 192241 43082 192247
rect 43030 192183 43082 192189
rect 42658 188168 42974 188196
rect 42166 187135 42218 187141
rect 42166 187077 42218 187083
rect 42454 187135 42506 187141
rect 42454 187077 42506 187083
rect 42178 186776 42206 187077
rect 42658 186549 42686 188168
rect 42742 187875 42794 187881
rect 42742 187817 42794 187823
rect 42070 186543 42122 186549
rect 42070 186485 42122 186491
rect 42646 186543 42698 186549
rect 42646 186485 42698 186491
rect 42082 186184 42110 186485
rect 41780 185990 41836 185999
rect 41780 185925 41836 185934
rect 41794 185592 41822 185925
rect 41780 184214 41836 184223
rect 41780 184149 41836 184158
rect 41794 183742 41822 184149
rect 41780 183622 41836 183631
rect 41780 183557 41836 183566
rect 41794 183121 41822 183557
rect 41780 182882 41836 182891
rect 41780 182817 41836 182826
rect 41794 182484 41822 182817
rect 42754 177119 42782 187817
rect 144020 184510 144076 184519
rect 144020 184445 144076 184454
rect 144034 184403 144062 184445
rect 144022 184397 144074 184403
rect 144022 184339 144074 184345
rect 144020 181846 144076 181855
rect 144020 181781 144076 181790
rect 144034 181517 144062 181781
rect 144022 181511 144074 181517
rect 144022 181453 144074 181459
rect 144116 180514 144172 180523
rect 144116 180449 144172 180458
rect 144130 178705 144158 180449
rect 144118 178699 144170 178705
rect 144118 178641 144170 178647
rect 144022 178625 144074 178631
rect 144020 178590 144022 178599
rect 144074 178590 144076 178599
rect 144020 178525 144076 178534
rect 42740 177110 42796 177119
rect 42740 177045 42796 177054
rect 144020 176814 144076 176823
rect 144020 176749 144076 176758
rect 144034 175745 144062 176749
rect 144022 175739 144074 175745
rect 144022 175681 144074 175687
rect 144020 173410 144076 173419
rect 144020 173345 144076 173354
rect 144034 172859 144062 173345
rect 144022 172853 144074 172859
rect 144022 172795 144074 172801
rect 144020 171338 144076 171347
rect 144020 171273 144076 171282
rect 144034 170417 144062 171273
rect 144022 170411 144074 170417
rect 144022 170353 144074 170359
rect 144116 168378 144172 168387
rect 144116 168313 144172 168322
rect 144020 167638 144076 167647
rect 144020 167573 144076 167582
rect 144034 167161 144062 167573
rect 144022 167155 144074 167161
rect 144022 167097 144074 167103
rect 144130 167087 144158 168313
rect 144118 167081 144170 167087
rect 144118 167023 144170 167029
rect 144020 166602 144076 166611
rect 144020 166537 144076 166546
rect 144034 164201 144062 166537
rect 144022 164195 144074 164201
rect 144022 164137 144074 164143
rect 144116 163642 144172 163651
rect 144116 163577 144172 163586
rect 144020 162902 144076 162911
rect 144020 162837 144076 162846
rect 144034 161389 144062 162837
rect 144022 161383 144074 161389
rect 144022 161325 144074 161331
rect 144130 161315 144158 163577
rect 144118 161309 144170 161315
rect 144118 161251 144170 161257
rect 144500 159942 144556 159951
rect 144500 159877 144556 159886
rect 144020 159350 144076 159359
rect 144020 159285 144076 159294
rect 144034 158503 144062 159285
rect 144022 158497 144074 158503
rect 144022 158439 144074 158445
rect 144308 158166 144364 158175
rect 144308 158101 144364 158110
rect 144212 156390 144268 156399
rect 144212 156325 144268 156334
rect 144020 155650 144076 155659
rect 144020 155585 144022 155594
rect 144074 155585 144076 155594
rect 144022 155553 144074 155559
rect 144116 154466 144172 154475
rect 144116 154401 144172 154410
rect 144020 152986 144076 152995
rect 144020 152921 144076 152930
rect 144034 152805 144062 152921
rect 144022 152799 144074 152805
rect 144022 152741 144074 152747
rect 144130 152731 144158 154401
rect 144118 152725 144170 152731
rect 144118 152667 144170 152673
rect 144116 151654 144172 151663
rect 144116 151589 144172 151598
rect 144020 150914 144076 150923
rect 144020 150849 144076 150858
rect 144034 149845 144062 150849
rect 144130 149919 144158 151589
rect 144118 149913 144170 149919
rect 144118 149855 144170 149861
rect 144022 149839 144074 149845
rect 144022 149781 144074 149787
rect 144226 149728 144254 156325
rect 144130 149700 144254 149728
rect 144022 149691 144074 149697
rect 144022 149633 144074 149639
rect 144034 147280 144062 149633
rect 143938 147252 144062 147280
rect 143938 146904 143966 147252
rect 144020 147214 144076 147223
rect 144020 147149 144076 147158
rect 144034 147033 144062 147149
rect 144022 147027 144074 147033
rect 144022 146969 144074 146975
rect 143938 146876 144062 146904
rect 141524 137594 141580 137603
rect 141524 137529 141580 137538
rect 141538 121027 141566 137529
rect 143926 134151 143978 134157
rect 143926 134093 143978 134099
rect 143938 132455 143966 134093
rect 143926 132449 143978 132455
rect 143926 132391 143978 132397
rect 141524 121018 141580 121027
rect 141524 120953 141580 120962
rect 141044 118650 141100 118659
rect 141044 118585 141100 118594
rect 141058 118363 141086 118585
rect 141044 118354 141100 118363
rect 141044 118289 141100 118298
rect 143926 106771 143978 106777
rect 143926 106713 143978 106719
rect 143938 106407 143966 106713
rect 144034 106555 144062 146876
rect 144022 106549 144074 106555
rect 144022 106491 144074 106497
rect 143926 106401 143978 106407
rect 143926 106343 143978 106349
rect 144130 106037 144158 149700
rect 144322 149697 144350 158101
rect 144310 149691 144362 149697
rect 144310 149633 144362 149639
rect 144514 149549 144542 159877
rect 144310 149543 144362 149549
rect 144310 149485 144362 149491
rect 144502 149543 144554 149549
rect 144502 149485 144554 149491
rect 144212 147954 144268 147963
rect 144212 147889 144268 147898
rect 144226 146959 144254 147889
rect 144214 146953 144266 146959
rect 144214 146895 144266 146901
rect 144212 146030 144268 146039
rect 144212 145965 144268 145974
rect 144226 144073 144254 145965
rect 144214 144067 144266 144073
rect 144214 144009 144266 144015
rect 144212 142478 144268 142487
rect 144212 142413 144268 142422
rect 144226 141187 144254 142413
rect 144214 141181 144266 141187
rect 144214 141123 144266 141129
rect 144214 141033 144266 141039
rect 144214 140975 144266 140981
rect 144226 138597 144254 140975
rect 144214 138591 144266 138597
rect 144214 138533 144266 138539
rect 144212 138482 144268 138491
rect 144212 138417 144268 138426
rect 144226 138375 144254 138417
rect 144214 138369 144266 138375
rect 144214 138311 144266 138317
rect 144212 132858 144268 132867
rect 144212 132793 144268 132802
rect 144226 132529 144254 132793
rect 144214 132523 144266 132529
rect 144214 132465 144266 132471
rect 144212 131082 144268 131091
rect 144212 131017 144268 131026
rect 144226 130161 144254 131017
rect 144214 130155 144266 130161
rect 144214 130097 144266 130103
rect 144212 130046 144268 130055
rect 144212 129981 144268 129990
rect 144226 129643 144254 129981
rect 144214 129637 144266 129643
rect 144214 129579 144266 129585
rect 144214 129489 144266 129495
rect 144214 129431 144266 129437
rect 144118 106031 144170 106037
rect 144118 105973 144170 105979
rect 144116 105922 144172 105931
rect 144116 105857 144172 105866
rect 144020 104886 144076 104895
rect 144020 104821 144076 104830
rect 144034 104409 144062 104821
rect 144022 104403 144074 104409
rect 144022 104345 144074 104351
rect 144022 104255 144074 104261
rect 144022 104197 144074 104203
rect 144034 104007 144062 104197
rect 144020 103998 144076 104007
rect 144020 103933 144076 103942
rect 144130 103743 144158 105857
rect 144118 103737 144170 103743
rect 144118 103679 144170 103685
rect 144116 102814 144172 102823
rect 144116 102749 144172 102758
rect 144020 101334 144076 101343
rect 144020 101269 144076 101278
rect 144034 100931 144062 101269
rect 144022 100925 144074 100931
rect 144022 100867 144074 100873
rect 144130 100857 144158 102749
rect 144118 100851 144170 100857
rect 144118 100793 144170 100799
rect 144020 99854 144076 99863
rect 144020 99789 144076 99798
rect 144034 98341 144062 99789
rect 144116 99114 144172 99123
rect 144116 99049 144172 99058
rect 144022 98335 144074 98341
rect 144022 98277 144074 98283
rect 144020 98078 144076 98087
rect 144020 98013 144022 98022
rect 144074 98013 144076 98022
rect 144022 97981 144074 97987
rect 144130 97971 144158 99049
rect 144118 97965 144170 97971
rect 144118 97907 144170 97913
rect 144020 96302 144076 96311
rect 144020 96237 144076 96246
rect 144034 95085 144062 96237
rect 144022 95079 144074 95085
rect 144022 95021 144074 95027
rect 144116 94378 144172 94387
rect 144116 94313 144172 94322
rect 144020 92750 144076 92759
rect 144020 92685 144076 92694
rect 144034 92199 144062 92685
rect 144130 92273 144158 94313
rect 144118 92267 144170 92273
rect 144118 92209 144170 92215
rect 144022 92193 144074 92199
rect 144022 92135 144074 92141
rect 144118 91231 144170 91237
rect 144118 91173 144170 91179
rect 144130 90960 144158 91173
rect 144226 91108 144254 129431
rect 144322 106523 144350 149485
rect 144500 149138 144556 149147
rect 144500 149073 144556 149082
rect 144404 143218 144460 143227
rect 144404 143153 144460 143162
rect 144418 141261 144446 143153
rect 144406 141255 144458 141261
rect 144406 141197 144458 141203
rect 144404 139518 144460 139527
rect 144404 139453 144460 139462
rect 144418 138301 144446 139453
rect 144406 138295 144458 138301
rect 144406 138237 144458 138243
rect 144406 138147 144458 138153
rect 144406 138089 144458 138095
rect 144418 136692 144446 138089
rect 144514 136821 144542 149073
rect 144502 136815 144554 136821
rect 144502 136757 144554 136763
rect 144418 136664 144542 136692
rect 144406 136297 144458 136303
rect 144406 136239 144458 136245
rect 144418 134157 144446 136239
rect 144514 135489 144542 136664
rect 144610 136229 144638 194805
rect 144694 144363 144746 144369
rect 144694 144305 144746 144311
rect 144706 141409 144734 144305
rect 144694 141403 144746 141409
rect 144694 141345 144746 141351
rect 144692 141294 144748 141303
rect 144692 141229 144748 141238
rect 144706 136303 144734 141229
rect 144694 136297 144746 136303
rect 144694 136239 144746 136245
rect 144598 136223 144650 136229
rect 144598 136165 144650 136171
rect 144598 136001 144650 136007
rect 144598 135943 144650 135949
rect 144692 135966 144748 135975
rect 144502 135483 144554 135489
rect 144502 135425 144554 135431
rect 144500 135078 144556 135087
rect 144500 135013 144556 135022
rect 144406 134151 144458 134157
rect 144406 134093 144458 134099
rect 144404 134042 144460 134051
rect 144404 133977 144460 133986
rect 144418 132603 144446 133977
rect 144514 132751 144542 135013
rect 144502 132745 144554 132751
rect 144502 132687 144554 132693
rect 144406 132597 144458 132603
rect 144406 132539 144458 132545
rect 144502 132449 144554 132455
rect 144502 132391 144554 132397
rect 144404 121018 144460 121027
rect 144404 120953 144460 120962
rect 144308 106514 144364 106523
rect 144308 106449 144364 106458
rect 144310 106401 144362 106407
rect 144310 106343 144362 106349
rect 144322 100709 144350 106343
rect 144310 100703 144362 100709
rect 144310 100645 144362 100651
rect 144418 95548 144446 120953
rect 144322 95520 144446 95548
rect 144322 91237 144350 95520
rect 144406 95449 144458 95455
rect 144406 95391 144458 95397
rect 144310 91231 144362 91237
rect 144310 91173 144362 91179
rect 144226 91080 144350 91108
rect 144130 90932 144254 90960
rect 144116 90826 144172 90835
rect 144116 90761 144172 90770
rect 144020 89642 144076 89651
rect 144020 89577 144076 89586
rect 144034 89461 144062 89577
rect 144022 89455 144074 89461
rect 144022 89397 144074 89403
rect 144130 89387 144158 90761
rect 144118 89381 144170 89387
rect 144118 89323 144170 89329
rect 144118 89233 144170 89239
rect 144118 89175 144170 89181
rect 144020 87866 144076 87875
rect 144020 87801 144076 87810
rect 144034 86501 144062 87801
rect 144022 86495 144074 86501
rect 144022 86437 144074 86443
rect 144020 85942 144076 85951
rect 144020 85877 144076 85886
rect 144034 85021 144062 85877
rect 144022 85015 144074 85021
rect 144022 84957 144074 84963
rect 144020 82390 144076 82399
rect 144020 82325 144076 82334
rect 144034 82135 144062 82325
rect 144022 82129 144074 82135
rect 144022 82071 144074 82077
rect 144020 81206 144076 81215
rect 144020 81141 144076 81150
rect 144034 80803 144062 81141
rect 144022 80797 144074 80803
rect 144022 80739 144074 80745
rect 144130 80729 144158 89175
rect 144118 80723 144170 80729
rect 144118 80665 144170 80671
rect 144116 79430 144172 79439
rect 144116 79365 144172 79374
rect 144020 78690 144076 78699
rect 144020 78625 144076 78634
rect 144034 77917 144062 78625
rect 144022 77911 144074 77917
rect 144022 77853 144074 77859
rect 144130 77843 144158 79365
rect 144118 77837 144170 77843
rect 144118 77779 144170 77785
rect 144118 76579 144170 76585
rect 144118 76521 144170 76527
rect 144130 75864 144158 76521
rect 144226 76363 144254 90932
rect 144214 76357 144266 76363
rect 144214 76299 144266 76305
rect 144130 75836 144254 75864
rect 144116 75730 144172 75739
rect 144116 75665 144172 75674
rect 144020 75138 144076 75147
rect 144020 75073 144076 75082
rect 144034 74957 144062 75073
rect 144130 75031 144158 75665
rect 144118 75025 144170 75031
rect 144118 74967 144170 74973
rect 144022 74951 144074 74957
rect 144022 74893 144074 74899
rect 144118 74877 144170 74883
rect 144118 74819 144170 74825
rect 144020 73954 144076 73963
rect 144020 73889 144076 73898
rect 144034 72071 144062 73889
rect 144130 72779 144158 74819
rect 144116 72770 144172 72779
rect 144116 72705 144172 72714
rect 144118 72657 144170 72663
rect 144118 72599 144170 72605
rect 144022 72065 144074 72071
rect 144022 72007 144074 72013
rect 144020 70994 144076 71003
rect 144020 70929 144076 70938
rect 144034 70295 144062 70929
rect 144022 70289 144074 70295
rect 144022 70231 144074 70237
rect 144020 69810 144076 69819
rect 144020 69745 144076 69754
rect 144034 69185 144062 69745
rect 144022 69179 144074 69185
rect 144022 69121 144074 69127
rect 144020 67590 144076 67599
rect 144020 67525 144076 67534
rect 144034 67039 144062 67525
rect 144022 67033 144074 67039
rect 144022 66975 144074 66981
rect 144020 66406 144076 66415
rect 144020 66341 144076 66350
rect 144034 66299 144062 66341
rect 144022 66293 144074 66299
rect 144022 66235 144074 66241
rect 144022 64813 144074 64819
rect 144020 64778 144022 64787
rect 144074 64778 144076 64787
rect 144020 64713 144076 64722
rect 144020 62706 144076 62715
rect 144020 62641 144076 62650
rect 144034 62229 144062 62641
rect 144022 62223 144074 62229
rect 144022 62165 144074 62171
rect 144022 59041 144074 59047
rect 144022 58983 144074 58989
rect 144034 58719 144062 58983
rect 144020 58710 144076 58719
rect 144130 58677 144158 72599
rect 144226 69407 144254 75836
rect 144322 72663 144350 91080
rect 144418 76511 144446 95391
rect 144406 76505 144458 76511
rect 144406 76447 144458 76453
rect 144406 76357 144458 76363
rect 144406 76299 144458 76305
rect 144310 72657 144362 72663
rect 144310 72599 144362 72605
rect 144310 72509 144362 72515
rect 144310 72451 144362 72457
rect 144214 69401 144266 69407
rect 144214 69343 144266 69349
rect 144212 69070 144268 69079
rect 144212 69005 144268 69014
rect 144226 66595 144254 69005
rect 144214 66589 144266 66595
rect 144214 66531 144266 66537
rect 144214 66219 144266 66225
rect 144214 66161 144266 66167
rect 144020 58645 144076 58654
rect 144118 58671 144170 58677
rect 144118 58613 144170 58619
rect 144226 58548 144254 66161
rect 144034 58520 144254 58548
rect 144034 57660 144062 58520
rect 144214 58449 144266 58455
rect 144214 58391 144266 58397
rect 143938 57632 144062 57660
rect 143938 57216 143966 57632
rect 144022 57561 144074 57567
rect 144022 57503 144074 57509
rect 144034 57387 144062 57503
rect 144118 57487 144170 57493
rect 144118 57429 144170 57435
rect 144020 57378 144076 57387
rect 144020 57313 144076 57322
rect 143938 57188 144062 57216
rect 144034 56328 144062 57188
rect 144130 56499 144158 57429
rect 144116 56490 144172 56499
rect 144116 56425 144172 56434
rect 144034 56300 144158 56328
rect 144020 54714 144076 54723
rect 144020 54649 144022 54658
rect 144074 54649 144076 54658
rect 144022 54617 144074 54623
rect 144022 54157 144074 54163
rect 144022 54099 144074 54105
rect 144034 53835 144062 54099
rect 144020 53826 144076 53835
rect 144020 53761 144076 53770
rect 144130 50537 144158 56300
rect 144118 50531 144170 50537
rect 144118 50473 144170 50479
rect 144226 50167 144254 58391
rect 144214 50161 144266 50167
rect 144214 50103 144266 50109
rect 144322 49797 144350 72451
rect 144418 50093 144446 76299
rect 144406 50087 144458 50093
rect 144406 50029 144458 50035
rect 144514 50019 144542 132391
rect 144610 124537 144638 135943
rect 144692 135901 144748 135910
rect 144706 129495 144734 135901
rect 144694 129489 144746 129495
rect 144694 129431 144746 129437
rect 144694 129341 144746 129347
rect 144694 129283 144746 129289
rect 144598 124531 144650 124537
rect 144598 124473 144650 124479
rect 144596 124422 144652 124431
rect 144596 124357 144652 124366
rect 144610 124019 144638 124357
rect 144598 124013 144650 124019
rect 144598 123955 144650 123961
rect 144596 121610 144652 121619
rect 144596 121545 144652 121554
rect 144610 121207 144638 121545
rect 144598 121201 144650 121207
rect 144598 121143 144650 121149
rect 144596 120870 144652 120879
rect 144596 120805 144652 120814
rect 144610 118617 144638 120805
rect 144598 118611 144650 118617
rect 144598 118553 144650 118559
rect 144596 118354 144652 118363
rect 144596 118289 144598 118298
rect 144650 118289 144652 118298
rect 144598 118257 144650 118263
rect 144596 116726 144652 116735
rect 144596 116661 144652 116670
rect 144610 115287 144638 116661
rect 144598 115281 144650 115287
rect 144598 115223 144650 115229
rect 144596 114210 144652 114219
rect 144596 114145 144652 114154
rect 144610 112549 144638 114145
rect 144598 112543 144650 112549
rect 144598 112485 144650 112491
rect 144596 112434 144652 112443
rect 144596 112369 144598 112378
rect 144650 112369 144652 112378
rect 144598 112337 144650 112343
rect 144596 109770 144652 109779
rect 144596 109705 144652 109714
rect 144610 109515 144638 109705
rect 144598 109509 144650 109515
rect 144598 109451 144650 109457
rect 144596 107550 144652 107559
rect 144596 107485 144598 107494
rect 144650 107485 144652 107494
rect 144598 107453 144650 107459
rect 144706 106671 144734 129283
rect 144802 125351 144830 196581
rect 144884 174446 144940 174455
rect 144884 174381 144940 174390
rect 144898 157171 144926 174381
rect 145076 172078 145132 172087
rect 145076 172013 145132 172022
rect 144980 161422 145036 161431
rect 144980 161357 145036 161366
rect 144886 157165 144938 157171
rect 144886 157107 144938 157113
rect 144886 157017 144938 157023
rect 144886 156959 144938 156965
rect 144898 144369 144926 156959
rect 144886 144363 144938 144369
rect 144886 144305 144938 144311
rect 144884 144254 144940 144263
rect 144884 144189 144940 144198
rect 144898 136969 144926 144189
rect 144886 136963 144938 136969
rect 144886 136905 144938 136911
rect 144886 136815 144938 136821
rect 144886 136757 144938 136763
rect 144790 125345 144842 125351
rect 144790 125287 144842 125293
rect 144788 125162 144844 125171
rect 144788 125097 144844 125106
rect 144802 123945 144830 125097
rect 144790 123939 144842 123945
rect 144790 123881 144842 123887
rect 144788 122646 144844 122655
rect 144788 122581 144844 122590
rect 144802 121059 144830 122581
rect 144790 121053 144842 121059
rect 144790 120995 144842 121001
rect 144788 119094 144844 119103
rect 144788 119029 144844 119038
rect 144802 118173 144830 119029
rect 144790 118167 144842 118173
rect 144790 118109 144842 118115
rect 144790 118019 144842 118025
rect 144790 117961 144842 117967
rect 144802 113289 144830 117961
rect 144790 113283 144842 113289
rect 144790 113225 144842 113231
rect 144788 113174 144844 113183
rect 144788 113109 144844 113118
rect 144802 112475 144830 113109
rect 144790 112469 144842 112475
rect 144790 112411 144842 112417
rect 144788 111250 144844 111259
rect 144788 111185 144844 111194
rect 144802 109589 144830 111185
rect 144790 109583 144842 109589
rect 144790 109525 144842 109531
rect 144790 109435 144842 109441
rect 144790 109377 144842 109383
rect 144802 106777 144830 109377
rect 144790 106771 144842 106777
rect 144790 106713 144842 106719
rect 144692 106662 144748 106671
rect 144692 106597 144748 106606
rect 144790 106623 144842 106629
rect 144790 106565 144842 106571
rect 144596 106366 144652 106375
rect 144596 106301 144652 106310
rect 144610 94715 144638 106301
rect 144802 103595 144830 106565
rect 144790 103589 144842 103595
rect 144790 103531 144842 103537
rect 144692 100890 144748 100899
rect 144692 100825 144748 100834
rect 144706 100691 144734 100825
rect 144706 100663 144830 100691
rect 144598 94709 144650 94715
rect 144598 94651 144650 94657
rect 144802 89239 144830 100663
rect 144790 89233 144842 89239
rect 144790 89175 144842 89181
rect 144788 87126 144844 87135
rect 144788 87061 144844 87070
rect 144598 86421 144650 86427
rect 144598 86363 144650 86369
rect 144610 76585 144638 86363
rect 144694 80723 144746 80729
rect 144694 80665 144746 80671
rect 144598 76579 144650 76585
rect 144598 76521 144650 76527
rect 144598 76357 144650 76363
rect 144598 76299 144650 76305
rect 144502 50013 144554 50019
rect 144502 49955 144554 49961
rect 144310 49791 144362 49797
rect 144310 49733 144362 49739
rect 144610 49649 144638 76299
rect 144706 66225 144734 80665
rect 144802 76289 144830 87061
rect 144898 86427 144926 136757
rect 144886 86421 144938 86427
rect 144886 86363 144938 86369
rect 144790 76283 144842 76289
rect 144790 76225 144842 76231
rect 144790 72731 144842 72737
rect 144790 72673 144842 72679
rect 144694 66219 144746 66225
rect 144694 66161 144746 66167
rect 144598 49643 144650 49649
rect 144598 49585 144650 49591
rect 144802 49575 144830 72673
rect 144886 66367 144938 66373
rect 144886 66309 144938 66315
rect 144898 50463 144926 66309
rect 144994 51425 145022 161357
rect 144982 51419 145034 51425
rect 144982 51361 145034 51367
rect 145090 50907 145118 172013
rect 145268 170154 145324 170163
rect 145268 170089 145324 170098
rect 145172 164826 145228 164835
rect 145172 164761 145228 164770
rect 145186 76363 145214 164761
rect 145174 76357 145226 76363
rect 145174 76299 145226 76305
rect 145174 76209 145226 76215
rect 145174 76151 145226 76157
rect 145186 72219 145214 76151
rect 145174 72213 145226 72219
rect 145174 72155 145226 72161
rect 145174 69549 145226 69555
rect 145174 69491 145226 69497
rect 145078 50901 145130 50907
rect 145078 50843 145130 50849
rect 144886 50457 144938 50463
rect 144886 50399 144938 50405
rect 145186 49945 145214 69491
rect 145282 50759 145310 170089
rect 145378 72737 145406 214489
rect 145460 210558 145516 210567
rect 145460 210493 145516 210502
rect 145366 72731 145418 72737
rect 145366 72673 145418 72679
rect 145366 72583 145418 72589
rect 145366 72525 145418 72531
rect 145270 50753 145322 50759
rect 145270 50695 145322 50701
rect 145378 50611 145406 72525
rect 145474 51351 145502 210493
rect 145556 208042 145612 208051
rect 145556 207977 145612 207986
rect 145570 69555 145598 207977
rect 145652 205674 145708 205683
rect 145652 205609 145708 205618
rect 145558 69549 145610 69555
rect 145558 69491 145610 69497
rect 145558 69401 145610 69407
rect 145558 69343 145610 69349
rect 145570 66373 145598 69343
rect 145558 66367 145610 66373
rect 145558 66309 145610 66315
rect 145558 66071 145610 66077
rect 145558 66013 145610 66019
rect 145462 51345 145514 51351
rect 145462 51287 145514 51293
rect 145366 50605 145418 50611
rect 145366 50547 145418 50553
rect 145174 49939 145226 49945
rect 145174 49881 145226 49887
rect 145570 49871 145598 66013
rect 145666 51277 145694 205609
rect 145844 205082 145900 205091
rect 145844 205017 145900 205026
rect 145748 201382 145804 201391
rect 145748 201317 145804 201326
rect 145762 51647 145790 201317
rect 145858 66077 145886 205017
rect 145940 190134 145996 190143
rect 145940 190069 145996 190078
rect 145954 83689 145982 190069
rect 146050 140521 146078 240537
rect 146530 239071 146558 259153
rect 149590 244041 149642 244047
rect 149590 243983 149642 243989
rect 149602 240463 149630 243983
rect 149588 240454 149644 240463
rect 149588 240389 149644 240398
rect 146530 239043 146846 239071
rect 146228 236902 146284 236911
rect 146228 236837 146284 236846
rect 146132 186434 146188 186443
rect 146132 186369 146188 186378
rect 146038 140515 146090 140521
rect 146038 140457 146090 140463
rect 146038 124531 146090 124537
rect 146038 124473 146090 124479
rect 146050 109441 146078 124473
rect 146038 109435 146090 109441
rect 146038 109377 146090 109383
rect 146036 108290 146092 108299
rect 146036 108225 146092 108234
rect 146050 106629 146078 108225
rect 146038 106623 146090 106629
rect 146038 106565 146090 106571
rect 146038 106031 146090 106037
rect 146038 105973 146090 105979
rect 146050 92051 146078 105973
rect 146038 92045 146090 92051
rect 146038 91987 146090 91993
rect 145942 83683 145994 83689
rect 145942 83625 145994 83631
rect 145940 83574 145996 83583
rect 145940 83509 145996 83518
rect 145846 66071 145898 66077
rect 145846 66013 145898 66019
rect 145954 65948 145982 83509
rect 146038 76283 146090 76289
rect 146038 76225 146090 76231
rect 145858 65920 145982 65948
rect 145750 51641 145802 51647
rect 145750 51583 145802 51589
rect 145654 51271 145706 51277
rect 145654 51213 145706 51219
rect 145858 50241 145886 65920
rect 146050 65800 146078 76225
rect 145954 65772 146078 65800
rect 145954 50389 145982 65772
rect 146038 65627 146090 65633
rect 146038 65569 146090 65575
rect 145942 50383 145994 50389
rect 145942 50325 145994 50331
rect 146050 50315 146078 65569
rect 146146 51203 146174 186369
rect 146242 116693 146270 236837
rect 146420 235126 146476 235135
rect 146420 235061 146476 235070
rect 146434 221773 146462 235061
rect 146818 224437 146846 239043
rect 146902 230129 146954 230135
rect 146900 230094 146902 230103
rect 146954 230094 146956 230103
rect 146900 230029 146956 230038
rect 146806 224431 146858 224437
rect 146806 224373 146858 224379
rect 149698 224363 149726 267811
rect 150274 264101 150302 275650
rect 151426 267875 151454 275650
rect 152674 270243 152702 275650
rect 152662 270237 152714 270243
rect 152662 270179 152714 270185
rect 153826 270095 153854 275650
rect 153814 270089 153866 270095
rect 153814 270031 153866 270037
rect 151414 267869 151466 267875
rect 151414 267811 151466 267817
rect 152566 267869 152618 267875
rect 152566 267811 152618 267817
rect 151126 265131 151178 265137
rect 151126 265073 151178 265079
rect 151138 264989 151166 265073
rect 151126 264983 151178 264989
rect 151126 264925 151178 264931
rect 150262 264095 150314 264101
rect 150262 264037 150314 264043
rect 152470 243967 152522 243973
rect 152470 243909 152522 243915
rect 152482 241901 152510 243909
rect 152470 241895 152522 241901
rect 152470 241837 152522 241843
rect 151126 230573 151178 230579
rect 151126 230515 151178 230521
rect 149686 224357 149738 224363
rect 149686 224299 149738 224305
rect 146422 221767 146474 221773
rect 146422 221709 146474 221715
rect 146710 221767 146762 221773
rect 146710 221709 146762 221715
rect 146722 207343 146750 221709
rect 148246 210297 148298 210303
rect 148246 210239 148298 210245
rect 146422 207337 146474 207343
rect 146422 207279 146474 207285
rect 146710 207337 146762 207343
rect 146710 207279 146762 207285
rect 146434 201627 146462 207279
rect 146804 202122 146860 202131
rect 146804 202057 146860 202066
rect 146818 201719 146846 202057
rect 146806 201713 146858 201719
rect 146806 201655 146858 201661
rect 146434 201599 146558 201627
rect 146324 185250 146380 185259
rect 146324 185185 146380 185194
rect 146230 116687 146282 116693
rect 146230 116629 146282 116635
rect 146230 115651 146282 115657
rect 146230 115593 146282 115599
rect 146242 110995 146270 115593
rect 146230 110989 146282 110995
rect 146230 110931 146282 110937
rect 146230 110841 146282 110847
rect 146230 110783 146282 110789
rect 146242 106703 146270 110783
rect 146230 106697 146282 106703
rect 146230 106639 146282 106645
rect 146230 106549 146282 106555
rect 146230 106491 146282 106497
rect 146242 92125 146270 106491
rect 146230 92119 146282 92125
rect 146230 92061 146282 92067
rect 146228 91418 146284 91427
rect 146228 91353 146284 91362
rect 146242 89313 146270 91353
rect 146230 89307 146282 89313
rect 146230 89249 146282 89255
rect 146230 83683 146282 83689
rect 146230 83625 146282 83631
rect 146242 72515 146270 83625
rect 146230 72509 146282 72515
rect 146230 72451 146282 72457
rect 146230 72361 146282 72367
rect 146230 72303 146282 72309
rect 146242 65633 146270 72303
rect 146230 65627 146282 65633
rect 146230 65569 146282 65575
rect 146228 65518 146284 65527
rect 146228 65453 146284 65462
rect 146242 64893 146270 65453
rect 146230 64887 146282 64893
rect 146230 64829 146282 64835
rect 146134 51197 146186 51203
rect 146134 51139 146186 51145
rect 146338 51055 146366 185185
rect 146420 183326 146476 183335
rect 146420 183261 146476 183270
rect 146434 51129 146462 183261
rect 146530 141113 146558 201599
rect 146708 199606 146764 199615
rect 146708 199541 146764 199550
rect 146722 198759 146750 199541
rect 146804 199014 146860 199023
rect 146804 198949 146806 198958
rect 146858 198949 146860 198958
rect 146806 198917 146858 198923
rect 146710 198753 146762 198759
rect 146710 198695 146762 198701
rect 146804 197830 146860 197839
rect 146804 197765 146860 197774
rect 146818 195873 146846 197765
rect 146806 195867 146858 195873
rect 146806 195809 146858 195815
rect 146804 193686 146860 193695
rect 146804 193621 146860 193630
rect 146818 193061 146846 193621
rect 146806 193055 146858 193061
rect 146806 192997 146858 193003
rect 146804 192946 146860 192955
rect 146804 192881 146860 192890
rect 146708 191762 146764 191771
rect 146708 191697 146764 191706
rect 146722 190249 146750 191697
rect 146710 190243 146762 190249
rect 146710 190185 146762 190191
rect 146818 190175 146846 192881
rect 146806 190169 146858 190175
rect 146806 190111 146858 190117
rect 146708 189394 146764 189403
rect 146708 189329 146764 189338
rect 146722 187363 146750 189329
rect 146804 188210 146860 188219
rect 146804 188145 146860 188154
rect 146710 187357 146762 187363
rect 146710 187299 146762 187305
rect 146818 187289 146846 188145
rect 146806 187283 146858 187289
rect 146806 187225 146858 187231
rect 146804 179774 146860 179783
rect 146804 179709 146860 179718
rect 146612 176074 146668 176083
rect 146612 176009 146668 176018
rect 146626 157023 146654 176009
rect 146818 157287 146846 179709
rect 146804 157278 146860 157287
rect 146804 157213 146860 157222
rect 146806 157165 146858 157171
rect 146806 157107 146858 157113
rect 146614 157017 146666 157023
rect 146614 156959 146666 156965
rect 146612 156834 146668 156843
rect 146612 156769 146668 156778
rect 146518 141107 146570 141113
rect 146518 141049 146570 141055
rect 146518 136667 146570 136673
rect 146518 136609 146570 136615
rect 146530 129421 146558 136609
rect 146518 129415 146570 129421
rect 146518 129357 146570 129363
rect 146516 129306 146572 129315
rect 146516 129241 146572 129250
rect 146530 126757 146558 129241
rect 146518 126751 146570 126757
rect 146518 126693 146570 126699
rect 146626 126628 146654 156769
rect 146710 140515 146762 140521
rect 146710 140457 146762 140463
rect 146722 134157 146750 140457
rect 146710 134151 146762 134157
rect 146710 134093 146762 134099
rect 146530 126600 146654 126628
rect 146530 114325 146558 126600
rect 146614 125345 146666 125351
rect 146614 125287 146666 125293
rect 146626 118025 146654 125287
rect 146614 118019 146666 118025
rect 146614 117961 146666 117967
rect 146614 116687 146666 116693
rect 146614 116629 146666 116635
rect 146518 114319 146570 114325
rect 146518 114261 146570 114267
rect 146518 114171 146570 114177
rect 146518 114113 146570 114119
rect 146530 111143 146558 114113
rect 146518 111137 146570 111143
rect 146518 111079 146570 111085
rect 146518 110989 146570 110995
rect 146518 110931 146570 110937
rect 146530 103521 146558 110931
rect 146626 103669 146654 116629
rect 146708 115394 146764 115403
rect 146708 115329 146710 115338
rect 146762 115329 146764 115338
rect 146710 115297 146762 115303
rect 146708 115246 146764 115255
rect 146708 115181 146764 115190
rect 146614 103663 146666 103669
rect 146614 103605 146666 103611
rect 146722 103540 146750 115181
rect 146518 103515 146570 103521
rect 146518 103457 146570 103463
rect 146626 103512 146750 103540
rect 146516 95562 146572 95571
rect 146516 95497 146572 95506
rect 146530 95159 146558 95497
rect 146626 95455 146654 103512
rect 146710 103441 146762 103447
rect 146710 103383 146762 103389
rect 146614 95449 146666 95455
rect 146614 95391 146666 95397
rect 146518 95153 146570 95159
rect 146518 95095 146570 95101
rect 146516 84166 146572 84175
rect 146516 84101 146572 84110
rect 146530 72367 146558 84101
rect 146518 72361 146570 72367
rect 146518 72303 146570 72309
rect 146518 72213 146570 72219
rect 146518 72155 146570 72161
rect 146530 60435 146558 72155
rect 146722 64912 146750 103383
rect 146818 72589 146846 157107
rect 147190 141033 147242 141039
rect 147190 140975 147242 140981
rect 147094 135483 147146 135489
rect 147094 135425 147146 135431
rect 146998 134151 147050 134157
rect 146998 134093 147050 134099
rect 146900 127530 146956 127539
rect 146900 127465 146956 127474
rect 146914 127053 146942 127465
rect 146902 127047 146954 127053
rect 146902 126989 146954 126995
rect 146900 126938 146956 126947
rect 146900 126873 146956 126882
rect 146914 126831 146942 126873
rect 146902 126825 146954 126831
rect 146902 126767 146954 126773
rect 146902 126677 146954 126683
rect 146902 126619 146954 126625
rect 146914 115435 146942 126619
rect 146902 115429 146954 115435
rect 146902 115371 146954 115377
rect 147010 115232 147038 134093
rect 147106 115255 147134 135425
rect 147202 126683 147230 140975
rect 148150 127047 148202 127053
rect 148150 126989 148202 126995
rect 148054 126825 148106 126831
rect 148054 126767 148106 126773
rect 147190 126677 147242 126683
rect 147190 126619 147242 126625
rect 146914 115204 147038 115232
rect 147092 115246 147148 115255
rect 146914 114917 146942 115204
rect 147092 115181 147148 115190
rect 146902 114911 146954 114917
rect 146902 114853 146954 114859
rect 146998 114319 147050 114325
rect 146998 114261 147050 114267
rect 146902 113283 146954 113289
rect 146902 113225 146954 113231
rect 146914 100709 146942 113225
rect 147010 103447 147038 114261
rect 146998 103441 147050 103447
rect 146998 103383 147050 103389
rect 146902 100703 146954 100709
rect 146902 100645 146954 100651
rect 146900 77506 146956 77515
rect 146900 77441 146956 77450
rect 146806 72583 146858 72589
rect 146806 72525 146858 72531
rect 146914 71997 146942 77441
rect 146902 71991 146954 71997
rect 146902 71933 146954 71939
rect 146722 64884 146942 64912
rect 146914 64616 146942 64884
rect 146818 64588 146942 64616
rect 146530 60407 146750 60435
rect 146518 60299 146570 60305
rect 146518 60241 146570 60247
rect 146530 59607 146558 60241
rect 146516 59598 146572 59607
rect 146516 59533 146572 59542
rect 146422 51123 146474 51129
rect 146422 51065 146474 51071
rect 146326 51049 146378 51055
rect 146326 50991 146378 50997
rect 146722 50685 146750 60407
rect 146818 57660 146846 64588
rect 146902 63407 146954 63413
rect 146902 63349 146954 63355
rect 146914 62419 146942 63349
rect 146900 62410 146956 62419
rect 146900 62345 146956 62354
rect 147958 60817 148010 60823
rect 146900 60782 146956 60791
rect 147958 60759 148010 60765
rect 146900 60717 146956 60726
rect 146914 60453 146942 60717
rect 146902 60447 146954 60453
rect 146902 60389 146954 60395
rect 146818 57632 146942 57660
rect 146914 57216 146942 57632
rect 146818 57188 146942 57216
rect 146818 50981 146846 57188
rect 146806 50975 146858 50981
rect 146806 50917 146858 50923
rect 146710 50679 146762 50685
rect 146710 50621 146762 50627
rect 146038 50309 146090 50315
rect 146038 50251 146090 50257
rect 145846 50235 145898 50241
rect 145846 50177 145898 50183
rect 145558 49865 145610 49871
rect 145558 49807 145610 49813
rect 144790 49569 144842 49575
rect 144790 49511 144842 49517
rect 147970 46171 147998 60759
rect 148066 47651 148094 126767
rect 148162 47725 148190 126989
rect 148258 60823 148286 210239
rect 148342 193055 148394 193061
rect 148342 192997 148394 193003
rect 148246 60817 148298 60823
rect 148246 60759 148298 60765
rect 148354 60731 148382 192997
rect 148438 190243 148490 190249
rect 148438 190185 148490 190191
rect 148258 60703 148382 60731
rect 148150 47719 148202 47725
rect 148150 47661 148202 47667
rect 148054 47645 148106 47651
rect 148054 47587 148106 47593
rect 148258 46393 148286 60703
rect 148450 60620 148478 190185
rect 148534 187357 148586 187363
rect 148534 187299 148586 187305
rect 148354 60592 148478 60620
rect 148354 46689 148382 60592
rect 148438 60521 148490 60527
rect 148438 60463 148490 60469
rect 148450 54163 148478 60463
rect 148438 54157 148490 54163
rect 148438 54099 148490 54105
rect 148342 46683 148394 46689
rect 148342 46625 148394 46631
rect 148546 46615 148574 187299
rect 148630 178699 148682 178705
rect 148630 178641 148682 178647
rect 148642 46763 148670 178641
rect 148726 167081 148778 167087
rect 148726 167023 148778 167029
rect 148630 46757 148682 46763
rect 148630 46699 148682 46705
rect 148534 46609 148586 46615
rect 148534 46551 148586 46557
rect 148738 46541 148766 167023
rect 148822 164195 148874 164201
rect 148822 164137 148874 164143
rect 148834 48391 148862 164137
rect 148918 161383 148970 161389
rect 148918 161325 148970 161331
rect 148822 48385 148874 48391
rect 148822 48327 148874 48333
rect 148930 46837 148958 161325
rect 149206 158497 149258 158503
rect 149206 158439 149258 158445
rect 149014 100925 149066 100931
rect 149014 100867 149066 100873
rect 149026 77769 149054 100867
rect 149014 77763 149066 77769
rect 149014 77705 149066 77711
rect 149218 47429 149246 158439
rect 149302 155611 149354 155617
rect 149302 155553 149354 155559
rect 149314 48317 149342 155553
rect 149398 149913 149450 149919
rect 149398 149855 149450 149861
rect 149302 48311 149354 48317
rect 149302 48253 149354 48259
rect 149410 48243 149438 149855
rect 149494 147027 149546 147033
rect 149494 146969 149546 146975
rect 149398 48237 149450 48243
rect 149398 48179 149450 48185
rect 149506 48169 149534 146969
rect 149590 141255 149642 141261
rect 149590 141197 149642 141203
rect 149494 48163 149546 48169
rect 149494 48105 149546 48111
rect 149602 48095 149630 141197
rect 149686 138369 149738 138375
rect 149686 138311 149738 138317
rect 149590 48089 149642 48095
rect 149590 48031 149642 48037
rect 149698 48021 149726 138311
rect 151138 100635 151166 230515
rect 152578 224289 152606 267811
rect 152566 224283 152618 224289
rect 152566 224225 152618 224231
rect 155458 221773 155486 275784
rect 155542 269941 155594 269947
rect 155542 269883 155594 269889
rect 155554 269207 155582 269883
rect 155542 269201 155594 269207
rect 155542 269143 155594 269149
rect 156226 264249 156254 275650
rect 156214 264243 156266 264249
rect 156214 264185 156266 264191
rect 157474 264175 157502 275650
rect 158626 267875 158654 275650
rect 160162 270613 160190 275784
rect 160150 270607 160202 270613
rect 160150 270549 160202 270555
rect 161026 270169 161054 275650
rect 161014 270163 161066 270169
rect 161014 270105 161066 270111
rect 162178 267875 162206 275650
rect 158614 267869 158666 267875
rect 158614 267811 158666 267817
rect 161206 267869 161258 267875
rect 161206 267811 161258 267817
rect 162166 267869 162218 267875
rect 162166 267811 162218 267817
rect 157462 264169 157514 264175
rect 157462 264111 157514 264117
rect 158422 245077 158474 245083
rect 158420 245042 158422 245051
rect 158474 245042 158476 245051
rect 158420 244977 158476 244986
rect 156886 225689 156938 225695
rect 156886 225631 156938 225637
rect 155446 221767 155498 221773
rect 155446 221709 155498 221715
rect 154006 216735 154058 216741
rect 154006 216677 154058 216683
rect 151222 184397 151274 184403
rect 151222 184339 151274 184345
rect 151126 100629 151178 100635
rect 151126 100571 151178 100577
rect 151234 91977 151262 184339
rect 151318 130155 151370 130161
rect 151318 130097 151370 130103
rect 151222 91971 151274 91977
rect 151222 91913 151274 91919
rect 151126 89455 151178 89461
rect 151126 89397 151178 89403
rect 151138 71923 151166 89397
rect 151330 83541 151358 130097
rect 154018 97527 154046 216677
rect 154102 144067 154154 144073
rect 154102 144009 154154 144015
rect 154006 97521 154058 97527
rect 154006 97463 154058 97469
rect 154006 92267 154058 92273
rect 154006 92209 154058 92215
rect 151318 83535 151370 83541
rect 151318 83477 151370 83483
rect 154018 74809 154046 92209
rect 154114 86427 154142 144009
rect 156898 97823 156926 225631
rect 161218 221699 161246 267811
rect 163426 264323 163454 275650
rect 164086 267869 164138 267875
rect 164086 267811 164138 267817
rect 163414 264317 163466 264323
rect 163414 264259 163466 264265
rect 162646 230499 162698 230505
rect 162646 230441 162698 230447
rect 161206 221693 161258 221699
rect 161206 221635 161258 221641
rect 159766 198975 159818 198981
rect 159766 198917 159818 198923
rect 156982 167155 157034 167161
rect 156982 167097 157034 167103
rect 156886 97817 156938 97823
rect 156886 97759 156938 97765
rect 156994 89239 157022 167097
rect 157078 104255 157130 104261
rect 157078 104197 157130 104203
rect 156982 89233 157034 89239
rect 156982 89175 157034 89181
rect 154102 86421 154154 86427
rect 154102 86363 154154 86369
rect 157090 77695 157118 104197
rect 159778 100561 159806 198917
rect 159862 170411 159914 170417
rect 159862 170353 159914 170359
rect 159766 100555 159818 100561
rect 159766 100497 159818 100503
rect 159874 89165 159902 170353
rect 160150 107511 160202 107517
rect 160150 107453 160202 107459
rect 159958 104403 160010 104409
rect 159958 104345 160010 104351
rect 159862 89159 159914 89165
rect 159862 89101 159914 89107
rect 157078 77689 157130 77695
rect 157078 77631 157130 77637
rect 155542 74951 155594 74957
rect 155542 74893 155594 74899
rect 154006 74803 154058 74809
rect 154006 74745 154058 74751
rect 154102 72065 154154 72071
rect 154102 72007 154154 72013
rect 151126 71917 151178 71923
rect 151126 71859 151178 71865
rect 149782 70289 149834 70295
rect 149782 70231 149834 70237
rect 149794 69037 149822 70231
rect 149782 69031 149834 69037
rect 149782 68973 149834 68979
rect 154114 68963 154142 72007
rect 154102 68957 154154 68963
rect 154102 68899 154154 68905
rect 155554 68889 155582 74893
rect 155542 68883 155594 68889
rect 155542 68825 155594 68831
rect 152662 67033 152714 67039
rect 152662 66975 152714 66981
rect 152674 66151 152702 66975
rect 158326 66589 158378 66595
rect 158326 66531 158378 66537
rect 152662 66145 152714 66151
rect 152662 66087 152714 66093
rect 158338 66077 158366 66531
rect 158326 66071 158378 66077
rect 158326 66013 158378 66019
rect 151414 62223 151466 62229
rect 151414 62165 151466 62171
rect 151426 60379 151454 62165
rect 152470 60595 152522 60601
rect 152470 60537 152522 60543
rect 151414 60373 151466 60379
rect 151414 60315 151466 60321
rect 152482 54681 152510 60537
rect 159168 55708 159422 55736
rect 152470 54675 152522 54681
rect 152470 54617 152522 54623
rect 155520 51416 155582 51444
rect 149686 48015 149738 48021
rect 149686 47957 149738 47963
rect 149206 47423 149258 47429
rect 149206 47365 149258 47371
rect 148918 46831 148970 46837
rect 148918 46773 148970 46779
rect 148726 46535 148778 46541
rect 148726 46477 148778 46483
rect 148246 46387 148298 46393
rect 148246 46329 148298 46335
rect 147958 46165 148010 46171
rect 147958 46107 148010 46113
rect 155554 44691 155582 51416
rect 159394 50833 159422 55708
rect 159970 52017 159998 104345
rect 160054 98335 160106 98341
rect 160054 98277 160106 98283
rect 160066 52165 160094 98277
rect 160162 77621 160190 107453
rect 160150 77615 160202 77621
rect 160150 77557 160202 77563
rect 160150 75025 160202 75031
rect 160150 74967 160202 74973
rect 160162 68815 160190 74967
rect 160150 68809 160202 68815
rect 160150 68751 160202 68757
rect 160054 52159 160106 52165
rect 160054 52101 160106 52107
rect 159958 52011 160010 52017
rect 159958 51953 160010 51959
rect 159382 50827 159434 50833
rect 159382 50769 159434 50775
rect 162658 47915 162686 230441
rect 164098 221625 164126 267811
rect 164578 264397 164606 275650
rect 165826 267875 165854 275650
rect 166882 269947 166910 275650
rect 168130 270391 168158 275650
rect 169296 275636 169886 275664
rect 168118 270385 168170 270391
rect 168118 270327 168170 270333
rect 166870 269941 166922 269947
rect 166870 269883 166922 269889
rect 165814 267869 165866 267875
rect 165814 267811 165866 267817
rect 166966 267869 167018 267875
rect 166966 267811 167018 267817
rect 164566 264391 164618 264397
rect 164566 264333 164618 264339
rect 165526 236271 165578 236277
rect 165526 236213 165578 236219
rect 164086 221619 164138 221625
rect 164086 221561 164138 221567
rect 162742 207485 162794 207491
rect 162742 207427 162794 207433
rect 162754 94937 162782 207427
rect 162934 132745 162986 132751
rect 162934 132687 162986 132693
rect 162838 109583 162890 109589
rect 162838 109525 162890 109531
rect 162742 94931 162794 94937
rect 162742 94873 162794 94879
rect 162742 86495 162794 86501
rect 162742 86437 162794 86443
rect 162754 51943 162782 86437
rect 162850 52461 162878 109525
rect 162946 83467 162974 132687
rect 163126 89381 163178 89387
rect 163126 89323 163178 89329
rect 162934 83461 162986 83467
rect 162934 83403 162986 83409
rect 163030 80797 163082 80803
rect 163030 80739 163082 80745
rect 162838 52455 162890 52461
rect 162838 52397 162890 52403
rect 163042 52091 163070 80739
rect 163138 71849 163166 89323
rect 163126 71843 163178 71849
rect 163126 71785 163178 71791
rect 164182 60669 164234 60675
rect 164182 60611 164234 60617
rect 164194 57493 164222 60611
rect 164182 57487 164234 57493
rect 164182 57429 164234 57435
rect 163030 52085 163082 52091
rect 163030 52027 163082 52033
rect 162742 51937 162794 51943
rect 162742 51879 162794 51885
rect 162644 47906 162700 47915
rect 162644 47841 162700 47850
rect 165538 47619 165566 236213
rect 166868 230094 166924 230103
rect 166868 230029 166870 230038
rect 166922 230029 166924 230038
rect 166870 229997 166922 230003
rect 166978 221551 167006 267811
rect 168310 264983 168362 264989
rect 168310 264925 168362 264931
rect 168406 264983 168458 264989
rect 168406 264925 168458 264931
rect 168322 264712 168350 264925
rect 168418 264841 168446 264925
rect 168406 264835 168458 264841
rect 168406 264777 168458 264783
rect 168502 264835 168554 264841
rect 168502 264777 168554 264783
rect 168514 264712 168542 264777
rect 168322 264684 168542 264712
rect 168502 245077 168554 245083
rect 168502 245019 168554 245025
rect 168514 244903 168542 245019
rect 168500 244894 168556 244903
rect 168500 244829 168556 244838
rect 168406 236197 168458 236203
rect 168406 236139 168458 236145
rect 166966 221545 167018 221551
rect 166966 221487 167018 221493
rect 165622 207411 165674 207417
rect 165622 207353 165674 207359
rect 165634 94863 165662 207353
rect 165718 138295 165770 138301
rect 165718 138237 165770 138243
rect 165622 94857 165674 94863
rect 165622 94799 165674 94805
rect 165730 83393 165758 138237
rect 165814 89307 165866 89313
rect 165814 89249 165866 89255
rect 165718 83387 165770 83393
rect 165718 83329 165770 83335
rect 165622 77911 165674 77917
rect 165622 77853 165674 77859
rect 165634 52609 165662 77853
rect 165826 71775 165854 89249
rect 165814 71769 165866 71775
rect 165814 71711 165866 71717
rect 167062 60743 167114 60749
rect 167062 60685 167114 60691
rect 167074 57567 167102 60685
rect 167062 57561 167114 57567
rect 167062 57503 167114 57509
rect 165622 52603 165674 52609
rect 165622 52545 165674 52551
rect 168418 48655 168446 236139
rect 169858 221477 169886 275636
rect 170530 264471 170558 275650
rect 171682 264545 171710 275650
rect 172930 270539 172958 275650
rect 172918 270533 172970 270539
rect 172918 270475 172970 270481
rect 174082 270465 174110 275650
rect 174070 270459 174122 270465
rect 174070 270401 174122 270407
rect 175522 268837 175550 275784
rect 176482 270613 176510 275650
rect 176470 270607 176522 270613
rect 176470 270549 176522 270555
rect 175606 270533 175658 270539
rect 175606 270475 175658 270481
rect 175510 268831 175562 268837
rect 175510 268773 175562 268779
rect 171670 264539 171722 264545
rect 171670 264481 171722 264487
rect 170518 264465 170570 264471
rect 170518 264407 170570 264413
rect 174166 239083 174218 239089
rect 174166 239025 174218 239031
rect 171286 233311 171338 233317
rect 171286 233253 171338 233259
rect 169846 221471 169898 221477
rect 169846 221413 169898 221419
rect 168502 213257 168554 213263
rect 168502 213199 168554 213205
rect 168514 97749 168542 213199
rect 168598 141181 168650 141187
rect 168598 141123 168650 141129
rect 168502 97743 168554 97749
rect 168502 97685 168554 97691
rect 168502 92193 168554 92199
rect 168502 92135 168554 92141
rect 168514 71701 168542 92135
rect 168610 83319 168638 141123
rect 168598 83313 168650 83319
rect 168598 83255 168650 83261
rect 168502 71695 168554 71701
rect 168502 71637 168554 71643
rect 169942 60817 169994 60823
rect 169942 60759 169994 60765
rect 169954 60305 169982 60759
rect 169942 60299 169994 60305
rect 169942 60241 169994 60247
rect 168404 48646 168460 48655
rect 168404 48581 168460 48590
rect 171298 48507 171326 233253
rect 172726 230203 172778 230209
rect 172726 230145 172778 230151
rect 172738 230061 172766 230145
rect 172726 230055 172778 230061
rect 172726 229997 172778 230003
rect 171382 213183 171434 213189
rect 171382 213125 171434 213131
rect 171394 97675 171422 213125
rect 171478 146953 171530 146959
rect 171478 146895 171530 146901
rect 171382 97669 171434 97675
rect 171382 97611 171434 97617
rect 171490 86353 171518 146895
rect 171574 95153 171626 95159
rect 171574 95095 171626 95101
rect 171478 86347 171530 86353
rect 171478 86289 171530 86295
rect 171586 74735 171614 95095
rect 171574 74729 171626 74735
rect 171574 74671 171626 74677
rect 171284 48498 171340 48507
rect 171284 48433 171340 48442
rect 174178 48359 174206 239025
rect 174262 218955 174314 218961
rect 174262 218897 174314 218903
rect 174274 97601 174302 218897
rect 175618 218813 175646 270475
rect 177634 264619 177662 275650
rect 178486 270607 178538 270613
rect 178486 270549 178538 270555
rect 177622 264613 177674 264619
rect 177622 264555 177674 264561
rect 177046 221915 177098 221921
rect 177046 221857 177098 221863
rect 175606 218807 175658 218813
rect 175606 218749 175658 218755
rect 174358 149839 174410 149845
rect 174358 149781 174410 149787
rect 174262 97595 174314 97601
rect 174262 97537 174314 97543
rect 174370 86279 174398 149781
rect 174454 95079 174506 95085
rect 174454 95021 174506 95027
rect 174358 86273 174410 86279
rect 174358 86215 174410 86221
rect 174466 74661 174494 95021
rect 174454 74655 174506 74661
rect 174454 74597 174506 74603
rect 174164 48350 174220 48359
rect 174164 48285 174220 48294
rect 177058 47651 177086 221857
rect 178498 218739 178526 270549
rect 178882 264693 178910 275650
rect 180034 270613 180062 275650
rect 180022 270607 180074 270613
rect 180022 270549 180074 270555
rect 181282 269133 181310 275650
rect 182448 275636 182750 275664
rect 183600 275636 184286 275664
rect 181366 275047 181418 275053
rect 181366 274989 181418 274995
rect 181378 270780 181406 274989
rect 181378 270752 181502 270780
rect 181366 270607 181418 270613
rect 181366 270549 181418 270555
rect 181270 269127 181322 269133
rect 181270 269069 181322 269075
rect 178870 264687 178922 264693
rect 178870 264629 178922 264635
rect 178582 230277 178634 230283
rect 178582 230219 178634 230225
rect 178594 230191 178622 230219
rect 178678 230203 178730 230209
rect 178594 230163 178678 230191
rect 178678 230145 178730 230151
rect 179926 224727 179978 224733
rect 179926 224669 179978 224675
rect 178486 218733 178538 218739
rect 178486 218675 178538 218681
rect 177142 152799 177194 152805
rect 177142 152741 177194 152747
rect 177154 86205 177182 152741
rect 177238 98039 177290 98045
rect 177238 97981 177290 97987
rect 177142 86199 177194 86205
rect 177142 86141 177194 86147
rect 177250 74587 177278 97981
rect 177238 74581 177290 74587
rect 177238 74523 177290 74529
rect 177046 47645 177098 47651
rect 165524 47610 165580 47619
rect 177046 47587 177098 47593
rect 165524 47545 165580 47554
rect 179938 46467 179966 224669
rect 181378 218665 181406 270549
rect 181474 267801 181502 270752
rect 182422 270459 182474 270465
rect 182422 270401 182474 270407
rect 182434 269947 182462 270401
rect 182422 269941 182474 269947
rect 182422 269883 182474 269889
rect 182518 269941 182570 269947
rect 182518 269883 182570 269889
rect 182530 269207 182558 269883
rect 182722 269207 182750 275636
rect 182518 269201 182570 269207
rect 182518 269143 182570 269149
rect 182710 269201 182762 269207
rect 182710 269143 182762 269149
rect 181462 267795 181514 267801
rect 181462 267737 181514 267743
rect 181462 265131 181514 265137
rect 181462 265073 181514 265079
rect 181474 264841 181502 265073
rect 181462 264835 181514 264841
rect 181462 264777 181514 264783
rect 181366 218659 181418 218665
rect 181366 218601 181418 218607
rect 184258 218591 184286 275636
rect 184738 268985 184766 275650
rect 185986 269059 186014 275650
rect 187030 270533 187082 270539
rect 187030 270475 187082 270481
rect 185974 269053 186026 269059
rect 185974 268995 186026 269001
rect 184726 268979 184778 268985
rect 184726 268921 184778 268927
rect 187042 268837 187070 270475
rect 187030 268831 187082 268837
rect 187030 268773 187082 268779
rect 184246 218585 184298 218591
rect 184246 218527 184298 218533
rect 187138 215705 187166 275650
rect 188386 264767 188414 275650
rect 189538 266987 189566 275650
rect 191074 267875 191102 275784
rect 191062 267869 191114 267875
rect 191062 267811 191114 267817
rect 191254 267795 191306 267801
rect 191254 267737 191306 267743
rect 189526 266981 189578 266987
rect 189526 266923 189578 266929
rect 188374 264761 188426 264767
rect 188374 264703 188426 264709
rect 191266 263435 191294 267737
rect 191938 267061 191966 275650
rect 192886 267869 192938 267875
rect 192886 267811 192938 267817
rect 191926 267055 191978 267061
rect 191926 266997 191978 267003
rect 191542 265131 191594 265137
rect 191542 265073 191594 265079
rect 191554 264915 191582 265073
rect 191542 264909 191594 264915
rect 191542 264851 191594 264857
rect 191254 263429 191306 263435
rect 191254 263371 191306 263377
rect 188566 227761 188618 227767
rect 188566 227703 188618 227709
rect 187126 215699 187178 215705
rect 187126 215641 187178 215647
rect 185686 201713 185738 201719
rect 185686 201655 185738 201661
rect 182806 195867 182858 195873
rect 182806 195809 182858 195815
rect 180022 152725 180074 152731
rect 180022 152667 180074 152673
rect 180034 86131 180062 152667
rect 180118 97965 180170 97971
rect 180118 97907 180170 97913
rect 180022 86125 180074 86131
rect 180022 86067 180074 86073
rect 180130 74513 180158 97907
rect 180118 74507 180170 74513
rect 180118 74449 180170 74455
rect 182818 48465 182846 195809
rect 182902 172853 182954 172859
rect 182902 172795 182954 172801
rect 182914 89091 182942 172795
rect 182998 109509 183050 109515
rect 182998 109451 183050 109457
rect 182902 89085 182954 89091
rect 182902 89027 182954 89033
rect 183010 77547 183038 109451
rect 185698 100487 185726 201655
rect 185782 181511 185834 181517
rect 185782 181453 185834 181459
rect 185686 100481 185738 100487
rect 185686 100423 185738 100429
rect 185794 91903 185822 181453
rect 185878 118315 185930 118321
rect 185878 118257 185930 118263
rect 185782 91897 185834 91903
rect 185782 91839 185834 91845
rect 185890 80655 185918 118257
rect 185878 80649 185930 80655
rect 185878 80591 185930 80597
rect 185686 77837 185738 77843
rect 185686 77779 185738 77785
rect 182998 77541 183050 77547
rect 182998 77483 183050 77489
rect 185698 77473 185726 77779
rect 185686 77467 185738 77473
rect 185686 77409 185738 77415
rect 182806 48459 182858 48465
rect 182806 48401 182858 48407
rect 188578 48211 188606 227703
rect 192898 215631 192926 267811
rect 193090 266469 193118 275650
rect 193078 266463 193130 266469
rect 193078 266405 193130 266411
rect 194338 266321 194366 275650
rect 194326 266315 194378 266321
rect 194326 266257 194378 266263
rect 195490 263509 195518 275650
rect 195874 270613 196094 270632
rect 195862 270607 196094 270613
rect 195914 270604 196094 270607
rect 195862 270549 195914 270555
rect 195874 270465 195998 270484
rect 196066 270465 196094 270604
rect 195862 270459 195998 270465
rect 195914 270456 195998 270459
rect 195862 270401 195914 270407
rect 195970 270317 195998 270456
rect 196054 270459 196106 270465
rect 196054 270401 196106 270407
rect 195862 270311 195914 270317
rect 195862 270253 195914 270259
rect 195958 270311 196010 270317
rect 195958 270253 196010 270259
rect 195874 270188 195902 270253
rect 195874 270160 195998 270188
rect 195970 269947 195998 270160
rect 195862 269941 195914 269947
rect 195862 269883 195914 269889
rect 195958 269941 196010 269947
rect 195958 269883 196010 269889
rect 195874 268837 195902 269883
rect 195862 268831 195914 268837
rect 195862 268773 195914 268779
rect 196738 266617 196766 275650
rect 196726 266611 196778 266617
rect 196726 266553 196778 266559
rect 197890 266543 197918 275650
rect 197878 266537 197930 266543
rect 197878 266479 197930 266485
rect 195478 263503 195530 263509
rect 195478 263445 195530 263451
rect 198742 263429 198794 263435
rect 198742 263371 198794 263377
rect 198754 250633 198782 263371
rect 199138 263361 199166 275650
rect 200194 266765 200222 275650
rect 200182 266759 200234 266765
rect 200182 266701 200234 266707
rect 201442 266691 201470 275650
rect 201430 266685 201482 266691
rect 201430 266627 201482 266633
rect 202594 264989 202622 275650
rect 203842 266913 203870 275650
rect 203830 266907 203882 266913
rect 203830 266849 203882 266855
rect 204994 266839 205022 275650
rect 206530 270613 206558 275784
rect 221506 275784 221616 275812
rect 237168 275784 237470 275812
rect 206518 270607 206570 270613
rect 206518 270549 206570 270555
rect 207394 267283 207422 275650
rect 207382 267277 207434 267283
rect 207382 267219 207434 267225
rect 204982 266833 205034 266839
rect 204982 266775 205034 266781
rect 208546 266247 208574 275650
rect 209794 269947 209822 275650
rect 209686 269941 209738 269947
rect 209686 269883 209738 269889
rect 209782 269941 209834 269947
rect 209782 269883 209834 269889
rect 209698 268319 209726 269883
rect 209686 268313 209738 268319
rect 209686 268255 209738 268261
rect 210946 267653 210974 275650
rect 212194 268689 212222 275650
rect 213346 270317 213374 275650
rect 213238 270311 213290 270317
rect 213238 270253 213290 270259
rect 213334 270311 213386 270317
rect 213334 270253 213386 270259
rect 213250 268763 213278 270253
rect 213238 268757 213290 268763
rect 213238 268699 213290 268705
rect 212182 268683 212234 268689
rect 212182 268625 212234 268631
rect 210934 267647 210986 267653
rect 210934 267589 210986 267595
rect 208534 266241 208586 266247
rect 208534 266183 208586 266189
rect 214594 265655 214622 275650
rect 215746 267135 215774 275650
rect 216790 270755 216842 270761
rect 216790 270697 216842 270703
rect 216802 270539 216830 270697
rect 216898 270539 216926 275650
rect 217462 270607 217514 270613
rect 217462 270549 217514 270555
rect 216790 270533 216842 270539
rect 216790 270475 216842 270481
rect 216886 270533 216938 270539
rect 216886 270475 216938 270481
rect 217474 268615 217502 270549
rect 217462 268609 217514 268615
rect 217462 268551 217514 268557
rect 215734 267129 215786 267135
rect 215734 267071 215786 267077
rect 217654 267055 217706 267061
rect 217654 266997 217706 267003
rect 214582 265649 214634 265655
rect 214582 265591 214634 265597
rect 202582 264983 202634 264989
rect 202582 264925 202634 264931
rect 216694 264909 216746 264915
rect 216694 264851 216746 264857
rect 216022 264835 216074 264841
rect 216022 264777 216074 264783
rect 199126 263355 199178 263361
rect 199126 263297 199178 263303
rect 216034 258630 216062 264777
rect 216596 263542 216652 263551
rect 216596 263477 216652 263486
rect 216610 258644 216638 263477
rect 216384 258616 216638 258644
rect 216706 258644 216734 264851
rect 216706 258616 216864 258644
rect 217666 258630 217694 266997
rect 218050 265951 218078 275650
rect 219298 268837 219326 275650
rect 220464 275636 220958 275664
rect 220630 270681 220682 270687
rect 220726 270681 220778 270687
rect 220682 270629 220726 270632
rect 220630 270623 220778 270629
rect 220642 270604 220766 270623
rect 220534 270533 220586 270539
rect 220534 270475 220586 270481
rect 220342 270311 220394 270317
rect 220342 270253 220394 270259
rect 219862 269941 219914 269947
rect 219862 269883 219914 269889
rect 219958 269941 220010 269947
rect 219958 269883 220010 269889
rect 218806 268831 218858 268837
rect 218806 268773 218858 268779
rect 219286 268831 219338 268837
rect 219286 268773 219338 268779
rect 218818 268467 218846 268773
rect 219382 268609 219434 268615
rect 219382 268551 219434 268557
rect 218806 268461 218858 268467
rect 218806 268403 218858 268409
rect 218038 265945 218090 265951
rect 218038 265887 218090 265893
rect 218902 264983 218954 264989
rect 218902 264925 218954 264931
rect 218134 263503 218186 263509
rect 218134 263445 218186 263451
rect 218146 258630 218174 263445
rect 218326 263355 218378 263361
rect 218326 263297 218378 263303
rect 218338 258644 218366 263297
rect 218914 258644 218942 264925
rect 218338 258616 218592 258644
rect 218914 258616 219072 258644
rect 219394 258630 219422 268551
rect 219874 258630 219902 269883
rect 219970 268763 219998 269883
rect 219958 268757 220010 268763
rect 219958 268699 220010 268705
rect 220354 258630 220382 270253
rect 220546 258644 220574 270475
rect 220930 258644 220958 275636
rect 221506 265803 221534 275784
rect 222550 267943 222602 267949
rect 222550 267885 222602 267891
rect 222070 267869 222122 267875
rect 222070 267811 222122 267817
rect 221494 265797 221546 265803
rect 221494 265739 221546 265745
rect 221590 262171 221642 262177
rect 221590 262113 221642 262119
rect 220546 258616 220800 258644
rect 220930 258616 221184 258644
rect 221602 258630 221630 262113
rect 222082 258630 222110 267811
rect 222562 258630 222590 267885
rect 222850 267061 222878 275650
rect 223606 268535 223658 268541
rect 223606 268477 223658 268483
rect 222838 267055 222890 267061
rect 222838 266997 222890 267003
rect 223030 266981 223082 266987
rect 223030 266923 223082 266929
rect 223042 264915 223070 266923
rect 223030 264909 223082 264915
rect 223030 264851 223082 264857
rect 223126 263059 223178 263065
rect 223126 263001 223178 263007
rect 223138 258644 223166 263001
rect 223618 258644 223646 268477
rect 223798 263503 223850 263509
rect 223798 263445 223850 263451
rect 222912 258616 223166 258644
rect 223392 258616 223646 258644
rect 223810 258630 223838 263445
rect 224002 262177 224030 275650
rect 224182 268387 224234 268393
rect 224182 268329 224234 268335
rect 223990 262171 224042 262177
rect 223990 262113 224042 262119
rect 224194 258630 224222 268329
rect 225250 265729 225278 275650
rect 226402 268763 226430 275650
rect 227446 271717 227498 271723
rect 227446 271659 227498 271665
rect 226390 268757 226442 268763
rect 226390 268699 226442 268705
rect 225334 267203 225386 267209
rect 225334 267145 225386 267151
rect 225238 265723 225290 265729
rect 225238 265665 225290 265671
rect 224662 263429 224714 263435
rect 224662 263371 224714 263377
rect 224674 258630 224702 263371
rect 225346 258644 225374 267145
rect 225814 261061 225866 261067
rect 225814 261003 225866 261009
rect 225826 258644 225854 261003
rect 225910 260987 225962 260993
rect 225910 260929 225962 260935
rect 225120 258616 225374 258644
rect 225600 258616 225854 258644
rect 225922 258630 225950 260929
rect 226390 260765 226442 260771
rect 226390 260707 226442 260713
rect 226402 258630 226430 260707
rect 226870 260321 226922 260327
rect 226870 260263 226922 260269
rect 226882 258630 226910 260263
rect 227458 258644 227486 271659
rect 227650 267875 227678 275650
rect 228118 272087 228170 272093
rect 228118 272029 228170 272035
rect 227926 271939 227978 271945
rect 227926 271881 227978 271887
rect 227638 267869 227690 267875
rect 227638 267811 227690 267817
rect 227638 264835 227690 264841
rect 227638 264777 227690 264783
rect 227650 263435 227678 264777
rect 227638 263429 227690 263435
rect 227638 263371 227690 263377
rect 227938 258644 227966 271881
rect 227328 258616 227486 258644
rect 227712 258616 227966 258644
rect 228130 258630 228158 272029
rect 228802 265581 228830 275650
rect 229078 272827 229130 272833
rect 229078 272769 229130 272775
rect 228886 270755 228938 270761
rect 228886 270697 228938 270703
rect 228898 270539 228926 270697
rect 228886 270533 228938 270539
rect 228886 270475 228938 270481
rect 228790 265575 228842 265581
rect 228790 265517 228842 265523
rect 228598 260469 228650 260475
rect 228598 260411 228650 260417
rect 228610 258630 228638 260411
rect 229090 258630 229118 272769
rect 230050 270761 230078 275650
rect 230134 272753 230186 272759
rect 230134 272695 230186 272701
rect 230038 270755 230090 270761
rect 230038 270697 230090 270703
rect 229654 261357 229706 261363
rect 229654 261299 229706 261305
rect 229666 258644 229694 261299
rect 230146 258644 230174 272695
rect 230806 272679 230858 272685
rect 230806 272621 230858 272627
rect 230326 261283 230378 261289
rect 230326 261225 230378 261231
rect 229440 258616 229694 258644
rect 229920 258616 230174 258644
rect 230338 258630 230366 261225
rect 230818 258630 230846 272621
rect 231202 267949 231230 275650
rect 231862 272605 231914 272611
rect 231862 272547 231914 272553
rect 231190 267943 231242 267949
rect 231190 267885 231242 267891
rect 231190 261209 231242 261215
rect 231190 261151 231242 261157
rect 231202 258630 231230 261151
rect 231874 258644 231902 272547
rect 232450 265507 232478 275650
rect 232726 272457 232778 272463
rect 232726 272399 232778 272405
rect 232438 265501 232490 265507
rect 232438 265443 232490 265449
rect 232342 261135 232394 261141
rect 232342 261077 232394 261083
rect 232354 258644 232382 261077
rect 232738 258644 232766 272399
rect 233398 272383 233450 272389
rect 233398 272325 233450 272331
rect 232918 260913 232970 260919
rect 232918 260855 232970 260861
rect 231648 258616 231902 258644
rect 232128 258616 232382 258644
rect 232512 258616 232766 258644
rect 232930 258630 232958 260855
rect 233410 258630 233438 272325
rect 233506 259957 233534 275650
rect 234454 272309 234506 272315
rect 234454 272251 234506 272257
rect 234070 260839 234122 260845
rect 234070 260781 234122 260787
rect 233494 259951 233546 259957
rect 233494 259893 233546 259899
rect 234082 258644 234110 260781
rect 234466 258644 234494 272251
rect 234754 263065 234782 275650
rect 235126 271421 235178 271427
rect 235126 271363 235178 271369
rect 234742 263059 234794 263065
rect 234742 263001 234794 263007
rect 234934 260691 234986 260697
rect 234934 260633 234986 260639
rect 234946 258644 234974 260633
rect 233856 258616 234110 258644
rect 234240 258616 234494 258644
rect 234720 258616 234974 258644
rect 235138 258630 235166 271363
rect 235906 265359 235934 275650
rect 237142 271791 237194 271797
rect 237142 271733 237194 271739
rect 235990 271569 236042 271575
rect 235990 271511 236042 271517
rect 235894 265353 235946 265359
rect 235894 265295 235946 265301
rect 235606 260025 235658 260031
rect 235606 259967 235658 259973
rect 235618 258630 235646 259967
rect 236002 258630 236030 271511
rect 236086 270459 236138 270465
rect 236086 270401 236138 270407
rect 236098 269947 236126 270401
rect 236086 269941 236138 269947
rect 236086 269883 236138 269889
rect 236662 260173 236714 260179
rect 236662 260115 236714 260121
rect 236674 258644 236702 260115
rect 237154 258644 237182 271733
rect 237442 271279 237470 275784
rect 252226 275784 252528 275812
rect 265776 275784 266078 275812
rect 268080 275784 268382 275812
rect 237718 271865 237770 271871
rect 237718 271807 237770 271813
rect 237430 271273 237482 271279
rect 237430 271215 237482 271221
rect 237622 270311 237674 270317
rect 237622 270253 237674 270259
rect 237526 269941 237578 269947
rect 237526 269883 237578 269889
rect 237538 268467 237566 269883
rect 237526 268461 237578 268467
rect 237526 268403 237578 268409
rect 237634 268319 237662 270253
rect 237622 268313 237674 268319
rect 237622 268255 237674 268261
rect 237334 260247 237386 260253
rect 237334 260189 237386 260195
rect 236448 258616 236702 258644
rect 236928 258616 237182 258644
rect 237346 258630 237374 260189
rect 237730 258630 237758 271807
rect 238306 268541 238334 275650
rect 238870 272013 238922 272019
rect 238870 271955 238922 271961
rect 238294 268535 238346 268541
rect 238294 268477 238346 268483
rect 238198 260395 238250 260401
rect 238198 260337 238250 260343
rect 238210 258630 238238 260337
rect 238882 258644 238910 271955
rect 239458 265285 239486 275650
rect 239734 273567 239786 273573
rect 239734 273509 239786 273515
rect 239446 265279 239498 265285
rect 239446 265221 239498 265227
rect 239350 260543 239402 260549
rect 239350 260485 239402 260491
rect 239362 258644 239390 260485
rect 239746 258644 239774 273509
rect 240406 273493 240458 273499
rect 240406 273435 240458 273441
rect 239926 261505 239978 261511
rect 239926 261447 239978 261453
rect 238656 258616 238910 258644
rect 239136 258616 239390 258644
rect 239472 258616 239774 258644
rect 239938 258630 239966 261447
rect 240418 258630 240446 273435
rect 240706 268541 240734 275650
rect 241462 273419 241514 273425
rect 241462 273361 241514 273367
rect 240694 268535 240746 268541
rect 240694 268477 240746 268483
rect 240982 260617 241034 260623
rect 240982 260559 241034 260565
rect 240994 258644 241022 260559
rect 241474 258644 241502 273361
rect 241858 263509 241886 275650
rect 242134 273345 242186 273351
rect 242134 273287 242186 273293
rect 241846 263503 241898 263509
rect 241846 263445 241898 263451
rect 241654 259285 241706 259291
rect 241654 259227 241706 259233
rect 240768 258616 241022 258644
rect 241248 258616 241502 258644
rect 241666 258630 241694 259227
rect 242146 258630 242174 273287
rect 243106 265433 243134 275650
rect 243190 273271 243242 273277
rect 243190 273213 243242 273219
rect 243094 265427 243146 265433
rect 243094 265369 243146 265375
rect 242518 259359 242570 259365
rect 242518 259301 242570 259307
rect 242530 258630 242558 259301
rect 243202 258644 243230 273213
rect 243862 273197 243914 273203
rect 243862 273139 243914 273145
rect 243670 261875 243722 261881
rect 243670 261817 243722 261823
rect 243682 258644 243710 261817
rect 242976 258616 243230 258644
rect 243456 258616 243710 258644
rect 243874 258630 243902 273139
rect 244258 262029 244286 275650
rect 244726 273123 244778 273129
rect 244726 273065 244778 273071
rect 244246 262023 244298 262029
rect 244246 261965 244298 261971
rect 244246 261801 244298 261807
rect 244246 261743 244298 261749
rect 244258 258630 244286 261743
rect 244738 258630 244766 273065
rect 245506 268393 245534 275650
rect 245878 273049 245930 273055
rect 245878 272991 245930 272997
rect 245494 268387 245546 268393
rect 245494 268329 245546 268335
rect 245398 261727 245450 261733
rect 245398 261669 245450 261675
rect 245410 258644 245438 261669
rect 245890 258644 245918 272991
rect 246454 272975 246506 272981
rect 246454 272917 246506 272923
rect 245974 261653 246026 261659
rect 245974 261595 246026 261601
rect 245184 258616 245438 258644
rect 245664 258616 245918 258644
rect 245986 258630 246014 261595
rect 246466 258630 246494 272917
rect 246658 265211 246686 275650
rect 247606 272901 247658 272907
rect 247606 272843 247658 272849
rect 246646 265205 246698 265211
rect 246646 265147 246698 265153
rect 246934 261579 246986 261585
rect 246934 261521 246986 261527
rect 246946 258630 246974 261521
rect 247618 258644 247646 272843
rect 247906 270909 247934 275650
rect 247894 270903 247946 270909
rect 247894 270845 247946 270851
rect 247702 268609 247754 268615
rect 247702 268551 247754 268557
rect 247714 267209 247742 268551
rect 247702 267203 247754 267209
rect 247702 267145 247754 267151
rect 249058 264841 249086 275650
rect 250006 266463 250058 266469
rect 250006 266405 250058 266411
rect 250102 266463 250154 266469
rect 250102 266405 250154 266411
rect 250018 266247 250046 266405
rect 250006 266241 250058 266247
rect 250006 266183 250058 266189
rect 249334 266019 249386 266025
rect 249334 265961 249386 265967
rect 249046 264835 249098 264841
rect 249046 264777 249098 264783
rect 248182 262911 248234 262917
rect 248182 262853 248234 262859
rect 247990 262171 248042 262177
rect 247990 262113 248042 262119
rect 248002 258644 248030 262113
rect 247392 258616 247646 258644
rect 247776 258616 248030 258644
rect 248194 258630 248222 262853
rect 248662 262837 248714 262843
rect 248662 262779 248714 262785
rect 248674 258630 248702 262779
rect 249346 258644 249374 265961
rect 249718 265871 249770 265877
rect 249718 265813 249770 265819
rect 249730 258644 249758 265813
rect 250114 258644 250142 266405
rect 250210 265137 250238 275650
rect 250486 267795 250538 267801
rect 250486 267737 250538 267743
rect 250198 265131 250250 265137
rect 250198 265073 250250 265079
rect 250390 264835 250442 264841
rect 250390 264777 250442 264783
rect 250402 262177 250430 264777
rect 250390 262171 250442 262177
rect 250390 262113 250442 262119
rect 250498 258644 250526 267737
rect 250774 267721 250826 267727
rect 250774 267663 250826 267669
rect 249072 258616 249374 258644
rect 249504 258616 249758 258644
rect 249984 258616 250142 258644
rect 250416 258616 250526 258644
rect 250786 258630 250814 267663
rect 251254 267573 251306 267579
rect 251254 267515 251306 267521
rect 251266 258630 251294 267515
rect 251362 262103 251390 275650
rect 252226 268615 252254 275784
rect 253776 275636 254078 275664
rect 252214 268609 252266 268615
rect 252214 268551 252266 268557
rect 251926 267499 251978 267505
rect 251926 267441 251978 267447
rect 251350 262097 251402 262103
rect 251350 262039 251402 262045
rect 251938 258644 251966 267441
rect 252406 267425 252458 267431
rect 252406 267367 252458 267373
rect 252020 266946 252076 266955
rect 252020 266881 252022 266890
rect 252074 266881 252076 266890
rect 252022 266849 252074 266855
rect 252418 258644 252446 267367
rect 252982 267203 253034 267209
rect 252982 267145 253034 267151
rect 252502 263281 252554 263287
rect 252502 263223 252554 263229
rect 251712 258616 251966 258644
rect 252192 258616 252446 258644
rect 252514 258630 252542 263223
rect 252994 258630 253022 267145
rect 253654 267129 253706 267135
rect 253654 267071 253706 267077
rect 253750 267129 253802 267135
rect 253750 267071 253802 267077
rect 253366 267055 253418 267061
rect 253366 266997 253418 267003
rect 253378 264989 253406 266997
rect 253366 264983 253418 264989
rect 253366 264925 253418 264931
rect 253666 263435 253694 267071
rect 253654 263429 253706 263435
rect 253654 263371 253706 263377
rect 253762 258644 253790 267071
rect 253846 266685 253898 266691
rect 253846 266627 253898 266633
rect 253858 263139 253886 266627
rect 254050 265063 254078 275636
rect 254134 267055 254186 267061
rect 254134 266997 254186 267003
rect 254038 265057 254090 265063
rect 254038 264999 254090 265005
rect 253846 263133 253898 263139
rect 253846 263075 253898 263081
rect 254146 258644 254174 266997
rect 254518 266981 254570 266987
rect 254518 266923 254570 266929
rect 254422 266389 254474 266395
rect 254422 266331 254474 266337
rect 254434 263213 254462 266331
rect 254422 263207 254474 263213
rect 254422 263149 254474 263155
rect 254530 258644 254558 266923
rect 254710 266685 254762 266691
rect 254710 266627 254762 266633
rect 253488 258616 253790 258644
rect 253920 258616 254174 258644
rect 254304 258616 254558 258644
rect 254722 258630 254750 266627
rect 254914 266099 254942 275650
rect 255874 275636 256176 275664
rect 257328 275636 257630 275664
rect 255766 266537 255818 266543
rect 255766 266479 255818 266485
rect 255190 266463 255242 266469
rect 255190 266405 255242 266411
rect 254902 266093 254954 266099
rect 254902 266035 254954 266041
rect 255202 258630 255230 266405
rect 255668 266058 255724 266067
rect 255668 265993 255724 266002
rect 255682 258630 255710 265993
rect 255778 263361 255806 266479
rect 255766 263355 255818 263361
rect 255766 263297 255818 263303
rect 255874 261067 255902 275636
rect 256148 267834 256204 267843
rect 257602 267820 257630 275636
rect 258562 267875 258590 275650
rect 259222 268905 259274 268911
rect 259222 268847 259274 268853
rect 259234 268245 259262 268847
rect 259222 268239 259274 268245
rect 259222 268181 259274 268187
rect 258550 267869 258602 267875
rect 257602 267792 257726 267820
rect 258550 267811 258602 267817
rect 256148 267769 256204 267778
rect 255862 261061 255914 261067
rect 255862 261003 255914 261009
rect 256162 258644 256190 267769
rect 256916 267390 256972 267399
rect 256916 267325 256972 267334
rect 256532 266946 256588 266955
rect 256532 266881 256534 266890
rect 256586 266881 256588 266890
rect 256534 266849 256586 266855
rect 256246 266833 256298 266839
rect 256246 266775 256298 266781
rect 256258 262177 256286 266775
rect 256724 266206 256780 266215
rect 256724 266141 256780 266150
rect 256342 266093 256394 266099
rect 256342 266035 256394 266041
rect 256438 266093 256490 266099
rect 256438 266035 256490 266041
rect 256354 263509 256382 266035
rect 256450 265877 256478 266035
rect 256438 265871 256490 265877
rect 256438 265813 256490 265819
rect 256342 263503 256394 263509
rect 256342 263445 256394 263451
rect 256246 262171 256298 262177
rect 256246 262113 256298 262119
rect 256738 258644 256766 266141
rect 256032 258616 256190 258644
rect 256512 258616 256766 258644
rect 256930 258630 256958 267325
rect 257300 267242 257356 267251
rect 257300 267177 257356 267186
rect 257314 258630 257342 267177
rect 257494 266167 257546 266173
rect 257494 266109 257546 266115
rect 257590 266167 257642 266173
rect 257590 266109 257642 266115
rect 257506 263065 257534 266109
rect 257602 265433 257630 266109
rect 257590 265427 257642 265433
rect 257590 265369 257642 265375
rect 257494 263059 257546 263065
rect 257494 263001 257546 263007
rect 257698 262769 257726 267792
rect 259126 267795 259178 267801
rect 259126 267737 259178 267743
rect 258838 267721 258890 267727
rect 258838 267663 258890 267669
rect 258850 267579 258878 267663
rect 258838 267573 258890 267579
rect 258838 267515 258890 267521
rect 258358 267277 258410 267283
rect 258550 267277 258602 267283
rect 258410 267225 258550 267228
rect 258358 267219 258602 267225
rect 258370 267200 258590 267219
rect 258646 267203 258698 267209
rect 258646 267145 258698 267151
rect 258262 267129 258314 267135
rect 257780 267094 257836 267103
rect 258454 267129 258506 267135
rect 258314 267077 258454 267080
rect 258262 267071 258506 267077
rect 258274 267052 258494 267071
rect 257780 267029 257836 267038
rect 257686 262763 257738 262769
rect 257686 262705 257738 262711
rect 257794 258630 257822 267029
rect 258452 266946 258508 266955
rect 258452 266881 258508 266890
rect 258466 258644 258494 266881
rect 258658 263287 258686 267145
rect 258932 266798 258988 266807
rect 258932 266733 258988 266742
rect 258646 263281 258698 263287
rect 258646 263223 258698 263229
rect 258946 258644 258974 266733
rect 259028 266650 259084 266659
rect 259028 266585 259084 266594
rect 258240 258616 258494 258644
rect 258720 258616 258974 258644
rect 259042 258630 259070 266585
rect 259138 266395 259166 267737
rect 259508 266502 259564 266511
rect 259508 266437 259564 266446
rect 259126 266389 259178 266395
rect 259126 266331 259178 266337
rect 259522 258630 259550 266437
rect 259714 260993 259742 275650
rect 259988 266354 260044 266363
rect 259988 266289 260044 266298
rect 259702 260987 259754 260993
rect 259702 260929 259754 260935
rect 260002 258630 260030 266289
rect 260962 262695 260990 275650
rect 262114 273721 262142 275650
rect 262102 273715 262154 273721
rect 262102 273657 262154 273663
rect 261046 272531 261098 272537
rect 261046 272473 261098 272479
rect 260950 262689 261002 262695
rect 260950 262631 261002 262637
rect 260662 261061 260714 261067
rect 260662 261003 260714 261009
rect 260674 258644 260702 261003
rect 261058 258644 261086 272473
rect 261238 262985 261290 262991
rect 261238 262927 261290 262933
rect 260448 258616 260702 258644
rect 260832 258616 261086 258644
rect 261250 258630 261278 262927
rect 263362 261955 263390 275650
rect 264514 268393 264542 275650
rect 264502 268387 264554 268393
rect 264502 268329 264554 268335
rect 266050 266469 266078 275784
rect 266518 272235 266570 272241
rect 266518 272177 266570 272183
rect 266038 266463 266090 266469
rect 266038 266405 266090 266411
rect 263444 262062 263500 262071
rect 263444 261997 263500 262006
rect 262102 261949 262154 261955
rect 262102 261891 262154 261897
rect 263350 261949 263402 261955
rect 263350 261891 263402 261897
rect 261718 260987 261770 260993
rect 261718 260929 261770 260935
rect 261730 258630 261758 260929
rect 262114 260771 262142 261891
rect 262102 260765 262154 260771
rect 262102 260707 262154 260713
rect 262198 260765 262250 260771
rect 262198 260707 262250 260713
rect 262210 258630 262238 260707
rect 263252 260434 263308 260443
rect 263252 260369 263308 260378
rect 262772 260286 262828 260295
rect 262772 260221 262828 260230
rect 262786 258644 262814 260221
rect 263266 258644 263294 260369
rect 262560 258616 262814 258644
rect 263040 258616 263294 258644
rect 263458 258630 263486 261997
rect 263924 261766 263980 261775
rect 263924 261701 263980 261710
rect 263938 258630 263966 261701
rect 264308 261470 264364 261479
rect 264308 261405 264364 261414
rect 264322 258630 264350 261405
rect 264884 261322 264940 261331
rect 264884 261257 264940 261266
rect 264898 258644 264926 261257
rect 265460 261174 265516 261183
rect 265460 261109 265516 261118
rect 265474 258644 265502 261109
rect 265844 261026 265900 261035
rect 265844 260961 265900 260970
rect 265858 258644 265886 260961
rect 266036 260878 266092 260887
rect 266036 260813 266092 260822
rect 264768 258616 264926 258644
rect 265248 258616 265502 258644
rect 265632 258616 265886 258644
rect 266050 258630 266078 260813
rect 266530 258630 266558 272177
rect 266818 260327 266846 275650
rect 268244 273606 268300 273615
rect 268244 273541 268300 273550
rect 267764 273458 267820 273467
rect 267764 273393 267820 273402
rect 267190 272161 267242 272167
rect 267190 272103 267242 272109
rect 266806 260321 266858 260327
rect 266806 260263 266858 260269
rect 267202 258644 267230 272103
rect 267572 271978 267628 271987
rect 267572 271913 267628 271922
rect 267586 258644 267614 271913
rect 267778 258792 267806 273393
rect 267862 268535 267914 268541
rect 267862 268477 267914 268483
rect 267874 265877 267902 268477
rect 267862 265871 267914 265877
rect 267862 265813 267914 265819
rect 267778 258764 267854 258792
rect 266976 258616 267230 258644
rect 267360 258616 267614 258644
rect 267826 258630 267854 258764
rect 268258 258630 268286 273541
rect 268354 262621 268382 275784
rect 280834 275784 281136 275812
rect 283536 275784 283838 275812
rect 296688 275784 296798 275812
rect 268724 273310 268780 273319
rect 268724 273245 268780 273254
rect 268342 262615 268394 262621
rect 268342 262557 268394 262563
rect 268738 258630 268766 273245
rect 269108 273162 269164 273171
rect 269108 273097 269164 273106
rect 269122 258630 269150 273097
rect 269218 268615 269246 275650
rect 269780 273014 269836 273023
rect 269780 272949 269836 272958
rect 269206 268609 269258 268615
rect 269206 268551 269258 268557
rect 269794 258644 269822 272949
rect 270260 272866 270316 272875
rect 270260 272801 270316 272810
rect 270274 258644 270302 272801
rect 270370 271723 270398 275650
rect 270452 272718 270508 272727
rect 270452 272653 270508 272662
rect 270358 271717 270410 271723
rect 270358 271659 270410 271665
rect 269568 258616 269822 258644
rect 270048 258616 270302 258644
rect 270466 258630 270494 272653
rect 270836 272570 270892 272579
rect 270836 272505 270892 272514
rect 270850 258630 270878 272505
rect 271316 272422 271372 272431
rect 271316 272357 271372 272366
rect 271330 258630 271358 272357
rect 271618 268319 271646 275650
rect 272564 272274 272620 272283
rect 272564 272209 272620 272218
rect 271606 268313 271658 268319
rect 271606 268255 271658 268261
rect 271988 260730 272044 260739
rect 271988 260665 272044 260674
rect 272002 258644 272030 260665
rect 272372 260582 272428 260591
rect 272372 260517 272428 260526
rect 272386 258644 272414 260517
rect 271776 258616 272030 258644
rect 272160 258616 272414 258644
rect 272578 258630 272606 272209
rect 272770 268541 272798 275650
rect 273044 272126 273100 272135
rect 273044 272061 273100 272070
rect 272758 268535 272810 268541
rect 272758 268477 272810 268483
rect 272854 266241 272906 266247
rect 272854 266183 272906 266189
rect 272662 266167 272714 266173
rect 272662 266109 272714 266115
rect 272674 265581 272702 266109
rect 272662 265575 272714 265581
rect 272662 265517 272714 265523
rect 272866 262843 272894 266183
rect 272854 262837 272906 262843
rect 272854 262779 272906 262785
rect 273058 258630 273086 272061
rect 274018 271945 274046 275650
rect 274006 271939 274058 271945
rect 274006 271881 274058 271887
rect 274774 266907 274826 266913
rect 274774 266849 274826 266855
rect 274198 266759 274250 266765
rect 274198 266701 274250 266707
rect 273622 266611 273674 266617
rect 273622 266553 273674 266559
rect 273526 266167 273578 266173
rect 273526 266109 273578 266115
rect 273538 258630 273566 266109
rect 273634 258644 273662 266553
rect 274102 266167 274154 266173
rect 274102 266109 274154 266115
rect 274114 262917 274142 266109
rect 274102 262911 274154 262917
rect 274102 262853 274154 262859
rect 274210 258644 274238 266701
rect 273634 258616 273888 258644
rect 274210 258616 274368 258644
rect 274786 258630 274814 266849
rect 275170 262695 275198 275650
rect 275926 267869 275978 267875
rect 275926 267811 275978 267817
rect 275638 267647 275690 267653
rect 275638 267589 275690 267595
rect 275254 267277 275306 267283
rect 275254 267219 275306 267225
rect 275158 262689 275210 262695
rect 275158 262631 275210 262637
rect 275266 258630 275294 267219
rect 275650 258630 275678 267589
rect 275938 265655 275966 267811
rect 276418 266913 276446 275650
rect 277570 272093 277598 275650
rect 277558 272087 277610 272093
rect 277558 272029 277610 272035
rect 278818 267875 278846 275650
rect 279970 268467 279998 275650
rect 279958 268461 280010 268467
rect 279958 268403 280010 268409
rect 279286 268239 279338 268245
rect 279286 268181 279338 268187
rect 278806 267869 278858 267875
rect 278806 267811 278858 267817
rect 276406 266907 276458 266913
rect 276406 266849 276458 266855
rect 276502 265945 276554 265951
rect 276502 265887 276554 265893
rect 275830 265649 275882 265655
rect 275830 265591 275882 265597
rect 275926 265649 275978 265655
rect 275926 265591 275978 265597
rect 275842 258644 275870 265591
rect 276514 258644 276542 265887
rect 276982 265797 277034 265803
rect 276982 265739 277034 265745
rect 275842 258616 276096 258644
rect 276514 258616 276576 258644
rect 276994 258630 277022 265739
rect 277366 265723 277418 265729
rect 277366 265665 277418 265671
rect 277378 258630 277406 265665
rect 277846 265501 277898 265507
rect 277846 265443 277898 265449
rect 277858 258630 277886 265443
rect 278038 265427 278090 265433
rect 278038 265369 278090 265375
rect 278050 258644 278078 265369
rect 278518 265353 278570 265359
rect 278518 265295 278570 265301
rect 278530 258644 278558 265295
rect 279094 265279 279146 265285
rect 279094 265221 279146 265227
rect 278050 258616 278304 258644
rect 278530 258616 278784 258644
rect 279106 258630 279134 265221
rect 279298 263107 279326 268181
rect 279574 265575 279626 265581
rect 279574 265517 279626 265523
rect 279284 263098 279340 263107
rect 279284 263033 279340 263042
rect 279586 258630 279614 265517
rect 280054 265205 280106 265211
rect 280054 265147 280106 265153
rect 280066 258630 280094 265147
rect 280150 265131 280202 265137
rect 280150 265073 280202 265079
rect 280162 258644 280190 265073
rect 280630 265057 280682 265063
rect 280630 264999 280682 265005
rect 280642 258644 280670 264999
rect 280834 260475 280862 275784
rect 282166 268387 282218 268393
rect 282166 268329 282218 268335
rect 281302 262763 281354 262769
rect 281302 262705 281354 262711
rect 280822 260469 280874 260475
rect 280822 260411 280874 260417
rect 280162 258616 280416 258644
rect 280642 258616 280896 258644
rect 281314 258630 281342 262705
rect 281782 262467 281834 262473
rect 281782 262409 281834 262415
rect 281794 258630 281822 262409
rect 282178 258630 282206 268329
rect 282370 262769 282398 275650
rect 283810 268911 283838 275784
rect 284674 272833 284702 275650
rect 284662 272827 284714 272833
rect 284662 272769 284714 272775
rect 283798 268905 283850 268911
rect 283798 268847 283850 268853
rect 282838 268313 282890 268319
rect 282838 268255 282890 268261
rect 282358 262763 282410 262769
rect 282358 262705 282410 262711
rect 282358 262615 282410 262621
rect 282358 262557 282410 262563
rect 282370 258644 282398 262557
rect 282850 258644 282878 268255
rect 283894 267869 283946 267875
rect 283894 267811 283946 267817
rect 285622 267869 285674 267875
rect 285622 267811 285674 267817
rect 283510 262689 283562 262695
rect 283510 262631 283562 262637
rect 282370 258616 282624 258644
rect 282850 258616 283104 258644
rect 283522 258630 283550 262631
rect 283906 258630 283934 267811
rect 285526 262911 285578 262917
rect 285526 262853 285578 262859
rect 284374 262763 284426 262769
rect 284374 262705 284426 262711
rect 284386 258630 284414 262705
rect 285046 262615 285098 262621
rect 285046 262557 285098 262563
rect 285058 258644 285086 262557
rect 285538 258644 285566 262853
rect 284832 258616 285086 258644
rect 285312 258616 285566 258644
rect 285634 258630 285662 267811
rect 285826 262621 285854 275650
rect 286102 268387 286154 268393
rect 286102 268329 286154 268335
rect 285814 262615 285866 262621
rect 285814 262557 285866 262563
rect 286114 258630 286142 268329
rect 287074 268171 287102 275650
rect 287062 268165 287114 268171
rect 287062 268107 287114 268113
rect 287638 268091 287690 268097
rect 287638 268033 287690 268039
rect 286582 263281 286634 263287
rect 286582 263223 286634 263229
rect 286594 258630 286622 263223
rect 287254 262689 287306 262695
rect 287254 262631 287306 262637
rect 287266 258644 287294 262631
rect 287650 258644 287678 268033
rect 287830 262541 287882 262547
rect 287830 262483 287882 262489
rect 287040 258616 287294 258644
rect 287424 258616 287678 258644
rect 287842 258630 287870 262483
rect 288226 261363 288254 275650
rect 288310 266759 288362 266765
rect 288310 266701 288362 266707
rect 288214 261357 288266 261363
rect 288214 261299 288266 261305
rect 288322 258630 288350 266701
rect 289366 266611 289418 266617
rect 289366 266553 289418 266559
rect 288694 266389 288746 266395
rect 288694 266331 288746 266337
rect 288706 258630 288734 266331
rect 289378 258644 289406 266553
rect 289474 262917 289502 275650
rect 290640 275636 290846 275664
rect 290818 267820 290846 275636
rect 291874 272759 291902 275650
rect 291862 272753 291914 272759
rect 291862 272695 291914 272701
rect 293026 267875 293054 275650
rect 294274 268245 294302 275650
rect 294838 271199 294890 271205
rect 294838 271141 294890 271147
rect 294262 268239 294314 268245
rect 294262 268181 294314 268187
rect 293014 267869 293066 267875
rect 290818 267792 291038 267820
rect 293014 267811 293066 267817
rect 289846 267277 289898 267283
rect 289846 267219 289898 267225
rect 289462 262911 289514 262917
rect 289462 262853 289514 262859
rect 289858 258644 289886 267219
rect 290422 265205 290474 265211
rect 290422 265147 290474 265153
rect 290038 265057 290090 265063
rect 290038 264999 290090 265005
rect 289152 258616 289406 258644
rect 289632 258616 289886 258644
rect 290050 258630 290078 264999
rect 290434 258630 290462 265147
rect 291010 262917 291038 267792
rect 294166 266907 294218 266913
rect 294166 266849 294218 266855
rect 294070 265797 294122 265803
rect 294070 265739 294122 265745
rect 293686 265723 293738 265729
rect 293686 265665 293738 265671
rect 293110 265575 293162 265581
rect 293110 265517 293162 265523
rect 292630 265501 292682 265507
rect 292630 265443 292682 265449
rect 292150 265427 292202 265433
rect 292150 265369 292202 265375
rect 292054 265353 292106 265359
rect 292054 265295 292106 265301
rect 291574 265279 291626 265285
rect 291574 265221 291626 265227
rect 291190 265131 291242 265137
rect 291190 265073 291242 265079
rect 290998 262911 291050 262917
rect 290998 262853 291050 262859
rect 291202 258644 291230 265073
rect 291586 258644 291614 265221
rect 292066 258644 292094 265295
rect 290928 258616 291230 258644
rect 291360 258616 291614 258644
rect 291840 258616 292094 258644
rect 292162 258630 292190 265369
rect 292642 258630 292670 265443
rect 293122 258630 293150 265517
rect 293698 258644 293726 265665
rect 294082 258644 294110 265739
rect 294178 262843 294206 266849
rect 294166 262837 294218 262843
rect 294166 262779 294218 262785
rect 294358 259507 294410 259513
rect 294358 259449 294410 259455
rect 293568 258616 293726 258644
rect 293952 258616 294110 258644
rect 294370 258630 294398 259449
rect 294850 258630 294878 271141
rect 295426 261289 295454 275650
rect 296566 271125 296618 271131
rect 296566 271067 296618 271073
rect 295894 271051 295946 271057
rect 295894 270993 295946 270999
rect 295414 261283 295466 261289
rect 295414 261225 295466 261231
rect 295318 259581 295370 259587
rect 295318 259523 295370 259529
rect 295330 258630 295358 259523
rect 295906 258644 295934 270993
rect 296374 259655 296426 259661
rect 296374 259597 296426 259603
rect 296386 258644 296414 259597
rect 295680 258616 295934 258644
rect 296160 258616 296414 258644
rect 296578 258630 296606 271067
rect 296770 268393 296798 275784
rect 297430 270977 297482 270983
rect 297430 270919 297482 270925
rect 296758 268387 296810 268393
rect 296758 268329 296810 268335
rect 296950 259729 297002 259735
rect 296950 259671 297002 259677
rect 296962 258630 296990 259671
rect 297442 258630 297470 270919
rect 297826 262769 297854 275650
rect 298978 272685 299006 275650
rect 298966 272679 299018 272685
rect 298966 272621 299018 272627
rect 299158 271643 299210 271649
rect 299158 271585 299210 271591
rect 298486 271347 298538 271353
rect 298486 271289 298538 271295
rect 297814 262763 297866 262769
rect 297814 262705 297866 262711
rect 298006 261209 298058 261215
rect 298006 261151 298058 261157
rect 298018 260919 298046 261151
rect 298006 260913 298058 260919
rect 298006 260855 298058 260861
rect 298102 259803 298154 259809
rect 298102 259745 298154 259751
rect 298114 258644 298142 259745
rect 298498 258644 298526 271289
rect 298582 268387 298634 268393
rect 298582 268329 298634 268335
rect 298594 268171 298622 268329
rect 298582 268165 298634 268171
rect 298582 268107 298634 268113
rect 298966 259951 299018 259957
rect 298966 259893 299018 259899
rect 298978 258644 299006 259893
rect 297888 258616 298142 258644
rect 298368 258616 298526 258644
rect 298752 258616 299006 258644
rect 299170 258630 299198 271585
rect 299542 266463 299594 266469
rect 299542 266405 299594 266411
rect 299554 262621 299582 266405
rect 300130 263287 300158 275650
rect 300310 271717 300362 271723
rect 300310 271659 300362 271665
rect 300118 263281 300170 263287
rect 300118 263223 300170 263229
rect 299542 262615 299594 262621
rect 299542 262557 299594 262563
rect 299638 260099 299690 260105
rect 299638 260041 299690 260047
rect 299650 258630 299678 260041
rect 300322 258644 300350 271659
rect 301282 268245 301310 275650
rect 302230 272087 302282 272093
rect 302230 272029 302282 272035
rect 301366 271939 301418 271945
rect 301366 271881 301418 271887
rect 301270 268239 301322 268245
rect 301270 268181 301322 268187
rect 300694 265945 300746 265951
rect 300694 265887 300746 265893
rect 300706 258644 300734 265887
rect 301174 260321 301226 260327
rect 301174 260263 301226 260269
rect 301186 258644 301214 260263
rect 300096 258616 300350 258644
rect 300480 258616 300734 258644
rect 300960 258616 301214 258644
rect 301378 258630 301406 271881
rect 301846 260469 301898 260475
rect 301846 260411 301898 260417
rect 301858 258630 301886 260411
rect 302242 258630 302270 272029
rect 302530 261289 302558 275650
rect 302902 273789 302954 273795
rect 302902 273731 302954 273737
rect 302518 261283 302570 261289
rect 302518 261225 302570 261231
rect 302914 258644 302942 273731
rect 303394 258644 303422 276321
rect 397558 276305 397610 276311
rect 397558 276247 397610 276253
rect 386326 276157 386378 276163
rect 386326 276099 386378 276105
rect 303574 276009 303626 276015
rect 303574 275951 303626 275957
rect 302688 258616 302942 258644
rect 303168 258616 303422 258644
rect 303586 258630 303614 275951
rect 303958 275935 304010 275941
rect 303958 275877 304010 275883
rect 303682 262695 303710 275650
rect 303670 262689 303722 262695
rect 303670 262631 303722 262637
rect 303970 258630 303998 275877
rect 304438 275861 304490 275867
rect 304438 275803 304490 275809
rect 304450 258630 304478 275803
rect 305110 275787 305162 275793
rect 312144 275784 312446 275812
rect 305110 275729 305162 275735
rect 304930 262695 304958 275650
rect 304918 262689 304970 262695
rect 304918 262631 304970 262637
rect 305122 258644 305150 275729
rect 305206 275713 305258 275719
rect 305206 275655 305258 275661
rect 304896 258616 305150 258644
rect 305218 258644 305246 275655
rect 306082 272611 306110 275650
rect 306646 275565 306698 275571
rect 306646 275507 306698 275513
rect 306166 273641 306218 273647
rect 306166 273583 306218 273589
rect 306070 272605 306122 272611
rect 306070 272547 306122 272553
rect 305686 260913 305738 260919
rect 305686 260855 305738 260861
rect 305218 258616 305280 258644
rect 305698 258630 305726 260855
rect 306178 258630 306206 273583
rect 306658 258630 306686 275507
rect 307222 275491 307274 275497
rect 307222 275433 307274 275439
rect 307234 258644 307262 275433
rect 307330 268097 307358 275650
rect 307702 275417 307754 275423
rect 307702 275359 307754 275365
rect 307318 268091 307370 268097
rect 307318 268033 307370 268039
rect 307714 258644 307742 275359
rect 307894 275343 307946 275349
rect 307894 275285 307946 275291
rect 307008 258616 307262 258644
rect 307488 258616 307742 258644
rect 307906 258630 307934 275285
rect 308374 275269 308426 275275
rect 308374 275211 308426 275217
rect 308182 261283 308234 261289
rect 308182 261225 308234 261231
rect 308194 259883 308222 261225
rect 308086 259877 308138 259883
rect 308086 259819 308138 259825
rect 308182 259877 308234 259883
rect 308182 259819 308234 259825
rect 308098 259439 308126 259819
rect 308086 259433 308138 259439
rect 308086 259375 308138 259381
rect 308386 258630 308414 275211
rect 308482 268171 308510 275650
rect 308758 275195 308810 275201
rect 308758 275137 308810 275143
rect 308470 268165 308522 268171
rect 308470 268107 308522 268113
rect 308770 258630 308798 275137
rect 309430 275121 309482 275127
rect 309430 275063 309482 275069
rect 309442 258644 309470 275063
rect 309730 261141 309758 275650
rect 309910 275047 309962 275053
rect 309910 274989 309962 274995
rect 309718 261135 309770 261141
rect 309718 261077 309770 261083
rect 309922 258644 309950 274989
rect 310102 274973 310154 274979
rect 310102 274915 310154 274921
rect 309216 258616 309470 258644
rect 309696 258616 309950 258644
rect 310114 258630 310142 274915
rect 310486 274899 310538 274905
rect 310486 274841 310538 274847
rect 310498 258630 310526 274841
rect 310882 262547 310910 275650
rect 311638 274825 311690 274831
rect 311638 274767 311690 274773
rect 310966 274751 311018 274757
rect 310966 274693 311018 274699
rect 310870 262541 310922 262547
rect 310870 262483 310922 262489
rect 310978 258630 311006 274693
rect 311650 258644 311678 274767
rect 312118 274677 312170 274683
rect 312118 274619 312170 274625
rect 312130 258644 312158 274619
rect 312214 274603 312266 274609
rect 312214 274545 312266 274551
rect 311424 258616 311678 258644
rect 311904 258616 312158 258644
rect 312226 258630 312254 274545
rect 312418 262547 312446 275784
rect 327202 275784 327504 275812
rect 342754 275784 342960 275812
rect 345058 275784 345360 275812
rect 358114 275784 358416 275812
rect 373570 275784 373872 275812
rect 375970 275784 376272 275812
rect 312694 274529 312746 274535
rect 312694 274471 312746 274477
rect 312406 262541 312458 262547
rect 312406 262483 312458 262489
rect 312706 258630 312734 274471
rect 313174 274455 313226 274461
rect 313174 274397 313226 274403
rect 313186 258630 313214 274397
rect 313282 272463 313310 275650
rect 313750 274381 313802 274387
rect 313750 274323 313802 274329
rect 313270 272457 313322 272463
rect 313270 272399 313322 272405
rect 313762 258644 313790 274323
rect 313942 268683 313994 268689
rect 313942 268625 313994 268631
rect 313954 262473 313982 268625
rect 314434 266765 314462 275650
rect 314710 274307 314762 274313
rect 314710 274249 314762 274255
rect 314422 266759 314474 266765
rect 314422 266701 314474 266707
rect 314230 266389 314282 266395
rect 314230 266331 314282 266337
rect 313942 262467 313994 262473
rect 313942 262409 313994 262415
rect 314242 258644 314270 266331
rect 314722 258644 314750 274249
rect 314902 274233 314954 274239
rect 314902 274175 314954 274181
rect 313536 258616 313790 258644
rect 314016 258616 314270 258644
rect 314448 258616 314750 258644
rect 314914 258630 314942 274175
rect 315286 274159 315338 274165
rect 315286 274101 315338 274107
rect 315298 258630 315326 274101
rect 315682 268097 315710 275650
rect 315958 274085 316010 274091
rect 315958 274027 316010 274033
rect 315670 268091 315722 268097
rect 315670 268033 315722 268039
rect 315970 258644 315998 274027
rect 316438 274011 316490 274017
rect 316438 273953 316490 273959
rect 316450 258644 316478 273953
rect 316630 273937 316682 273943
rect 316630 273879 316682 273885
rect 315744 258616 315998 258644
rect 316224 258616 316478 258644
rect 316642 258630 316670 273879
rect 316738 261215 316766 275650
rect 317494 267647 317546 267653
rect 317494 267589 317546 267595
rect 317014 262393 317066 262399
rect 317014 262335 317066 262341
rect 316726 261209 316778 261215
rect 316726 261151 316778 261157
rect 317026 258630 317054 262335
rect 317506 258630 317534 267589
rect 317986 266469 318014 275650
rect 319138 267949 319166 275650
rect 320386 272389 320414 275650
rect 320374 272383 320426 272389
rect 320374 272325 320426 272331
rect 320950 270829 321002 270835
rect 320950 270771 321002 270777
rect 319126 267943 319178 267949
rect 319126 267885 319178 267891
rect 319220 267686 319276 267695
rect 319220 267621 319276 267630
rect 318070 266907 318122 266913
rect 318070 266849 318122 266855
rect 317974 266463 318026 266469
rect 317974 266405 318026 266411
rect 318082 262048 318110 266849
rect 318646 266759 318698 266765
rect 318646 266701 318698 266707
rect 318166 265205 318218 265211
rect 318218 265153 318398 265156
rect 318166 265147 318398 265153
rect 318178 265137 318398 265147
rect 318178 265131 318410 265137
rect 318178 265128 318358 265131
rect 318358 265073 318410 265079
rect 317986 262020 318110 262048
rect 317986 258496 318014 262020
rect 318358 261283 318410 261289
rect 318358 261225 318410 261231
rect 318070 261135 318122 261141
rect 318070 261077 318122 261083
rect 318082 260031 318110 261077
rect 318262 260913 318314 260919
rect 318262 260855 318314 260861
rect 318166 260691 318218 260697
rect 318166 260633 318218 260639
rect 318178 260031 318206 260633
rect 318070 260025 318122 260031
rect 318070 259967 318122 259973
rect 318166 260025 318218 260031
rect 318166 259967 318218 259973
rect 318274 259439 318302 260855
rect 318370 260697 318398 261225
rect 318358 260691 318410 260697
rect 318358 260633 318410 260639
rect 318262 259433 318314 259439
rect 318262 259375 318314 259381
rect 318658 258644 318686 266701
rect 318742 266463 318794 266469
rect 318742 266405 318794 266411
rect 318432 258616 318686 258644
rect 318754 258630 318782 266405
rect 319234 258630 319262 267621
rect 320276 267538 320332 267547
rect 320276 267473 320332 267482
rect 319606 266389 319658 266395
rect 319606 266331 319658 266337
rect 319702 266389 319754 266395
rect 319702 266331 319754 266337
rect 319618 265919 319646 266331
rect 319604 265910 319660 265919
rect 319604 265845 319660 265854
rect 319714 258630 319742 266331
rect 320290 258644 320318 267473
rect 320758 261431 320810 261437
rect 320758 261373 320810 261379
rect 320770 258644 320798 261373
rect 320064 258616 320318 258644
rect 320544 258616 320798 258644
rect 320962 258630 320990 270771
rect 321538 266617 321566 275650
rect 322102 272827 322154 272833
rect 322102 272769 322154 272775
rect 321814 267647 321866 267653
rect 321814 267589 321866 267595
rect 321910 267647 321962 267653
rect 321910 267589 321962 267595
rect 321826 266913 321854 267589
rect 321718 266907 321770 266913
rect 321718 266849 321770 266855
rect 321814 266907 321866 266913
rect 321814 266849 321866 266855
rect 321730 266765 321758 266849
rect 321622 266759 321674 266765
rect 321622 266701 321674 266707
rect 321718 266759 321770 266765
rect 321718 266701 321770 266707
rect 321634 266617 321662 266701
rect 321526 266611 321578 266617
rect 321526 266553 321578 266559
rect 321622 266611 321674 266617
rect 321622 266553 321674 266559
rect 321922 265919 321950 267589
rect 321908 265910 321964 265919
rect 321908 265845 321964 265854
rect 321430 261357 321482 261363
rect 321430 261299 321482 261305
rect 321442 258630 321470 261299
rect 322114 258644 322142 272769
rect 322786 268023 322814 275650
rect 322966 272753 323018 272759
rect 322966 272695 323018 272701
rect 322774 268017 322826 268023
rect 322774 267959 322826 267965
rect 322486 261283 322538 261289
rect 322486 261225 322538 261231
rect 322498 258644 322526 261225
rect 322978 258644 323006 272695
rect 323542 272679 323594 272685
rect 323542 272621 323594 272627
rect 323158 261209 323210 261215
rect 323158 261151 323210 261157
rect 321840 258616 322142 258644
rect 322272 258616 322526 258644
rect 322752 258616 323006 258644
rect 323170 258630 323198 261151
rect 323554 258630 323582 272621
rect 323938 260845 323966 275650
rect 324694 272605 324746 272611
rect 324694 272547 324746 272553
rect 324406 268757 324458 268763
rect 324406 268699 324458 268705
rect 324418 267875 324446 268699
rect 324406 267869 324458 267875
rect 324406 267811 324458 267817
rect 324022 261949 324074 261955
rect 324022 261891 324074 261897
rect 323926 260839 323978 260845
rect 323926 260781 323978 260787
rect 324034 258630 324062 261891
rect 324706 258644 324734 272547
rect 325186 267283 325214 275650
rect 326352 275636 327038 275664
rect 325270 272457 325322 272463
rect 325270 272399 325322 272405
rect 325174 267277 325226 267283
rect 325174 267219 325226 267225
rect 325174 260913 325226 260919
rect 325174 260855 325226 260861
rect 325186 258644 325214 260855
rect 324480 258616 324734 258644
rect 324960 258616 325214 258644
rect 325282 258630 325310 272399
rect 326230 272383 326282 272389
rect 326230 272325 326282 272331
rect 325462 267277 325514 267283
rect 325462 267219 325514 267225
rect 325474 262399 325502 267219
rect 325462 262393 325514 262399
rect 325462 262335 325514 262341
rect 325750 260839 325802 260845
rect 325750 260781 325802 260787
rect 325762 258630 325790 260781
rect 326242 258630 326270 272325
rect 326804 268722 326860 268731
rect 326804 268657 326860 268666
rect 326818 262991 326846 268657
rect 327010 262991 327038 275636
rect 327202 272315 327230 275784
rect 327862 272827 327914 272833
rect 327862 272769 327914 272775
rect 327394 272537 327614 272556
rect 327382 272531 327626 272537
rect 327434 272528 327574 272531
rect 327382 272473 327434 272479
rect 327574 272473 327626 272479
rect 327190 272309 327242 272315
rect 327190 272251 327242 272257
rect 327286 271495 327338 271501
rect 327286 271437 327338 271443
rect 327094 270681 327146 270687
rect 327094 270623 327146 270629
rect 326806 262985 326858 262991
rect 326806 262927 326858 262933
rect 326998 262985 327050 262991
rect 326998 262927 327050 262933
rect 327106 262399 327134 270623
rect 327094 262393 327146 262399
rect 327094 262335 327146 262341
rect 326900 261914 326956 261923
rect 326900 261849 326956 261858
rect 326914 258644 326942 261849
rect 327298 258644 327326 271437
rect 327766 270903 327818 270909
rect 327766 270845 327818 270851
rect 327778 263287 327806 270845
rect 327874 270835 327902 272769
rect 327862 270829 327914 270835
rect 327862 270771 327914 270777
rect 327958 270829 328010 270835
rect 327958 270771 328010 270777
rect 327766 263281 327818 263287
rect 327766 263223 327818 263229
rect 327476 261618 327532 261627
rect 327476 261553 327532 261562
rect 326688 258616 326942 258644
rect 327072 258616 327326 258644
rect 327490 258630 327518 261553
rect 327970 258630 327998 270771
rect 328738 265063 328766 275650
rect 328918 270903 328970 270909
rect 328918 270845 328970 270851
rect 328726 265057 328778 265063
rect 328726 264999 328778 265005
rect 328246 260691 328298 260697
rect 328246 260633 328298 260639
rect 328342 260691 328394 260697
rect 328342 260633 328394 260639
rect 328258 259883 328286 260633
rect 328246 259877 328298 259883
rect 328246 259819 328298 259825
rect 328354 258630 328382 260633
rect 328930 258644 328958 270845
rect 329890 270687 329918 275650
rect 331030 271273 331082 271279
rect 331030 271215 331082 271221
rect 329878 270681 329930 270687
rect 329878 270623 329930 270629
rect 330166 267869 330218 267875
rect 330166 267811 330218 267817
rect 329014 266315 329066 266321
rect 329014 266257 329066 266263
rect 328800 258616 328958 258644
rect 329026 258644 329054 266257
rect 329686 263355 329738 263361
rect 329686 263297 329738 263303
rect 329026 258616 329280 258644
rect 329698 258630 329726 263297
rect 330178 263139 330206 267811
rect 330070 263133 330122 263139
rect 330070 263075 330122 263081
rect 330166 263133 330218 263139
rect 330166 263075 330218 263081
rect 330082 258630 330110 263075
rect 331042 263065 331070 271215
rect 330742 263059 330794 263065
rect 330742 263001 330794 263007
rect 331030 263059 331082 263065
rect 331030 263001 331082 263007
rect 330550 262171 330602 262177
rect 330550 262113 330602 262119
rect 330562 258630 330590 262113
rect 330754 258644 330782 263001
rect 331138 260031 331166 275650
rect 331990 268683 332042 268689
rect 331990 268625 332042 268631
rect 331222 268609 331274 268615
rect 331222 268551 331274 268557
rect 331234 263361 331262 268551
rect 331606 263429 331658 263435
rect 331606 263371 331658 263377
rect 331222 263355 331274 263361
rect 331222 263297 331274 263303
rect 331222 262467 331274 262473
rect 331222 262409 331274 262415
rect 331126 260025 331178 260031
rect 331126 259967 331178 259973
rect 331234 258644 331262 262409
rect 331618 258644 331646 263371
rect 332002 258644 332030 268625
rect 332290 265137 332318 275650
rect 333334 270755 333386 270761
rect 333334 270697 333386 270703
rect 332278 265131 332330 265137
rect 332278 265073 332330 265079
rect 332758 264983 332810 264989
rect 332758 264925 332810 264931
rect 330754 258616 331008 258644
rect 331234 258616 331488 258644
rect 331618 258616 331872 258644
rect 332002 258616 332304 258644
rect 332770 258630 332798 264925
rect 332950 263133 333002 263139
rect 332950 263075 333002 263081
rect 332962 258644 332990 263075
rect 333346 258644 333374 270697
rect 333442 264989 333470 275650
rect 334594 271427 334622 275650
rect 334582 271421 334634 271427
rect 334582 271363 334634 271369
rect 334102 268535 334154 268541
rect 334102 268477 334154 268483
rect 334114 264989 334142 268477
rect 334198 268461 334250 268467
rect 334198 268403 334250 268409
rect 333430 264983 333482 264989
rect 333430 264925 333482 264931
rect 334102 264983 334154 264989
rect 334102 264925 334154 264931
rect 334210 263435 334238 268403
rect 334966 265871 335018 265877
rect 334966 265813 335018 265819
rect 334198 263429 334250 263435
rect 334198 263371 334250 263377
rect 334486 263059 334538 263065
rect 334486 263001 334538 263007
rect 334006 259877 334058 259883
rect 334006 259819 334058 259825
rect 334018 258644 334046 259819
rect 332962 258616 333216 258644
rect 333346 258616 333600 258644
rect 334018 258616 334080 258644
rect 334498 258630 334526 263001
rect 334978 258630 335006 265813
rect 335842 265211 335870 275650
rect 336994 268467 337022 275650
rect 337558 273715 337610 273721
rect 337558 273657 337610 273663
rect 337090 270613 337406 270632
rect 337078 270607 337406 270613
rect 337130 270604 337406 270607
rect 337078 270549 337130 270555
rect 337090 270465 337310 270484
rect 337078 270459 337310 270465
rect 337130 270456 337310 270459
rect 337078 270401 337130 270407
rect 337078 270311 337130 270317
rect 337078 270253 337130 270259
rect 337090 270040 337118 270253
rect 337090 270012 337214 270040
rect 337078 269941 337130 269947
rect 337078 269883 337130 269889
rect 337090 268911 337118 269883
rect 337078 268905 337130 268911
rect 337078 268847 337130 268853
rect 337186 268763 337214 270012
rect 337174 268757 337226 268763
rect 337174 268699 337226 268705
rect 337282 268615 337310 270456
rect 337378 269947 337406 270604
rect 337366 269941 337418 269947
rect 337366 269883 337418 269889
rect 337270 268609 337322 268615
rect 337270 268551 337322 268557
rect 336982 268461 337034 268467
rect 336982 268403 337034 268409
rect 337078 265649 337130 265655
rect 337078 265591 337130 265597
rect 335830 265205 335882 265211
rect 335830 265147 335882 265153
rect 336598 263503 336650 263509
rect 336598 263445 336650 263451
rect 335542 263281 335594 263287
rect 335542 263223 335594 263229
rect 335350 262171 335402 262177
rect 335350 262113 335402 262119
rect 335362 258630 335390 262113
rect 335554 258644 335582 263223
rect 336022 262245 336074 262251
rect 336022 262187 336074 262193
rect 336034 258644 336062 262187
rect 335554 258616 335808 258644
rect 336034 258616 336288 258644
rect 336610 258630 336638 263445
rect 337090 258630 337118 265591
rect 337570 258630 337598 273657
rect 338134 263355 338186 263361
rect 338134 263297 338186 263303
rect 337750 262615 337802 262621
rect 337750 262557 337802 262563
rect 337762 258644 337790 262557
rect 338146 258644 338174 263297
rect 338242 261141 338270 275650
rect 339106 275636 339408 275664
rect 338710 268387 338762 268393
rect 338710 268329 338762 268335
rect 338722 263065 338750 268329
rect 339106 265285 339134 275636
rect 339862 268683 339914 268689
rect 339862 268625 339914 268631
rect 339382 268313 339434 268319
rect 339382 268255 339434 268261
rect 339094 265279 339146 265285
rect 339094 265221 339146 265227
rect 338806 264983 338858 264989
rect 338806 264925 338858 264931
rect 338710 263059 338762 263065
rect 338710 263001 338762 263007
rect 338230 261135 338282 261141
rect 338230 261077 338282 261083
rect 337762 258616 338016 258644
rect 338146 258616 338400 258644
rect 338818 258630 338846 264925
rect 339394 262843 339422 268255
rect 339670 268239 339722 268245
rect 339670 268181 339722 268187
rect 339682 263139 339710 268181
rect 339766 263429 339818 263435
rect 339766 263371 339818 263377
rect 339670 263133 339722 263139
rect 339670 263075 339722 263081
rect 339286 262837 339338 262843
rect 339286 262779 339338 262785
rect 339382 262837 339434 262843
rect 339382 262779 339434 262785
rect 339298 258630 339326 262779
rect 339778 258630 339806 263371
rect 339874 258644 339902 268625
rect 340642 263361 340670 275650
rect 341794 271575 341822 275650
rect 341782 271569 341834 271575
rect 341782 271511 341834 271517
rect 341974 268091 342026 268097
rect 341974 268033 342026 268039
rect 341590 267943 341642 267949
rect 341590 267885 341642 267891
rect 340630 263355 340682 263361
rect 340630 263297 340682 263303
rect 340342 263059 340394 263065
rect 340342 263001 340394 263007
rect 340354 258644 340382 263001
rect 341014 262911 341066 262917
rect 341014 262853 341066 262859
rect 339874 258616 340128 258644
rect 340354 258616 340608 258644
rect 341026 258630 341054 262853
rect 341602 262843 341630 267885
rect 341494 262837 341546 262843
rect 341494 262779 341546 262785
rect 341590 262837 341642 262843
rect 341590 262779 341642 262785
rect 341506 258630 341534 262779
rect 341986 262769 342014 268033
rect 342754 265359 342782 275784
rect 343222 268165 343274 268171
rect 343222 268107 343274 268113
rect 342742 265353 342794 265359
rect 342742 265295 342794 265301
rect 342070 263133 342122 263139
rect 342070 263075 342122 263081
rect 341878 262763 341930 262769
rect 341878 262705 341930 262711
rect 341974 262763 342026 262769
rect 341974 262705 342026 262711
rect 341890 258630 341918 262705
rect 342082 258644 342110 263075
rect 342742 262689 342794 262695
rect 342742 262631 342794 262637
rect 342754 258644 342782 262631
rect 342082 258616 342336 258644
rect 342754 258616 342816 258644
rect 343234 258630 343262 268107
rect 344194 267875 344222 275650
rect 344662 268017 344714 268023
rect 344662 267959 344714 267965
rect 344182 267869 344234 267875
rect 344182 267811 344234 267817
rect 344278 262837 344330 262843
rect 344278 262779 344330 262785
rect 344086 262763 344138 262769
rect 344086 262705 344138 262711
rect 343606 262541 343658 262547
rect 343606 262483 343658 262489
rect 343618 258630 343646 262483
rect 344098 258630 344126 262705
rect 344290 258644 344318 262779
rect 344674 258644 344702 267959
rect 345058 260179 345086 275784
rect 345814 270681 345866 270687
rect 345814 270623 345866 270629
rect 345334 262985 345386 262991
rect 345334 262927 345386 262933
rect 345046 260173 345098 260179
rect 345046 260115 345098 260121
rect 344290 258616 344544 258644
rect 344674 258616 344928 258644
rect 345346 258630 345374 262927
rect 345826 258630 345854 270623
rect 346390 268461 346442 268467
rect 346390 268403 346442 268409
rect 346294 264983 346346 264989
rect 346294 264925 346346 264931
rect 346306 258630 346334 264925
rect 346402 258644 346430 268403
rect 346594 265433 346622 275650
rect 347542 267869 347594 267875
rect 347542 267811 347594 267817
rect 346582 265427 346634 265433
rect 346582 265369 346634 265375
rect 346870 263355 346922 263361
rect 346870 263297 346922 263303
rect 346882 258644 346910 263297
rect 346966 261949 347018 261955
rect 346966 261891 347018 261897
rect 346978 261141 347006 261891
rect 346966 261135 347018 261141
rect 346966 261077 347018 261083
rect 346402 258616 346656 258644
rect 346882 258616 347136 258644
rect 347554 258630 347582 267811
rect 347746 258644 347774 275650
rect 348994 271797 349022 275650
rect 348982 271791 349034 271797
rect 348982 271733 349034 271739
rect 349558 268831 349610 268837
rect 349558 268773 349610 268779
rect 348406 264983 348458 264989
rect 348406 264925 348458 264931
rect 347746 258616 348048 258644
rect 348418 258630 348446 264925
rect 349078 263355 349130 263361
rect 349078 263297 349130 263303
rect 349090 258644 349118 263297
rect 349570 258644 349598 268773
rect 350050 265507 350078 275650
rect 351190 270681 351242 270687
rect 351190 270623 351242 270629
rect 350134 268757 350186 268763
rect 350134 268699 350186 268705
rect 350038 265501 350090 265507
rect 350038 265443 350090 265449
rect 349750 263133 349802 263139
rect 349750 263075 349802 263081
rect 348864 258616 349118 258644
rect 349344 258616 349598 258644
rect 349762 258630 349790 263075
rect 350146 258630 350174 268699
rect 350902 265057 350954 265063
rect 350902 264999 350954 265005
rect 350914 258644 350942 264999
rect 351202 258644 351230 270623
rect 351298 264989 351326 275650
rect 351286 264983 351338 264989
rect 351286 264925 351338 264931
rect 351862 262985 351914 262991
rect 351862 262927 351914 262933
rect 351766 262319 351818 262325
rect 351766 262261 351818 262267
rect 351778 258644 351806 262261
rect 350640 258616 350942 258644
rect 351072 258616 351230 258644
rect 351552 258616 351806 258644
rect 351874 258630 351902 262927
rect 352342 262911 352394 262917
rect 352342 262853 352394 262859
rect 352354 258630 352382 262853
rect 352450 260253 352478 275650
rect 353698 265581 353726 275650
rect 353686 265575 353738 265581
rect 353686 265517 353738 265523
rect 354550 265427 354602 265433
rect 354550 265369 354602 265375
rect 353398 263503 353450 263509
rect 353398 263445 353450 263451
rect 352822 262171 352874 262177
rect 352822 262113 352874 262119
rect 352438 260247 352490 260253
rect 352438 260189 352490 260195
rect 352834 258630 352862 262113
rect 353410 258644 353438 263445
rect 353878 263429 353930 263435
rect 353878 263371 353930 263377
rect 353890 258644 353918 263371
rect 354070 263059 354122 263065
rect 354070 263001 354122 263007
rect 353184 258616 353438 258644
rect 353664 258616 353918 258644
rect 354082 258630 354110 263001
rect 354562 258630 354590 265369
rect 354850 263361 354878 275650
rect 356098 271871 356126 275650
rect 356086 271865 356138 271871
rect 356086 271807 356138 271813
rect 356278 271791 356330 271797
rect 356278 271733 356330 271739
rect 356086 265871 356138 265877
rect 356086 265813 356138 265819
rect 355606 265649 355658 265655
rect 355606 265591 355658 265597
rect 354934 265575 354986 265581
rect 354934 265517 354986 265523
rect 354838 263355 354890 263361
rect 354838 263297 354890 263303
rect 354946 258630 354974 265517
rect 355030 263355 355082 263361
rect 355030 263297 355082 263303
rect 355042 262991 355070 263297
rect 355030 262985 355082 262991
rect 355030 262927 355082 262933
rect 355618 258644 355646 265591
rect 356098 258644 356126 265813
rect 355392 258616 355646 258644
rect 355872 258616 356126 258644
rect 356290 258630 356318 271733
rect 356770 270613 357086 270632
rect 356770 270607 357098 270613
rect 356770 270604 357046 270607
rect 356770 269947 356798 270604
rect 357046 270549 357098 270555
rect 356866 270465 357086 270484
rect 356866 270459 357098 270465
rect 356866 270456 357046 270459
rect 356758 269941 356810 269947
rect 356758 269883 356810 269889
rect 356866 268615 356894 270456
rect 357046 270401 357098 270407
rect 357046 270311 357098 270317
rect 357046 270253 357098 270259
rect 357058 270188 357086 270253
rect 356962 270160 357086 270188
rect 356962 268689 356990 270160
rect 357046 269941 357098 269947
rect 357046 269883 357098 269889
rect 357058 268911 357086 269883
rect 357046 268905 357098 268911
rect 357046 268847 357098 268853
rect 356950 268683 357002 268689
rect 356950 268625 357002 268631
rect 356854 268609 356906 268615
rect 356854 268551 356906 268557
rect 357250 265729 357278 275650
rect 358114 268837 358142 275784
rect 358294 273863 358346 273869
rect 358294 273805 358346 273811
rect 358102 268831 358154 268837
rect 358102 268773 358154 268779
rect 357238 265723 357290 265729
rect 357238 265665 357290 265671
rect 357142 265353 357194 265359
rect 357142 265295 357194 265301
rect 357046 262097 357098 262103
rect 357046 262039 357098 262045
rect 357058 258644 357086 262039
rect 356688 258616 357086 258644
rect 357154 258630 357182 265295
rect 357814 263281 357866 263287
rect 357814 263223 357866 263229
rect 357826 258644 357854 263223
rect 358306 258644 358334 273805
rect 358390 273715 358442 273721
rect 358390 273657 358442 273663
rect 357600 258616 357854 258644
rect 358080 258616 358334 258644
rect 358402 258630 358430 273657
rect 358870 265279 358922 265285
rect 358870 265221 358922 265227
rect 358882 258630 358910 265221
rect 359350 262245 359402 262251
rect 359350 262187 359402 262193
rect 359362 258630 359390 262187
rect 359650 260401 359678 275650
rect 360598 267943 360650 267949
rect 360598 267885 360650 267891
rect 359926 267869 359978 267875
rect 359926 267811 359978 267817
rect 359638 260395 359690 260401
rect 359638 260337 359690 260343
rect 359938 258644 359966 267811
rect 360406 262467 360458 262473
rect 360406 262409 360458 262415
rect 360418 258644 360446 262409
rect 359808 258616 359966 258644
rect 360192 258616 360446 258644
rect 360610 258630 360638 267885
rect 360802 265803 360830 275650
rect 361462 268017 361514 268023
rect 361462 267959 361514 267965
rect 360790 265797 360842 265803
rect 360790 265739 360842 265745
rect 361078 262615 361130 262621
rect 361078 262557 361130 262563
rect 361090 258630 361118 262557
rect 361474 258630 361502 267959
rect 362050 263139 362078 275650
rect 363202 272019 363230 275650
rect 363190 272013 363242 272019
rect 363190 271955 363242 271961
rect 362806 271569 362858 271575
rect 362806 271511 362858 271517
rect 362614 268091 362666 268097
rect 362614 268033 362666 268039
rect 362134 265797 362186 265803
rect 362134 265739 362186 265745
rect 362038 263133 362090 263139
rect 362038 263075 362090 263081
rect 362146 263065 362174 265739
rect 362134 263059 362186 263065
rect 362134 263001 362186 263007
rect 362134 262689 362186 262695
rect 362134 262631 362186 262637
rect 362146 258644 362174 262631
rect 362626 258644 362654 268033
rect 362818 262917 362846 271511
rect 364342 268239 364394 268245
rect 364342 268181 364394 268187
rect 363190 268165 363242 268171
rect 363190 268107 363242 268113
rect 362806 262911 362858 262917
rect 362806 262853 362858 262859
rect 362710 262763 362762 262769
rect 362710 262705 362762 262711
rect 361920 258616 362174 258644
rect 362400 258616 362654 258644
rect 362722 258644 362750 262705
rect 362806 262171 362858 262177
rect 362806 262113 362858 262119
rect 362818 261955 362846 262113
rect 362806 261949 362858 261955
rect 362806 261891 362858 261897
rect 362722 258616 362832 258644
rect 363202 258630 363230 268107
rect 363670 262837 363722 262843
rect 363670 262779 363722 262785
rect 363682 258630 363710 262779
rect 364354 258644 364382 268181
rect 364450 259513 364478 275650
rect 364630 272013 364682 272019
rect 364630 271955 364682 271961
rect 364642 263287 364670 271955
rect 365602 268763 365630 275650
rect 365590 268757 365642 268763
rect 365590 268699 365642 268705
rect 365878 268387 365930 268393
rect 365878 268329 365930 268335
rect 365206 268313 365258 268319
rect 365206 268255 365258 268261
rect 364630 263281 364682 263287
rect 364630 263223 364682 263229
rect 364822 262911 364874 262917
rect 364822 262853 364874 262859
rect 364438 259507 364490 259513
rect 364438 259449 364490 259455
rect 364834 258644 364862 262853
rect 365218 258644 365246 268255
rect 365686 265057 365738 265063
rect 365686 264999 365738 265005
rect 365698 263361 365726 264999
rect 365686 263355 365738 263361
rect 365686 263297 365738 263303
rect 365398 262985 365450 262991
rect 365398 262927 365450 262933
rect 364128 258616 364382 258644
rect 364608 258616 364862 258644
rect 364992 258616 365246 258644
rect 365410 258630 365438 262927
rect 365890 258630 365918 268329
rect 366550 263059 366602 263065
rect 366550 263001 366602 263007
rect 366562 258644 366590 263001
rect 366754 260549 366782 275650
rect 367906 271205 367934 275650
rect 367894 271199 367946 271205
rect 367894 271141 367946 271147
rect 367990 269719 368042 269725
rect 367990 269661 368042 269667
rect 367606 268535 367658 268541
rect 367606 268477 367658 268483
rect 366934 268461 366986 268467
rect 366934 268403 366986 268409
rect 366742 260543 366794 260549
rect 366742 260485 366794 260491
rect 366946 258644 366974 268403
rect 367222 265501 367274 265507
rect 367222 265443 367274 265449
rect 367126 265205 367178 265211
rect 367126 265147 367178 265153
rect 367138 263509 367166 265147
rect 367126 263503 367178 263509
rect 367126 263445 367178 263451
rect 367234 263435 367262 265443
rect 367222 263429 367274 263435
rect 367222 263371 367274 263377
rect 367414 263133 367466 263139
rect 367414 263075 367466 263081
rect 367426 258644 367454 263075
rect 366336 258616 366590 258644
rect 366720 258616 366974 258644
rect 367200 258616 367454 258644
rect 367618 258630 367646 268477
rect 368002 262959 368030 269661
rect 368470 268609 368522 268615
rect 368470 268551 368522 268557
rect 367988 262950 368044 262959
rect 367988 262885 368044 262894
rect 367990 262541 368042 262547
rect 367990 262483 368042 262489
rect 368002 258630 368030 262483
rect 368482 258630 368510 268551
rect 369154 264989 369182 275650
rect 370306 273573 370334 275650
rect 370294 273567 370346 273573
rect 370294 273509 370346 273515
rect 371350 268831 371402 268837
rect 371350 268773 371402 268779
rect 370198 268757 370250 268763
rect 370198 268699 370250 268705
rect 369622 265131 369674 265137
rect 369622 265073 369674 265079
rect 369142 264983 369194 264989
rect 369142 264925 369194 264931
rect 369142 263281 369194 263287
rect 369142 263223 369194 263229
rect 369154 258644 369182 263223
rect 369634 258644 369662 265073
rect 369718 263355 369770 263361
rect 369718 263297 369770 263303
rect 368928 258616 369182 258644
rect 369408 258616 369662 258644
rect 369730 258630 369758 263297
rect 370210 258630 370238 268699
rect 370678 263429 370730 263435
rect 370678 263371 370730 263377
rect 370690 258630 370718 263371
rect 371362 258644 371390 268773
rect 371446 263503 371498 263509
rect 371446 263445 371498 263451
rect 371136 258616 371390 258644
rect 371458 258644 371486 263445
rect 371554 259587 371582 275650
rect 372706 270687 372734 275650
rect 372694 270681 372746 270687
rect 372694 270623 372746 270629
rect 371926 268905 371978 268911
rect 371926 268847 371978 268853
rect 371542 259581 371594 259587
rect 371542 259523 371594 259529
rect 371458 258616 371520 258644
rect 371938 258630 371966 268847
rect 373174 268683 373226 268689
rect 373174 268625 373226 268631
rect 372886 266315 372938 266321
rect 372886 266257 372938 266263
rect 372406 264983 372458 264989
rect 372406 264925 372458 264931
rect 372418 258630 372446 264925
rect 372898 258630 372926 266257
rect 373186 265137 373214 268625
rect 373462 265723 373514 265729
rect 373462 265665 373514 265671
rect 373174 265131 373226 265137
rect 373174 265073 373226 265079
rect 373474 258644 373502 265665
rect 373570 261511 373598 275784
rect 374134 271865 374186 271871
rect 374134 271807 374186 271813
rect 373558 261505 373610 261511
rect 373558 261447 373610 261453
rect 373942 260395 373994 260401
rect 373942 260337 373994 260343
rect 373954 258644 373982 260337
rect 373248 258616 373502 258644
rect 373728 258616 373982 258644
rect 374146 258630 374174 271807
rect 375106 271057 375134 275650
rect 375670 273567 375722 273573
rect 375670 273509 375722 273515
rect 375094 271051 375146 271057
rect 375094 270993 375146 270999
rect 374422 270681 374474 270687
rect 374422 270623 374474 270629
rect 374434 265285 374462 270623
rect 374422 265279 374474 265285
rect 374422 265221 374474 265227
rect 374998 265279 375050 265285
rect 374998 265221 375050 265227
rect 374614 261505 374666 261511
rect 374614 261447 374666 261453
rect 374626 258630 374654 261447
rect 375010 258630 375038 265221
rect 375682 258644 375710 273509
rect 375970 262325 375998 275784
rect 377506 273499 377534 275650
rect 377494 273493 377546 273499
rect 377494 273435 377546 273441
rect 378454 271421 378506 271427
rect 378454 271363 378506 271369
rect 376246 271273 376298 271279
rect 376246 271215 376298 271221
rect 376054 269349 376106 269355
rect 376054 269291 376106 269297
rect 376066 262325 376094 269291
rect 375958 262319 376010 262325
rect 375958 262261 376010 262267
rect 376054 262319 376106 262325
rect 376054 262261 376106 262267
rect 376150 260247 376202 260253
rect 376150 260189 376202 260195
rect 376162 258644 376190 260189
rect 375456 258616 375710 258644
rect 375936 258616 376190 258644
rect 376258 258630 376286 271215
rect 377206 271199 377258 271205
rect 377206 271141 377258 271147
rect 376726 260173 376778 260179
rect 376726 260115 376778 260121
rect 376738 258630 376766 260115
rect 377218 258630 377246 271141
rect 377878 265131 377930 265137
rect 377878 265073 377930 265079
rect 377890 258644 377918 265073
rect 378262 260025 378314 260031
rect 378262 259967 378314 259973
rect 378274 258644 378302 259967
rect 377664 258616 377918 258644
rect 378048 258616 378302 258644
rect 378466 258630 378494 271363
rect 378658 259661 378686 275650
rect 379414 271051 379466 271057
rect 379414 270993 379466 270999
rect 378934 260543 378986 260549
rect 378934 260485 378986 260491
rect 378646 259655 378698 259661
rect 378646 259597 378698 259603
rect 378946 258630 378974 260485
rect 379426 258630 379454 270993
rect 379906 265063 379934 275650
rect 380662 273493 380714 273499
rect 380662 273435 380714 273441
rect 380386 270456 380606 270484
rect 380386 270317 380414 270456
rect 380374 270311 380426 270317
rect 380374 270253 380426 270259
rect 380470 270311 380522 270317
rect 380470 270253 380522 270259
rect 380182 270015 380234 270021
rect 380182 269957 380234 269963
rect 380086 269941 380138 269947
rect 380086 269883 380138 269889
rect 380098 269725 380126 269883
rect 380086 269719 380138 269725
rect 380086 269661 380138 269667
rect 380194 269355 380222 269957
rect 380182 269349 380234 269355
rect 380182 269291 380234 269297
rect 380482 269133 380510 270253
rect 380578 269873 380606 270456
rect 380566 269867 380618 269873
rect 380566 269809 380618 269815
rect 380470 269127 380522 269133
rect 380470 269069 380522 269075
rect 380084 265318 380140 265327
rect 380084 265253 380140 265262
rect 380098 265137 380126 265253
rect 380086 265131 380138 265137
rect 380086 265073 380138 265079
rect 380470 265131 380522 265137
rect 380470 265073 380522 265079
rect 379894 265057 379946 265063
rect 379894 264999 379946 265005
rect 379990 259877 380042 259883
rect 379990 259819 380042 259825
rect 380002 258644 380030 259819
rect 380482 258644 380510 265073
rect 379776 258616 380030 258644
rect 380256 258616 380510 258644
rect 380674 258630 380702 273435
rect 381058 260623 381086 275650
rect 382306 271131 382334 275650
rect 383362 271575 383390 275650
rect 384610 273425 384638 275650
rect 385570 275636 385776 275664
rect 384598 273419 384650 273425
rect 384598 273361 384650 273367
rect 383350 271569 383402 271575
rect 383350 271511 383402 271517
rect 382294 271125 382346 271131
rect 382294 271067 382346 271073
rect 382198 270755 382250 270761
rect 382198 270697 382250 270703
rect 381142 265057 381194 265063
rect 381142 264999 381194 265005
rect 381046 260617 381098 260623
rect 381046 260559 381098 260565
rect 381154 258630 381182 264999
rect 381526 260617 381578 260623
rect 381526 260559 381578 260565
rect 381538 258630 381566 260559
rect 382210 258644 382238 270697
rect 382294 269941 382346 269947
rect 382294 269883 382346 269889
rect 382306 265359 382334 269883
rect 383158 269793 383210 269799
rect 383158 269735 383210 269741
rect 383254 269793 383306 269799
rect 383254 269735 383306 269741
rect 382774 269719 382826 269725
rect 382774 269661 382826 269667
rect 382870 269719 382922 269725
rect 382870 269661 382922 269667
rect 382786 269133 382814 269661
rect 382774 269127 382826 269133
rect 382774 269069 382826 269075
rect 382294 265353 382346 265359
rect 382390 265353 382442 265359
rect 382294 265295 382346 265301
rect 382388 265318 382390 265327
rect 382442 265318 382444 265327
rect 382388 265253 382444 265262
rect 382580 262210 382636 262219
rect 382580 262145 382636 262154
rect 382594 262029 382622 262145
rect 382582 262023 382634 262029
rect 382582 261965 382634 261971
rect 382678 262023 382730 262029
rect 382678 261965 382730 261971
rect 382690 258644 382718 261965
rect 381984 258616 382238 258644
rect 382464 258616 382718 258644
rect 382882 258630 382910 269661
rect 382966 269423 383018 269429
rect 382966 269365 383018 269371
rect 382978 262177 383006 269365
rect 383170 269355 383198 269735
rect 383158 269349 383210 269355
rect 383158 269291 383210 269297
rect 382966 262171 383018 262177
rect 382966 262113 383018 262119
rect 383266 258630 383294 269735
rect 383638 269423 383690 269429
rect 383638 269365 383690 269371
rect 383734 269423 383786 269429
rect 383734 269365 383786 269371
rect 383650 268583 383678 269365
rect 383636 268574 383692 268583
rect 383636 268509 383692 268518
rect 383746 258630 383774 269365
rect 384788 269018 384844 269027
rect 384788 268953 384844 268962
rect 384406 262245 384458 262251
rect 384406 262187 384458 262193
rect 384418 258644 384446 262187
rect 384802 258644 384830 268953
rect 385460 262802 385516 262811
rect 385460 262737 385516 262746
rect 384982 262319 385034 262325
rect 384982 262261 385034 262267
rect 384192 258616 384446 258644
rect 384576 258616 384830 258644
rect 384994 258630 385022 262261
rect 385474 258630 385502 262737
rect 385570 259735 385598 275636
rect 386038 269571 386090 269577
rect 386038 269513 386090 269519
rect 385654 269497 385706 269503
rect 385654 269439 385706 269445
rect 385666 262325 385694 269439
rect 385942 269349 385994 269355
rect 385942 269291 385994 269297
rect 385750 269275 385802 269281
rect 385750 269217 385802 269223
rect 385654 262319 385706 262325
rect 385654 262261 385706 262267
rect 385762 262048 385790 269217
rect 385954 265008 385982 269291
rect 386050 265063 386078 269513
rect 386132 269462 386188 269471
rect 386132 269397 386188 269406
rect 385858 264980 385982 265008
rect 386038 265057 386090 265063
rect 386038 264999 386090 265005
rect 385858 262251 385886 264980
rect 386146 262251 386174 269397
rect 385846 262245 385898 262251
rect 385846 262187 385898 262193
rect 386134 262245 386186 262251
rect 386134 262187 386186 262193
rect 385762 262020 385982 262048
rect 385558 259729 385610 259735
rect 385558 259671 385610 259677
rect 385954 258630 385982 262020
rect 386338 258496 386366 276099
rect 396790 276083 396842 276089
rect 396790 276025 396842 276031
rect 389026 275784 389328 275812
rect 386722 275636 387024 275664
rect 386516 262950 386572 262959
rect 386516 262885 386572 262894
rect 386530 258644 386558 262885
rect 386722 262219 386750 275636
rect 387490 271945 387710 271964
rect 387478 271939 387722 271945
rect 387530 271936 387670 271939
rect 387478 271881 387530 271887
rect 387670 271881 387722 271887
rect 387382 271865 387434 271871
rect 387382 271807 387434 271813
rect 387286 271569 387338 271575
rect 387286 271511 387338 271517
rect 387298 271205 387326 271511
rect 387394 271205 387422 271807
rect 387286 271199 387338 271205
rect 387286 271141 387338 271147
rect 387382 271199 387434 271205
rect 387382 271141 387434 271147
rect 387106 270752 387422 270780
rect 387106 270021 387134 270752
rect 387394 270687 387422 270752
rect 387286 270681 387338 270687
rect 387286 270623 387338 270629
rect 387382 270681 387434 270687
rect 387382 270623 387434 270629
rect 387298 270465 387326 270623
rect 387190 270459 387242 270465
rect 387190 270401 387242 270407
rect 387286 270459 387338 270465
rect 387286 270401 387338 270407
rect 387202 270188 387230 270401
rect 387202 270160 387422 270188
rect 387094 270015 387146 270021
rect 387094 269957 387146 269963
rect 387286 270015 387338 270021
rect 387286 269957 387338 269963
rect 387298 268985 387326 269957
rect 387394 268985 387422 270160
rect 387668 269314 387724 269323
rect 387668 269249 387724 269258
rect 387286 268979 387338 268985
rect 387286 268921 387338 268927
rect 387382 268979 387434 268985
rect 387382 268921 387434 268927
rect 387190 263577 387242 263583
rect 387190 263519 387242 263525
rect 386708 262210 386764 262219
rect 386708 262145 386764 262154
rect 386530 258616 386784 258644
rect 387202 258630 387230 263519
rect 387682 258630 387710 269249
rect 388054 262171 388106 262177
rect 388054 262113 388106 262119
rect 388066 258630 388094 262113
rect 388162 259291 388190 275650
rect 389026 270983 389054 275784
rect 389014 270977 389066 270983
rect 389014 270919 389066 270925
rect 390358 270681 390410 270687
rect 390358 270623 390410 270629
rect 389012 270054 389068 270063
rect 389012 269989 389068 269998
rect 388822 269867 388874 269873
rect 388822 269809 388874 269815
rect 388630 269645 388682 269651
rect 388630 269587 388682 269593
rect 388532 269314 388588 269323
rect 388532 269249 388588 269258
rect 388546 269133 388574 269249
rect 388534 269127 388586 269133
rect 388534 269069 388586 269075
rect 388642 262325 388670 269587
rect 388834 269503 388862 269809
rect 388918 269645 388970 269651
rect 388918 269587 388970 269593
rect 388726 269497 388778 269503
rect 388726 269439 388778 269445
rect 388822 269497 388874 269503
rect 388822 269439 388874 269445
rect 388738 263583 388766 269439
rect 388822 269127 388874 269133
rect 388822 269069 388874 269075
rect 388834 266025 388862 269069
rect 388822 266019 388874 266025
rect 388822 265961 388874 265967
rect 388930 265137 388958 269587
rect 388918 265131 388970 265137
rect 388918 265073 388970 265079
rect 388820 263838 388876 263847
rect 388820 263773 388876 263782
rect 388726 263577 388778 263583
rect 388726 263519 388778 263525
rect 388246 262319 388298 262325
rect 388246 262261 388298 262267
rect 388630 262319 388682 262325
rect 388630 262261 388682 262267
rect 388150 259285 388202 259291
rect 388150 259227 388202 259233
rect 388258 258644 388286 262261
rect 388834 258644 388862 263773
rect 389026 262177 389054 269989
rect 389396 264134 389452 264143
rect 389396 264069 389452 264078
rect 389014 262171 389066 262177
rect 389014 262113 389066 262119
rect 388258 258616 388512 258644
rect 388834 258616 388992 258644
rect 389410 258630 389438 264069
rect 389780 263986 389836 263995
rect 389780 263921 389836 263930
rect 389794 258630 389822 263921
rect 390370 263583 390398 270623
rect 390562 265211 390590 275650
rect 391714 273351 391742 275650
rect 391702 273345 391754 273351
rect 391702 273287 391754 273293
rect 392180 270646 392236 270655
rect 392180 270581 392236 270590
rect 390644 270350 390700 270359
rect 390644 270285 390700 270294
rect 390550 265205 390602 265211
rect 390550 265147 390602 265153
rect 390262 263577 390314 263583
rect 390262 263519 390314 263525
rect 390358 263577 390410 263583
rect 390358 263519 390410 263525
rect 390274 258630 390302 263519
rect 390658 262251 390686 270285
rect 391702 269867 391754 269873
rect 391702 269809 391754 269815
rect 391604 269758 391660 269767
rect 391604 269693 391660 269702
rect 391414 269275 391466 269281
rect 391414 269217 391466 269223
rect 391426 262325 391454 269217
rect 391618 264860 391646 269693
rect 391714 265359 391742 269809
rect 391796 269314 391852 269323
rect 391796 269249 391798 269258
rect 391850 269249 391852 269258
rect 391798 269217 391850 269223
rect 391702 265353 391754 265359
rect 391702 265295 391754 265301
rect 391618 264832 392126 264860
rect 391988 264282 392044 264291
rect 391988 264217 392044 264226
rect 391510 263651 391562 263657
rect 391510 263593 391562 263599
rect 390934 262319 390986 262325
rect 390934 262261 390986 262267
rect 391414 262319 391466 262325
rect 391414 262261 391466 262267
rect 390454 262245 390506 262251
rect 390454 262187 390506 262193
rect 390646 262245 390698 262251
rect 390646 262187 390698 262193
rect 390466 258644 390494 262187
rect 390946 258644 390974 262261
rect 390466 258616 390720 258644
rect 390946 258616 391200 258644
rect 391522 258630 391550 263593
rect 392002 258630 392030 264217
rect 392098 258644 392126 264832
rect 392194 264143 392222 270581
rect 392564 269610 392620 269619
rect 392564 269545 392620 269554
rect 392180 264134 392236 264143
rect 392180 264069 392236 264078
rect 392578 258644 392606 269545
rect 392962 259809 392990 275650
rect 393046 272013 393098 272019
rect 393046 271955 393098 271961
rect 393058 271871 393086 271955
rect 393046 271865 393098 271871
rect 393046 271807 393098 271813
rect 394114 265507 394142 275650
rect 395170 275636 395376 275664
rect 394774 271569 394826 271575
rect 394774 271511 394826 271517
rect 394786 271057 394814 271511
rect 394678 271051 394730 271057
rect 394678 270993 394730 270999
rect 394774 271051 394826 271057
rect 394774 270993 394826 270999
rect 394690 270761 394718 270993
rect 394678 270755 394730 270761
rect 394678 270697 394730 270703
rect 394870 270237 394922 270243
rect 394870 270179 394922 270185
rect 394594 269568 394814 269596
rect 394594 269503 394622 269568
rect 394582 269497 394634 269503
rect 394582 269439 394634 269445
rect 394678 269497 394730 269503
rect 394678 269439 394730 269445
rect 394486 269275 394538 269281
rect 394486 269217 394538 269223
rect 394582 269275 394634 269281
rect 394582 269217 394634 269223
rect 394102 265501 394154 265507
rect 394102 265443 394154 265449
rect 393044 264578 393100 264587
rect 393044 264513 393100 264522
rect 392950 259803 393002 259809
rect 392950 259745 393002 259751
rect 393058 258644 393086 264513
rect 393716 264430 393772 264439
rect 393716 264365 393772 264374
rect 392098 258616 392496 258644
rect 392578 258616 392832 258644
rect 393058 258616 393312 258644
rect 393730 258630 393758 264365
rect 394294 263577 394346 263583
rect 394294 263519 394346 263525
rect 394306 262177 394334 263519
rect 394498 262367 394526 269217
rect 394594 266099 394622 269217
rect 394582 266093 394634 266099
rect 394582 266035 394634 266041
rect 394484 262358 394540 262367
rect 394484 262293 394540 262302
rect 394198 262171 394250 262177
rect 394198 262113 394250 262119
rect 394294 262171 394346 262177
rect 394294 262113 394346 262119
rect 394210 258630 394238 262113
rect 394690 262029 394718 269439
rect 394786 266099 394814 269568
rect 394774 266093 394826 266099
rect 394774 266035 394826 266041
rect 394772 264726 394828 264735
rect 394772 264661 394828 264670
rect 394678 262023 394730 262029
rect 394678 261965 394730 261971
rect 394678 259803 394730 259809
rect 394678 259745 394730 259751
rect 394690 258644 394718 259745
rect 394608 258616 394718 258644
rect 394786 258644 394814 264661
rect 394882 263583 394910 270179
rect 395060 269906 395116 269915
rect 395060 269841 395116 269850
rect 394966 266093 395018 266099
rect 394966 266035 395018 266041
rect 394978 263657 395006 266035
rect 394966 263651 395018 263657
rect 394966 263593 395018 263599
rect 394870 263577 394922 263583
rect 394870 263519 394922 263525
rect 395074 259809 395102 269841
rect 395062 259803 395114 259809
rect 395062 259745 395114 259751
rect 395170 259365 395198 275636
rect 396514 271353 396542 275650
rect 396502 271347 396554 271353
rect 396502 271289 396554 271295
rect 395924 270202 395980 270211
rect 395924 270137 395980 270146
rect 395348 268574 395404 268583
rect 395348 268509 395404 268518
rect 395362 263731 395390 268509
rect 395254 263725 395306 263731
rect 395254 263667 395306 263673
rect 395350 263725 395402 263731
rect 395350 263667 395402 263673
rect 395158 259359 395210 259365
rect 395158 259301 395210 259307
rect 395266 258644 395294 263667
rect 394786 258616 395040 258644
rect 395266 258616 395520 258644
rect 395938 258630 395966 270137
rect 396502 263725 396554 263731
rect 396502 263667 396554 263673
rect 396310 262245 396362 262251
rect 396310 262187 396362 262193
rect 396322 258630 396350 262187
rect 396514 262177 396542 263667
rect 396502 262171 396554 262177
rect 396502 262113 396554 262119
rect 396802 258630 396830 276025
rect 397378 270752 397502 270780
rect 397378 270613 397406 270752
rect 397474 270613 397502 270752
rect 397366 270607 397418 270613
rect 397366 270549 397418 270555
rect 397462 270607 397514 270613
rect 397462 270549 397514 270555
rect 397076 262358 397132 262367
rect 396982 262319 397034 262325
rect 397076 262293 397078 262302
rect 396982 262261 397034 262267
rect 397130 262293 397132 262302
rect 397078 262261 397130 262267
rect 396994 258644 397022 262261
rect 397570 258644 397598 276247
rect 398518 276231 398570 276237
rect 398518 276173 398570 276179
rect 397762 265803 397790 275650
rect 397750 265797 397802 265803
rect 397750 265739 397802 265745
rect 397844 264874 397900 264883
rect 397844 264809 397900 264818
rect 397858 258644 397886 264809
rect 396994 258616 397248 258644
rect 397570 258616 397728 258644
rect 397858 258616 398112 258644
rect 398530 258630 398558 276173
rect 439030 276009 439082 276015
rect 439082 275957 439344 275960
rect 439030 275951 439344 275957
rect 439042 275932 439344 275951
rect 442594 275941 442896 275960
rect 442582 275935 442896 275941
rect 442634 275932 442896 275935
rect 442582 275877 442634 275883
rect 446326 275861 446378 275867
rect 404482 275784 404784 275812
rect 419938 275784 420240 275812
rect 446378 275809 446544 275812
rect 446326 275803 446544 275809
rect 446338 275784 446544 275803
rect 449698 275793 450000 275812
rect 449686 275787 450000 275793
rect 398914 273277 398942 275650
rect 398902 273271 398954 273277
rect 398902 273213 398954 273219
rect 398996 270498 399052 270507
rect 398996 270433 399052 270442
rect 398612 268870 398668 268879
rect 398612 268805 398668 268814
rect 398626 263731 398654 268805
rect 398614 263725 398666 263731
rect 398614 263667 398666 263673
rect 399010 258630 399038 270433
rect 399572 263394 399628 263403
rect 399572 263329 399628 263338
rect 399190 262393 399242 262399
rect 399190 262335 399242 262341
rect 399202 258644 399230 262335
rect 399586 258644 399614 263329
rect 400066 259957 400094 275650
rect 400342 270607 400394 270613
rect 400342 270549 400394 270555
rect 400246 270237 400298 270243
rect 400246 270179 400298 270185
rect 400150 268979 400202 268985
rect 400150 268921 400202 268927
rect 400162 262399 400190 268921
rect 400258 265285 400286 270179
rect 400246 265279 400298 265285
rect 400246 265221 400298 265227
rect 400150 262393 400202 262399
rect 400150 262335 400202 262341
rect 400354 262251 400382 270549
rect 401218 265433 401246 275650
rect 402166 270311 402218 270317
rect 402166 270253 402218 270259
rect 402358 270311 402410 270317
rect 402358 270253 402410 270259
rect 401206 265427 401258 265433
rect 401206 265369 401258 265375
rect 400724 264134 400780 264143
rect 400724 264069 400780 264078
rect 400150 262245 400202 262251
rect 400150 262187 400202 262193
rect 400342 262245 400394 262251
rect 400342 262187 400394 262193
rect 400054 259951 400106 259957
rect 400054 259893 400106 259899
rect 399202 258616 399456 258644
rect 399586 258616 399840 258644
rect 317952 258468 318014 258496
rect 386304 258468 386366 258496
rect 400162 258496 400190 262187
rect 400738 258630 400766 264069
rect 401590 263799 401642 263805
rect 401590 263741 401642 263747
rect 401108 263098 401164 263107
rect 401108 263033 401164 263042
rect 401122 258630 401150 263033
rect 401602 258630 401630 263741
rect 402178 262325 402206 270253
rect 402260 269166 402316 269175
rect 402260 269101 402316 269110
rect 401782 262319 401834 262325
rect 401782 262261 401834 262267
rect 402166 262319 402218 262325
rect 402166 262261 402218 262267
rect 401794 258644 401822 262261
rect 402274 258644 402302 269101
rect 402370 265729 402398 270253
rect 402358 265723 402410 265729
rect 402358 265665 402410 265671
rect 402466 261881 402494 275650
rect 403618 271649 403646 275650
rect 403606 271643 403658 271649
rect 403606 271585 403658 271591
rect 403126 270755 403178 270761
rect 403126 270697 403178 270703
rect 403138 270613 403166 270697
rect 403126 270607 403178 270613
rect 403126 270549 403178 270555
rect 403894 270163 403946 270169
rect 403894 270105 403946 270111
rect 403222 270089 403274 270095
rect 403222 270031 403274 270037
rect 403030 270015 403082 270021
rect 403030 269957 403082 269963
rect 403042 263805 403070 269957
rect 403234 265655 403262 270031
rect 403222 265649 403274 265655
rect 403222 265591 403274 265597
rect 403030 263799 403082 263805
rect 403030 263741 403082 263747
rect 403316 263246 403372 263255
rect 402838 263207 402890 263213
rect 403316 263181 403372 263190
rect 402838 263149 402890 263155
rect 402454 261875 402506 261881
rect 402454 261817 402506 261823
rect 401794 258616 402048 258644
rect 402274 258616 402528 258644
rect 402850 258630 402878 263149
rect 403330 258630 403358 263181
rect 403906 262177 403934 270105
rect 404482 265581 404510 275784
rect 406018 273203 406046 275650
rect 406006 273197 406058 273203
rect 406006 273139 406058 273145
rect 405910 270533 405962 270539
rect 405910 270475 405962 270481
rect 405718 270385 405770 270391
rect 405718 270327 405770 270333
rect 405142 270015 405194 270021
rect 405142 269957 405194 269963
rect 404470 265575 404522 265581
rect 404470 265517 404522 265523
rect 404374 263947 404426 263953
rect 404374 263889 404426 263895
rect 403990 263725 404042 263731
rect 403990 263667 404042 263673
rect 403798 262171 403850 262177
rect 403798 262113 403850 262119
rect 403894 262171 403946 262177
rect 403894 262113 403946 262119
rect 403810 258630 403838 262113
rect 404002 258644 404030 263667
rect 404386 258644 404414 263889
rect 405154 263879 405182 269957
rect 405622 269201 405674 269207
rect 405622 269143 405674 269149
rect 405526 264021 405578 264027
rect 405526 263963 405578 263969
rect 405046 263873 405098 263879
rect 405046 263815 405098 263821
rect 405142 263873 405194 263879
rect 405142 263815 405194 263821
rect 404002 258616 404256 258644
rect 404386 258616 404640 258644
rect 405058 258630 405086 263815
rect 405538 258630 405566 263963
rect 405634 263731 405662 269143
rect 405730 264027 405758 270327
rect 405814 269127 405866 269133
rect 405814 269069 405866 269075
rect 405718 264021 405770 264027
rect 405718 263963 405770 263969
rect 405622 263725 405674 263731
rect 405622 263667 405674 263673
rect 405826 259883 405854 269069
rect 405922 263953 405950 270475
rect 406102 270015 406154 270021
rect 406102 269957 406154 269963
rect 406114 265877 406142 269957
rect 406678 268979 406730 268985
rect 406678 268921 406730 268927
rect 406102 265871 406154 265877
rect 406102 265813 406154 265819
rect 406006 264095 406058 264101
rect 406006 264037 406058 264043
rect 405910 263947 405962 263953
rect 405910 263889 405962 263895
rect 405814 259877 405866 259883
rect 405814 259819 405866 259825
rect 406018 258630 406046 264037
rect 406582 263873 406634 263879
rect 406582 263815 406634 263821
rect 406102 263577 406154 263583
rect 406102 263519 406154 263525
rect 406114 258644 406142 263519
rect 406594 258644 406622 263815
rect 406690 263213 406718 268921
rect 406678 263207 406730 263213
rect 406678 263149 406730 263155
rect 407170 260105 407198 275650
rect 407350 271421 407402 271427
rect 407350 271363 407402 271369
rect 407362 270539 407390 271363
rect 407350 270533 407402 270539
rect 407350 270475 407402 270481
rect 408418 270095 408446 275650
rect 408982 270163 409034 270169
rect 408982 270105 409034 270111
rect 408406 270089 408458 270095
rect 408406 270031 408458 270037
rect 408994 269947 409022 270105
rect 409078 270015 409130 270021
rect 409078 269957 409130 269963
rect 408982 269941 409034 269947
rect 408982 269883 409034 269889
rect 407542 269793 407594 269799
rect 407542 269735 407594 269741
rect 407638 269793 407690 269799
rect 407638 269735 407690 269741
rect 407554 269429 407582 269735
rect 407542 269423 407594 269429
rect 407542 269365 407594 269371
rect 407650 269133 407678 269735
rect 407638 269127 407690 269133
rect 407638 269069 407690 269075
rect 408982 264317 409034 264323
rect 408982 264259 409034 264265
rect 407254 264243 407306 264249
rect 407254 264185 407306 264191
rect 407158 260099 407210 260105
rect 407158 260041 407210 260047
rect 406114 258616 406368 258644
rect 406594 258616 406848 258644
rect 407266 258630 407294 264185
rect 407734 264169 407786 264175
rect 407734 264111 407786 264117
rect 407746 258630 407774 264111
rect 408118 263651 408170 263657
rect 408118 263593 408170 263599
rect 408130 258630 408158 263593
rect 408310 262171 408362 262177
rect 408310 262113 408362 262119
rect 408322 258644 408350 262113
rect 408994 258644 409022 264259
rect 409090 260179 409118 269957
rect 409174 269941 409226 269947
rect 409174 269883 409226 269889
rect 409078 260173 409130 260179
rect 409078 260115 409130 260121
rect 409186 260031 409214 269883
rect 409366 264391 409418 264397
rect 409366 264333 409418 264339
rect 409174 260025 409226 260031
rect 409174 259967 409226 259973
rect 408322 258616 408576 258644
rect 408994 258616 409056 258644
rect 409378 258630 409406 264333
rect 409570 261807 409598 275650
rect 410818 271723 410846 275650
rect 410806 271717 410858 271723
rect 410806 271659 410858 271665
rect 411970 270095 411998 275650
rect 413218 273129 413246 275650
rect 413206 273123 413258 273129
rect 413206 273065 413258 273071
rect 411958 270089 412010 270095
rect 411958 270031 412010 270037
rect 414370 265951 414398 275650
rect 415618 271797 415646 275650
rect 415606 271791 415658 271797
rect 415606 271733 415658 271739
rect 414358 265945 414410 265951
rect 414358 265887 414410 265893
rect 415318 264909 415370 264915
rect 415318 264851 415370 264857
rect 414838 264761 414890 264767
rect 414838 264703 414890 264709
rect 412630 264687 412682 264693
rect 412630 264629 412682 264635
rect 412534 264613 412586 264619
rect 412534 264555 412586 264561
rect 410902 264539 410954 264545
rect 410902 264481 410954 264487
rect 410518 264465 410570 264471
rect 410518 264407 410570 264413
rect 410326 264021 410378 264027
rect 410326 263963 410378 263969
rect 409846 262393 409898 262399
rect 409846 262335 409898 262341
rect 409558 261801 409610 261807
rect 409558 261743 409610 261749
rect 409858 258630 409886 262335
rect 410338 258630 410366 263963
rect 410530 258644 410558 264407
rect 410914 258644 410942 264481
rect 412054 263947 412106 263953
rect 412054 263889 412106 263895
rect 411574 262245 411626 262251
rect 411574 262187 411626 262193
rect 410530 258616 410784 258644
rect 410914 258616 411168 258644
rect 411586 258630 411614 262187
rect 412066 258630 412094 263889
rect 412546 258630 412574 264555
rect 412642 258644 412670 264629
rect 414262 263799 414314 263805
rect 414262 263741 414314 263747
rect 413782 263725 413834 263731
rect 413782 263667 413834 263673
rect 413110 262319 413162 262325
rect 413110 262261 413162 262267
rect 413122 258644 413150 262261
rect 412642 258616 412896 258644
rect 413122 258616 413376 258644
rect 413794 258630 413822 263667
rect 414274 258630 414302 263741
rect 414646 263207 414698 263213
rect 414646 263149 414698 263155
rect 414658 258630 414686 263149
rect 414850 258644 414878 264703
rect 415330 258644 415358 264851
rect 416674 261733 416702 275650
rect 416662 261727 416714 261733
rect 416662 261669 416714 261675
rect 417922 260327 417950 275650
rect 419074 261955 419102 275650
rect 419938 273055 419966 275784
rect 449738 275784 450000 275787
rect 450850 275784 451152 275812
rect 453250 275784 453552 275812
rect 455650 275784 455952 275812
rect 466704 275784 466814 275812
rect 449686 275729 449738 275735
rect 419926 273049 419978 273055
rect 419926 272991 419978 272997
rect 421474 271945 421502 275650
rect 421846 275639 421898 275645
rect 421846 275581 421898 275587
rect 421462 271939 421514 271945
rect 421462 271881 421514 271887
rect 419062 261949 419114 261955
rect 419062 261891 419114 261897
rect 417910 260321 417962 260327
rect 417910 260263 417962 260269
rect 414850 258616 415104 258644
rect 415330 258616 415584 258644
rect 400162 258468 400320 258496
rect 210164 256438 210220 256447
rect 210164 256373 210220 256382
rect 198742 250627 198794 250633
rect 198742 250569 198794 250575
rect 207286 250553 207338 250559
rect 207286 250495 207338 250501
rect 204982 246557 205034 246563
rect 204982 246499 205034 246505
rect 204886 246483 204938 246489
rect 204886 246425 204938 246431
rect 204502 246409 204554 246415
rect 204502 246351 204554 246357
rect 204514 244935 204542 246351
rect 204790 246261 204842 246267
rect 204790 246203 204842 246209
rect 204502 244929 204554 244935
rect 204502 244871 204554 244877
rect 204694 243893 204746 243899
rect 204694 243835 204746 243841
rect 204598 243819 204650 243825
rect 204598 243761 204650 243767
rect 204502 243671 204554 243677
rect 204502 243613 204554 243619
rect 204514 233169 204542 243613
rect 204502 233163 204554 233169
rect 204502 233105 204554 233111
rect 204610 232799 204638 243761
rect 204706 233095 204734 243835
rect 204694 233089 204746 233095
rect 204694 233031 204746 233037
rect 204598 232793 204650 232799
rect 204598 232735 204650 232741
rect 204802 230547 204830 246203
rect 204788 230538 204844 230547
rect 204788 230473 204844 230482
rect 201814 230425 201866 230431
rect 201814 230367 201866 230373
rect 201622 230351 201674 230357
rect 201622 230293 201674 230299
rect 201634 228475 201662 230293
rect 201718 230203 201770 230209
rect 201718 230145 201770 230151
rect 201730 229511 201758 230145
rect 201716 229502 201772 229511
rect 201716 229437 201772 229446
rect 201620 228466 201676 228475
rect 201620 228401 201676 228410
rect 201826 227883 201854 230367
rect 204898 230103 204926 246425
rect 204994 233243 205022 246499
rect 207190 246335 207242 246341
rect 207190 246277 207242 246283
rect 205174 244929 205226 244935
rect 205174 244871 205226 244877
rect 204982 233237 205034 233243
rect 204982 233179 205034 233185
rect 204884 230094 204940 230103
rect 204884 230029 204940 230038
rect 201812 227874 201868 227883
rect 201812 227809 201868 227818
rect 194326 227687 194378 227693
rect 194326 227629 194378 227635
rect 192886 215625 192938 215631
rect 192886 215567 192938 215573
rect 191446 198753 191498 198759
rect 191446 198695 191498 198701
rect 188662 175739 188714 175745
rect 188662 175681 188714 175687
rect 188674 89017 188702 175681
rect 188758 112543 188810 112549
rect 188758 112485 188810 112491
rect 188662 89011 188714 89017
rect 188662 88953 188714 88959
rect 188770 77399 188798 112485
rect 188758 77393 188810 77399
rect 188758 77335 188810 77341
rect 191458 48539 191486 198695
rect 191542 178625 191594 178631
rect 191542 178567 191594 178573
rect 191554 88943 191582 178567
rect 191638 118611 191690 118617
rect 191638 118553 191690 118559
rect 191542 88937 191594 88943
rect 191542 88879 191594 88885
rect 191650 80581 191678 118553
rect 193942 106623 193994 106629
rect 193942 106565 193994 106571
rect 193954 94123 193982 106565
rect 193942 94117 193994 94123
rect 193942 94059 193994 94065
rect 191638 80575 191690 80581
rect 191638 80517 191690 80523
rect 193750 64813 193802 64819
rect 193750 64755 193802 64761
rect 193762 64195 193790 64755
rect 193748 64186 193804 64195
rect 193748 64121 193804 64130
rect 194132 62558 194188 62567
rect 194132 62493 194188 62502
rect 194146 60749 194174 62493
rect 194134 60743 194186 60749
rect 194134 60685 194186 60691
rect 191446 48533 191498 48539
rect 191446 48475 191498 48481
rect 188564 48202 188620 48211
rect 188564 48137 188620 48146
rect 194338 48063 194366 227629
rect 197206 227613 197258 227619
rect 197206 227555 197258 227561
rect 194422 187283 194474 187289
rect 194422 187225 194474 187231
rect 194434 90835 194462 187225
rect 194518 124013 194570 124019
rect 194518 123955 194570 123961
rect 194420 90826 194476 90835
rect 194420 90761 194476 90770
rect 194530 79735 194558 123955
rect 194614 83535 194666 83541
rect 194614 83477 194666 83483
rect 194626 81363 194654 83477
rect 194612 81354 194668 81363
rect 194612 81289 194668 81298
rect 194516 79726 194572 79735
rect 194516 79661 194572 79670
rect 195574 77615 195626 77621
rect 195574 77557 195626 77563
rect 195586 76479 195614 77557
rect 195572 76470 195628 76479
rect 195572 76405 195628 76414
rect 194708 69070 194764 69079
rect 194708 69005 194764 69014
rect 194722 68815 194750 69005
rect 194710 68809 194762 68815
rect 194710 68751 194762 68757
rect 194324 48054 194380 48063
rect 194324 47989 194380 47998
rect 197218 46911 197246 227555
rect 201814 227539 201866 227545
rect 201814 227481 201866 227487
rect 197590 227465 197642 227471
rect 197590 227407 197642 227413
rect 197602 225663 197630 227407
rect 201718 227391 201770 227397
rect 201718 227333 201770 227339
rect 201526 227317 201578 227323
rect 201730 227291 201758 227333
rect 201526 227259 201578 227265
rect 201716 227282 201772 227291
rect 197588 225654 197644 225663
rect 197588 225589 197644 225598
rect 201538 225219 201566 227259
rect 201622 227243 201674 227249
rect 201716 227217 201772 227226
rect 201622 227185 201674 227191
rect 201634 226255 201662 227185
rect 201826 226847 201854 227481
rect 201812 226838 201868 226847
rect 201812 226773 201868 226782
rect 201620 226246 201676 226255
rect 201620 226181 201676 226190
rect 201524 225210 201580 225219
rect 201524 225145 201580 225154
rect 201526 224653 201578 224659
rect 201526 224595 201578 224601
rect 201716 224618 201772 224627
rect 201538 222407 201566 224595
rect 201716 224553 201718 224562
rect 201770 224553 201772 224562
rect 201718 224521 201770 224527
rect 201622 224505 201674 224511
rect 201622 224447 201674 224453
rect 201634 224035 201662 224447
rect 201718 224431 201770 224437
rect 201718 224373 201770 224379
rect 201620 224026 201676 224035
rect 201620 223961 201676 223970
rect 201730 223591 201758 224373
rect 201814 224357 201866 224363
rect 201814 224299 201866 224305
rect 201716 223582 201772 223591
rect 201716 223517 201772 223526
rect 201826 222999 201854 224299
rect 201812 222990 201868 222999
rect 201812 222925 201868 222934
rect 201524 222398 201580 222407
rect 201524 222333 201580 222342
rect 202966 221841 203018 221847
rect 202966 221783 203018 221789
rect 198646 221767 198698 221773
rect 198646 221709 198698 221715
rect 198658 221371 198686 221709
rect 201718 221693 201770 221699
rect 201718 221635 201770 221641
rect 201622 221545 201674 221551
rect 201622 221487 201674 221493
rect 198644 221362 198700 221371
rect 198644 221297 198700 221306
rect 201634 219743 201662 221487
rect 201730 220779 201758 221635
rect 201814 221471 201866 221477
rect 201814 221413 201866 221419
rect 201716 220770 201772 220779
rect 201716 220705 201772 220714
rect 201620 219734 201676 219743
rect 201620 219669 201676 219678
rect 201826 219151 201854 221413
rect 201812 219142 201868 219151
rect 201812 219077 201868 219086
rect 197590 218881 197642 218887
rect 197590 218823 197642 218829
rect 197602 216487 197630 218823
rect 201718 218733 201770 218739
rect 201718 218675 201770 218681
rect 198166 218659 198218 218665
rect 198166 218601 198218 218607
rect 198178 217523 198206 218601
rect 201730 218115 201758 218675
rect 201716 218106 201772 218115
rect 201716 218041 201772 218050
rect 198164 217514 198220 217523
rect 198164 217449 198220 217458
rect 197588 216478 197644 216487
rect 197588 216413 197644 216422
rect 201622 215995 201674 216001
rect 201622 215937 201674 215943
rect 201238 215773 201290 215779
rect 201238 215715 201290 215721
rect 201250 214267 201278 215715
rect 201634 214859 201662 215937
rect 201716 215886 201772 215895
rect 201716 215821 201772 215830
rect 201814 215847 201866 215853
rect 201730 215705 201758 215821
rect 201814 215789 201866 215795
rect 201718 215699 201770 215705
rect 201718 215641 201770 215647
rect 201620 214850 201676 214859
rect 201620 214785 201676 214794
rect 201236 214258 201292 214267
rect 201236 214193 201292 214202
rect 201826 213231 201854 215789
rect 201812 213222 201868 213231
rect 201812 213157 201868 213166
rect 201622 213109 201674 213115
rect 201622 213051 201674 213057
rect 201634 211603 201662 213051
rect 201718 213035 201770 213041
rect 201718 212977 201770 212983
rect 201730 212639 201758 212977
rect 201716 212630 201772 212639
rect 201716 212565 201772 212574
rect 201620 211594 201676 211603
rect 201620 211529 201676 211538
rect 200086 201639 200138 201645
rect 200086 201581 200138 201587
rect 197302 161309 197354 161315
rect 197302 161251 197354 161257
rect 197314 93351 197342 161251
rect 197398 123939 197450 123945
rect 197398 123881 197450 123887
rect 197300 93342 197356 93351
rect 197300 93277 197356 93286
rect 197410 79883 197438 123881
rect 199990 103589 200042 103595
rect 199990 103531 200042 103537
rect 200002 102231 200030 103531
rect 199988 102222 200044 102231
rect 199988 102157 200044 102166
rect 197686 92045 197738 92051
rect 197686 91987 197738 91993
rect 197698 91723 197726 91987
rect 197684 91714 197740 91723
rect 197684 91649 197740 91658
rect 198742 89011 198794 89017
rect 198742 88953 198794 88959
rect 198754 88615 198782 88953
rect 198740 88606 198796 88615
rect 198740 88541 198796 88550
rect 197782 82129 197834 82135
rect 197780 82094 197782 82103
rect 197834 82094 197836 82103
rect 197780 82029 197836 82038
rect 197396 79874 197452 79883
rect 197396 79809 197452 79818
rect 198358 74655 198410 74661
rect 198358 74597 198410 74603
rect 198370 73371 198398 74597
rect 198356 73362 198412 73371
rect 198356 73297 198412 73306
rect 199316 61374 199372 61383
rect 199316 61309 199372 61318
rect 199330 60527 199358 61309
rect 199318 60521 199370 60527
rect 199318 60463 199370 60469
rect 200098 48465 200126 201581
rect 200182 190169 200234 190175
rect 200182 190111 200234 190117
rect 200194 93499 200222 190111
rect 200278 126751 200330 126757
rect 200278 126693 200330 126699
rect 200180 93490 200236 93499
rect 200180 93425 200236 93434
rect 200290 80475 200318 126693
rect 201718 103663 201770 103669
rect 201718 103605 201770 103611
rect 201730 101639 201758 103605
rect 201716 101630 201772 101639
rect 201716 101565 201772 101574
rect 201814 100777 201866 100783
rect 201814 100719 201866 100725
rect 201622 100703 201674 100709
rect 201622 100645 201674 100651
rect 201634 98975 201662 100645
rect 201718 100629 201770 100635
rect 201716 100594 201718 100603
rect 201770 100594 201772 100603
rect 201716 100529 201772 100538
rect 201718 100481 201770 100487
rect 201718 100423 201770 100429
rect 201730 100011 201758 100423
rect 201716 100002 201772 100011
rect 201716 99937 201772 99946
rect 201620 98966 201676 98975
rect 201620 98901 201676 98910
rect 201826 98383 201854 100719
rect 201812 98374 201868 98383
rect 201812 98309 201868 98318
rect 201814 97743 201866 97749
rect 201814 97685 201866 97691
rect 201622 97669 201674 97675
rect 201622 97611 201674 97617
rect 201634 95719 201662 97611
rect 201718 97595 201770 97601
rect 201718 97537 201770 97543
rect 201730 96755 201758 97537
rect 201716 96746 201772 96755
rect 201716 96681 201772 96690
rect 201620 95710 201676 95719
rect 201620 95645 201676 95654
rect 201826 95127 201854 97685
rect 202978 97347 203006 221783
rect 203062 121201 203114 121207
rect 203062 121143 203114 121149
rect 202964 97338 203020 97347
rect 202964 97273 203020 97282
rect 201812 95118 201868 95127
rect 201812 95053 201868 95062
rect 201718 94931 201770 94937
rect 201718 94873 201770 94879
rect 201622 94709 201674 94715
rect 201622 94651 201674 94657
rect 201634 92463 201662 94651
rect 201730 94091 201758 94873
rect 201716 94082 201772 94091
rect 201716 94017 201772 94026
rect 201620 92454 201676 92463
rect 201620 92389 201676 92398
rect 201718 92119 201770 92125
rect 201718 92061 201770 92067
rect 201622 91971 201674 91977
rect 201622 91913 201674 91919
rect 201634 90243 201662 91913
rect 201730 91871 201758 92061
rect 201814 91897 201866 91903
rect 201716 91862 201772 91871
rect 201814 91839 201866 91845
rect 201716 91797 201772 91806
rect 201620 90234 201676 90243
rect 201620 90169 201676 90178
rect 201826 89651 201854 91839
rect 201812 89642 201868 89651
rect 201812 89577 201868 89586
rect 201814 89233 201866 89239
rect 201716 89198 201772 89207
rect 201622 89159 201674 89165
rect 201814 89175 201866 89181
rect 201716 89133 201772 89142
rect 201622 89101 201674 89107
rect 201526 89085 201578 89091
rect 201526 89027 201578 89033
rect 201538 88023 201566 89027
rect 201524 88014 201580 88023
rect 201524 87949 201580 87958
rect 201634 87579 201662 89101
rect 201730 88943 201758 89133
rect 201718 88937 201770 88943
rect 201718 88879 201770 88885
rect 201620 87570 201676 87579
rect 201620 87505 201676 87514
rect 201826 86987 201854 89175
rect 201812 86978 201868 86987
rect 201812 86913 201868 86922
rect 201910 86421 201962 86427
rect 201716 86386 201772 86395
rect 201526 86347 201578 86353
rect 201910 86363 201962 86369
rect 201716 86321 201772 86330
rect 201526 86289 201578 86295
rect 201538 84323 201566 86289
rect 201622 86199 201674 86205
rect 201622 86141 201674 86147
rect 201634 85359 201662 86141
rect 201730 86131 201758 86321
rect 201814 86273 201866 86279
rect 201814 86215 201866 86221
rect 201718 86125 201770 86131
rect 201718 86067 201770 86073
rect 201716 85942 201772 85951
rect 201716 85877 201772 85886
rect 201620 85350 201676 85359
rect 201620 85285 201676 85294
rect 201730 85021 201758 85877
rect 201718 85015 201770 85021
rect 201718 84957 201770 84963
rect 201826 84767 201854 86215
rect 201812 84758 201868 84767
rect 201812 84693 201868 84702
rect 201524 84314 201580 84323
rect 201524 84249 201580 84258
rect 201922 83731 201950 86363
rect 201908 83722 201964 83731
rect 201908 83657 201964 83666
rect 201622 83461 201674 83467
rect 201622 83403 201674 83409
rect 201046 83313 201098 83319
rect 201046 83255 201098 83261
rect 201058 83139 201086 83255
rect 201044 83130 201100 83139
rect 201044 83065 201100 83074
rect 201634 81511 201662 83403
rect 201718 83387 201770 83393
rect 201718 83329 201770 83335
rect 201730 82695 201758 83329
rect 201716 82686 201772 82695
rect 201716 82621 201772 82630
rect 201620 81502 201676 81511
rect 201620 81437 201676 81446
rect 201718 80649 201770 80655
rect 201718 80591 201770 80597
rect 200374 80575 200426 80581
rect 200374 80517 200426 80523
rect 200276 80466 200332 80475
rect 200276 80401 200332 80410
rect 200386 78847 200414 80517
rect 200372 78838 200428 78847
rect 200372 78773 200428 78782
rect 201730 78255 201758 80591
rect 201716 78246 201772 78255
rect 201716 78181 201772 78190
rect 201526 77763 201578 77769
rect 201526 77705 201578 77711
rect 201538 74999 201566 77705
rect 201814 77689 201866 77695
rect 201814 77631 201866 77637
rect 201622 77541 201674 77547
rect 201622 77483 201674 77489
rect 201634 76627 201662 77483
rect 201718 77467 201770 77473
rect 201718 77409 201770 77415
rect 201730 77219 201758 77409
rect 201716 77210 201772 77219
rect 201716 77145 201772 77154
rect 201620 76618 201676 76627
rect 201620 76553 201676 76562
rect 201826 75591 201854 77631
rect 201812 75582 201868 75591
rect 201812 75517 201868 75526
rect 201524 74990 201580 74999
rect 201524 74925 201580 74934
rect 201718 74803 201770 74809
rect 201718 74745 201770 74751
rect 200950 74729 201002 74735
rect 200950 74671 201002 74677
rect 200962 73223 200990 74671
rect 201046 74581 201098 74587
rect 201046 74523 201098 74529
rect 201058 73963 201086 74523
rect 201044 73954 201100 73963
rect 201044 73889 201100 73898
rect 200948 73214 201004 73223
rect 200948 73149 201004 73158
rect 201730 72335 201758 74745
rect 201716 72326 201772 72335
rect 201716 72261 201772 72270
rect 200470 71991 200522 71997
rect 200470 71933 200522 71939
rect 200482 69523 200510 71933
rect 201814 71917 201866 71923
rect 201814 71859 201866 71865
rect 201622 71843 201674 71849
rect 201622 71785 201674 71791
rect 201634 70707 201662 71785
rect 201716 71734 201772 71743
rect 201716 71669 201718 71678
rect 201770 71669 201772 71678
rect 201718 71637 201770 71643
rect 201620 70698 201676 70707
rect 201620 70633 201676 70642
rect 201826 70115 201854 71859
rect 201812 70106 201868 70115
rect 201812 70041 201868 70050
rect 200468 69514 200524 69523
rect 200468 69449 200524 69458
rect 201526 69105 201578 69111
rect 201526 69047 201578 69053
rect 201538 66859 201566 69047
rect 201814 69031 201866 69037
rect 201814 68973 201866 68979
rect 201622 68957 201674 68963
rect 201622 68899 201674 68905
rect 201634 67895 201662 68899
rect 201718 68883 201770 68889
rect 201718 68825 201770 68831
rect 201730 68487 201758 68825
rect 201716 68478 201772 68487
rect 201716 68413 201772 68422
rect 201620 67886 201676 67895
rect 201620 67821 201676 67830
rect 201826 67451 201854 68973
rect 201812 67442 201868 67451
rect 201812 67377 201868 67386
rect 201524 66850 201580 66859
rect 201524 66785 201580 66794
rect 201620 66258 201676 66267
rect 200182 66219 200234 66225
rect 201620 66193 201676 66202
rect 200182 66161 200234 66167
rect 200194 65231 200222 66161
rect 201634 66077 201662 66193
rect 201718 66145 201770 66151
rect 201718 66087 201770 66093
rect 201622 66071 201674 66077
rect 201622 66013 201674 66019
rect 201730 65823 201758 66087
rect 201716 65814 201772 65823
rect 201716 65749 201772 65758
rect 200180 65222 200236 65231
rect 200180 65157 200236 65166
rect 201718 64887 201770 64893
rect 201718 64829 201770 64835
rect 201730 64639 201758 64829
rect 201716 64630 201772 64639
rect 201716 64565 201772 64574
rect 201716 63594 201772 63603
rect 201716 63529 201772 63538
rect 201730 63413 201758 63529
rect 201718 63407 201770 63413
rect 201718 63349 201770 63355
rect 201716 63002 201772 63011
rect 201716 62937 201772 62946
rect 201620 61966 201676 61975
rect 201620 61901 201676 61910
rect 201634 60601 201662 61901
rect 201730 60823 201758 62937
rect 201718 60817 201770 60823
rect 201718 60759 201770 60765
rect 201622 60595 201674 60601
rect 201622 60537 201674 60543
rect 201718 60447 201770 60453
rect 201718 60389 201770 60395
rect 201620 60338 201676 60347
rect 201620 60273 201676 60282
rect 201634 59047 201662 60273
rect 201730 59755 201758 60389
rect 201716 59746 201772 59755
rect 201716 59681 201772 59690
rect 201622 59041 201674 59047
rect 201622 58983 201674 58989
rect 203074 48613 203102 121143
rect 203158 112469 203210 112475
rect 203158 112411 203210 112417
rect 203170 54279 203198 112411
rect 203156 54270 203212 54279
rect 203156 54205 203212 54214
rect 203062 48607 203114 48613
rect 203062 48549 203114 48555
rect 199222 48459 199274 48465
rect 199222 48401 199274 48407
rect 200086 48459 200138 48465
rect 200086 48401 200138 48407
rect 199234 47873 199262 48401
rect 199222 47867 199274 47873
rect 199222 47809 199274 47815
rect 205186 47767 205214 244871
rect 206518 243745 206570 243751
rect 206518 243687 206570 243693
rect 206530 241975 206558 243687
rect 206422 241969 206474 241975
rect 206422 241911 206474 241917
rect 206518 241969 206570 241975
rect 206518 241911 206570 241917
rect 207094 241969 207146 241975
rect 207094 241911 207146 241917
rect 206434 202871 206462 241911
rect 206806 233237 206858 233243
rect 206806 233179 206858 233185
rect 206710 233089 206762 233095
rect 206710 233031 206762 233037
rect 206614 232793 206666 232799
rect 206614 232735 206666 232741
rect 206626 231139 206654 232735
rect 206722 231731 206750 233031
rect 206818 232767 206846 233179
rect 206902 233163 206954 233169
rect 206902 233105 206954 233111
rect 206804 232758 206860 232767
rect 206804 232693 206860 232702
rect 206708 231722 206764 231731
rect 206708 231657 206764 231666
rect 206612 231130 206668 231139
rect 206612 231065 206668 231074
rect 206516 230094 206572 230103
rect 206516 230029 206572 230038
rect 206420 202862 206476 202871
rect 206420 202797 206476 202806
rect 206434 53793 206462 202797
rect 206530 54163 206558 230029
rect 206626 54237 206654 231065
rect 206614 54231 206666 54237
rect 206614 54173 206666 54179
rect 206518 54157 206570 54163
rect 206518 54099 206570 54105
rect 206422 53787 206474 53793
rect 206422 53729 206474 53735
rect 206722 53349 206750 231657
rect 206710 53343 206762 53349
rect 206710 53285 206762 53291
rect 206818 53275 206846 232693
rect 206914 232175 206942 233105
rect 206900 232166 206956 232175
rect 206900 232101 206956 232110
rect 206914 53941 206942 232101
rect 206996 230538 207052 230547
rect 206996 230473 207052 230482
rect 207010 54015 207038 230473
rect 206998 54009 207050 54015
rect 206998 53951 207050 53957
rect 206902 53935 206954 53941
rect 206902 53877 206954 53883
rect 206806 53269 206858 53275
rect 206806 53211 206858 53217
rect 207106 52979 207134 241911
rect 207202 233761 207230 246277
rect 207298 241943 207326 250495
rect 210178 244121 210206 256373
rect 215540 252146 215596 252155
rect 215540 252081 215596 252090
rect 214102 244929 214154 244935
rect 214102 244871 214154 244877
rect 210166 244115 210218 244121
rect 210166 244057 210218 244063
rect 212374 243597 212426 243603
rect 212374 243539 212426 243545
rect 211894 243449 211946 243455
rect 211894 243391 211946 243397
rect 209972 242230 210028 242239
rect 209972 242165 210028 242174
rect 208340 242082 208396 242091
rect 208340 242017 208396 242026
rect 207284 241934 207340 241943
rect 207284 241869 207340 241878
rect 207190 233755 207242 233761
rect 207190 233697 207242 233703
rect 207094 52973 207146 52979
rect 207094 52915 207146 52921
rect 207202 48803 207230 233697
rect 208246 62001 208298 62007
rect 208246 61943 208298 61949
rect 208150 61853 208202 61859
rect 208150 61795 208202 61801
rect 207284 55602 207340 55611
rect 207284 55537 207340 55546
rect 207188 48794 207244 48803
rect 207188 48729 207244 48738
rect 205172 47758 205228 47767
rect 205172 47693 205228 47702
rect 197206 46905 197258 46911
rect 197206 46847 197258 46853
rect 179926 46461 179978 46467
rect 179926 46403 179978 46409
rect 141814 44685 141866 44691
rect 141814 44627 141866 44633
rect 155542 44685 155594 44691
rect 155542 44627 155594 44633
rect 141826 40367 141854 44627
rect 207298 42175 207326 55537
rect 208054 48089 208106 48095
rect 208054 48031 208106 48037
rect 208066 47577 208094 48031
rect 208162 48021 208190 61795
rect 208258 48095 208286 61943
rect 208354 51795 208382 242017
rect 208724 241934 208780 241943
rect 208724 241869 208780 241878
rect 208738 239871 208766 241869
rect 208916 240454 208972 240463
rect 208916 240389 208972 240398
rect 208724 239862 208780 239871
rect 208450 239820 208724 239848
rect 208342 51789 208394 51795
rect 208342 51731 208394 51737
rect 208450 51721 208478 239820
rect 208724 239797 208780 239806
rect 208930 239723 208958 240389
rect 208916 239714 208972 239723
rect 208916 239649 208972 239658
rect 209876 239714 209932 239723
rect 209876 239649 209932 239658
rect 208726 239083 208778 239089
rect 208726 239025 208778 239031
rect 208738 74883 208766 239025
rect 209782 223247 209834 223253
rect 209782 223189 209834 223195
rect 209794 208527 209822 223189
rect 209782 208521 209834 208527
rect 209782 208463 209834 208469
rect 209890 169899 209918 239649
rect 209986 227268 210014 242165
rect 211508 237198 211564 237207
rect 211508 237133 211564 237142
rect 210070 234791 210122 234797
rect 210070 234733 210122 234739
rect 210082 228919 210110 234733
rect 211522 233803 211550 237133
rect 211906 234099 211934 243391
rect 212278 243375 212330 243381
rect 212278 243317 212330 243323
rect 211892 234090 211948 234099
rect 211892 234025 211948 234034
rect 211508 233794 211564 233803
rect 211508 233729 211564 233738
rect 210166 233681 210218 233687
rect 211316 233646 211372 233655
rect 210166 233623 210218 233629
rect 210068 228910 210124 228919
rect 210068 228845 210124 228854
rect 209986 227240 210110 227268
rect 209974 224283 210026 224289
rect 209974 224225 210026 224231
rect 209986 221889 210014 224225
rect 209972 221880 210028 221889
rect 209972 221815 210028 221824
rect 209974 221619 210026 221625
rect 209974 221561 210026 221567
rect 209986 220261 210014 221561
rect 209972 220252 210028 220261
rect 209972 220187 210028 220196
rect 209974 218807 210026 218813
rect 209974 218749 210026 218755
rect 209986 218633 210014 218749
rect 209972 218624 210028 218633
rect 209972 218559 210028 218568
rect 209974 215625 210026 215631
rect 209974 215567 210026 215573
rect 209986 215377 210014 215567
rect 209972 215368 210028 215377
rect 209972 215303 210028 215312
rect 209974 212961 210026 212967
rect 209974 212903 210026 212909
rect 209986 212121 210014 212903
rect 209972 212112 210028 212121
rect 209972 212047 210028 212056
rect 209974 169967 210026 169973
rect 209974 169909 210026 169915
rect 209878 169893 209930 169899
rect 209878 169835 209930 169841
rect 209986 169825 210014 169909
rect 209782 169819 209834 169825
rect 209782 169761 209834 169767
rect 209974 169819 210026 169825
rect 209974 169761 210026 169767
rect 209794 149845 209822 169761
rect 209878 169745 209930 169751
rect 209878 169687 209930 169693
rect 209782 149839 209834 149845
rect 209782 149781 209834 149787
rect 208822 132597 208874 132603
rect 208822 132539 208874 132545
rect 208726 74877 208778 74883
rect 208726 74819 208778 74825
rect 208630 71991 208682 71997
rect 208630 71933 208682 71939
rect 208534 61927 208586 61933
rect 208534 61869 208586 61875
rect 208438 51715 208490 51721
rect 208438 51657 208490 51663
rect 208546 48169 208574 61869
rect 208642 59195 208670 71933
rect 208726 63111 208778 63117
rect 208726 63053 208778 63059
rect 208630 59189 208682 59195
rect 208630 59131 208682 59137
rect 208738 53423 208766 63053
rect 208834 61859 208862 132539
rect 208918 132523 208970 132529
rect 208918 132465 208970 132471
rect 208930 62007 208958 132465
rect 209014 129637 209066 129643
rect 209014 129579 209066 129585
rect 208918 62001 208970 62007
rect 208918 61943 208970 61949
rect 209026 61933 209054 129579
rect 209110 121053 209162 121059
rect 209110 120995 209162 121001
rect 209014 61927 209066 61933
rect 209014 61869 209066 61875
rect 208822 61853 208874 61859
rect 208822 61795 208874 61801
rect 209122 59288 209150 120995
rect 209206 118167 209258 118173
rect 209206 118109 209258 118115
rect 209218 71997 209246 118109
rect 209302 115355 209354 115361
rect 209302 115297 209354 115303
rect 209206 71991 209258 71997
rect 209206 71933 209258 71939
rect 208834 59260 209150 59288
rect 208726 53417 208778 53423
rect 208726 53359 208778 53365
rect 208630 48977 208682 48983
rect 208630 48919 208682 48925
rect 208642 48243 208670 48919
rect 208834 48613 208862 59260
rect 209014 59189 209066 59195
rect 209014 59131 209066 59137
rect 209026 48687 209054 59131
rect 209314 48835 209342 115297
rect 209398 115281 209450 115287
rect 209398 115223 209450 115229
rect 209410 53719 209438 115223
rect 209494 112395 209546 112401
rect 209494 112337 209546 112343
rect 209506 54089 209534 112337
rect 209590 103737 209642 103743
rect 209590 103679 209642 103685
rect 209602 94216 209630 103679
rect 209686 100851 209738 100857
rect 209686 100793 209738 100799
rect 209698 94364 209726 100793
rect 209698 94336 209822 94364
rect 209602 94188 209726 94216
rect 209590 94117 209642 94123
rect 209590 94059 209642 94065
rect 209602 63117 209630 94059
rect 209590 63111 209642 63117
rect 209590 63053 209642 63059
rect 209698 62988 209726 94188
rect 209602 62960 209726 62988
rect 209494 54083 209546 54089
rect 209494 54025 209546 54031
rect 209398 53713 209450 53719
rect 209398 53655 209450 53661
rect 209602 53497 209630 62960
rect 209686 62889 209738 62895
rect 209686 62831 209738 62837
rect 209590 53491 209642 53497
rect 209590 53433 209642 53439
rect 209698 53391 209726 62831
rect 209794 54311 209822 94336
rect 209782 54305 209834 54311
rect 209782 54247 209834 54253
rect 209684 53382 209740 53391
rect 209684 53317 209740 53326
rect 209890 51869 209918 169687
rect 209974 149839 210026 149845
rect 209974 149781 210026 149787
rect 209986 148291 210014 149781
rect 209974 148285 210026 148291
rect 209974 148227 210026 148233
rect 210082 147033 210110 227240
rect 210178 223253 210206 233623
rect 210262 233607 210314 233613
rect 211200 233604 211316 233632
rect 211522 233618 211550 233729
rect 211906 233618 211934 234025
rect 212290 233951 212318 243317
rect 212276 233942 212332 233951
rect 212276 233877 212332 233886
rect 212290 233618 212318 233877
rect 212386 233687 212414 243539
rect 212758 243523 212810 243529
rect 212758 243465 212810 243471
rect 212374 233681 212426 233687
rect 212770 233632 212798 243465
rect 213142 241969 213194 241975
rect 213142 241911 213194 241917
rect 213154 233632 213182 241911
rect 213526 233755 213578 233761
rect 213526 233697 213578 233703
rect 213538 233632 213566 233697
rect 212426 233629 212640 233632
rect 212374 233623 212640 233629
rect 211316 233581 211372 233590
rect 212386 233604 212640 233623
rect 212770 233613 213024 233632
rect 212758 233607 213024 233613
rect 212386 233558 212414 233604
rect 210262 233549 210314 233555
rect 212810 233604 213024 233607
rect 213154 233604 213408 233632
rect 213538 233604 213744 233632
rect 214114 233618 214142 244871
rect 214486 244855 214538 244861
rect 214486 244797 214538 244803
rect 214196 233646 214252 233655
rect 214498 233632 214526 244797
rect 215554 243423 215582 252081
rect 215636 248594 215692 248603
rect 215636 248529 215692 248538
rect 215540 243414 215596 243423
rect 215540 243349 215596 243358
rect 215060 241786 215116 241795
rect 215060 241721 215116 241730
rect 215074 233632 215102 241721
rect 215444 239714 215500 239723
rect 215444 239649 215500 239658
rect 215458 233632 215486 239649
rect 215650 239089 215678 248529
rect 216034 244163 216062 246938
rect 216384 246924 216638 246952
rect 216864 246924 217118 246952
rect 216020 244154 216076 244163
rect 216020 244089 216076 244098
rect 215828 240602 215884 240611
rect 215828 240537 215884 240546
rect 215638 239083 215690 239089
rect 215638 239025 215690 239031
rect 215842 233632 215870 240537
rect 215924 240454 215980 240463
rect 215924 240389 215980 240398
rect 214252 233618 214526 233632
rect 214252 233604 214512 233618
rect 214848 233604 215102 233632
rect 215232 233604 215486 233632
rect 215616 233604 215870 233632
rect 215938 233618 215966 240389
rect 216610 239237 216638 246924
rect 216694 241747 216746 241753
rect 216694 241689 216746 241695
rect 216598 239231 216650 239237
rect 216598 239173 216650 239179
rect 216706 233803 216734 241689
rect 217090 237947 217118 246924
rect 217282 241309 217310 246938
rect 217558 244707 217610 244713
rect 217558 244649 217610 244655
rect 217270 241303 217322 241309
rect 217270 241245 217322 241251
rect 217270 238565 217322 238571
rect 217270 238507 217322 238513
rect 217076 237938 217132 237947
rect 217076 237873 217132 237882
rect 216692 233794 216748 233803
rect 216692 233729 216748 233738
rect 216336 233613 216542 233632
rect 216706 233618 216734 233729
rect 217282 233632 217310 238507
rect 217570 233632 217598 244649
rect 217666 243571 217694 246938
rect 217652 243562 217708 243571
rect 217652 243497 217708 243506
rect 218146 239977 218174 246938
rect 218592 246924 218846 246952
rect 218422 244337 218474 244343
rect 218422 244279 218474 244285
rect 218134 239971 218186 239977
rect 218134 239913 218186 239919
rect 218038 238343 218090 238349
rect 218038 238285 218090 238291
rect 218050 233632 218078 238285
rect 218434 233632 218462 244279
rect 218518 238269 218570 238275
rect 218518 238211 218570 238217
rect 216336 233607 216554 233613
rect 216336 233604 216502 233607
rect 214196 233581 214252 233590
rect 212758 233549 212810 233555
rect 217056 233604 217310 233632
rect 217440 233604 217598 233632
rect 217824 233604 218078 233632
rect 218160 233604 218462 233632
rect 218530 233618 218558 238211
rect 218818 237799 218846 246924
rect 219010 246924 219072 246952
rect 219202 246924 219408 246952
rect 219888 246924 220190 246952
rect 218804 237790 218860 237799
rect 218804 237725 218860 237734
rect 219010 237651 219038 246924
rect 218996 237642 219052 237651
rect 218996 237577 219052 237586
rect 219202 233780 219230 246924
rect 219478 244041 219530 244047
rect 219478 243983 219530 243989
rect 219106 233752 219230 233780
rect 219106 233632 219134 233752
rect 219490 233632 219518 243983
rect 219862 238417 219914 238423
rect 219862 238359 219914 238365
rect 219874 233632 219902 238359
rect 220162 233761 220190 246924
rect 220354 241161 220382 246938
rect 220800 246924 221054 246952
rect 221184 246924 221438 246952
rect 220726 243893 220778 243899
rect 220726 243835 220778 243841
rect 220342 241155 220394 241161
rect 220342 241097 220394 241103
rect 220246 239749 220298 239755
rect 220246 239691 220298 239697
rect 220150 233755 220202 233761
rect 220150 233697 220202 233703
rect 220258 233632 220286 239691
rect 220342 238195 220394 238201
rect 220342 238137 220394 238143
rect 218928 233604 219134 233632
rect 219264 233604 219518 233632
rect 219648 233604 219902 233632
rect 220032 233604 220286 233632
rect 220354 233618 220382 238137
rect 220738 233618 220766 243835
rect 221026 238391 221054 246924
rect 221410 241901 221438 246924
rect 221602 243719 221630 246938
rect 221588 243710 221644 243719
rect 221588 243645 221644 243654
rect 221398 241895 221450 241901
rect 221398 241837 221450 241843
rect 221686 240711 221738 240717
rect 221686 240653 221738 240659
rect 221110 240637 221162 240643
rect 221110 240579 221162 240585
rect 221012 238382 221068 238391
rect 221012 238317 221068 238326
rect 221122 233618 221150 240579
rect 221698 233632 221726 240653
rect 222082 240273 222110 246938
rect 222576 246924 222782 246952
rect 222912 246924 223166 246952
rect 223392 246924 223646 246952
rect 222550 240785 222602 240791
rect 222550 240727 222602 240733
rect 222070 240267 222122 240273
rect 222070 240209 222122 240215
rect 222070 239675 222122 239681
rect 222070 239617 222122 239623
rect 222082 233632 222110 239617
rect 222166 239083 222218 239089
rect 222166 239025 222218 239031
rect 221472 233604 221726 233632
rect 221856 233604 222110 233632
rect 222178 233632 222206 239025
rect 222178 233604 222240 233632
rect 222562 233618 222590 240727
rect 222754 238539 222782 246924
rect 223138 241827 223166 246924
rect 223618 244015 223646 246924
rect 223604 244006 223660 244015
rect 223604 243941 223660 243950
rect 223126 241821 223178 241827
rect 223126 241763 223178 241769
rect 223318 241007 223370 241013
rect 223318 240949 223370 240955
rect 222934 239305 222986 239311
rect 222934 239247 222986 239253
rect 222740 238530 222796 238539
rect 222740 238465 222796 238474
rect 222946 233618 222974 239247
rect 223330 233618 223358 240949
rect 223810 239533 223838 246938
rect 223894 240859 223946 240865
rect 223894 240801 223946 240807
rect 223798 239527 223850 239533
rect 223798 239469 223850 239475
rect 223906 233632 223934 240801
rect 224194 238095 224222 246938
rect 224468 245338 224524 245347
rect 224468 245273 224524 245282
rect 224482 244755 224510 245273
rect 224674 244755 224702 246938
rect 225120 246924 225374 246952
rect 225600 246924 225854 246952
rect 224468 244746 224524 244755
rect 224468 244681 224524 244690
rect 224660 244746 224716 244755
rect 224660 244681 224716 244690
rect 225346 241383 225374 246924
rect 225334 241377 225386 241383
rect 225334 241319 225386 241325
rect 224566 240933 224618 240939
rect 224566 240875 224618 240881
rect 224278 240415 224330 240421
rect 224278 240357 224330 240363
rect 224180 238086 224236 238095
rect 224180 238021 224236 238030
rect 224290 233632 224318 240357
rect 224578 233632 224606 240875
rect 225526 240563 225578 240569
rect 225526 240505 225578 240511
rect 225142 239971 225194 239977
rect 225142 239913 225194 239919
rect 224758 239601 224810 239607
rect 224758 239543 224810 239549
rect 223680 233604 223934 233632
rect 224064 233604 224318 233632
rect 224448 233604 224606 233632
rect 224770 233618 224798 239543
rect 225154 233618 225182 239913
rect 225538 233618 225566 240505
rect 225826 238243 225854 246924
rect 225922 241457 225950 246938
rect 226402 243867 226430 246938
rect 226388 243858 226444 243867
rect 226388 243793 226444 243802
rect 226882 241679 226910 246938
rect 227328 246924 227486 246952
rect 227712 246924 227966 246952
rect 226870 241673 226922 241679
rect 226870 241615 226922 241621
rect 225910 241451 225962 241457
rect 225910 241393 225962 241399
rect 226486 241081 226538 241087
rect 226486 241023 226538 241029
rect 226102 240489 226154 240495
rect 226102 240431 226154 240437
rect 225812 238234 225868 238243
rect 225812 238169 225868 238178
rect 226114 233632 226142 240431
rect 226498 233632 226526 241023
rect 226870 240193 226922 240199
rect 226870 240135 226922 240141
rect 226882 233632 226910 240135
rect 226966 240045 227018 240051
rect 226966 239987 227018 239993
rect 225888 233604 226142 233632
rect 226272 233604 226526 233632
rect 226656 233604 226910 233632
rect 226978 233618 227006 239987
rect 227350 239971 227402 239977
rect 227350 239913 227402 239919
rect 227362 233618 227390 239913
rect 227458 238687 227486 246924
rect 227542 241599 227594 241605
rect 227542 241541 227594 241547
rect 227554 240421 227582 241541
rect 227542 240415 227594 240421
rect 227542 240357 227594 240363
rect 227938 240125 227966 246924
rect 228130 244607 228158 246938
rect 228116 244598 228172 244607
rect 228116 244533 228172 244542
rect 228502 241525 228554 241531
rect 228502 241467 228554 241473
rect 228310 240267 228362 240273
rect 228310 240209 228362 240215
rect 227926 240119 227978 240125
rect 227926 240061 227978 240067
rect 227734 239083 227786 239089
rect 227734 239025 227786 239031
rect 227444 238678 227500 238687
rect 227444 238613 227500 238622
rect 227746 233618 227774 239025
rect 228322 233632 228350 240209
rect 228514 240199 228542 241467
rect 228502 240193 228554 240199
rect 228502 240135 228554 240141
rect 228610 239163 228638 246938
rect 228886 241747 228938 241753
rect 228886 241689 228938 241695
rect 228898 240569 228926 241689
rect 228886 240563 228938 240569
rect 228886 240505 228938 240511
rect 228982 240563 229034 240569
rect 228982 240505 229034 240511
rect 228694 240193 228746 240199
rect 228694 240135 228746 240141
rect 228598 239157 228650 239163
rect 228598 239099 228650 239105
rect 228706 233632 228734 240135
rect 228994 240051 229022 240505
rect 229090 240051 229118 246938
rect 229440 246924 229694 246952
rect 229920 246924 230174 246952
rect 229666 244459 229694 246924
rect 229652 244450 229708 244459
rect 229652 244385 229708 244394
rect 229174 241303 229226 241309
rect 229174 241245 229226 241251
rect 228982 240045 229034 240051
rect 228982 239987 229034 239993
rect 229078 240045 229130 240051
rect 229078 239987 229130 239993
rect 229078 239823 229130 239829
rect 229078 239765 229130 239771
rect 229090 233632 229118 239765
rect 228096 233604 228350 233632
rect 228480 233604 228734 233632
rect 228864 233604 229118 233632
rect 229186 233618 229214 241245
rect 229942 241155 229994 241161
rect 229942 241097 229994 241103
rect 229954 240495 229982 241097
rect 229942 240489 229994 240495
rect 229942 240431 229994 240437
rect 230038 240489 230090 240495
rect 230038 240431 230090 240437
rect 230050 239977 230078 240431
rect 230146 239977 230174 246924
rect 230242 246924 230352 246952
rect 230434 246924 230832 246952
rect 230038 239971 230090 239977
rect 230038 239913 230090 239919
rect 230134 239971 230186 239977
rect 230134 239913 230186 239919
rect 229558 239897 229610 239903
rect 229558 239839 229610 239845
rect 229570 233618 229598 239839
rect 229942 239305 229994 239311
rect 229942 239247 229994 239253
rect 229954 233618 229982 239247
rect 230242 238835 230270 246924
rect 230434 239108 230462 246924
rect 231202 243127 231230 246938
rect 231394 246924 231648 246952
rect 231188 243118 231244 243127
rect 231188 243053 231244 243062
rect 230806 240045 230858 240051
rect 230806 239987 230858 239993
rect 230518 239971 230570 239977
rect 230518 239913 230570 239919
rect 230338 239080 230462 239108
rect 230228 238826 230284 238835
rect 230228 238761 230284 238770
rect 230338 233632 230366 239080
rect 230304 233604 230366 233632
rect 230530 233632 230558 239913
rect 230818 233632 230846 239987
rect 231394 239311 231422 246924
rect 232114 246656 232142 246938
rect 232066 246628 232142 246656
rect 232258 246924 232512 246952
rect 231766 240119 231818 240125
rect 231766 240061 231818 240067
rect 231382 239305 231434 239311
rect 231382 239247 231434 239253
rect 231382 239157 231434 239163
rect 231382 239099 231434 239105
rect 230530 233604 230688 233632
rect 230818 233604 231072 233632
rect 231394 233618 231422 239099
rect 231778 233618 231806 240061
rect 232066 238983 232094 246628
rect 232150 241673 232202 241679
rect 232150 241615 232202 241621
rect 232052 238974 232108 238983
rect 232052 238909 232108 238918
rect 232162 233618 232190 241615
rect 232258 239903 232286 246924
rect 232930 244311 232958 246938
rect 232916 244302 232972 244311
rect 232916 244237 232972 244246
rect 232342 241451 232394 241457
rect 232342 241393 232394 241399
rect 232246 239897 232298 239903
rect 232246 239839 232298 239845
rect 232354 233632 232382 241393
rect 232630 241377 232682 241383
rect 232630 241319 232682 241325
rect 232642 233632 232670 241319
rect 233206 239231 233258 239237
rect 233206 239173 233258 239179
rect 233218 233632 233246 239173
rect 233410 237609 233438 246938
rect 233602 246924 233856 246952
rect 234240 246924 234398 246952
rect 233602 239829 233630 246924
rect 234370 242979 234398 246924
rect 234466 246924 234720 246952
rect 234356 242970 234412 242979
rect 234356 242905 234412 242914
rect 233974 241821 234026 241827
rect 233974 241763 234026 241769
rect 233590 239823 233642 239829
rect 233590 239765 233642 239771
rect 233590 239527 233642 239533
rect 233590 239469 233642 239475
rect 233398 237603 233450 237609
rect 233398 237545 233450 237551
rect 232354 233604 232512 233632
rect 232642 233604 232896 233632
rect 233218 233604 233280 233632
rect 233602 233618 233630 239469
rect 233986 233618 234014 241763
rect 234358 240341 234410 240347
rect 234358 240283 234410 240289
rect 234370 233618 234398 240283
rect 234466 240199 234494 246924
rect 234550 241895 234602 241901
rect 234550 241837 234602 241843
rect 234454 240193 234506 240199
rect 234454 240135 234506 240141
rect 234562 233632 234590 241837
rect 235138 237503 235166 246938
rect 235318 241377 235370 241383
rect 235318 241319 235370 241325
rect 235330 241013 235358 241319
rect 235318 241007 235370 241013
rect 235318 240949 235370 240955
rect 235618 240273 235646 246938
rect 236002 243275 236030 246938
rect 236194 246924 236448 246952
rect 236928 246924 237086 246952
rect 235988 243266 236044 243275
rect 235988 243201 236044 243210
rect 235606 240267 235658 240273
rect 235606 240209 235658 240215
rect 236194 239089 236222 246924
rect 236470 244559 236522 244565
rect 236470 244501 236522 244507
rect 236278 241303 236330 241309
rect 236278 241245 236330 241251
rect 236290 240865 236318 241245
rect 236278 240859 236330 240865
rect 236278 240801 236330 240807
rect 236182 239083 236234 239089
rect 236182 239025 236234 239031
rect 235318 238935 235370 238941
rect 235318 238877 235370 238883
rect 235124 237494 235180 237503
rect 235124 237429 235180 237438
rect 235330 233632 235358 238877
rect 235798 238787 235850 238793
rect 235798 238729 235850 238735
rect 235702 237011 235754 237017
rect 235702 236953 235754 236959
rect 235714 233632 235742 236953
rect 234562 233604 234720 233632
rect 235104 233604 235358 233632
rect 235488 233604 235742 233632
rect 235810 233618 235838 238729
rect 236482 233632 236510 244501
rect 236662 241599 236714 241605
rect 236662 241541 236714 241547
rect 236566 241451 236618 241457
rect 236566 241393 236618 241399
rect 236578 239089 236606 241393
rect 236674 239681 236702 241541
rect 236662 239675 236714 239681
rect 236662 239617 236714 239623
rect 236758 239675 236810 239681
rect 236758 239617 236810 239623
rect 236566 239083 236618 239089
rect 236566 239025 236618 239031
rect 236770 233632 236798 239617
rect 237058 238497 237086 246924
rect 237238 241451 237290 241457
rect 237238 241393 237290 241399
rect 237250 240791 237278 241393
rect 237238 240785 237290 240791
rect 237238 240727 237290 240733
rect 237346 240495 237374 246938
rect 237442 246924 237744 246952
rect 237442 240569 237470 246924
rect 237622 240785 237674 240791
rect 237622 240727 237674 240733
rect 237430 240563 237482 240569
rect 237430 240505 237482 240511
rect 237334 240489 237386 240495
rect 237334 240431 237386 240437
rect 237142 239157 237194 239163
rect 237142 239099 237194 239105
rect 237046 238491 237098 238497
rect 237046 238433 237098 238439
rect 237154 233632 237182 239099
rect 237634 233780 237662 240727
rect 237910 240563 237962 240569
rect 237910 240505 237962 240511
rect 237538 233752 237662 233780
rect 237538 233632 237566 233752
rect 237922 233632 237950 240505
rect 238006 240489 238058 240495
rect 238006 240431 238058 240437
rect 236208 233604 236510 233632
rect 236592 233604 236798 233632
rect 236928 233604 237182 233632
rect 237312 233604 237566 233632
rect 237696 233604 237950 233632
rect 238018 233618 238046 240431
rect 238210 237355 238238 246938
rect 238402 246924 238656 246952
rect 239136 246924 239390 246952
rect 238402 241531 238430 246924
rect 239362 243455 239390 246924
rect 239350 243449 239402 243455
rect 239350 243391 239402 243397
rect 238390 241525 238442 241531
rect 238390 241467 238442 241473
rect 238774 241525 238826 241531
rect 238774 241467 238826 241473
rect 238390 239083 238442 239089
rect 238390 239025 238442 239031
rect 238196 237346 238252 237355
rect 238196 237281 238252 237290
rect 238402 233618 238430 239025
rect 238786 233618 238814 241467
rect 239350 241229 239402 241235
rect 239350 241171 239402 241177
rect 238966 240711 239018 240717
rect 238966 240653 239018 240659
rect 238978 239163 239006 240653
rect 238966 239157 239018 239163
rect 238966 239099 239018 239105
rect 239362 233632 239390 241171
rect 239458 241087 239486 246938
rect 239734 241821 239786 241827
rect 239734 241763 239786 241769
rect 239446 241081 239498 241087
rect 239446 241023 239498 241029
rect 239746 233632 239774 241763
rect 239938 237683 239966 246938
rect 240214 241895 240266 241901
rect 240214 241837 240266 241843
rect 240118 240267 240170 240273
rect 240118 240209 240170 240215
rect 239926 237677 239978 237683
rect 239926 237619 239978 237625
rect 240130 233632 240158 240209
rect 239136 233604 239390 233632
rect 239520 233604 239774 233632
rect 239904 233604 240158 233632
rect 240226 233618 240254 241837
rect 240418 241161 240446 246938
rect 240768 246924 241022 246952
rect 240994 243529 241022 246924
rect 241090 246924 241248 246952
rect 240982 243523 241034 243529
rect 240982 243465 241034 243471
rect 240596 241934 240652 241943
rect 240596 241869 240652 241878
rect 240406 241155 240458 241161
rect 240406 241097 240458 241103
rect 240502 241155 240554 241161
rect 240502 241097 240554 241103
rect 240514 240495 240542 241097
rect 240502 240489 240554 240495
rect 240502 240431 240554 240437
rect 240610 233618 240638 241869
rect 241090 241753 241118 246924
rect 241078 241747 241130 241753
rect 241078 241689 241130 241695
rect 241556 240898 241612 240907
rect 241556 240833 241612 240842
rect 240980 240750 241036 240759
rect 240980 240685 241036 240694
rect 240994 233618 241022 240685
rect 241570 233632 241598 240833
rect 241666 237831 241694 246938
rect 242146 243381 242174 246938
rect 242134 243375 242186 243381
rect 242134 243317 242186 243323
rect 242420 241342 242476 241351
rect 242420 241277 242476 241286
rect 242324 241194 242380 241203
rect 242324 241129 242380 241138
rect 241844 240158 241900 240167
rect 241844 240093 241900 240102
rect 241654 237825 241706 237831
rect 241654 237767 241706 237773
rect 241858 233632 241886 240093
rect 242338 233632 242366 241129
rect 241344 233604 241598 233632
rect 241728 233604 241886 233632
rect 242112 233604 242366 233632
rect 242434 233618 242462 241277
rect 242530 239607 242558 246938
rect 242976 246924 243134 246952
rect 242804 241490 242860 241499
rect 242804 241425 242860 241434
rect 242518 239601 242570 239607
rect 242518 239543 242570 239549
rect 242818 233618 242846 241425
rect 243106 237905 243134 246924
rect 243202 246924 243456 246952
rect 243202 241013 243230 246924
rect 243874 243307 243902 246938
rect 243862 243301 243914 243307
rect 243862 243243 243914 243249
rect 244258 241679 244286 246938
rect 244630 241969 244682 241975
rect 244630 241911 244682 241917
rect 244246 241673 244298 241679
rect 243380 241638 243436 241647
rect 244246 241615 244298 241621
rect 243380 241573 243436 241582
rect 243190 241007 243242 241013
rect 243190 240949 243242 240955
rect 243286 241007 243338 241013
rect 243286 240949 243338 240955
rect 243298 240569 243326 240949
rect 243286 240563 243338 240569
rect 243286 240505 243338 240511
rect 243094 237899 243146 237905
rect 243094 237841 243146 237847
rect 243394 233632 243422 241573
rect 244534 240563 244586 240569
rect 244534 240505 244586 240511
rect 243766 239601 243818 239607
rect 243766 239543 243818 239549
rect 243778 233632 243806 239543
rect 243910 233903 243962 233909
rect 243910 233845 243962 233851
rect 243216 233604 243422 233632
rect 243552 233604 243806 233632
rect 243922 233618 243950 233845
rect 244546 233632 244574 240505
rect 244320 233604 244574 233632
rect 244642 233618 244670 241911
rect 244738 237757 244766 246938
rect 244930 246924 245184 246952
rect 245664 246924 245918 246952
rect 244930 241309 244958 246924
rect 245890 243603 245918 246924
rect 245878 243597 245930 243603
rect 245878 243539 245930 243545
rect 245398 241821 245450 241827
rect 245398 241763 245450 241769
rect 244918 241303 244970 241309
rect 244918 241245 244970 241251
rect 245014 239379 245066 239385
rect 245014 239321 245066 239327
rect 244726 237751 244778 237757
rect 244726 237693 244778 237699
rect 245026 233618 245054 239321
rect 245410 233618 245438 241763
rect 245986 241383 246014 246938
rect 246358 245151 246410 245157
rect 246358 245093 246410 245099
rect 245974 241377 246026 241383
rect 245974 241319 246026 241325
rect 245974 234273 246026 234279
rect 245974 234215 246026 234221
rect 245986 233632 246014 234215
rect 246370 233632 246398 245093
rect 246466 239533 246494 246938
rect 246838 245225 246890 245231
rect 246838 245167 246890 245173
rect 246454 239527 246506 239533
rect 246454 239469 246506 239475
rect 246742 234347 246794 234353
rect 246742 234289 246794 234295
rect 246754 233632 246782 234289
rect 245760 233604 246014 233632
rect 246144 233604 246398 233632
rect 246528 233604 246782 233632
rect 246850 233618 246878 245167
rect 246946 243751 246974 246938
rect 247138 246924 247392 246952
rect 247776 246924 248030 246952
rect 246934 243745 246986 243751
rect 246934 243687 246986 243693
rect 247138 241457 247166 246924
rect 247606 245373 247658 245379
rect 247606 245315 247658 245321
rect 247318 241525 247370 241531
rect 247318 241467 247370 241473
rect 247126 241451 247178 241457
rect 247126 241393 247178 241399
rect 247330 241235 247358 241467
rect 247318 241229 247370 241235
rect 247318 241171 247370 241177
rect 247414 241081 247466 241087
rect 247414 241023 247466 241029
rect 247426 239681 247454 241023
rect 247414 239675 247466 239681
rect 247414 239617 247466 239623
rect 247222 234421 247274 234427
rect 247222 234363 247274 234369
rect 247234 233618 247262 234363
rect 247618 233618 247646 245315
rect 248002 238645 248030 246924
rect 248194 243973 248222 246938
rect 248566 245595 248618 245601
rect 248566 245537 248618 245543
rect 248182 243967 248234 243973
rect 248182 243909 248234 243915
rect 247990 238639 248042 238645
rect 247990 238581 248042 238587
rect 248182 234569 248234 234575
rect 248182 234511 248234 234517
rect 248194 233632 248222 234511
rect 248578 233632 248606 245537
rect 248674 241605 248702 246938
rect 248662 241599 248714 241605
rect 248662 241541 248714 241547
rect 249058 238053 249086 246938
rect 249250 246924 249504 246952
rect 249984 246924 250238 246952
rect 249250 240939 249278 246924
rect 249814 245669 249866 245675
rect 249814 245611 249866 245617
rect 249334 245521 249386 245527
rect 249334 245463 249386 245469
rect 249238 240933 249290 240939
rect 249238 240875 249290 240881
rect 249046 238047 249098 238053
rect 249046 237989 249098 237995
rect 248950 235679 249002 235685
rect 248950 235621 249002 235627
rect 248962 233632 248990 235621
rect 249346 233632 249374 245463
rect 249430 234717 249482 234723
rect 249430 234659 249482 234665
rect 247968 233604 248222 233632
rect 248352 233604 248606 233632
rect 248736 233604 248990 233632
rect 249072 233604 249374 233632
rect 249442 233618 249470 234659
rect 249826 233618 249854 245611
rect 250210 244343 250238 246924
rect 250198 244337 250250 244343
rect 250198 244279 250250 244285
rect 250402 240865 250430 246938
rect 250486 245743 250538 245749
rect 250486 245685 250538 245691
rect 250390 240859 250442 240865
rect 250390 240801 250442 240807
rect 250390 234865 250442 234871
rect 250390 234807 250442 234813
rect 250402 233632 250430 234807
rect 250498 233928 250526 245685
rect 250786 243899 250814 246938
rect 251266 244121 251294 246938
rect 251458 246924 251712 246952
rect 252192 246924 252446 246952
rect 251254 244115 251306 244121
rect 251254 244057 251306 244063
rect 250774 243893 250826 243899
rect 250774 243835 250826 243841
rect 251458 238201 251486 246924
rect 251542 245891 251594 245897
rect 251542 245833 251594 245839
rect 251446 238195 251498 238201
rect 251446 238137 251498 238143
rect 251158 235013 251210 235019
rect 251158 234955 251210 234961
rect 250498 233900 250574 233928
rect 250176 233604 250430 233632
rect 250546 233618 250574 233900
rect 251170 233632 251198 234955
rect 251554 233632 251582 245833
rect 252022 245817 252074 245823
rect 252022 245759 252074 245765
rect 251638 235161 251690 235167
rect 251638 235103 251690 235109
rect 250944 233604 251198 233632
rect 251280 233604 251582 233632
rect 251650 233618 251678 235103
rect 252034 233618 252062 245759
rect 252418 238127 252446 246924
rect 252514 240643 252542 246938
rect 252886 246705 252938 246711
rect 252886 246647 252938 246653
rect 252502 240637 252554 240643
rect 252502 240579 252554 240585
rect 252406 238121 252458 238127
rect 252406 238063 252458 238069
rect 252598 235235 252650 235241
rect 252598 235177 252650 235183
rect 252610 233632 252638 235177
rect 252898 233632 252926 246647
rect 252994 243899 253022 246938
rect 252982 243893 253034 243899
rect 252982 243835 253034 243841
rect 253474 238423 253502 246938
rect 253920 246924 253982 246952
rect 253750 246039 253802 246045
rect 253750 245981 253802 245987
rect 253462 238417 253514 238423
rect 253462 238359 253514 238365
rect 253366 235309 253418 235315
rect 253366 235251 253418 235257
rect 253378 233632 253406 235251
rect 253762 233632 253790 245981
rect 253954 238201 253982 246924
rect 254050 246924 254304 246952
rect 254050 244047 254078 246924
rect 254230 246261 254282 246267
rect 254230 246203 254282 246209
rect 254038 244041 254090 244047
rect 254038 243983 254090 243989
rect 253942 238195 253994 238201
rect 253942 238137 253994 238143
rect 253846 235383 253898 235389
rect 253846 235325 253898 235331
rect 252384 233604 252638 233632
rect 252768 233604 252926 233632
rect 253152 233604 253406 233632
rect 253488 233604 253790 233632
rect 253858 233618 253886 235325
rect 254242 233618 254270 246203
rect 254722 244195 254750 246938
rect 255094 246335 255146 246341
rect 255094 246277 255146 246283
rect 254710 244189 254762 244195
rect 254710 244131 254762 244137
rect 254326 243671 254378 243677
rect 254326 243613 254378 243619
rect 254338 243381 254366 243613
rect 254326 243375 254378 243381
rect 254326 243317 254378 243323
rect 254806 235457 254858 235463
rect 254806 235399 254858 235405
rect 254818 233632 254846 235399
rect 255106 233632 255134 246277
rect 255202 238423 255230 246938
rect 255190 238417 255242 238423
rect 255190 238359 255242 238365
rect 255682 238275 255710 246938
rect 256032 246924 256286 246952
rect 255958 246409 256010 246415
rect 255958 246351 256010 246357
rect 255670 238269 255722 238275
rect 255670 238211 255722 238217
rect 255574 235531 255626 235537
rect 255574 235473 255626 235479
rect 255586 233632 255614 235473
rect 255970 233632 255998 246351
rect 256258 244047 256286 246924
rect 256354 246924 256512 246952
rect 256354 244639 256382 246924
rect 256438 246483 256490 246489
rect 256438 246425 256490 246431
rect 256342 244633 256394 244639
rect 256342 244575 256394 244581
rect 256246 244041 256298 244047
rect 256246 243983 256298 243989
rect 256054 235605 256106 235611
rect 256054 235547 256106 235553
rect 254592 233604 254846 233632
rect 254976 233604 255134 233632
rect 255360 233604 255614 233632
rect 255696 233604 255998 233632
rect 256066 233618 256094 235547
rect 256450 233618 256478 246425
rect 256930 238719 256958 246938
rect 257014 246853 257066 246859
rect 257014 246795 257066 246801
rect 256918 238713 256970 238719
rect 256918 238655 256970 238661
rect 257026 233632 257054 246795
rect 257314 238349 257342 246938
rect 257590 246557 257642 246563
rect 257590 246499 257642 246505
rect 257302 238343 257354 238349
rect 257302 238285 257354 238291
rect 257398 235753 257450 235759
rect 257398 235695 257450 235701
rect 257410 233632 257438 235695
rect 257602 233928 257630 246499
rect 257686 238491 257738 238497
rect 257686 238433 257738 238439
rect 257698 237905 257726 238433
rect 257686 237899 257738 237905
rect 257686 237841 257738 237847
rect 257794 235093 257822 246938
rect 257986 246924 258240 246952
rect 258720 246924 258974 246952
rect 257986 244713 258014 246924
rect 258262 246631 258314 246637
rect 258262 246573 258314 246579
rect 257974 244707 258026 244713
rect 257974 244649 258026 244655
rect 257878 235827 257930 235833
rect 257878 235769 257930 235775
rect 257782 235087 257834 235093
rect 257782 235029 257834 235035
rect 256800 233604 257054 233632
rect 257184 233604 257438 233632
rect 257554 233900 257630 233928
rect 257554 233618 257582 233900
rect 257890 233618 257918 235769
rect 258274 233618 258302 246573
rect 258838 244337 258890 244343
rect 258838 244279 258890 244285
rect 258850 243677 258878 244279
rect 258838 243671 258890 243677
rect 258838 243613 258890 243619
rect 258946 234945 258974 246924
rect 259042 238571 259070 246938
rect 259220 245190 259276 245199
rect 259220 245125 259276 245134
rect 259234 245051 259262 245125
rect 259220 245042 259276 245051
rect 259220 244977 259276 244986
rect 259522 241901 259550 246938
rect 259894 244929 259946 244935
rect 259894 244871 259946 244877
rect 259606 244855 259658 244861
rect 259606 244797 259658 244803
rect 259510 241895 259562 241901
rect 259510 241837 259562 241843
rect 259030 238565 259082 238571
rect 259030 238507 259082 238513
rect 258934 234939 258986 234945
rect 258934 234881 258986 234887
rect 258982 233829 259034 233835
rect 258982 233771 259034 233777
rect 258838 233755 258890 233761
rect 258838 233697 258890 233703
rect 258850 233632 258878 233697
rect 258672 233604 258878 233632
rect 258994 233618 259022 233771
rect 259618 233632 259646 244797
rect 259906 233632 259934 244871
rect 260002 238497 260030 246938
rect 260194 246924 260448 246952
rect 260832 246924 261086 246952
rect 260194 240273 260222 246924
rect 260470 245003 260522 245009
rect 260470 244945 260522 244951
rect 260182 240267 260234 240273
rect 260182 240209 260234 240215
rect 259990 238491 260042 238497
rect 259990 238433 260042 238439
rect 260086 234051 260138 234057
rect 260086 233993 260138 233999
rect 259392 233604 259646 233632
rect 259776 233604 259934 233632
rect 260098 233618 260126 233993
rect 260482 233618 260510 244945
rect 261058 244417 261086 246924
rect 261046 244411 261098 244417
rect 261046 244353 261098 244359
rect 261250 241753 261278 246938
rect 261430 245077 261482 245083
rect 261430 245019 261482 245025
rect 261238 241747 261290 241753
rect 261238 241689 261290 241695
rect 260854 233977 260906 233983
rect 260854 233919 260906 233925
rect 260866 233618 260894 233919
rect 261442 233632 261470 245019
rect 261730 238645 261758 246938
rect 262006 246779 262058 246785
rect 262006 246721 262058 246727
rect 261718 238639 261770 238645
rect 261718 238581 261770 238587
rect 261814 234125 261866 234131
rect 261814 234067 261866 234073
rect 261826 233632 261854 234067
rect 262018 233928 262046 246721
rect 262210 241531 262238 246938
rect 262560 246924 262814 246952
rect 262678 245299 262730 245305
rect 262678 245241 262730 245247
rect 262198 241525 262250 241531
rect 262198 241467 262250 241473
rect 262294 234199 262346 234205
rect 262294 234141 262346 234147
rect 261216 233604 261470 233632
rect 261600 233604 261854 233632
rect 261970 233900 262046 233928
rect 261970 233618 261998 233900
rect 262306 233618 262334 234141
rect 262690 233618 262718 245241
rect 262786 242863 262814 246924
rect 262882 246924 263040 246952
rect 262774 242857 262826 242863
rect 262774 242799 262826 242805
rect 262882 241383 262910 246924
rect 263062 245447 263114 245453
rect 263062 245389 263114 245395
rect 262870 241377 262922 241383
rect 262870 241319 262922 241325
rect 263074 233618 263102 245389
rect 263458 238349 263486 246938
rect 263938 242789 263966 246938
rect 263926 242783 263978 242789
rect 263926 242725 263978 242731
rect 264322 241161 264350 246938
rect 264768 246924 264926 246952
rect 264790 243301 264842 243307
rect 264790 243243 264842 243249
rect 264406 241525 264458 241531
rect 264406 241467 264458 241473
rect 264310 241155 264362 241161
rect 264310 241097 264362 241103
rect 264214 238565 264266 238571
rect 264214 238507 264266 238513
rect 263446 238343 263498 238349
rect 263446 238285 263498 238291
rect 264226 238127 264254 238507
rect 264214 238121 264266 238127
rect 264214 238063 264266 238069
rect 264022 234643 264074 234649
rect 264022 234585 264074 234591
rect 263638 234495 263690 234501
rect 263638 234437 263690 234443
rect 263650 233632 263678 234437
rect 264034 233632 264062 234585
rect 264418 233632 264446 241467
rect 264502 239009 264554 239015
rect 264502 238951 264554 238957
rect 263424 233604 263678 233632
rect 263808 233604 264062 233632
rect 264192 233604 264446 233632
rect 264514 233618 264542 238951
rect 264802 233632 264830 243243
rect 264898 238571 264926 246924
rect 264994 246924 265248 246952
rect 265632 246924 265886 246952
rect 264994 241013 265022 246924
rect 265750 243227 265802 243233
rect 265750 243169 265802 243175
rect 264982 241007 265034 241013
rect 264982 240949 265034 240955
rect 264886 238565 264938 238571
rect 264886 238507 264938 238513
rect 265270 236937 265322 236943
rect 265270 236879 265322 236885
rect 264802 233604 264912 233632
rect 265282 233618 265310 236879
rect 265762 233632 265790 243169
rect 265858 242937 265886 246924
rect 265846 242931 265898 242937
rect 265846 242873 265898 242879
rect 266050 240791 266078 246938
rect 266038 240785 266090 240791
rect 266038 240727 266090 240733
rect 266530 238867 266558 246938
rect 266722 246924 266976 246952
rect 267360 246924 267614 246952
rect 266614 243153 266666 243159
rect 266614 243095 266666 243101
rect 266518 238861 266570 238867
rect 266518 238803 266570 238809
rect 266230 237381 266282 237387
rect 266230 237323 266282 237329
rect 266242 233632 266270 237323
rect 266626 233632 266654 243095
rect 266722 240717 266750 246924
rect 267586 244713 267614 246924
rect 267826 246656 267854 246938
rect 267778 246628 267854 246656
rect 267574 244707 267626 244713
rect 267574 244649 267626 244655
rect 267778 241087 267806 246628
rect 268258 244565 268286 246938
rect 268738 244787 268766 246938
rect 268726 244781 268778 244787
rect 268726 244723 268778 244729
rect 268246 244559 268298 244565
rect 268246 244501 268298 244507
rect 268054 243079 268106 243085
rect 268054 243021 268106 243027
rect 267766 241081 267818 241087
rect 267766 241023 267818 241029
rect 266710 240711 266762 240717
rect 266710 240653 266762 240659
rect 266710 237455 266762 237461
rect 266710 237397 266762 237403
rect 265632 233604 265790 233632
rect 266016 233604 266270 233632
rect 266400 233604 266654 233632
rect 266722 233618 266750 237397
rect 267094 237307 267146 237313
rect 267094 237249 267146 237255
rect 267106 233618 267134 237249
rect 267478 237233 267530 237239
rect 267478 237175 267530 237181
rect 267490 233618 267518 237175
rect 268066 233632 268094 243021
rect 268822 243005 268874 243011
rect 268822 242947 268874 242953
rect 268438 239897 268490 239903
rect 268438 239839 268490 239845
rect 268450 233632 268478 239839
rect 268834 233632 268862 242947
rect 268918 242339 268970 242345
rect 268918 242281 268970 242287
rect 267840 233604 268094 233632
rect 268224 233604 268478 233632
rect 268608 233604 268862 233632
rect 268930 233618 268958 242281
rect 269122 238793 269150 246938
rect 269568 246924 269726 246952
rect 269110 238787 269162 238793
rect 269110 238729 269162 238735
rect 269302 237159 269354 237165
rect 269302 237101 269354 237107
rect 269314 233618 269342 237101
rect 269698 237091 269726 246924
rect 269794 246924 270048 246952
rect 269686 237085 269738 237091
rect 269686 237027 269738 237033
rect 269794 237017 269822 246924
rect 270466 244565 270494 246938
rect 270454 244559 270506 244565
rect 270454 244501 270506 244507
rect 270262 242709 270314 242715
rect 270262 242651 270314 242657
rect 269878 242487 269930 242493
rect 269878 242429 269930 242435
rect 269782 237011 269834 237017
rect 269782 236953 269834 236959
rect 269890 233632 269918 242429
rect 270274 233632 270302 242651
rect 270850 238941 270878 246938
rect 271030 241747 271082 241753
rect 271030 241689 271082 241695
rect 270838 238935 270890 238941
rect 270838 238877 270890 238883
rect 270646 236863 270698 236869
rect 270646 236805 270698 236811
rect 270658 233632 270686 236805
rect 271042 233632 271070 241689
rect 271126 241377 271178 241383
rect 271126 241319 271178 241325
rect 269712 233604 269918 233632
rect 270048 233604 270302 233632
rect 270432 233604 270686 233632
rect 270816 233604 271070 233632
rect 271138 233618 271166 241319
rect 271330 238941 271358 246938
rect 271776 246924 272030 246952
rect 272160 246924 272414 246952
rect 271894 241895 271946 241901
rect 271894 241837 271946 241843
rect 271510 240933 271562 240939
rect 271510 240875 271562 240881
rect 271318 238935 271370 238941
rect 271318 238877 271370 238883
rect 271522 233618 271550 240875
rect 271906 233618 271934 241837
rect 272002 241605 272030 246924
rect 271990 241599 272042 241605
rect 271990 241541 272042 241547
rect 272386 233803 272414 246924
rect 272578 241309 272606 246938
rect 272566 241303 272618 241309
rect 272566 241245 272618 241251
rect 272854 241007 272906 241013
rect 272854 240949 272906 240955
rect 272470 240045 272522 240051
rect 272470 239987 272522 239993
rect 272372 233794 272428 233803
rect 272372 233729 272428 233738
rect 272482 233632 272510 239987
rect 272866 233632 272894 240949
rect 273058 239977 273086 246938
rect 273238 245965 273290 245971
rect 273238 245907 273290 245913
rect 273250 241827 273278 245907
rect 273238 241821 273290 241827
rect 273238 241763 273290 241769
rect 273538 241235 273566 246938
rect 273634 246924 273888 246952
rect 274368 246924 274622 246952
rect 273526 241229 273578 241235
rect 273526 241171 273578 241177
rect 273238 240637 273290 240643
rect 273238 240579 273290 240585
rect 273046 239971 273098 239977
rect 273046 239913 273098 239919
rect 273250 233632 273278 240579
rect 273334 240563 273386 240569
rect 273334 240505 273386 240511
rect 272256 233604 272510 233632
rect 272640 233604 272894 233632
rect 273024 233604 273278 233632
rect 273346 233618 273374 240505
rect 273634 240051 273662 246924
rect 273718 241451 273770 241457
rect 273718 241393 273770 241399
rect 273622 240045 273674 240051
rect 273622 239987 273674 239993
rect 273526 239379 273578 239385
rect 273526 239321 273578 239327
rect 273538 236129 273566 239321
rect 273526 236123 273578 236129
rect 273526 236065 273578 236071
rect 273730 233618 273758 241393
rect 274102 239379 274154 239385
rect 274102 239321 274154 239327
rect 274114 233618 274142 239321
rect 274594 237017 274622 246924
rect 274786 239903 274814 246938
rect 275266 242567 275294 246938
rect 275254 242561 275306 242567
rect 275254 242503 275306 242509
rect 275446 241821 275498 241827
rect 275446 241763 275498 241769
rect 274774 239897 274826 239903
rect 274774 239839 274826 239845
rect 275062 239305 275114 239311
rect 275062 239247 275114 239253
rect 274678 239157 274730 239163
rect 274678 239099 274730 239105
rect 274582 237011 274634 237017
rect 274582 236953 274634 236959
rect 274690 233632 274718 239099
rect 275074 233632 275102 239247
rect 275458 233632 275486 241763
rect 275650 241531 275678 246938
rect 276096 246924 276254 246952
rect 276576 246924 276830 246952
rect 275638 241525 275690 241531
rect 275638 241467 275690 241473
rect 275926 241155 275978 241161
rect 275926 241097 275978 241103
rect 275542 240341 275594 240347
rect 275542 240283 275594 240289
rect 274464 233604 274718 233632
rect 274848 233604 275102 233632
rect 275232 233604 275486 233632
rect 275554 233618 275582 240283
rect 275938 233618 275966 241097
rect 276226 239681 276254 246924
rect 276406 246113 276458 246119
rect 276406 246055 276458 246061
rect 276418 240791 276446 246055
rect 276406 240785 276458 240791
rect 276406 240727 276458 240733
rect 276802 240495 276830 246924
rect 276886 240859 276938 240865
rect 276886 240801 276938 240807
rect 276790 240489 276842 240495
rect 276790 240431 276842 240437
rect 276310 239971 276362 239977
rect 276310 239913 276362 239919
rect 276214 239675 276266 239681
rect 276214 239617 276266 239623
rect 276322 233618 276350 239913
rect 276502 238713 276554 238719
rect 276502 238655 276554 238661
rect 276514 238349 276542 238655
rect 276502 238343 276554 238349
rect 276502 238285 276554 238291
rect 276898 233632 276926 240801
rect 276994 239533 277022 246938
rect 277378 241087 277406 246938
rect 277558 246187 277610 246193
rect 277558 246129 277610 246135
rect 277366 241081 277418 241087
rect 277366 241023 277418 241029
rect 277570 239755 277598 246129
rect 277750 240267 277802 240273
rect 277750 240209 277802 240215
rect 277558 239749 277610 239755
rect 277558 239691 277610 239697
rect 277270 239601 277322 239607
rect 277270 239543 277322 239549
rect 276982 239527 277034 239533
rect 276982 239469 277034 239475
rect 277282 233632 277310 239543
rect 277654 239083 277706 239089
rect 277654 239025 277706 239031
rect 277666 233632 277694 239025
rect 276672 233604 276926 233632
rect 277056 233604 277310 233632
rect 277440 233604 277694 233632
rect 277762 233618 277790 240209
rect 277858 239237 277886 246938
rect 278304 246924 278558 246952
rect 278784 246924 279038 246952
rect 278134 244707 278186 244713
rect 278134 244649 278186 244655
rect 278038 244633 278090 244639
rect 278038 244575 278090 244581
rect 277942 244337 277994 244343
rect 277942 244279 277994 244285
rect 277954 242789 277982 244279
rect 278050 242863 278078 244575
rect 278146 242937 278174 244649
rect 278134 242931 278186 242937
rect 278134 242873 278186 242879
rect 278038 242857 278090 242863
rect 278038 242799 278090 242805
rect 277942 242783 277994 242789
rect 277942 242725 277994 242731
rect 278530 240791 278558 246924
rect 278518 240785 278570 240791
rect 278518 240727 278570 240733
rect 278518 240193 278570 240199
rect 278518 240135 278570 240141
rect 278134 239749 278186 239755
rect 278134 239691 278186 239697
rect 277846 239231 277898 239237
rect 277846 239173 277898 239179
rect 277846 238787 277898 238793
rect 277846 238729 277898 238735
rect 277858 238349 277886 238729
rect 277846 238343 277898 238349
rect 277846 238285 277898 238291
rect 277846 237529 277898 237535
rect 277846 237471 277898 237477
rect 277858 236943 277886 237471
rect 277846 236937 277898 236943
rect 277846 236879 277898 236885
rect 278146 233618 278174 239691
rect 278530 233618 278558 240135
rect 279010 240051 279038 246924
rect 279106 240421 279134 246938
rect 279600 246924 279902 246952
rect 279284 245190 279340 245199
rect 279284 245125 279340 245134
rect 279298 244903 279326 245125
rect 279284 244894 279340 244903
rect 279284 244829 279340 244838
rect 279094 240415 279146 240421
rect 279094 240357 279146 240363
rect 279094 240119 279146 240125
rect 279094 240061 279146 240067
rect 278998 240045 279050 240051
rect 278998 239987 279050 239993
rect 278710 238787 278762 238793
rect 278710 238729 278762 238735
rect 278722 237091 278750 238729
rect 278710 237085 278762 237091
rect 278710 237027 278762 237033
rect 279106 233632 279134 240061
rect 279874 239977 279902 246924
rect 280066 240717 280094 246938
rect 280416 246924 280478 246952
rect 280054 240711 280106 240717
rect 280054 240653 280106 240659
rect 280450 240495 280478 246924
rect 280546 246924 280896 246952
rect 280342 240489 280394 240495
rect 280342 240431 280394 240437
rect 280438 240489 280490 240495
rect 280438 240431 280490 240437
rect 279862 239971 279914 239977
rect 279862 239913 279914 239919
rect 279286 239897 279338 239903
rect 279286 239839 279338 239845
rect 279298 233780 279326 239839
rect 279862 239823 279914 239829
rect 279862 239765 279914 239771
rect 278880 233604 279134 233632
rect 279250 233752 279326 233780
rect 279250 233618 279278 233752
rect 279874 233632 279902 239765
rect 280354 239552 280382 240431
rect 280354 239524 280478 239552
rect 280450 239459 280478 239524
rect 280438 239453 280490 239459
rect 280438 239395 280490 239401
rect 280546 234224 280574 246924
rect 281314 241679 281342 246938
rect 281506 246924 281808 246952
rect 281302 241673 281354 241679
rect 281302 241615 281354 241621
rect 280822 240045 280874 240051
rect 280822 239987 280874 239993
rect 280630 239971 280682 239977
rect 280630 239913 280682 239919
rect 280258 234196 280574 234224
rect 280258 233632 280286 234196
rect 280340 233794 280396 233803
rect 280340 233729 280396 233738
rect 279648 233604 279902 233632
rect 279984 233604 280286 233632
rect 280354 233618 280382 233729
rect 280642 233632 280670 239913
rect 280834 233632 280862 239987
rect 281506 239829 281534 246924
rect 282070 242931 282122 242937
rect 282070 242873 282122 242879
rect 281686 240933 281738 240939
rect 281686 240875 281738 240881
rect 281698 240569 281726 240875
rect 281590 240563 281642 240569
rect 281590 240505 281642 240511
rect 281686 240563 281738 240569
rect 281686 240505 281738 240511
rect 281602 239829 281630 240505
rect 281494 239823 281546 239829
rect 281494 239765 281546 239771
rect 281590 239823 281642 239829
rect 281590 239765 281642 239771
rect 281590 239527 281642 239533
rect 281590 239469 281642 239475
rect 281206 239231 281258 239237
rect 281206 239173 281258 239179
rect 281218 233632 281246 239173
rect 281602 233632 281630 239469
rect 282082 233632 282110 242873
rect 282178 239533 282206 246938
rect 282370 246924 282624 246952
rect 283104 246924 283358 246952
rect 282370 239903 282398 246924
rect 282934 242635 282986 242641
rect 282934 242577 282986 242583
rect 282358 239897 282410 239903
rect 282358 239839 282410 239845
rect 282166 239527 282218 239533
rect 282166 239469 282218 239475
rect 282550 239231 282602 239237
rect 282550 239173 282602 239179
rect 280642 233604 280752 233632
rect 280834 233604 281088 233632
rect 281218 233604 281472 233632
rect 281602 233604 281856 233632
rect 282082 233604 282192 233632
rect 282562 233618 282590 239173
rect 282946 233618 282974 242577
rect 283330 241531 283358 246924
rect 283414 242857 283466 242863
rect 283414 242799 283466 242805
rect 283318 241525 283370 241531
rect 283318 241467 283370 241473
rect 283426 233632 283454 242799
rect 283522 240125 283550 246938
rect 283798 242265 283850 242271
rect 283798 242207 283850 242213
rect 283510 240119 283562 240125
rect 283510 240061 283562 240067
rect 283810 233632 283838 242207
rect 283906 240939 283934 246938
rect 283894 240933 283946 240939
rect 283894 240875 283946 240881
rect 284386 240199 284414 246938
rect 284578 246924 284832 246952
rect 285312 246924 285566 246952
rect 284374 240193 284426 240199
rect 284374 240135 284426 240141
rect 284578 239755 284606 246924
rect 285428 241046 285484 241055
rect 285538 241013 285566 246924
rect 285428 240981 285430 240990
rect 285482 240981 285484 240990
rect 285526 241007 285578 241013
rect 285430 240949 285482 240955
rect 285526 240949 285578 240955
rect 284662 240637 284714 240643
rect 284662 240579 284714 240585
rect 284674 239755 284702 240579
rect 285634 240273 285662 246938
rect 286114 241901 286142 246938
rect 286102 241895 286154 241901
rect 286102 241837 286154 241843
rect 286486 241747 286538 241753
rect 286486 241689 286538 241695
rect 286102 241451 286154 241457
rect 286102 241393 286154 241399
rect 286114 241087 286142 241393
rect 286390 241377 286442 241383
rect 286390 241319 286442 241325
rect 286294 241303 286346 241309
rect 286294 241245 286346 241251
rect 286198 241229 286250 241235
rect 286198 241171 286250 241177
rect 286006 241081 286058 241087
rect 286006 241023 286058 241029
rect 286102 241081 286154 241087
rect 286102 241023 286154 241029
rect 285910 240785 285962 240791
rect 285910 240727 285962 240733
rect 285814 240711 285866 240717
rect 285814 240653 285866 240659
rect 285718 240563 285770 240569
rect 285718 240505 285770 240511
rect 285730 240315 285758 240505
rect 285716 240306 285772 240315
rect 285622 240267 285674 240273
rect 285716 240241 285772 240250
rect 285622 240209 285674 240215
rect 285826 239977 285854 240653
rect 285922 240199 285950 240727
rect 285910 240193 285962 240199
rect 285910 240135 285962 240141
rect 286018 240125 286046 241023
rect 286210 240347 286238 241171
rect 286198 240341 286250 240347
rect 286198 240283 286250 240289
rect 286006 240119 286058 240125
rect 286006 240061 286058 240067
rect 286306 240051 286334 241245
rect 286402 240643 286430 241319
rect 286498 241087 286526 241689
rect 286486 241081 286538 241087
rect 286486 241023 286538 241029
rect 286390 240637 286442 240643
rect 286390 240579 286442 240585
rect 286294 240045 286346 240051
rect 286294 239987 286346 239993
rect 285814 239971 285866 239977
rect 285814 239913 285866 239919
rect 285428 239862 285484 239871
rect 285428 239797 285484 239806
rect 284566 239749 284618 239755
rect 284566 239691 284618 239697
rect 284662 239749 284714 239755
rect 284662 239691 284714 239697
rect 285238 239675 285290 239681
rect 285238 239617 285290 239623
rect 284278 236863 284330 236869
rect 284278 236805 284330 236811
rect 284290 233632 284318 236805
rect 284758 236789 284810 236795
rect 284758 236731 284810 236737
rect 284374 236715 284426 236721
rect 284374 236657 284426 236663
rect 283296 233604 283454 233632
rect 283680 233604 283838 233632
rect 284064 233604 284318 233632
rect 284386 233618 284414 236657
rect 284770 233618 284798 236731
rect 285142 236641 285194 236647
rect 285142 236583 285194 236589
rect 285154 233618 285182 236583
rect 285250 233632 285278 239617
rect 285442 239385 285470 239797
rect 285430 239379 285482 239385
rect 285430 239321 285482 239327
rect 286594 239089 286622 246938
rect 287040 246924 287102 246952
rect 286774 242043 286826 242049
rect 286774 241985 286826 241991
rect 286678 241451 286730 241457
rect 286678 241393 286730 241399
rect 286690 241055 286718 241393
rect 286786 241309 286814 241985
rect 286774 241303 286826 241309
rect 286774 241245 286826 241251
rect 287074 241235 287102 246924
rect 287170 246924 287424 246952
rect 287062 241229 287114 241235
rect 287062 241171 287114 241177
rect 286676 241046 286732 241055
rect 286676 240981 286732 240990
rect 287170 239607 287198 246924
rect 287638 244263 287690 244269
rect 287638 244205 287690 244211
rect 287350 240859 287402 240865
rect 287350 240801 287402 240807
rect 287158 239601 287210 239607
rect 287158 239543 287210 239549
rect 286582 239083 286634 239089
rect 286582 239025 286634 239031
rect 286966 237085 287018 237091
rect 286966 237027 287018 237033
rect 286102 236567 286154 236573
rect 286102 236509 286154 236515
rect 286114 233632 286142 236509
rect 286582 236419 286634 236425
rect 286582 236361 286634 236367
rect 286486 236271 286538 236277
rect 286486 236213 286538 236219
rect 286498 233632 286526 236213
rect 285250 233604 285504 233632
rect 285888 233604 286142 233632
rect 286272 233604 286526 233632
rect 286594 233618 286622 236361
rect 286978 233618 287006 237027
rect 287362 233618 287390 240801
rect 287650 233928 287678 244205
rect 287734 242117 287786 242123
rect 287734 242059 287786 242065
rect 287746 239237 287774 242059
rect 287842 240791 287870 246938
rect 288118 241599 288170 241605
rect 288118 241541 288170 241547
rect 287830 240785 287882 240791
rect 287830 240727 287882 240733
rect 287734 239231 287786 239237
rect 287734 239173 287786 239179
rect 288022 239231 288074 239237
rect 288022 239173 288074 239179
rect 287926 239157 287978 239163
rect 288034 239145 288062 239173
rect 287978 239117 288062 239145
rect 287926 239099 287978 239105
rect 287650 233900 287726 233928
rect 287698 233618 287726 233900
rect 288130 233780 288158 241541
rect 288322 240717 288350 246938
rect 288310 240711 288362 240717
rect 288310 240653 288362 240659
rect 288502 240341 288554 240347
rect 288502 240283 288554 240289
rect 288598 240341 288650 240347
rect 288598 240283 288650 240289
rect 288514 239163 288542 240283
rect 288610 240199 288638 240283
rect 288706 240199 288734 246938
rect 289152 246924 289406 246952
rect 289270 240563 289322 240569
rect 289270 240505 289322 240511
rect 288598 240193 288650 240199
rect 288598 240135 288650 240141
rect 288694 240193 288746 240199
rect 288694 240135 288746 240141
rect 289282 239829 289310 240505
rect 289378 239829 289406 246924
rect 289474 246924 289632 246952
rect 289474 241383 289502 246924
rect 289846 241895 289898 241901
rect 289846 241837 289898 241843
rect 289942 241895 289994 241901
rect 289942 241837 289994 241843
rect 289750 241747 289802 241753
rect 289750 241689 289802 241695
rect 289762 241531 289790 241689
rect 289750 241525 289802 241531
rect 289750 241467 289802 241473
rect 289462 241377 289514 241383
rect 289462 241319 289514 241325
rect 289750 241377 289802 241383
rect 289750 241319 289802 241325
rect 289558 240711 289610 240717
rect 289558 240653 289610 240659
rect 289270 239823 289322 239829
rect 289270 239765 289322 239771
rect 289366 239823 289418 239829
rect 289366 239765 289418 239771
rect 288694 239601 288746 239607
rect 288694 239543 288746 239549
rect 288502 239157 288554 239163
rect 288502 239099 288554 239105
rect 288082 233752 288158 233780
rect 288082 233618 288110 233752
rect 288706 233632 288734 239543
rect 288790 239453 288842 239459
rect 288790 239395 288842 239401
rect 288480 233604 288734 233632
rect 288802 233618 288830 239395
rect 289570 233780 289598 240653
rect 289474 233752 289598 233780
rect 289474 233632 289502 233752
rect 289762 233632 289790 241319
rect 289858 241055 289886 241837
rect 289954 241679 289982 241837
rect 289942 241673 289994 241679
rect 289942 241615 289994 241621
rect 289844 241046 289900 241055
rect 289844 240981 289900 240990
rect 290050 239385 290078 246938
rect 290134 241673 290186 241679
rect 290134 241615 290186 241621
rect 290038 239379 290090 239385
rect 290038 239321 290090 239327
rect 290146 233632 290174 241615
rect 290434 239903 290462 246938
rect 290710 241525 290762 241531
rect 290710 241467 290762 241473
rect 290722 241013 290750 241467
rect 290710 241007 290762 241013
rect 290710 240949 290762 240955
rect 290806 241007 290858 241013
rect 290806 240949 290858 240955
rect 290818 240791 290846 240949
rect 290806 240785 290858 240791
rect 290806 240727 290858 240733
rect 290422 239897 290474 239903
rect 290422 239839 290474 239845
rect 290518 239897 290570 239903
rect 290518 239839 290570 239845
rect 290530 239459 290558 239839
rect 290914 239755 290942 246938
rect 291106 246924 291360 246952
rect 291840 246924 292094 246952
rect 291106 241827 291134 246924
rect 291094 241821 291146 241827
rect 291094 241763 291146 241769
rect 291286 241821 291338 241827
rect 291286 241763 291338 241769
rect 291298 241235 291326 241763
rect 291286 241229 291338 241235
rect 291286 241171 291338 241177
rect 291382 241229 291434 241235
rect 291382 241171 291434 241177
rect 290998 240785 291050 240791
rect 290998 240727 291050 240733
rect 290806 239749 290858 239755
rect 290806 239691 290858 239697
rect 290902 239749 290954 239755
rect 290902 239691 290954 239697
rect 290818 239459 290846 239691
rect 290518 239453 290570 239459
rect 290518 239395 290570 239401
rect 290806 239453 290858 239459
rect 290806 239395 290858 239401
rect 290518 236345 290570 236351
rect 290518 236287 290570 236293
rect 290530 233632 290558 236287
rect 290806 236197 290858 236203
rect 290806 236139 290858 236145
rect 290818 233632 290846 236139
rect 289200 233604 289502 233632
rect 289584 233604 289790 233632
rect 289920 233604 290174 233632
rect 290304 233604 290558 233632
rect 290688 233604 290846 233632
rect 291010 233618 291038 240727
rect 291394 233618 291422 241171
rect 292066 240125 292094 246924
rect 292054 240119 292106 240125
rect 292054 240061 292106 240067
rect 291862 240045 291914 240051
rect 291862 239987 291914 239993
rect 291874 239700 291902 239987
rect 291874 239672 291998 239700
rect 291970 239607 291998 239672
rect 291958 239601 292010 239607
rect 291958 239543 292010 239549
rect 291670 239527 291722 239533
rect 291670 239469 291722 239475
rect 291682 236592 291710 239469
rect 292162 239311 292190 246938
rect 292642 239903 292670 246938
rect 293014 242191 293066 242197
rect 293014 242133 293066 242139
rect 292726 242043 292778 242049
rect 292726 241985 292778 241991
rect 292246 239897 292298 239903
rect 292246 239839 292298 239845
rect 292630 239897 292682 239903
rect 292630 239839 292682 239845
rect 292258 239311 292286 239839
rect 292150 239305 292202 239311
rect 292150 239247 292202 239253
rect 292246 239305 292298 239311
rect 292246 239247 292298 239253
rect 291682 236564 291902 236592
rect 291766 236493 291818 236499
rect 291766 236435 291818 236441
rect 291778 233618 291806 236435
rect 291874 233632 291902 236564
rect 292738 233632 292766 241985
rect 293026 233632 293054 242133
rect 293122 239237 293150 246938
rect 293314 246924 293568 246952
rect 293952 246924 294206 246952
rect 293206 242413 293258 242419
rect 293206 242355 293258 242361
rect 293110 239231 293162 239237
rect 293110 239173 293162 239179
rect 291874 233604 292128 233632
rect 292512 233604 292766 233632
rect 292896 233604 293054 233632
rect 293218 233618 293246 242355
rect 293314 239871 293342 246924
rect 293590 242783 293642 242789
rect 293590 242725 293642 242731
rect 293300 239862 293356 239871
rect 293300 239797 293356 239806
rect 293602 233618 293630 242725
rect 294070 240341 294122 240347
rect 294070 240283 294122 240289
rect 293974 240045 294026 240051
rect 293974 239987 294026 239993
rect 293986 233618 294014 239987
rect 294082 233632 294110 240283
rect 294178 239237 294206 246924
rect 294370 241161 294398 246938
rect 294358 241155 294410 241161
rect 294358 241097 294410 241103
rect 294454 241155 294506 241161
rect 294454 241097 294506 241103
rect 294466 241055 294494 241097
rect 294452 241046 294508 241055
rect 294452 240981 294508 240990
rect 294454 240415 294506 240421
rect 294454 240357 294506 240363
rect 294166 239231 294218 239237
rect 294166 239173 294218 239179
rect 294466 233632 294494 240357
rect 294850 239089 294878 246938
rect 294934 244263 294986 244269
rect 294934 244205 294986 244211
rect 294946 243085 294974 244205
rect 294934 243079 294986 243085
rect 294934 243021 294986 243027
rect 295126 243005 295178 243011
rect 295126 242947 295178 242953
rect 295138 242715 295166 242947
rect 295126 242709 295178 242715
rect 295126 242651 295178 242657
rect 295330 240569 295358 246938
rect 295680 246924 295934 246952
rect 295798 241895 295850 241901
rect 295798 241837 295850 241843
rect 295318 240563 295370 240569
rect 295318 240505 295370 240511
rect 295414 240489 295466 240495
rect 295414 240431 295466 240437
rect 294934 239971 294986 239977
rect 294934 239913 294986 239919
rect 294838 239083 294890 239089
rect 294838 239025 294890 239031
rect 294946 233632 294974 239913
rect 294082 233604 294336 233632
rect 294466 233604 294720 233632
rect 294946 233604 295104 233632
rect 295426 233618 295454 240431
rect 295810 233618 295838 241837
rect 295906 240051 295934 246924
rect 296002 246924 296160 246952
rect 295894 240045 295946 240051
rect 295894 239987 295946 239993
rect 296002 239459 296030 246924
rect 296278 241747 296330 241753
rect 296278 241689 296330 241695
rect 296182 239675 296234 239681
rect 296182 239617 296234 239623
rect 295990 239453 296042 239459
rect 295990 239395 296042 239401
rect 296194 233618 296222 239617
rect 296290 233632 296318 241689
rect 296578 239977 296606 246938
rect 296660 245042 296716 245051
rect 296660 244977 296716 244986
rect 296674 244903 296702 244977
rect 296660 244894 296716 244903
rect 296660 244829 296716 244838
rect 296662 242783 296714 242789
rect 296662 242725 296714 242731
rect 296674 241975 296702 242725
rect 296662 241969 296714 241975
rect 296662 241911 296714 241917
rect 296962 241457 296990 246938
rect 296950 241451 297002 241457
rect 296950 241393 297002 241399
rect 296662 240933 296714 240939
rect 296662 240875 296714 240881
rect 296566 239971 296618 239977
rect 296566 239913 296618 239919
rect 296674 233632 296702 240875
rect 297442 239681 297470 246938
rect 297888 246924 298046 246952
rect 297622 241525 297674 241531
rect 297622 241467 297674 241473
rect 297430 239675 297482 239681
rect 297430 239617 297482 239623
rect 297046 239601 297098 239607
rect 297046 239543 297098 239549
rect 297058 233632 297086 239543
rect 296290 233604 296544 233632
rect 296674 233604 296928 233632
rect 297058 233604 297312 233632
rect 297634 233618 297662 241467
rect 297718 241155 297770 241161
rect 297718 241097 297770 241103
rect 297730 233632 297758 241097
rect 298018 239533 298046 246924
rect 298354 246656 298382 246938
rect 298752 246924 299006 246952
rect 298306 246628 298382 246656
rect 298102 242857 298154 242863
rect 298102 242799 298154 242805
rect 298114 242271 298142 242799
rect 298198 242783 298250 242789
rect 298198 242725 298250 242731
rect 298102 242265 298154 242271
rect 298102 242207 298154 242213
rect 298210 242123 298238 242725
rect 298198 242117 298250 242123
rect 298198 242059 298250 242065
rect 298306 241309 298334 246628
rect 298390 241821 298442 241827
rect 298390 241763 298442 241769
rect 298294 241303 298346 241309
rect 298294 241245 298346 241251
rect 298006 239527 298058 239533
rect 298006 239469 298058 239475
rect 297730 233604 298032 233632
rect 298402 233618 298430 241763
rect 298486 241007 298538 241013
rect 298486 240949 298538 240955
rect 298498 233632 298526 240949
rect 298978 240199 299006 246924
rect 299170 240315 299198 246938
rect 299156 240306 299212 240315
rect 299156 240241 299212 240250
rect 298870 240193 298922 240199
rect 298870 240135 298922 240141
rect 298966 240193 299018 240199
rect 298966 240135 299018 240141
rect 298882 233632 298910 240135
rect 299650 239829 299678 246938
rect 299842 246924 300096 246952
rect 300480 246924 300734 246952
rect 299842 240643 299870 246924
rect 300022 241377 300074 241383
rect 300022 241319 300074 241325
rect 300034 240717 300062 241319
rect 300022 240711 300074 240717
rect 300022 240653 300074 240659
rect 299830 240637 299882 240643
rect 299830 240579 299882 240585
rect 300706 240125 300734 246924
rect 300802 246924 300960 246952
rect 300802 241087 300830 246924
rect 301174 241303 301226 241309
rect 301174 241245 301226 241251
rect 301078 241155 301130 241161
rect 301078 241097 301130 241103
rect 300790 241081 300842 241087
rect 300790 241023 300842 241029
rect 300598 240119 300650 240125
rect 300598 240061 300650 240067
rect 300694 240119 300746 240125
rect 300694 240061 300746 240067
rect 299254 239823 299306 239829
rect 299254 239765 299306 239771
rect 299638 239823 299690 239829
rect 299638 239765 299690 239771
rect 299266 233632 299294 239765
rect 300214 239749 300266 239755
rect 300214 239691 300266 239697
rect 299830 239379 299882 239385
rect 299830 239321 299882 239327
rect 298498 233604 298752 233632
rect 298882 233604 299136 233632
rect 299266 233604 299520 233632
rect 299842 233618 299870 239321
rect 300226 233618 300254 239691
rect 300610 233618 300638 240061
rect 300694 239897 300746 239903
rect 300694 239839 300746 239845
rect 300706 233632 300734 239839
rect 301090 239607 301118 241097
rect 301078 239601 301130 239607
rect 301078 239543 301130 239549
rect 301186 239311 301214 241245
rect 301378 239903 301406 246938
rect 301366 239897 301418 239903
rect 301366 239839 301418 239845
rect 301174 239305 301226 239311
rect 301174 239247 301226 239253
rect 301462 239231 301514 239237
rect 301462 239173 301514 239179
rect 301078 239157 301130 239163
rect 301078 239099 301130 239105
rect 301090 233632 301118 239099
rect 301474 233632 301502 239173
rect 301858 236943 301886 246938
rect 302242 243011 302270 246938
rect 302688 246924 302942 246952
rect 302230 243005 302282 243011
rect 302230 242947 302282 242953
rect 302518 241081 302570 241087
rect 302518 241023 302570 241029
rect 302326 240341 302378 240347
rect 302146 240301 302326 240329
rect 302038 239083 302090 239089
rect 302038 239025 302090 239031
rect 301846 236937 301898 236943
rect 301846 236879 301898 236885
rect 300706 233604 300960 233632
rect 301090 233604 301344 233632
rect 301474 233604 301728 233632
rect 302050 233618 302078 239025
rect 302146 237091 302174 240301
rect 302326 240283 302378 240289
rect 302530 240273 302558 241023
rect 302518 240267 302570 240273
rect 302518 240209 302570 240215
rect 302422 240193 302474 240199
rect 302422 240135 302474 240141
rect 302134 237085 302186 237091
rect 302134 237027 302186 237033
rect 302434 236943 302462 240135
rect 302518 240045 302570 240051
rect 302518 239987 302570 239993
rect 302422 236937 302474 236943
rect 302422 236879 302474 236885
rect 302530 233632 302558 239987
rect 302914 239977 302942 246924
rect 303010 246924 303168 246952
rect 303010 242493 303038 246924
rect 302998 242487 303050 242493
rect 302998 242429 303050 242435
rect 303586 240051 303614 246938
rect 303574 240045 303626 240051
rect 303574 239987 303626 239993
rect 302806 239971 302858 239977
rect 302806 239913 302858 239919
rect 302902 239971 302954 239977
rect 302902 239913 302954 239919
rect 302448 233604 302558 233632
rect 302818 233618 302846 239913
rect 302902 239675 302954 239681
rect 302902 239617 302954 239623
rect 302914 233632 302942 239617
rect 303286 239527 303338 239533
rect 303286 239469 303338 239475
rect 303298 233632 303326 239469
rect 303970 237165 303998 246938
rect 304246 239823 304298 239829
rect 304246 239765 304298 239771
rect 303958 237159 304010 237165
rect 303958 237101 304010 237107
rect 303670 236937 303722 236943
rect 303670 236879 303722 236885
rect 303682 233632 303710 236879
rect 302914 233604 303168 233632
rect 303298 233604 303552 233632
rect 303682 233604 303936 233632
rect 304258 233618 304286 239765
rect 304450 239385 304478 246938
rect 304642 246924 304896 246952
rect 305218 246924 305280 246952
rect 304642 242345 304670 246924
rect 304630 242339 304682 242345
rect 304630 242281 304682 242287
rect 304630 240119 304682 240125
rect 304630 240061 304682 240067
rect 304438 239379 304490 239385
rect 304438 239321 304490 239327
rect 304642 233618 304670 240061
rect 305014 239897 305066 239903
rect 305014 239839 305066 239845
rect 305026 233618 305054 239839
rect 305218 239681 305246 246924
rect 305698 243085 305726 246938
rect 306192 246924 306590 246952
rect 306672 246924 306878 246952
rect 305686 243079 305738 243085
rect 305686 243021 305738 243027
rect 305878 240045 305930 240051
rect 305878 239987 305930 239993
rect 305494 239971 305546 239977
rect 305494 239913 305546 239919
rect 305206 239675 305258 239681
rect 305206 239617 305258 239623
rect 305398 237011 305450 237017
rect 305398 236953 305450 236959
rect 216502 233549 216554 233555
rect 210166 223247 210218 223253
rect 210166 223189 210218 223195
rect 210166 218585 210218 218591
rect 210166 218527 210218 218533
rect 210178 217005 210206 218527
rect 210164 216996 210220 217005
rect 210164 216931 210220 216940
rect 210166 215921 210218 215927
rect 210166 215863 210218 215869
rect 210178 213749 210206 215863
rect 210164 213740 210220 213749
rect 210164 213675 210220 213684
rect 210274 208620 210302 233549
rect 212770 233521 212798 233549
rect 305410 233484 305438 236953
rect 305506 233632 305534 239913
rect 305890 233632 305918 239987
rect 306454 239379 306506 239385
rect 306454 239321 306506 239327
rect 305506 233604 305760 233632
rect 305890 233604 306144 233632
rect 306466 233618 306494 239321
rect 306562 233803 306590 246924
rect 306646 239675 306698 239681
rect 306646 239617 306698 239623
rect 306548 233794 306604 233803
rect 306548 233729 306604 233738
rect 306658 233632 306686 239617
rect 306850 234076 306878 246924
rect 306994 246656 307022 246938
rect 307488 246924 307742 246952
rect 306946 246628 307022 246656
rect 306946 244269 306974 246628
rect 306934 244263 306986 244269
rect 306934 244205 306986 244211
rect 307030 244263 307082 244269
rect 307030 244205 307082 244211
rect 307042 241975 307070 244205
rect 307030 241969 307082 241975
rect 307030 241911 307082 241917
rect 306850 234048 307358 234076
rect 306932 233646 306988 233655
rect 306658 233604 306864 233632
rect 307330 233632 307358 234048
rect 307714 233632 307742 246924
rect 307906 237239 307934 246938
rect 307894 237233 307946 237239
rect 307894 237175 307946 237181
rect 308386 233928 308414 246938
rect 308770 237313 308798 246938
rect 308962 246924 309216 246952
rect 309538 246924 309696 246952
rect 309826 246924 310128 246952
rect 308758 237307 308810 237313
rect 308758 237249 308810 237255
rect 308338 233900 308414 233928
rect 306988 233604 307248 233632
rect 307330 233604 307584 233632
rect 307714 233604 307968 233632
rect 308338 233618 308366 233900
rect 308962 233632 308990 246924
rect 309430 242561 309482 242567
rect 309430 242503 309482 242509
rect 309334 239971 309386 239977
rect 309334 239913 309386 239919
rect 309346 233632 309374 239913
rect 308688 233604 308990 233632
rect 309072 233604 309374 233632
rect 309442 233618 309470 242503
rect 309538 237461 309566 246924
rect 309826 239977 309854 246924
rect 310498 243159 310526 246938
rect 310486 243153 310538 243159
rect 310486 243095 310538 243101
rect 310870 240045 310922 240051
rect 310870 239987 310922 239993
rect 309814 239971 309866 239977
rect 309814 239913 309866 239919
rect 310006 239971 310058 239977
rect 310006 239913 310058 239919
rect 309526 237455 309578 237461
rect 309526 237397 309578 237403
rect 310018 233632 310046 239913
rect 310774 239675 310826 239681
rect 310774 239617 310826 239623
rect 310390 239527 310442 239533
rect 310390 239469 310442 239475
rect 310402 233632 310430 239469
rect 310786 233632 310814 239617
rect 309792 233604 310046 233632
rect 310176 233604 310430 233632
rect 310560 233604 310814 233632
rect 310882 233618 310910 239987
rect 310978 237387 311006 246938
rect 311170 246924 311424 246952
rect 311650 246924 311904 246952
rect 311170 239977 311198 246924
rect 311650 243233 311678 246924
rect 311638 243227 311690 243233
rect 311638 243169 311690 243175
rect 311158 239971 311210 239977
rect 311158 239913 311210 239919
rect 311638 239971 311690 239977
rect 311638 239913 311690 239919
rect 311254 239823 311306 239829
rect 311254 239765 311306 239771
rect 310966 237381 311018 237387
rect 310966 237323 311018 237329
rect 311266 233618 311294 239765
rect 311650 233618 311678 239913
rect 312226 239533 312254 246938
rect 312214 239527 312266 239533
rect 312214 239469 312266 239475
rect 312706 237535 312734 246938
rect 312982 243079 313034 243085
rect 312982 243021 313034 243027
rect 312694 237529 312746 237535
rect 312694 237471 312746 237477
rect 312598 237011 312650 237017
rect 312598 236953 312650 236959
rect 312214 236937 312266 236943
rect 312214 236879 312266 236885
rect 312226 233632 312254 236879
rect 312610 233632 312638 236953
rect 312994 233632 313022 243021
rect 313186 239681 313214 246938
rect 313282 246924 313536 246952
rect 313954 246924 314016 246952
rect 313282 243307 313310 246924
rect 313270 243301 313322 243307
rect 313270 243243 313322 243249
rect 313462 242339 313514 242345
rect 313462 242281 313514 242287
rect 313174 239675 313226 239681
rect 313174 239617 313226 239623
rect 313078 237159 313130 237165
rect 313078 237101 313130 237107
rect 312000 233604 312254 233632
rect 312384 233604 312638 233632
rect 312768 233604 313022 233632
rect 313090 233618 313118 237101
rect 313474 233618 313502 242281
rect 313954 240051 313982 246924
rect 313942 240045 313994 240051
rect 313942 239987 313994 239993
rect 314434 239015 314462 246938
rect 314806 242265 314858 242271
rect 314806 242207 314858 242213
rect 314422 239009 314474 239015
rect 314422 238951 314474 238957
rect 313846 237307 313898 237313
rect 313846 237249 313898 237255
rect 313858 233618 313886 237249
rect 314422 237085 314474 237091
rect 314422 237027 314474 237033
rect 314434 233632 314462 237027
rect 314818 233632 314846 242207
rect 314914 239829 314942 246938
rect 315298 240865 315326 246938
rect 315490 246924 315744 246952
rect 315970 246924 316224 246952
rect 315490 241161 315518 246924
rect 315574 243227 315626 243233
rect 315574 243169 315626 243175
rect 315478 241155 315530 241161
rect 315478 241097 315530 241103
rect 315286 240859 315338 240865
rect 315286 240801 315338 240807
rect 314902 239823 314954 239829
rect 314902 239765 314954 239771
rect 315190 237381 315242 237387
rect 315190 237323 315242 237329
rect 315202 233632 315230 237323
rect 315586 233632 315614 243169
rect 315970 241087 315998 246924
rect 316534 243301 316586 243307
rect 316534 243243 316586 243249
rect 315958 241081 316010 241087
rect 315958 241023 316010 241029
rect 315670 240637 315722 240643
rect 315670 240579 315722 240585
rect 314208 233604 314462 233632
rect 314592 233604 314846 233632
rect 314976 233604 315230 233632
rect 315312 233604 315614 233632
rect 315682 233618 315710 240579
rect 316054 237529 316106 237535
rect 316054 237471 316106 237477
rect 316066 233618 316094 237471
rect 316546 233632 316574 243243
rect 316642 241309 316670 246938
rect 316726 242857 316778 242863
rect 316726 242799 316778 242805
rect 316738 242641 316766 242799
rect 316726 242635 316778 242641
rect 316726 242577 316778 242583
rect 316630 241303 316682 241309
rect 316630 241245 316682 241251
rect 316822 237455 316874 237461
rect 316822 237397 316874 237403
rect 316834 233780 316862 237397
rect 317026 236425 317054 246938
rect 317206 242857 317258 242863
rect 317206 242799 317258 242805
rect 317218 242641 317246 242799
rect 317206 242635 317258 242641
rect 317206 242577 317258 242583
rect 317506 240569 317534 246938
rect 317698 246924 317952 246952
rect 318370 246924 318432 246952
rect 317494 240563 317546 240569
rect 317494 240505 317546 240511
rect 317398 237233 317450 237239
rect 317398 237175 317450 237181
rect 317014 236419 317066 236425
rect 317014 236361 317066 236367
rect 316416 233604 316574 233632
rect 316786 233752 316862 233780
rect 316786 233618 316814 233752
rect 317410 233632 317438 237175
rect 317698 236277 317726 246924
rect 318262 244781 318314 244787
rect 318262 244723 318314 244729
rect 318070 244707 318122 244713
rect 318070 244649 318122 244655
rect 318082 242641 318110 244649
rect 318166 244559 318218 244565
rect 318166 244501 318218 244507
rect 318070 242635 318122 242641
rect 318070 242577 318122 242583
rect 318178 242419 318206 244501
rect 318274 242789 318302 244723
rect 318262 242783 318314 242789
rect 318262 242725 318314 242731
rect 318166 242413 318218 242419
rect 318166 242355 318218 242361
rect 318262 241747 318314 241753
rect 318262 241689 318314 241695
rect 317878 241525 317930 241531
rect 317878 241467 317930 241473
rect 317782 241081 317834 241087
rect 317782 241023 317834 241029
rect 317686 236271 317738 236277
rect 317686 236213 317738 236219
rect 317794 233632 317822 241023
rect 317184 233604 317438 233632
rect 317520 233604 317822 233632
rect 317890 233618 317918 241467
rect 318274 233618 318302 241689
rect 318370 240717 318398 246924
rect 318358 240711 318410 240717
rect 318358 240653 318410 240659
rect 318754 236573 318782 246938
rect 318838 241673 318890 241679
rect 318838 241615 318890 241621
rect 318742 236567 318794 236573
rect 318742 236509 318794 236515
rect 318850 233632 318878 241615
rect 319234 241013 319262 246938
rect 319222 241007 319274 241013
rect 319222 240949 319274 240955
rect 319222 240563 319274 240569
rect 319222 240505 319274 240511
rect 319234 233632 319262 240505
rect 319606 239305 319658 239311
rect 319606 239247 319658 239253
rect 319714 239256 319742 246938
rect 320050 246656 320078 246938
rect 320002 246628 320078 246656
rect 320290 246924 320544 246952
rect 319618 233632 319646 239247
rect 319714 239228 319934 239256
rect 319702 239157 319754 239163
rect 319702 239099 319754 239105
rect 318624 233604 318878 233632
rect 319008 233604 319262 233632
rect 319392 233604 319646 233632
rect 319714 233618 319742 239099
rect 319906 236351 319934 239228
rect 320002 236647 320030 246628
rect 320086 239601 320138 239607
rect 320086 239543 320138 239549
rect 319990 236641 320042 236647
rect 319990 236583 320042 236589
rect 319894 236345 319946 236351
rect 319894 236287 319946 236293
rect 320098 233618 320126 239543
rect 320290 236203 320318 246924
rect 320470 242117 320522 242123
rect 320470 242059 320522 242065
rect 320278 236197 320330 236203
rect 320278 236139 320330 236145
rect 320482 233618 320510 242059
rect 320962 236795 320990 246938
rect 321442 240791 321470 246938
rect 321538 246924 321840 246952
rect 322018 246924 322272 246952
rect 322594 246924 322752 246952
rect 321430 240785 321482 240791
rect 321430 240727 321482 240733
rect 321430 240415 321482 240421
rect 321430 240357 321482 240363
rect 321046 239675 321098 239681
rect 321046 239617 321098 239623
rect 320950 236789 321002 236795
rect 320950 236731 321002 236737
rect 321058 233632 321086 239617
rect 321442 233632 321470 240357
rect 321538 236721 321566 246924
rect 322018 240939 322046 246924
rect 322006 240933 322058 240939
rect 322006 240875 322058 240881
rect 321910 239897 321962 239903
rect 321910 239839 321962 239845
rect 321814 239749 321866 239755
rect 321814 239691 321866 239697
rect 321526 236715 321578 236721
rect 321526 236657 321578 236663
rect 321826 233632 321854 239691
rect 320832 233604 321086 233632
rect 321216 233604 321470 233632
rect 321600 233604 321854 233632
rect 321922 233618 321950 239839
rect 322294 239823 322346 239829
rect 322294 239765 322346 239771
rect 322306 233618 322334 239765
rect 322594 236869 322622 246924
rect 322678 239231 322730 239237
rect 322678 239173 322730 239179
rect 322582 236863 322634 236869
rect 322582 236805 322634 236811
rect 322690 233618 322718 239173
rect 323170 236499 323198 246938
rect 323554 242863 323582 246938
rect 323542 242857 323594 242863
rect 323542 242799 323594 242805
rect 324034 242715 324062 246938
rect 324226 246924 324480 246952
rect 324706 246924 324960 246952
rect 324022 242709 324074 242715
rect 324022 242651 324074 242657
rect 324226 242049 324254 246924
rect 324706 242567 324734 246924
rect 324694 242561 324746 242567
rect 324694 242503 324746 242509
rect 325282 242197 325310 246938
rect 325462 244559 325514 244565
rect 325462 244501 325514 244507
rect 325474 244436 325502 244501
rect 325378 244408 325502 244436
rect 325378 244269 325406 244408
rect 325366 244263 325418 244269
rect 325366 244205 325418 244211
rect 325462 244263 325514 244269
rect 325462 244205 325514 244211
rect 325270 242191 325322 242197
rect 325270 242133 325322 242139
rect 324214 242043 324266 242049
rect 324214 241985 324266 241991
rect 325474 241795 325502 244205
rect 325762 242937 325790 246938
rect 325750 242931 325802 242937
rect 325750 242873 325802 242879
rect 326242 242493 326270 246938
rect 326338 246924 326688 246952
rect 326818 246924 327072 246952
rect 326338 243011 326366 246924
rect 326818 244565 326846 246924
rect 326806 244559 326858 244565
rect 326806 244501 326858 244507
rect 326614 243153 326666 243159
rect 326614 243095 326666 243101
rect 326422 243079 326474 243085
rect 326474 243039 326558 243067
rect 326422 243021 326474 243027
rect 326530 243011 326558 243039
rect 326326 243005 326378 243011
rect 326326 242947 326378 242953
rect 326518 243005 326570 243011
rect 326518 242947 326570 242953
rect 326230 242487 326282 242493
rect 326230 242429 326282 242435
rect 326626 242345 326654 243095
rect 326710 243079 326762 243085
rect 326710 243021 326762 243027
rect 326614 242339 326666 242345
rect 326614 242281 326666 242287
rect 326722 242271 326750 243021
rect 326710 242265 326762 242271
rect 326710 242207 326762 242213
rect 325460 241786 325516 241795
rect 325460 241721 325516 241730
rect 324502 240859 324554 240865
rect 324502 240801 324554 240807
rect 323638 240637 323690 240643
rect 323638 240579 323690 240585
rect 323254 240045 323306 240051
rect 323254 239987 323306 239993
rect 323158 236493 323210 236499
rect 323158 236435 323210 236441
rect 323266 233632 323294 239987
rect 323650 233632 323678 240579
rect 324118 240489 324170 240495
rect 324118 240431 324170 240437
rect 324022 240119 324074 240125
rect 324022 240061 324074 240067
rect 324034 233632 324062 240061
rect 323040 233604 323294 233632
rect 323424 233604 323678 233632
rect 323808 233604 324062 233632
rect 324130 233618 324158 240431
rect 324514 233618 324542 240801
rect 326710 240711 326762 240717
rect 326710 240653 326762 240659
rect 326230 240341 326282 240347
rect 326230 240283 326282 240289
rect 324886 240267 324938 240273
rect 324886 240209 324938 240215
rect 324898 233618 324926 240209
rect 325846 240193 325898 240199
rect 325846 240135 325898 240141
rect 325460 239714 325516 239723
rect 325460 239649 325516 239658
rect 325366 239453 325418 239459
rect 325366 239395 325418 239401
rect 325378 233632 325406 239395
rect 325474 239015 325502 239649
rect 325462 239009 325514 239015
rect 325462 238951 325514 238957
rect 325858 233632 325886 240135
rect 326242 233632 326270 240283
rect 326326 239379 326378 239385
rect 326326 239321 326378 239327
rect 325248 233604 325406 233632
rect 325632 233604 325886 233632
rect 326016 233604 326270 233632
rect 326338 233618 326366 239321
rect 326722 233618 326750 240653
rect 327490 239977 327518 246938
rect 327970 246859 327998 246938
rect 327958 246853 328010 246859
rect 327958 246795 328010 246801
rect 327574 241303 327626 241309
rect 327574 241245 327626 241251
rect 327478 239971 327530 239977
rect 327478 239913 327530 239919
rect 327094 239083 327146 239089
rect 327094 239025 327146 239031
rect 327106 233618 327134 239025
rect 327586 233632 327614 241245
rect 328054 241229 328106 241235
rect 328054 241171 328106 241177
rect 327862 240785 327914 240791
rect 327862 240727 327914 240733
rect 327874 240569 327902 240727
rect 327766 240563 327818 240569
rect 327766 240505 327818 240511
rect 327862 240563 327914 240569
rect 327862 240505 327914 240511
rect 327778 240421 327806 240505
rect 327670 240415 327722 240421
rect 327670 240357 327722 240363
rect 327766 240415 327818 240421
rect 327766 240357 327818 240363
rect 327682 239903 327710 240357
rect 327670 239897 327722 239903
rect 327670 239839 327722 239845
rect 328066 233632 328094 241171
rect 328246 240785 328298 240791
rect 328246 240727 328298 240733
rect 328258 233928 328286 240727
rect 328354 239681 328382 246938
rect 328786 246711 328814 246938
rect 329026 246924 329280 246952
rect 328774 246705 328826 246711
rect 328774 246647 328826 246653
rect 328918 241821 328970 241827
rect 328918 241763 328970 241769
rect 328534 241451 328586 241457
rect 328534 241393 328586 241399
rect 328342 239675 328394 239681
rect 328342 239617 328394 239623
rect 327456 233604 327614 233632
rect 327840 233604 328094 233632
rect 328210 233900 328286 233928
rect 328210 233618 328238 233900
rect 328546 233618 328574 241393
rect 328930 239237 328958 241763
rect 329026 240273 329054 246924
rect 329014 240267 329066 240273
rect 329014 240209 329066 240215
rect 329206 240267 329258 240273
rect 329206 240209 329258 240215
rect 329110 239823 329162 239829
rect 329110 239765 329162 239771
rect 329122 239237 329150 239765
rect 328918 239231 328970 239237
rect 328918 239173 328970 239179
rect 329110 239231 329162 239237
rect 329110 239173 329162 239179
rect 329218 233632 329246 240209
rect 329302 239823 329354 239829
rect 329302 239765 329354 239771
rect 328944 233604 329246 233632
rect 329314 233618 329342 239765
rect 329698 235685 329726 246938
rect 329794 246924 330096 246952
rect 329794 240273 329822 246924
rect 330262 242709 330314 242715
rect 330262 242651 330314 242657
rect 329878 241377 329930 241383
rect 329878 241319 329930 241325
rect 329782 240267 329834 240273
rect 329782 240209 329834 240215
rect 329686 235679 329738 235685
rect 329686 235621 329738 235627
rect 329890 233632 329918 241319
rect 330274 233632 330302 242651
rect 330562 241901 330590 246938
rect 331008 246924 331166 246952
rect 330646 242931 330698 242937
rect 330646 242873 330698 242879
rect 330550 241895 330602 241901
rect 330550 241837 330602 241843
rect 330658 233632 330686 242873
rect 331030 242857 331082 242863
rect 331030 242799 331082 242805
rect 330742 242561 330794 242567
rect 330742 242503 330794 242509
rect 329664 233604 329918 233632
rect 330048 233604 330302 233632
rect 330432 233604 330686 233632
rect 330754 233618 330782 242503
rect 330934 239971 330986 239977
rect 330934 239913 330986 239919
rect 330946 239755 330974 239913
rect 330934 239749 330986 239755
rect 330934 239691 330986 239697
rect 331042 233632 331070 242799
rect 331138 239977 331166 246924
rect 331234 246924 331488 246952
rect 331234 241943 331262 246924
rect 331858 246785 331886 246938
rect 331846 246779 331898 246785
rect 331846 246721 331898 246727
rect 331220 241934 331276 241943
rect 331220 241869 331276 241878
rect 331318 241895 331370 241901
rect 331318 241837 331370 241843
rect 331330 240125 331358 241837
rect 332086 241155 332138 241161
rect 332086 241097 332138 241103
rect 331318 240119 331370 240125
rect 331318 240061 331370 240067
rect 331510 240045 331562 240051
rect 331510 239987 331562 239993
rect 331126 239971 331178 239977
rect 331126 239913 331178 239919
rect 331042 233604 331152 233632
rect 331522 233618 331550 239987
rect 332098 233632 332126 241097
rect 332290 240569 332318 246938
rect 332770 246637 332798 246938
rect 332962 246924 333216 246952
rect 333442 246924 333600 246952
rect 333826 246924 334080 246952
rect 332758 246631 332810 246637
rect 332758 246573 332810 246579
rect 332962 241087 332990 246924
rect 332950 241081 333002 241087
rect 332950 241023 333002 241029
rect 332470 241007 332522 241013
rect 332470 240949 332522 240955
rect 332278 240563 332330 240569
rect 332278 240505 332330 240511
rect 332482 233632 332510 240949
rect 332854 240563 332906 240569
rect 332854 240505 332906 240511
rect 332866 233632 332894 240505
rect 333334 240267 333386 240273
rect 333334 240209 333386 240215
rect 332950 239971 333002 239977
rect 332950 239913 333002 239919
rect 331872 233604 332126 233632
rect 332256 233604 332510 233632
rect 332640 233604 332894 233632
rect 332962 233618 332990 239913
rect 333346 233618 333374 240209
rect 333442 235833 333470 246924
rect 333826 241531 333854 246924
rect 334498 246563 334526 246938
rect 334486 246557 334538 246563
rect 334486 246499 334538 246505
rect 334978 241753 335006 246938
rect 335156 244154 335212 244163
rect 335156 244089 335212 244098
rect 334966 241747 335018 241753
rect 334966 241689 335018 241695
rect 334582 241599 334634 241605
rect 334582 241541 334634 241547
rect 333814 241525 333866 241531
rect 333814 241467 333866 241473
rect 333718 241007 333770 241013
rect 333718 240949 333770 240955
rect 333430 235827 333482 235833
rect 333430 235769 333482 235775
rect 333730 233618 333758 240949
rect 334594 240865 334622 241541
rect 335062 240933 335114 240939
rect 335062 240875 335114 240881
rect 334582 240859 334634 240865
rect 334582 240801 334634 240807
rect 334678 240859 334730 240865
rect 334678 240801 334730 240807
rect 334198 240489 334250 240495
rect 334198 240431 334250 240437
rect 334294 240489 334346 240495
rect 334294 240431 334346 240437
rect 334210 239977 334238 240431
rect 334198 239971 334250 239977
rect 334198 239913 334250 239919
rect 334306 233632 334334 240431
rect 334690 233632 334718 240801
rect 335074 233632 335102 240875
rect 334080 233604 334334 233632
rect 334464 233604 334718 233632
rect 334848 233604 335102 233632
rect 335170 233618 335198 244089
rect 335362 235759 335390 246938
rect 335554 246924 335808 246952
rect 336034 246924 336288 246952
rect 335554 241679 335582 246924
rect 335926 244411 335978 244417
rect 335926 244353 335978 244359
rect 335542 241673 335594 241679
rect 335542 241615 335594 241621
rect 335542 238491 335594 238497
rect 335542 238433 335594 238439
rect 335350 235753 335402 235759
rect 335350 235695 335402 235701
rect 335554 233618 335582 238433
rect 335938 233618 335966 244353
rect 336034 240421 336062 246924
rect 336610 246489 336638 246938
rect 336994 246924 337104 246952
rect 336598 246483 336650 246489
rect 336598 246425 336650 246431
rect 336406 244633 336458 244639
rect 336406 244575 336458 244581
rect 336022 240415 336074 240421
rect 336022 240357 336074 240363
rect 336022 238639 336074 238645
rect 336022 238581 336074 238587
rect 336034 233632 336062 238581
rect 336418 233632 336446 244575
rect 336994 239311 337022 246924
rect 337366 244337 337418 244343
rect 337366 244279 337418 244285
rect 337078 241747 337130 241753
rect 337078 241689 337130 241695
rect 337090 240643 337118 241689
rect 337078 240637 337130 240643
rect 337078 240579 337130 240585
rect 336982 239305 337034 239311
rect 336982 239247 337034 239253
rect 336982 238713 337034 238719
rect 336982 238655 337034 238661
rect 336994 233632 337022 238655
rect 336034 233604 336288 233632
rect 336418 233604 336672 233632
rect 336994 233604 337056 233632
rect 337378 233618 337406 244279
rect 337570 235611 337598 246938
rect 337762 246924 338016 246952
rect 338146 246924 338400 246952
rect 337762 239163 337790 246924
rect 338146 246415 338174 246924
rect 338134 246409 338186 246415
rect 338134 246351 338186 246357
rect 338710 244485 338762 244491
rect 338710 244427 338762 244433
rect 337846 242635 337898 242641
rect 337846 242577 337898 242583
rect 337750 239157 337802 239163
rect 337750 239099 337802 239105
rect 337750 238565 337802 238571
rect 337750 238507 337802 238513
rect 337558 235605 337610 235611
rect 337558 235547 337610 235553
rect 337762 233618 337790 238507
rect 337858 233632 337886 242577
rect 338146 242040 338366 242068
rect 338146 241827 338174 242040
rect 338338 241920 338366 242040
rect 338518 241969 338570 241975
rect 338230 241895 338282 241901
rect 338338 241892 338462 241920
rect 338518 241911 338570 241917
rect 338230 241837 338282 241843
rect 338134 241821 338186 241827
rect 338134 241763 338186 241769
rect 338134 241673 338186 241679
rect 338134 241615 338186 241621
rect 338038 241525 338090 241531
rect 338038 241467 338090 241473
rect 338050 241235 338078 241467
rect 338146 241309 338174 241615
rect 338134 241303 338186 241309
rect 338134 241245 338186 241251
rect 338038 241229 338090 241235
rect 338038 241171 338090 241177
rect 338134 240785 338186 240791
rect 338134 240727 338186 240733
rect 338146 240421 338174 240727
rect 338242 240717 338270 241837
rect 338434 241217 338462 241892
rect 338530 241309 338558 241911
rect 338518 241303 338570 241309
rect 338518 241245 338570 241251
rect 338614 241229 338666 241235
rect 338434 241189 338614 241217
rect 338614 241171 338666 241177
rect 338230 240711 338282 240717
rect 338230 240653 338282 240659
rect 338614 240711 338666 240717
rect 338614 240653 338666 240659
rect 338134 240415 338186 240421
rect 338134 240357 338186 240363
rect 338626 240273 338654 240653
rect 338614 240267 338666 240273
rect 338614 240209 338666 240215
rect 338518 240193 338570 240199
rect 338242 240141 338518 240144
rect 338242 240135 338570 240141
rect 338242 240125 338558 240135
rect 338230 240119 338558 240125
rect 338282 240116 338558 240119
rect 338230 240061 338282 240067
rect 338230 238861 338282 238867
rect 338230 238803 338282 238809
rect 338242 233632 338270 238803
rect 338722 233632 338750 244427
rect 338818 239607 338846 246938
rect 338902 241821 338954 241827
rect 338902 241763 338954 241769
rect 338806 239601 338858 239607
rect 338806 239543 338858 239549
rect 338914 239089 338942 241763
rect 338998 241081 339050 241087
rect 338998 241023 339050 241029
rect 339010 240051 339038 241023
rect 338998 240045 339050 240051
rect 338998 239987 339050 239993
rect 338902 239083 338954 239089
rect 338902 239025 338954 239031
rect 338996 238382 339052 238391
rect 338996 238317 339052 238326
rect 339010 233632 339038 238317
rect 339298 235537 339326 246938
rect 339490 246924 339792 246952
rect 339874 246924 340128 246952
rect 340546 246924 340608 246952
rect 339490 242123 339518 246924
rect 339874 246341 339902 246924
rect 339862 246335 339914 246341
rect 339862 246277 339914 246283
rect 339860 245190 339916 245199
rect 339860 245125 339916 245134
rect 339764 245042 339820 245051
rect 339874 245028 339902 245125
rect 339820 245000 339902 245028
rect 339764 244977 339820 244986
rect 339574 242783 339626 242789
rect 339574 242725 339626 242731
rect 339478 242117 339530 242123
rect 339478 242059 339530 242065
rect 339286 235531 339338 235537
rect 339286 235473 339338 235479
rect 337858 233604 338160 233632
rect 338242 233604 338496 233632
rect 338722 233604 338880 233632
rect 339010 233604 339264 233632
rect 339586 233618 339614 242725
rect 340342 242413 340394 242419
rect 340342 242355 340394 242361
rect 339958 238787 340010 238793
rect 339958 238729 340010 238735
rect 339970 233618 339998 238729
rect 340354 233618 340382 242355
rect 340438 238935 340490 238941
rect 340438 238877 340490 238883
rect 340450 233632 340478 238877
rect 340546 235463 340574 246924
rect 340820 243710 340876 243719
rect 340820 243645 340876 243654
rect 340534 235457 340586 235463
rect 340534 235399 340586 235405
rect 340834 233632 340862 243645
rect 341026 239903 341054 246938
rect 341506 246267 341534 246938
rect 341494 246261 341546 246267
rect 341494 246203 341546 246209
rect 341780 244006 341836 244015
rect 341780 243941 341836 243950
rect 341014 239897 341066 239903
rect 341014 239839 341066 239845
rect 341204 238530 341260 238539
rect 341204 238465 341260 238474
rect 341218 233632 341246 238465
rect 340450 233604 340704 233632
rect 340834 233604 341088 233632
rect 341218 233604 341472 233632
rect 341794 233618 341822 243941
rect 341890 239681 341918 246938
rect 342082 246924 342336 246952
rect 342754 246924 342816 246952
rect 341878 239675 341930 239681
rect 341878 239617 341930 239623
rect 342082 235389 342110 246924
rect 342548 244746 342604 244755
rect 342548 244681 342604 244690
rect 342164 238086 342220 238095
rect 342164 238021 342220 238030
rect 342070 235383 342122 235389
rect 342070 235325 342122 235331
rect 342178 233618 342206 238021
rect 342562 233618 342590 244681
rect 342754 240347 342782 246924
rect 343234 246045 343262 246938
rect 343222 246039 343274 246045
rect 343222 245981 343274 245987
rect 343028 243858 343084 243867
rect 343028 243793 343084 243802
rect 342742 240341 342794 240347
rect 342742 240283 342794 240289
rect 342836 240306 342892 240315
rect 342836 240241 342838 240250
rect 342890 240241 342892 240250
rect 342838 240209 342890 240215
rect 342742 240045 342794 240051
rect 342740 240010 342742 240019
rect 342794 240010 342796 240019
rect 342740 239945 342796 239954
rect 342740 238234 342796 238243
rect 342740 238169 342796 238178
rect 342754 233632 342782 238169
rect 343042 233632 343070 243793
rect 343126 240341 343178 240347
rect 343126 240283 343178 240289
rect 343138 239755 343166 240283
rect 343126 239749 343178 239755
rect 343126 239691 343178 239697
rect 343618 239237 343646 246938
rect 343988 244598 344044 244607
rect 343988 244533 344044 244542
rect 343606 239231 343658 239237
rect 343606 239173 343658 239179
rect 343412 238678 343468 238687
rect 343412 238613 343468 238622
rect 343426 233632 343454 238613
rect 342754 233604 342912 233632
rect 343042 233604 343296 233632
rect 343426 233604 343680 233632
rect 344002 233618 344030 244533
rect 344098 235315 344126 246938
rect 344290 246924 344544 246952
rect 344674 246924 344928 246952
rect 344290 241235 344318 246924
rect 344278 241229 344330 241235
rect 344278 241171 344330 241177
rect 344674 240125 344702 246924
rect 344756 244450 344812 244459
rect 344756 244385 344812 244394
rect 344662 240119 344714 240125
rect 344662 240061 344714 240067
rect 344372 237938 344428 237947
rect 344372 237873 344428 237882
rect 344086 235309 344138 235315
rect 344086 235251 344138 235257
rect 344386 233618 344414 237873
rect 344770 233618 344798 244385
rect 345236 243118 345292 243127
rect 345236 243053 345292 243062
rect 344852 238826 344908 238835
rect 344852 238761 344908 238770
rect 344866 233632 344894 238761
rect 345250 233632 345278 243053
rect 345346 235241 345374 246938
rect 345826 241753 345854 246938
rect 346306 245823 346334 246938
rect 346402 246924 346656 246952
rect 346882 246924 347136 246952
rect 346294 245817 346346 245823
rect 346294 245759 346346 245765
rect 346196 244302 346252 244311
rect 346196 244237 346252 244246
rect 345814 241747 345866 241753
rect 345814 241689 345866 241695
rect 345620 238974 345676 238983
rect 345620 238909 345676 238918
rect 345334 235235 345386 235241
rect 345334 235177 345386 235183
rect 345634 233632 345662 238909
rect 344866 233604 345120 233632
rect 345250 233604 345504 233632
rect 345634 233604 345888 233632
rect 346210 233618 346238 244237
rect 346402 241309 346430 246924
rect 346390 241303 346442 241309
rect 346390 241245 346442 241251
rect 346582 237603 346634 237609
rect 346582 237545 346634 237551
rect 346594 233618 346622 237545
rect 346882 235167 346910 246924
rect 347444 243266 347500 243275
rect 347444 243201 347500 243210
rect 346964 242970 347020 242979
rect 346964 242905 347020 242914
rect 346870 235161 346922 235167
rect 346870 235103 346922 235109
rect 346978 233618 347006 242905
rect 347060 237494 347116 237503
rect 347060 237429 347116 237438
rect 347074 233632 347102 237429
rect 347458 233632 347486 243201
rect 347554 239977 347582 246938
rect 348034 245897 348062 246938
rect 348130 246924 348432 246952
rect 348610 246924 348864 246952
rect 349090 246924 349344 246952
rect 348022 245891 348074 245897
rect 348022 245833 348074 245839
rect 348130 241605 348158 246924
rect 348502 244263 348554 244269
rect 348502 244205 348554 244211
rect 348514 243825 348542 244205
rect 348502 243819 348554 243825
rect 348502 243761 348554 243767
rect 348404 243562 348460 243571
rect 348404 243497 348460 243506
rect 348118 241599 348170 241605
rect 348118 241541 348170 241547
rect 348214 241599 348266 241605
rect 348214 241541 348266 241547
rect 347542 239971 347594 239977
rect 347542 239913 347594 239919
rect 348226 239829 348254 241541
rect 348214 239823 348266 239829
rect 348214 239765 348266 239771
rect 347830 237899 347882 237905
rect 347830 237841 347882 237847
rect 347842 233632 347870 237841
rect 347074 233604 347328 233632
rect 347458 233604 347712 233632
rect 347842 233604 348096 233632
rect 348418 233618 348446 243497
rect 348502 243227 348554 243233
rect 348502 243169 348554 243175
rect 348514 242789 348542 243169
rect 348502 242783 348554 242789
rect 348502 242725 348554 242731
rect 348610 235019 348638 246924
rect 349090 245749 349118 246924
rect 349078 245743 349130 245749
rect 349078 245685 349130 245691
rect 349654 243523 349706 243529
rect 349654 243465 349706 243471
rect 349174 243449 349226 243455
rect 349174 243391 349226 243397
rect 348788 237346 348844 237355
rect 348788 237281 348844 237290
rect 348598 235013 348650 235019
rect 348598 234955 348650 234961
rect 348802 233618 348830 237281
rect 349186 233618 349214 243391
rect 349270 237677 349322 237683
rect 349270 237619 349322 237625
rect 349282 233632 349310 237619
rect 349666 233632 349694 243465
rect 349762 239385 349790 246938
rect 349750 239379 349802 239385
rect 349750 239321 349802 239327
rect 350038 237825 350090 237831
rect 350038 237767 350090 237773
rect 350050 233632 350078 237767
rect 350146 234871 350174 246938
rect 350422 243597 350474 243603
rect 350422 243539 350474 243545
rect 350134 234865 350186 234871
rect 350134 234807 350186 234813
rect 350434 233632 350462 243539
rect 350626 240019 350654 246938
rect 350818 246924 351072 246952
rect 351394 246924 351552 246952
rect 351682 246924 351888 246952
rect 350818 245675 350846 246924
rect 350806 245669 350858 245675
rect 350806 245611 350858 245617
rect 351394 240315 351422 246924
rect 351478 243375 351530 243381
rect 351478 243317 351530 243323
rect 351380 240306 351436 240315
rect 351380 240241 351436 240250
rect 350612 240010 350668 240019
rect 350612 239945 350668 239954
rect 351490 238220 351518 243317
rect 351394 238192 351518 238220
rect 350998 237973 351050 237979
rect 350998 237915 351050 237921
rect 349282 233604 349536 233632
rect 349666 233604 349920 233632
rect 350050 233604 350304 233632
rect 350434 233604 350640 233632
rect 351010 233618 351038 237915
rect 351394 233618 351422 238192
rect 351478 237751 351530 237757
rect 351478 237693 351530 237699
rect 351490 233632 351518 237693
rect 351682 234723 351710 246924
rect 351862 243745 351914 243751
rect 351862 243687 351914 243693
rect 351670 234717 351722 234723
rect 351670 234659 351722 234665
rect 351874 233632 351902 243687
rect 352354 239311 352382 246938
rect 352834 245527 352862 246938
rect 352930 246924 353184 246952
rect 353410 246924 353664 246952
rect 352822 245521 352874 245527
rect 352822 245463 352874 245469
rect 352822 244263 352874 244269
rect 352822 244205 352874 244211
rect 352342 239305 352394 239311
rect 352342 239247 352394 239253
rect 352244 237790 352300 237799
rect 352244 237725 352300 237734
rect 352258 233632 352286 237725
rect 351490 233604 351744 233632
rect 351874 233604 352128 233632
rect 352258 233604 352512 233632
rect 352834 233618 352862 244205
rect 352930 241901 352958 246924
rect 352918 241895 352970 241901
rect 352918 241837 352970 241843
rect 353410 241827 353438 246924
rect 354082 245601 354110 246938
rect 354070 245595 354122 245601
rect 354070 245537 354122 245543
rect 353590 243967 353642 243973
rect 353590 243909 353642 243915
rect 353398 241821 353450 241827
rect 353398 241763 353450 241769
rect 353206 238121 353258 238127
rect 353206 238063 353258 238069
rect 353218 233618 353246 238063
rect 353602 233618 353630 243909
rect 354358 243671 354410 243677
rect 354358 243613 354410 243619
rect 353686 238047 353738 238053
rect 353686 237989 353738 237995
rect 353698 233632 353726 237989
rect 354370 233928 354398 243613
rect 354562 241753 354590 246938
rect 354550 241747 354602 241753
rect 354550 241689 354602 241695
rect 354452 237642 354508 237651
rect 354452 237577 354508 237586
rect 354322 233900 354398 233928
rect 353698 233604 353952 233632
rect 354322 233618 354350 233900
rect 354466 233632 354494 237577
rect 354946 234575 354974 246938
rect 355138 246924 355392 246952
rect 355618 246924 355872 246952
rect 355030 244115 355082 244121
rect 355030 244057 355082 244063
rect 354934 234569 354986 234575
rect 354934 234511 354986 234517
rect 354466 233604 354720 233632
rect 355042 233618 355070 244057
rect 355138 241531 355166 246924
rect 355618 245379 355646 246924
rect 355606 245373 355658 245379
rect 355606 245315 355658 245321
rect 355798 243893 355850 243899
rect 355798 243835 355850 243841
rect 355126 241525 355178 241531
rect 355126 241467 355178 241473
rect 355414 238195 355466 238201
rect 355414 238137 355466 238143
rect 355426 233618 355454 238137
rect 355810 233618 355838 243835
rect 356290 240421 356318 246938
rect 356482 246924 356688 246952
rect 356374 244189 356426 244195
rect 356374 244131 356426 244137
rect 356278 240415 356330 240421
rect 356278 240357 356330 240363
rect 355894 238269 355946 238275
rect 355894 238211 355946 238217
rect 355906 233632 355934 238211
rect 356386 233632 356414 244131
rect 356482 234427 356510 246924
rect 357154 241457 357182 246938
rect 357346 246924 357600 246952
rect 357826 246924 358080 246952
rect 357346 245231 357374 246924
rect 357334 245225 357386 245231
rect 357334 245167 357386 245173
rect 357238 244041 357290 244047
rect 357238 243983 357290 243989
rect 357142 241451 357194 241457
rect 357142 241393 357194 241399
rect 356662 238417 356714 238423
rect 356662 238359 356714 238365
rect 356470 234421 356522 234427
rect 356470 234363 356522 234369
rect 356674 233632 356702 238359
rect 355906 233604 356160 233632
rect 356386 233604 356544 233632
rect 356674 233604 356928 233632
rect 357250 233618 357278 243983
rect 357622 238343 357674 238349
rect 357622 238285 357674 238291
rect 357634 233618 357662 238285
rect 357826 234353 357854 246924
rect 358402 241605 358430 246938
rect 358882 245157 358910 246938
rect 358870 245151 358922 245157
rect 358870 245093 358922 245099
rect 358390 241599 358442 241605
rect 358390 241541 358442 241547
rect 359362 241383 359390 246938
rect 359554 246924 359808 246952
rect 360034 246924 360192 246952
rect 359350 241377 359402 241383
rect 359350 241319 359402 241325
rect 358868 239566 358924 239575
rect 358868 239501 358924 239510
rect 358006 235087 358058 235093
rect 358006 235029 358058 235035
rect 357814 234347 357866 234353
rect 357814 234289 357866 234295
rect 358018 233618 358046 235029
rect 358102 234939 358154 234945
rect 358102 234881 358154 234887
rect 358114 233632 358142 234881
rect 358486 233681 358538 233687
rect 358114 233604 358368 233632
rect 358882 233632 358910 239501
rect 359444 239418 359500 239427
rect 359444 239353 359500 239362
rect 358538 233629 358752 233632
rect 358486 233623 358752 233629
rect 358498 233604 358752 233623
rect 358882 233604 359136 233632
rect 359458 233618 359486 239353
rect 359554 234279 359582 246924
rect 360034 242715 360062 246924
rect 360610 245971 360638 246938
rect 360598 245965 360650 245971
rect 360598 245907 360650 245913
rect 360790 243819 360842 243825
rect 360790 243761 360842 243767
rect 360214 243745 360266 243751
rect 360214 243687 360266 243693
rect 360022 242709 360074 242715
rect 360022 242651 360074 242657
rect 359830 241081 359882 241087
rect 359830 241023 359882 241029
rect 359542 234273 359594 234279
rect 359542 234215 359594 234221
rect 359842 233618 359870 241023
rect 360226 233618 360254 243687
rect 360802 233632 360830 243761
rect 361090 242937 361118 246938
rect 361078 242931 361130 242937
rect 361078 242873 361130 242879
rect 361174 237899 361226 237905
rect 361174 237841 361226 237847
rect 361186 233632 361214 237841
rect 361474 236129 361502 246938
rect 361666 246924 361920 246952
rect 362146 246924 362400 246952
rect 361666 242567 361694 246924
rect 362038 243671 362090 243677
rect 362038 243613 362090 243619
rect 361942 243449 361994 243455
rect 361942 243391 361994 243397
rect 361654 242561 361706 242567
rect 361654 242503 361706 242509
rect 361558 237825 361610 237831
rect 361558 237767 361610 237773
rect 361462 236123 361514 236129
rect 361462 236065 361514 236071
rect 361570 233632 361598 237767
rect 361954 233632 361982 243391
rect 360576 233604 360830 233632
rect 360960 233604 361214 233632
rect 361344 233604 361598 233632
rect 361680 233604 361982 233632
rect 362050 233618 362078 243613
rect 362146 242863 362174 246924
rect 362818 246119 362846 246938
rect 362806 246113 362858 246119
rect 362806 246055 362858 246061
rect 362422 243597 362474 243603
rect 362422 243539 362474 243545
rect 362134 242857 362186 242863
rect 362134 242799 362186 242805
rect 362434 233618 362462 243539
rect 362806 241377 362858 241383
rect 362806 241319 362858 241325
rect 362818 233632 362846 241319
rect 363202 241235 363230 246938
rect 363190 241229 363242 241235
rect 363190 241171 363242 241177
rect 363382 237677 363434 237683
rect 363382 237619 363434 237625
rect 363394 233632 363422 237619
rect 363682 233909 363710 246938
rect 363970 246924 364128 246952
rect 364354 246924 364608 246952
rect 364738 246924 364992 246952
rect 363862 243523 363914 243529
rect 363862 243465 363914 243471
rect 363766 237751 363818 237757
rect 363766 237693 363818 237699
rect 363670 233903 363722 233909
rect 363670 233845 363722 233851
rect 363778 233632 363806 237693
rect 362784 233604 362846 233632
rect 363168 233604 363422 233632
rect 363552 233604 363806 233632
rect 363874 233618 363902 243465
rect 363970 241013 363998 246924
rect 364354 246193 364382 246924
rect 364342 246187 364394 246193
rect 364342 246129 364394 246135
rect 364630 243375 364682 243381
rect 364630 243317 364682 243323
rect 363958 241007 364010 241013
rect 363958 240949 364010 240955
rect 364246 237603 364298 237609
rect 364246 237545 364298 237551
rect 364258 233618 364286 237545
rect 364642 233618 364670 243317
rect 364738 240939 364766 246924
rect 365410 241647 365438 246938
rect 365684 241934 365740 241943
rect 365684 241869 365740 241878
rect 365588 241786 365644 241795
rect 365588 241721 365644 241730
rect 365396 241638 365452 241647
rect 365396 241573 365452 241582
rect 364726 240933 364778 240939
rect 364726 240875 364778 240881
rect 365204 240306 365260 240315
rect 365204 240241 365260 240250
rect 365218 233632 365246 240241
rect 365602 233632 365630 241721
rect 364992 233604 365246 233632
rect 365376 233604 365630 233632
rect 365698 233632 365726 241869
rect 365780 241638 365836 241647
rect 365780 241573 365836 241582
rect 365794 241203 365822 241573
rect 365780 241194 365836 241203
rect 365780 241129 365836 241138
rect 365890 240569 365918 246938
rect 366082 246924 366336 246952
rect 366466 246924 366720 246952
rect 366946 246924 367200 246952
rect 366082 241499 366110 246924
rect 366466 241499 366494 246924
rect 366068 241490 366124 241499
rect 366068 241425 366124 241434
rect 366452 241490 366508 241499
rect 366452 241425 366508 241434
rect 366452 241342 366508 241351
rect 366452 241277 366508 241286
rect 366068 241194 366124 241203
rect 366068 241129 366124 241138
rect 365878 240563 365930 240569
rect 365878 240505 365930 240511
rect 365698 233604 365760 233632
rect 366082 233618 366110 241129
rect 366466 233618 366494 241277
rect 366946 240717 366974 246924
rect 367618 241647 367646 246938
rect 367604 241638 367660 241647
rect 367604 241573 367660 241582
rect 367796 241638 367852 241647
rect 367796 241573 367852 241582
rect 367412 241046 367468 241055
rect 367412 240981 367468 240990
rect 366934 240711 366986 240717
rect 366934 240653 366986 240659
rect 366838 240193 366890 240199
rect 366838 240135 366890 240141
rect 366850 233618 366878 240135
rect 367426 233632 367454 240981
rect 367810 233632 367838 241573
rect 368002 240865 368030 246938
rect 368278 241895 368330 241901
rect 368278 241837 368330 241843
rect 367990 240859 368042 240865
rect 367990 240801 368042 240807
rect 368182 240119 368234 240125
rect 368182 240061 368234 240067
rect 368194 233632 368222 240061
rect 367200 233604 367454 233632
rect 367584 233604 367838 233632
rect 367968 233604 368222 233632
rect 368290 233618 368318 241837
rect 368482 240167 368510 246938
rect 368770 246924 368928 246952
rect 369154 246924 369408 246952
rect 368566 243227 368618 243233
rect 368566 243169 368618 243175
rect 368578 242789 368606 243169
rect 368566 242783 368618 242789
rect 368566 242725 368618 242731
rect 368770 240495 368798 246924
rect 369154 240907 369182 246924
rect 369140 240898 369196 240907
rect 369140 240833 369196 240842
rect 369730 240643 369758 246938
rect 370210 240759 370238 246938
rect 370486 241525 370538 241531
rect 370486 241467 370538 241473
rect 370196 240750 370252 240759
rect 370196 240685 370252 240694
rect 369718 240637 369770 240643
rect 369718 240579 369770 240585
rect 368758 240489 368810 240495
rect 368758 240431 368810 240437
rect 370006 240415 370058 240421
rect 370006 240357 370058 240363
rect 368468 240158 368524 240167
rect 368468 240093 368524 240102
rect 369622 239527 369674 239533
rect 369622 239469 369674 239475
rect 368662 239453 368714 239459
rect 368662 239395 368714 239401
rect 368674 233618 368702 239395
rect 369046 239379 369098 239385
rect 369046 239321 369098 239327
rect 369058 233618 369086 239321
rect 369634 233632 369662 239469
rect 370018 233632 370046 240357
rect 370390 239305 370442 239311
rect 370390 239247 370442 239253
rect 370402 233632 370430 239247
rect 369408 233604 369662 233632
rect 369792 233604 370046 233632
rect 370176 233604 370430 233632
rect 370498 233618 370526 241467
rect 370690 240791 370718 246938
rect 370978 246924 371136 246952
rect 371362 246924 371520 246952
rect 370678 240785 370730 240791
rect 370678 240727 370730 240733
rect 370870 239675 370922 239681
rect 370870 239617 370922 239623
rect 370882 233618 370910 239617
rect 370978 234649 371006 246924
rect 371254 239823 371306 239829
rect 371254 239765 371306 239771
rect 370966 234643 371018 234649
rect 370966 234585 371018 234591
rect 371266 233618 371294 239765
rect 371362 236943 371390 246924
rect 371830 239231 371882 239237
rect 371830 239173 371882 239179
rect 371350 236937 371402 236943
rect 371350 236879 371402 236885
rect 371842 233632 371870 239173
rect 371938 234501 371966 246938
rect 372214 241377 372266 241383
rect 372214 241319 372266 241325
rect 371926 234495 371978 234501
rect 371926 234437 371978 234443
rect 372226 233632 372254 241319
rect 372418 237017 372446 246938
rect 372898 245453 372926 246938
rect 372994 246924 373248 246952
rect 373474 246924 373728 246952
rect 372886 245447 372938 245453
rect 372886 245389 372938 245395
rect 372994 243011 373022 246924
rect 373474 245305 373502 246924
rect 373462 245299 373514 245305
rect 373462 245241 373514 245247
rect 372982 243005 373034 243011
rect 372982 242947 373034 242953
rect 372694 241821 372746 241827
rect 372694 241763 372746 241769
rect 372598 240711 372650 240717
rect 372598 240653 372650 240659
rect 372406 237011 372458 237017
rect 372406 236953 372458 236959
rect 372610 233632 372638 240653
rect 371616 233604 371870 233632
rect 372000 233604 372254 233632
rect 372384 233604 372638 233632
rect 372706 233618 372734 241763
rect 373078 241673 373130 241679
rect 373078 241615 373130 241621
rect 373090 233618 373118 241615
rect 373462 241229 373514 241235
rect 373462 241171 373514 241177
rect 373474 233618 373502 241171
rect 374038 240933 374090 240939
rect 374038 240875 374090 240881
rect 374050 233632 374078 240875
rect 374146 237165 374174 246938
rect 374326 240563 374378 240569
rect 374326 240505 374378 240511
rect 374134 237159 374186 237165
rect 374134 237101 374186 237107
rect 374338 233632 374366 240505
rect 374626 234205 374654 246938
rect 375010 243159 375038 246938
rect 375202 246924 375456 246952
rect 375778 246924 375936 246952
rect 376066 246924 376272 246952
rect 374998 243153 375050 243159
rect 374998 243095 375050 243101
rect 374902 241155 374954 241161
rect 374902 241097 374954 241103
rect 374806 239749 374858 239755
rect 374806 239691 374858 239697
rect 374614 234199 374666 234205
rect 374614 234141 374666 234147
rect 374818 233632 374846 239691
rect 373824 233604 374078 233632
rect 374208 233604 374366 233632
rect 374592 233604 374846 233632
rect 374914 233618 374942 241097
rect 375202 237313 375230 246924
rect 375670 241007 375722 241013
rect 375670 240949 375722 240955
rect 375286 240785 375338 240791
rect 375286 240727 375338 240733
rect 375190 237307 375242 237313
rect 375190 237249 375242 237255
rect 375298 233618 375326 240727
rect 375682 233618 375710 240949
rect 375778 234131 375806 246924
rect 376066 237091 376094 246924
rect 376738 245083 376766 246938
rect 376726 245077 376778 245083
rect 376726 245019 376778 245025
rect 377218 243085 377246 246938
rect 377410 246924 377664 246952
rect 377794 246924 378048 246952
rect 377206 243079 377258 243085
rect 377206 243021 377258 243027
rect 377108 240750 377164 240759
rect 377108 240685 377164 240694
rect 376630 240637 376682 240643
rect 376630 240579 376682 240585
rect 376246 240489 376298 240495
rect 376246 240431 376298 240437
rect 376054 237085 376106 237091
rect 376054 237027 376106 237033
rect 375766 234125 375818 234131
rect 375766 234067 375818 234073
rect 376258 233632 376286 240431
rect 376642 233632 376670 240579
rect 377012 239862 377068 239871
rect 377012 239797 377068 239806
rect 377026 233632 377054 239797
rect 376032 233604 376286 233632
rect 376416 233604 376670 233632
rect 376800 233604 377054 233632
rect 377122 233618 377150 240685
rect 377410 233983 377438 246924
rect 377492 240010 377548 240019
rect 377492 239945 377548 239954
rect 377398 233977 377450 233983
rect 377398 233919 377450 233925
rect 377506 233618 377534 239945
rect 377794 237387 377822 246924
rect 378466 245009 378494 246938
rect 378454 245003 378506 245009
rect 378454 244945 378506 244951
rect 378946 243233 378974 246938
rect 378934 243227 378986 243233
rect 378934 243169 378986 243175
rect 378550 241895 378602 241901
rect 378550 241837 378602 241843
rect 377878 241747 377930 241753
rect 377878 241689 377930 241695
rect 377890 240199 377918 241689
rect 377878 240193 377930 240199
rect 377878 240135 377930 240141
rect 378452 240158 378508 240167
rect 378562 240125 378590 241837
rect 379220 241490 379276 241499
rect 379220 241425 379276 241434
rect 378452 240093 378508 240102
rect 378550 240119 378602 240125
rect 377876 239714 377932 239723
rect 377876 239649 377932 239658
rect 377782 237381 377834 237387
rect 377782 237323 377834 237329
rect 377890 233618 377918 239649
rect 378466 233632 378494 240093
rect 378550 240061 378602 240067
rect 378838 240119 378890 240125
rect 378838 240061 378890 240067
rect 378850 233632 378878 240061
rect 379234 233632 379262 241425
rect 379316 240898 379372 240907
rect 379316 240833 379372 240842
rect 378240 233604 378494 233632
rect 378624 233604 378878 233632
rect 379008 233604 379262 233632
rect 379330 233618 379358 240833
rect 379426 234057 379454 246938
rect 379522 246924 379776 246952
rect 380194 246924 380256 246952
rect 379522 244935 379550 246924
rect 379510 244929 379562 244935
rect 379510 244871 379562 244877
rect 380086 240193 380138 240199
rect 380086 240135 380138 240141
rect 379702 239083 379754 239089
rect 379702 239025 379754 239031
rect 379414 234051 379466 234057
rect 379414 233993 379466 233999
rect 379714 233618 379742 239025
rect 380098 233618 380126 240135
rect 380194 237535 380222 246924
rect 380674 244861 380702 246938
rect 380662 244855 380714 244861
rect 380662 244797 380714 244803
rect 381154 243307 381182 246938
rect 381250 246924 381552 246952
rect 381730 246924 381984 246952
rect 382402 246924 382464 246952
rect 382594 246924 382896 246952
rect 381142 243301 381194 243307
rect 381142 243243 381194 243249
rect 380662 239601 380714 239607
rect 380662 239543 380714 239549
rect 380182 237529 380234 237535
rect 380182 237471 380234 237477
rect 380674 233632 380702 239543
rect 381046 239157 381098 239163
rect 381046 239099 381098 239105
rect 381058 233632 381086 239099
rect 381250 233835 381278 246924
rect 381430 241303 381482 241309
rect 381430 241245 381482 241251
rect 381238 233829 381290 233835
rect 381238 233771 381290 233777
rect 381442 233632 381470 241245
rect 381526 240341 381578 240347
rect 381526 240283 381578 240289
rect 380448 233604 380702 233632
rect 380832 233604 381086 233632
rect 381216 233604 381470 233632
rect 381538 233618 381566 240283
rect 381730 237461 381758 246924
rect 381910 240267 381962 240273
rect 381910 240209 381962 240215
rect 381718 237455 381770 237461
rect 381718 237397 381770 237403
rect 381922 233618 381950 240209
rect 382294 239971 382346 239977
rect 382294 239913 382346 239919
rect 382306 233618 382334 239913
rect 382402 233761 382430 246924
rect 382594 237239 382622 246924
rect 382870 240045 382922 240051
rect 382870 239987 382922 239993
rect 382582 237233 382634 237239
rect 382582 237175 382634 237181
rect 382390 233755 382442 233761
rect 382390 233697 382442 233703
rect 382882 233632 382910 239987
rect 382966 239897 383018 239903
rect 382966 239839 383018 239845
rect 382978 233928 383006 239839
rect 383062 239675 383114 239681
rect 383062 239617 383114 239623
rect 383074 239575 383102 239617
rect 383060 239566 383116 239575
rect 383060 239501 383116 239510
rect 383266 234797 383294 246938
rect 383542 241969 383594 241975
rect 383542 241911 383594 241917
rect 383554 241383 383582 241911
rect 383542 241377 383594 241383
rect 383542 241319 383594 241325
rect 383638 241377 383690 241383
rect 383638 241319 383690 241325
rect 383254 234791 383306 234797
rect 383254 234733 383306 234739
rect 382978 233900 383054 233928
rect 382656 233604 382910 233632
rect 383026 233618 383054 233900
rect 383650 233632 383678 241319
rect 383424 233604 383678 233632
rect 383746 233618 383774 246938
rect 384034 246924 384192 246952
rect 384514 246924 384576 246952
rect 384034 238941 384062 246924
rect 384514 241087 384542 246924
rect 384790 241673 384842 241679
rect 384790 241615 384842 241621
rect 384886 241673 384938 241679
rect 384886 241615 384938 241621
rect 384802 241235 384830 241615
rect 384694 241229 384746 241235
rect 384694 241171 384746 241177
rect 384790 241229 384842 241235
rect 384790 241171 384842 241177
rect 384502 241081 384554 241087
rect 384502 241023 384554 241029
rect 384706 241013 384734 241171
rect 384898 241032 384926 241615
rect 384994 241531 385022 246938
rect 385076 243414 385132 243423
rect 385076 243349 385132 243358
rect 384982 241525 385034 241531
rect 384982 241467 385034 241473
rect 384694 241007 384746 241013
rect 384694 240949 384746 240955
rect 384802 241004 384926 241032
rect 384802 240884 384830 241004
rect 384118 240859 384170 240865
rect 384118 240801 384170 240807
rect 384226 240856 384830 240884
rect 384022 238935 384074 238941
rect 384022 238877 384074 238883
rect 384130 233618 384158 240801
rect 384226 240717 384254 240856
rect 384214 240711 384266 240717
rect 384214 240653 384266 240659
rect 384310 240711 384362 240717
rect 384310 240653 384362 240659
rect 384322 233632 384350 240653
rect 384598 238935 384650 238941
rect 384598 238877 384650 238883
rect 384610 233632 384638 238877
rect 385090 233632 385118 243349
rect 385474 239977 385502 246938
rect 385654 241895 385706 241901
rect 385654 241837 385706 241843
rect 385666 241531 385694 241837
rect 385654 241525 385706 241531
rect 385654 241467 385706 241473
rect 385954 241457 385982 246938
rect 386050 246924 386304 246952
rect 386530 246924 386784 246952
rect 385942 241451 385994 241457
rect 385942 241393 385994 241399
rect 385462 239971 385514 239977
rect 385462 239913 385514 239919
rect 386050 239755 386078 246924
rect 386134 241821 386186 241827
rect 386134 241763 386186 241769
rect 386146 241457 386174 241763
rect 386134 241451 386186 241457
rect 386134 241393 386186 241399
rect 386530 240051 386558 246924
rect 387202 241753 387230 246938
rect 387286 241895 387338 241901
rect 387286 241837 387338 241843
rect 387298 241753 387326 241837
rect 387190 241747 387242 241753
rect 387190 241689 387242 241695
rect 387286 241747 387338 241753
rect 387286 241689 387338 241695
rect 386614 240415 386666 240421
rect 386614 240357 386666 240363
rect 386626 240051 386654 240357
rect 387682 240125 387710 246938
rect 387670 240119 387722 240125
rect 387670 240061 387722 240067
rect 386518 240045 386570 240051
rect 386518 239987 386570 239993
rect 386614 240045 386666 240051
rect 386614 239987 386666 239993
rect 388066 239903 388094 246938
rect 388258 246924 388512 246952
rect 388834 246924 388992 246952
rect 388258 241531 388286 246924
rect 388246 241525 388298 241531
rect 388246 241467 388298 241473
rect 388726 240119 388778 240125
rect 388726 240061 388778 240067
rect 388054 239897 388106 239903
rect 388054 239839 388106 239845
rect 388738 239829 388766 240061
rect 388726 239823 388778 239829
rect 388726 239765 388778 239771
rect 386038 239749 386090 239755
rect 386038 239691 386090 239697
rect 388834 239089 388862 246924
rect 389410 241383 389438 246938
rect 389794 241605 389822 246938
rect 389782 241599 389834 241605
rect 389782 241541 389834 241547
rect 389398 241377 389450 241383
rect 389398 241319 389450 241325
rect 390274 240199 390302 246938
rect 390466 246924 390720 246952
rect 390946 246924 391200 246952
rect 390262 240193 390314 240199
rect 390262 240135 390314 240141
rect 390466 239459 390494 246924
rect 390946 239607 390974 246924
rect 390934 239601 390986 239607
rect 390934 239543 390986 239549
rect 390454 239453 390506 239459
rect 390454 239395 390506 239401
rect 391522 239385 391550 246938
rect 391510 239379 391562 239385
rect 391510 239321 391562 239327
rect 392002 239163 392030 246938
rect 392482 239533 392510 246938
rect 392578 246924 392832 246952
rect 393058 246924 393312 246952
rect 392578 241309 392606 246924
rect 392566 241303 392618 241309
rect 392566 241245 392618 241251
rect 393058 240051 393086 246924
rect 393730 240347 393758 246938
rect 393718 240341 393770 240347
rect 393718 240283 393770 240289
rect 393046 240045 393098 240051
rect 393046 239987 393098 239993
rect 392470 239527 392522 239533
rect 392470 239469 392522 239475
rect 394210 239311 394238 246938
rect 394594 240273 394622 246938
rect 394786 246924 395040 246952
rect 395266 246924 395520 246952
rect 394786 240611 394814 246924
rect 394772 240602 394828 240611
rect 394772 240537 394828 240546
rect 394582 240267 394634 240273
rect 394582 240209 394634 240215
rect 395266 239575 395294 246924
rect 395938 243751 395966 246938
rect 395926 243745 395978 243751
rect 395926 243687 395978 243693
rect 396322 240125 396350 246938
rect 396310 240119 396362 240125
rect 396310 240061 396362 240067
rect 395252 239566 395308 239575
rect 395252 239501 395308 239510
rect 394198 239305 394250 239311
rect 394198 239247 394250 239253
rect 391990 239157 392042 239163
rect 391990 239099 392042 239105
rect 388822 239083 388874 239089
rect 388822 239025 388874 239031
rect 396802 239015 396830 246938
rect 396994 246924 397248 246952
rect 397474 246924 397728 246952
rect 397858 246924 398112 246952
rect 396994 239237 397022 246924
rect 397474 243825 397502 246924
rect 397462 243819 397514 243825
rect 397462 243761 397514 243767
rect 397858 241753 397886 246924
rect 398530 244491 398558 246938
rect 398518 244485 398570 244491
rect 398518 244427 398570 244433
rect 397846 241747 397898 241753
rect 397846 241689 397898 241695
rect 399010 241679 399038 246938
rect 399202 246924 399456 246952
rect 399586 246924 399840 246952
rect 398998 241673 399050 241679
rect 398998 241615 399050 241621
rect 396982 239231 397034 239237
rect 396982 239173 397034 239179
rect 396790 239009 396842 239015
rect 396790 238951 396842 238957
rect 399202 237905 399230 246924
rect 399586 241457 399614 246924
rect 400306 246656 400334 246938
rect 400258 246628 400334 246656
rect 399574 241451 399626 241457
rect 399574 241393 399626 241399
rect 399190 237899 399242 237905
rect 399190 237841 399242 237847
rect 400258 237831 400286 246628
rect 400738 241235 400766 246938
rect 401122 243455 401150 246938
rect 401110 243449 401162 243455
rect 401110 243391 401162 243397
rect 400726 241229 400778 241235
rect 400726 241171 400778 241177
rect 401602 241013 401630 246938
rect 401794 246924 402048 246952
rect 402274 246924 402528 246952
rect 401794 243677 401822 246924
rect 401782 243671 401834 243677
rect 401782 243613 401834 243619
rect 401590 241007 401642 241013
rect 401590 240949 401642 240955
rect 402274 240939 402302 246924
rect 402850 243603 402878 246938
rect 403028 245042 403084 245051
rect 403220 245042 403276 245051
rect 403084 245000 403220 245028
rect 403028 244977 403084 244986
rect 403220 244977 403276 244986
rect 402838 243597 402890 243603
rect 402838 243539 402890 243545
rect 402262 240933 402314 240939
rect 402262 240875 402314 240881
rect 403330 240569 403358 246938
rect 403318 240563 403370 240569
rect 403318 240505 403370 240511
rect 400246 237825 400298 237831
rect 400246 237767 400298 237773
rect 403810 237683 403838 246938
rect 404002 246924 404256 246952
rect 404386 246924 404640 246952
rect 404002 241161 404030 246924
rect 403990 241155 404042 241161
rect 403990 241097 404042 241103
rect 404386 237757 404414 246924
rect 405058 240791 405086 246938
rect 405538 243529 405566 246938
rect 405526 243523 405578 243529
rect 405526 243465 405578 243471
rect 406018 241087 406046 246938
rect 406114 246924 406368 246952
rect 406594 246924 406848 246952
rect 406006 241081 406058 241087
rect 406006 241023 406058 241029
rect 405046 240785 405098 240791
rect 405046 240727 405098 240733
rect 404374 237751 404426 237757
rect 404374 237693 404426 237699
rect 403798 237677 403850 237683
rect 403798 237619 403850 237625
rect 406114 237609 406142 246924
rect 406594 240495 406622 246924
rect 407266 243381 407294 246938
rect 407254 243375 407306 243381
rect 407254 243317 407306 243323
rect 407746 240643 407774 246938
rect 407734 240637 407786 240643
rect 407734 240579 407786 240585
rect 406582 240489 406634 240495
rect 406582 240431 406634 240437
rect 408130 240315 408158 246938
rect 408322 246924 408576 246952
rect 408994 246924 409056 246952
rect 408116 240306 408172 240315
rect 408116 240241 408172 240250
rect 408322 239871 408350 246924
rect 408994 241795 409022 246924
rect 408980 241786 409036 241795
rect 408980 241721 409036 241730
rect 409378 240759 409406 246938
rect 409858 241943 409886 246938
rect 409844 241934 409900 241943
rect 409844 241869 409900 241878
rect 409364 240750 409420 240759
rect 409364 240685 409420 240694
rect 410338 240019 410366 246938
rect 410530 246924 410784 246952
rect 410914 246924 411168 246952
rect 410530 241203 410558 246924
rect 410516 241194 410572 241203
rect 410516 241129 410572 241138
rect 410324 240010 410380 240019
rect 410324 239945 410380 239954
rect 408308 239862 408364 239871
rect 408308 239797 408364 239806
rect 410914 239723 410942 246924
rect 411586 241351 411614 246938
rect 411572 241342 411628 241351
rect 411572 241277 411628 241286
rect 412066 240167 412094 246938
rect 412546 241055 412574 246938
rect 412642 246924 412896 246952
rect 413122 246924 413376 246952
rect 412642 241499 412670 246924
rect 413122 241647 413150 246924
rect 413108 241638 413164 241647
rect 413108 241573 413164 241582
rect 412628 241490 412684 241499
rect 412628 241425 412684 241434
rect 412532 241046 412588 241055
rect 412532 240981 412588 240990
rect 413794 240907 413822 246938
rect 413780 240898 413836 240907
rect 414274 240865 414302 246938
rect 413780 240833 413836 240842
rect 414262 240859 414314 240865
rect 414262 240801 414314 240807
rect 414658 240717 414686 246938
rect 414850 246924 415104 246952
rect 415330 246924 415584 246952
rect 414646 240711 414698 240717
rect 414646 240653 414698 240659
rect 412052 240158 412108 240167
rect 412052 240093 412108 240102
rect 410900 239714 410956 239723
rect 410900 239649 410956 239658
rect 406102 237603 406154 237609
rect 406102 237545 406154 237551
rect 384322 233604 384528 233632
rect 384610 233604 384864 233632
rect 385090 233604 385248 233632
rect 414850 233613 414878 246924
rect 415330 240463 415358 246924
rect 420502 245003 420554 245009
rect 420502 244945 420554 244951
rect 420514 244903 420542 244945
rect 420500 244894 420556 244903
rect 420500 244829 420556 244838
rect 421858 242239 421886 275581
rect 422626 270169 422654 275650
rect 422614 270163 422666 270169
rect 422614 270105 422666 270111
rect 423874 261659 423902 275650
rect 423862 261653 423914 261659
rect 423862 261595 423914 261601
rect 425026 260475 425054 275650
rect 426274 271871 426302 275650
rect 427426 272981 427454 275650
rect 427414 272975 427466 272981
rect 427414 272917 427466 272923
rect 428674 272093 428702 275650
rect 429826 273869 429854 275650
rect 429814 273863 429866 273869
rect 429814 273805 429866 273811
rect 428662 272087 428714 272093
rect 428662 272029 428714 272035
rect 426262 271865 426314 271871
rect 426262 271807 426314 271813
rect 431074 261585 431102 275650
rect 432226 273795 432254 275650
rect 432214 273789 432266 273795
rect 432214 273731 432266 273737
rect 433378 273721 433406 275650
rect 433366 273715 433418 273721
rect 433366 273657 433418 273663
rect 434530 272907 434558 275650
rect 434518 272901 434570 272907
rect 434518 272843 434570 272849
rect 436930 270465 436958 275650
rect 436918 270459 436970 270465
rect 436918 270401 436970 270407
rect 438082 264841 438110 275650
rect 438070 264835 438122 264841
rect 438070 264777 438122 264783
rect 440482 262103 440510 275650
rect 441730 266173 441758 275650
rect 444130 267875 444158 275650
rect 444118 267869 444170 267875
rect 444118 267811 444170 267817
rect 445282 266247 445310 275650
rect 446230 270089 446282 270095
rect 446230 270031 446282 270037
rect 445270 266241 445322 266247
rect 445270 266183 445322 266189
rect 441718 266167 441770 266173
rect 441718 266109 441770 266115
rect 440470 262097 440522 262103
rect 440470 262039 440522 262045
rect 431062 261579 431114 261585
rect 431062 261521 431114 261527
rect 425014 260469 425066 260475
rect 425014 260411 425066 260417
rect 446242 260253 446270 270031
rect 447094 267795 447146 267801
rect 447094 267737 447146 267743
rect 447106 267579 447134 267737
rect 447190 267721 447242 267727
rect 447190 267663 447242 267669
rect 447202 267579 447230 267663
rect 447094 267573 447146 267579
rect 447094 267515 447146 267521
rect 447190 267573 447242 267579
rect 447190 267515 447242 267521
rect 447682 262473 447710 275650
rect 448930 268985 448958 275650
rect 448918 268979 448970 268985
rect 448918 268921 448970 268927
rect 450850 267949 450878 275784
rect 453250 275719 453278 275784
rect 453238 275713 453290 275719
rect 453238 275655 453290 275661
rect 452386 269133 452414 275650
rect 452374 269127 452426 269133
rect 452374 269069 452426 269075
rect 450838 267943 450890 267949
rect 450838 267885 450890 267891
rect 454786 262621 454814 275650
rect 455650 267875 455678 275784
rect 455638 267869 455690 267875
rect 455638 267811 455690 267817
rect 455062 267795 455114 267801
rect 455062 267737 455114 267743
rect 454774 262615 454826 262621
rect 454774 262557 454826 262563
rect 455074 262547 455102 267737
rect 455062 262541 455114 262547
rect 455062 262483 455114 262489
rect 447670 262467 447722 262473
rect 447670 262409 447722 262415
rect 446230 260247 446282 260253
rect 446230 260189 446282 260195
rect 457186 259439 457214 275650
rect 458338 268023 458366 275650
rect 458326 268017 458378 268023
rect 458326 267959 458378 267965
rect 459586 267579 459614 275650
rect 460738 273647 460766 275650
rect 460726 273641 460778 273647
rect 460726 273583 460778 273589
rect 459862 271273 459914 271279
rect 459862 271215 459914 271221
rect 459874 270465 459902 271215
rect 459862 270459 459914 270465
rect 459862 270401 459914 270407
rect 459574 267573 459626 267579
rect 459574 267515 459626 267521
rect 461986 262695 462014 275650
rect 463138 267727 463166 275650
rect 464386 275571 464414 275650
rect 464374 275565 464426 275571
rect 464374 275507 464426 275513
rect 465538 268097 465566 275650
rect 465526 268091 465578 268097
rect 465526 268033 465578 268039
rect 463126 267721 463178 267727
rect 463126 267663 463178 267669
rect 466786 267505 466814 275784
rect 481858 275784 482160 275812
rect 497314 275784 497616 275812
rect 512770 275784 513072 275812
rect 528226 275784 528528 275812
rect 543682 275784 543984 275812
rect 559138 275784 559440 275812
rect 574594 275784 574896 275812
rect 590050 275784 590352 275812
rect 605506 275784 605808 275812
rect 620962 275784 621264 275812
rect 636514 275784 636720 275812
rect 467842 275497 467870 275650
rect 467830 275491 467882 275497
rect 467830 275433 467882 275439
rect 466774 267499 466826 267505
rect 466774 267441 466826 267447
rect 468994 262769 469022 275650
rect 470242 267431 470270 275650
rect 471394 275423 471422 275650
rect 471382 275417 471434 275423
rect 471382 275359 471434 275365
rect 472342 271199 472394 271205
rect 472342 271141 472394 271147
rect 472354 269207 472382 271141
rect 472342 269201 472394 269207
rect 472342 269143 472394 269149
rect 472642 268171 472670 275650
rect 472630 268165 472682 268171
rect 472630 268107 472682 268113
rect 470230 267425 470282 267431
rect 470230 267367 470282 267373
rect 473794 267357 473822 275650
rect 475042 275349 475070 275650
rect 475030 275343 475082 275349
rect 475030 275285 475082 275291
rect 473782 267351 473834 267357
rect 473782 267293 473834 267299
rect 476194 262843 476222 275650
rect 477442 267209 477470 275650
rect 478594 275275 478622 275650
rect 478582 275269 478634 275275
rect 478582 275211 478634 275217
rect 478774 268979 478826 268985
rect 478774 268921 478826 268927
rect 477430 267203 477482 267209
rect 477430 267145 477482 267151
rect 476182 262837 476234 262843
rect 476182 262779 476234 262785
rect 468982 262763 469034 262769
rect 468982 262705 469034 262711
rect 461974 262689 462026 262695
rect 461974 262631 462026 262637
rect 478786 260401 478814 268921
rect 479842 268245 479870 275650
rect 479830 268239 479882 268245
rect 479830 268181 479882 268187
rect 480994 267061 481022 275650
rect 481858 275201 481886 275784
rect 481846 275195 481898 275201
rect 481846 275137 481898 275143
rect 480982 267055 481034 267061
rect 480982 266997 481034 267003
rect 483298 262917 483326 275650
rect 484450 267135 484478 275650
rect 485698 275127 485726 275650
rect 485686 275121 485738 275127
rect 485686 275063 485738 275069
rect 486850 268319 486878 275650
rect 487810 275636 488112 275664
rect 486838 268313 486890 268319
rect 486838 268255 486890 268261
rect 484438 267129 484490 267135
rect 484438 267071 484490 267077
rect 487810 266987 487838 275636
rect 489250 275053 489278 275650
rect 489238 275047 489290 275053
rect 489238 274989 489290 274995
rect 488086 273567 488138 273573
rect 488086 273509 488138 273515
rect 488098 269133 488126 273509
rect 488086 269127 488138 269133
rect 488086 269069 488138 269075
rect 487798 266981 487850 266987
rect 487798 266923 487850 266929
rect 490498 262991 490526 275650
rect 491650 266839 491678 275650
rect 492898 274979 492926 275650
rect 492886 274973 492938 274979
rect 492886 274915 492938 274921
rect 494050 268393 494078 275650
rect 494038 268387 494090 268393
rect 494038 268329 494090 268335
rect 491638 266833 491690 266839
rect 491638 266775 491690 266781
rect 495298 266691 495326 275650
rect 496450 274905 496478 275650
rect 496438 274899 496490 274905
rect 496438 274841 496490 274847
rect 495286 266685 495338 266691
rect 495286 266627 495338 266633
rect 497314 263065 497342 275784
rect 498850 266543 498878 275650
rect 499906 274757 499934 275650
rect 499894 274751 499946 274757
rect 499894 274693 499946 274699
rect 501154 268467 501182 275650
rect 501142 268461 501194 268467
rect 501142 268403 501194 268409
rect 498838 266537 498890 266543
rect 498838 266479 498890 266485
rect 502306 266067 502334 275650
rect 503554 274831 503582 275650
rect 503542 274825 503594 274831
rect 503542 274767 503594 274773
rect 502678 271051 502730 271057
rect 502678 270993 502730 270999
rect 502690 269059 502718 270993
rect 502678 269053 502730 269059
rect 502678 268995 502730 269001
rect 502292 266058 502348 266067
rect 502292 265993 502348 266002
rect 504706 263139 504734 275650
rect 505954 267843 505982 275650
rect 507106 274683 507134 275650
rect 507094 274677 507146 274683
rect 507094 274619 507146 274625
rect 508246 270385 508298 270391
rect 508246 270327 508298 270333
rect 505940 267834 505996 267843
rect 505940 267769 505996 267778
rect 504694 263133 504746 263139
rect 504694 263075 504746 263081
rect 497302 263059 497354 263065
rect 497302 263001 497354 263007
rect 490486 262985 490538 262991
rect 490486 262927 490538 262933
rect 483286 262911 483338 262917
rect 483286 262853 483338 262859
rect 508258 260549 508286 270327
rect 508354 268541 508382 275650
rect 508342 268535 508394 268541
rect 508342 268477 508394 268483
rect 509506 266215 509534 275650
rect 510754 274609 510782 275650
rect 510742 274603 510794 274609
rect 510742 274545 510794 274551
rect 511906 267801 511934 275650
rect 511894 267795 511946 267801
rect 511894 267737 511946 267743
rect 512770 267399 512798 275784
rect 514306 274535 514334 275650
rect 514294 274529 514346 274535
rect 514294 274471 514346 274477
rect 515458 268615 515486 275650
rect 515446 268609 515498 268615
rect 515446 268551 515498 268557
rect 512756 267390 512812 267399
rect 512756 267325 512812 267334
rect 516610 267251 516638 275650
rect 517762 274461 517790 275650
rect 517750 274455 517802 274461
rect 517750 274397 517802 274403
rect 516596 267242 516652 267251
rect 516596 267177 516652 267186
rect 509492 266206 509548 266215
rect 509492 266141 509548 266150
rect 519010 263287 519038 275650
rect 520162 267103 520190 275650
rect 521410 274387 521438 275650
rect 521398 274381 521450 274387
rect 521398 274323 521450 274329
rect 521782 270163 521834 270169
rect 521782 270105 521834 270111
rect 520148 267094 520204 267103
rect 520148 267029 520204 267038
rect 518998 263281 519050 263287
rect 518998 263223 519050 263229
rect 521302 261579 521354 261585
rect 521302 261521 521354 261527
rect 508246 260543 508298 260549
rect 508246 260485 508298 260491
rect 478774 260395 478826 260401
rect 478774 260337 478826 260343
rect 457174 259433 457226 259439
rect 457174 259375 457226 259381
rect 463604 245634 463660 245643
rect 463604 245569 463660 245578
rect 440564 245338 440620 245347
rect 440564 245273 440620 245282
rect 440578 245009 440606 245273
rect 463618 245199 463646 245569
rect 463604 245190 463660 245199
rect 463604 245125 463660 245134
rect 440566 245003 440618 245009
rect 440566 244945 440618 244951
rect 521314 243423 521342 261521
rect 521794 260623 521822 270105
rect 522562 268689 522590 275650
rect 522550 268683 522602 268689
rect 522550 268625 522602 268631
rect 523810 266955 523838 275650
rect 524962 267653 524990 275650
rect 524950 267647 525002 267653
rect 524950 267589 525002 267595
rect 523796 266946 523852 266955
rect 523796 266881 523852 266890
rect 526210 263361 526238 275650
rect 527362 266807 527390 275650
rect 528226 274313 528254 275784
rect 528214 274307 528266 274313
rect 528214 274249 528266 274255
rect 529762 268763 529790 275650
rect 529750 268757 529802 268763
rect 529750 268699 529802 268705
rect 527348 266798 527404 266807
rect 527348 266733 527404 266742
rect 530914 266659 530942 275650
rect 532162 274239 532190 275650
rect 532150 274233 532202 274239
rect 532150 274175 532202 274181
rect 530900 266650 530956 266659
rect 530900 266585 530956 266594
rect 533218 263435 533246 275650
rect 534466 266511 534494 275650
rect 535618 274165 535646 275650
rect 535606 274159 535658 274165
rect 535606 274101 535658 274107
rect 536866 268837 536894 275650
rect 536854 268831 536906 268837
rect 536854 268773 536906 268779
rect 534452 266502 534508 266511
rect 534452 266437 534508 266446
rect 538018 266363 538046 275650
rect 539266 274091 539294 275650
rect 539254 274085 539306 274091
rect 539254 274027 539306 274033
rect 538004 266354 538060 266363
rect 538004 266289 538060 266298
rect 540418 263509 540446 275650
rect 540406 263503 540458 263509
rect 540406 263445 540458 263451
rect 533206 263429 533258 263435
rect 533206 263371 533258 263377
rect 526198 263355 526250 263361
rect 526198 263297 526250 263303
rect 541666 261067 541694 275650
rect 542818 274017 542846 275650
rect 542806 274011 542858 274017
rect 542806 273953 542858 273959
rect 543682 268911 543710 275784
rect 545218 272537 545246 275650
rect 546370 273943 546398 275650
rect 546358 273937 546410 273943
rect 546358 273879 546410 273885
rect 545206 272531 545258 272537
rect 545206 272473 545258 272479
rect 543670 268905 543722 268911
rect 543670 268847 543722 268853
rect 547618 264989 547646 275650
rect 548770 268731 548798 275650
rect 548756 268722 548812 268731
rect 548756 268657 548812 268666
rect 549922 267283 549950 275650
rect 550102 273493 550154 273499
rect 550102 273435 550154 273441
rect 550114 268911 550142 273435
rect 550102 268905 550154 268911
rect 550102 268847 550154 268853
rect 549910 267277 549962 267283
rect 549910 267219 549962 267225
rect 548566 266537 548618 266543
rect 548566 266479 548618 266485
rect 547606 264983 547658 264989
rect 547606 264925 547658 264931
rect 548578 261585 548606 266479
rect 551074 266321 551102 275650
rect 551062 266315 551114 266321
rect 551062 266257 551114 266263
rect 548566 261579 548618 261585
rect 548566 261521 548618 261527
rect 541654 261061 541706 261067
rect 541654 261003 541706 261009
rect 552322 260993 552350 275650
rect 553474 266913 553502 275650
rect 554722 270317 554750 275650
rect 554710 270311 554762 270317
rect 554710 270253 554762 270259
rect 553462 266907 553514 266913
rect 553462 266849 553514 266855
rect 552310 260987 552362 260993
rect 552310 260929 552362 260935
rect 555874 260771 555902 275650
rect 557122 266765 557150 275650
rect 558274 268985 558302 275650
rect 558262 268979 558314 268985
rect 558262 268921 558314 268927
rect 557110 266759 557162 266765
rect 557110 266701 557162 266707
rect 555862 260765 555914 260771
rect 555862 260707 555914 260713
rect 521782 260617 521834 260623
rect 521782 260559 521834 260565
rect 559138 260295 559166 275784
rect 560674 266617 560702 275650
rect 561826 269207 561854 275650
rect 562198 270903 562250 270909
rect 562198 270845 562250 270851
rect 562210 270317 562238 270845
rect 562198 270311 562250 270317
rect 562198 270253 562250 270259
rect 561814 269201 561866 269207
rect 561814 269143 561866 269149
rect 560662 266611 560714 266617
rect 560662 266553 560714 266559
rect 563074 260443 563102 275650
rect 564226 266469 564254 275650
rect 564214 266463 564266 266469
rect 564214 266405 564266 266411
rect 565474 261511 565502 275650
rect 566530 262071 566558 275650
rect 567778 267695 567806 275650
rect 568930 270243 568958 275650
rect 568918 270237 568970 270243
rect 568918 270179 568970 270185
rect 567764 267686 567820 267695
rect 567764 267621 567820 267630
rect 566516 262062 566572 262071
rect 566516 261997 566572 262006
rect 570178 261775 570206 275650
rect 570262 270829 570314 270835
rect 570262 270771 570314 270777
rect 570274 269207 570302 270771
rect 570262 269201 570314 269207
rect 570262 269143 570314 269149
rect 571330 266395 571358 275650
rect 572578 269133 572606 275650
rect 573142 275047 573194 275053
rect 573142 274989 573194 274995
rect 572566 269127 572618 269133
rect 572566 269069 572618 269075
rect 573154 266543 573182 274989
rect 573142 266537 573194 266543
rect 573142 266479 573194 266485
rect 571318 266389 571370 266395
rect 571318 266331 571370 266337
rect 570164 261766 570220 261775
rect 570164 261701 570220 261710
rect 565462 261505 565514 261511
rect 573730 261479 573758 275650
rect 574594 267547 574622 275784
rect 576130 270095 576158 275650
rect 576118 270089 576170 270095
rect 576118 270031 576170 270037
rect 574580 267538 574636 267547
rect 574580 267473 574636 267482
rect 565462 261447 565514 261453
rect 573716 261470 573772 261479
rect 573716 261405 573772 261414
rect 577282 261331 577310 275650
rect 578530 261437 578558 275650
rect 579682 270465 579710 275650
rect 579670 270459 579722 270465
rect 579670 270401 579722 270407
rect 578518 261431 578570 261437
rect 578518 261373 578570 261379
rect 577268 261322 577324 261331
rect 577268 261257 577324 261266
rect 580930 261183 580958 275650
rect 582082 272833 582110 275650
rect 582070 272827 582122 272833
rect 582070 272769 582122 272775
rect 583234 270021 583262 275650
rect 583222 270015 583274 270021
rect 583222 269957 583274 269963
rect 580916 261174 580972 261183
rect 580916 261109 580972 261118
rect 584386 261035 584414 275650
rect 585634 261363 585662 275650
rect 586786 269059 586814 275650
rect 586774 269053 586826 269059
rect 586774 268995 586826 269001
rect 585622 261357 585674 261363
rect 585622 261299 585674 261305
rect 584372 261026 584428 261035
rect 584372 260961 584428 260970
rect 588034 260887 588062 275650
rect 589186 272759 589214 275650
rect 589174 272753 589226 272759
rect 589174 272695 589226 272701
rect 588886 271495 588938 271501
rect 588886 271437 588938 271443
rect 588898 270243 588926 271437
rect 588886 270237 588938 270243
rect 588886 270179 588938 270185
rect 590050 269873 590078 275784
rect 591586 272241 591614 275650
rect 591574 272235 591626 272241
rect 591574 272177 591626 272183
rect 590038 269867 590090 269873
rect 590038 269809 590090 269815
rect 592738 261289 592766 275650
rect 593986 269947 594014 275650
rect 595138 272167 595166 275650
rect 596386 272685 596414 275650
rect 596374 272679 596426 272685
rect 596374 272621 596426 272627
rect 595126 272161 595178 272167
rect 595126 272103 595178 272109
rect 597538 270539 597566 275650
rect 598786 271987 598814 275650
rect 598772 271978 598828 271987
rect 598772 271913 598828 271922
rect 597526 270533 597578 270539
rect 597526 270475 597578 270481
rect 593974 269941 594026 269947
rect 593974 269883 594026 269889
rect 592726 261283 592778 261289
rect 592726 261225 592778 261231
rect 599842 261215 599870 275650
rect 601090 270391 601118 275650
rect 602242 273467 602270 275650
rect 602228 273458 602284 273467
rect 602228 273393 602284 273402
rect 603490 272611 603518 275650
rect 603478 272605 603530 272611
rect 603478 272547 603530 272553
rect 604642 270613 604670 275650
rect 605506 273615 605534 275784
rect 605492 273606 605548 273615
rect 605492 273541 605548 273550
rect 604630 270607 604682 270613
rect 604630 270549 604682 270555
rect 601078 270385 601130 270391
rect 601078 270327 601130 270333
rect 599830 261209 599882 261215
rect 599830 261151 599882 261157
rect 607042 261141 607070 275650
rect 608194 269799 608222 275650
rect 609442 273319 609470 275650
rect 609428 273310 609484 273319
rect 609428 273245 609484 273254
rect 610594 272463 610622 275650
rect 610582 272457 610634 272463
rect 610582 272399 610634 272405
rect 608182 269793 608234 269799
rect 608182 269735 608234 269741
rect 611842 269651 611870 275650
rect 612994 273171 613022 275650
rect 612980 273162 613036 273171
rect 612980 273097 613036 273106
rect 611830 269645 611882 269651
rect 611830 269587 611882 269593
rect 607030 261135 607082 261141
rect 607030 261077 607082 261083
rect 614242 260919 614270 275650
rect 615394 268911 615422 275650
rect 616546 273023 616574 275650
rect 616532 273014 616588 273023
rect 616532 272949 616588 272958
rect 617698 272389 617726 275650
rect 617686 272383 617738 272389
rect 617686 272325 617738 272331
rect 618946 269577 618974 275650
rect 620098 272875 620126 275650
rect 620084 272866 620140 272875
rect 620084 272801 620140 272810
rect 618934 269571 618986 269577
rect 618934 269513 618986 269519
rect 615382 268905 615434 268911
rect 615382 268847 615434 268853
rect 614230 260913 614282 260919
rect 588020 260878 588076 260887
rect 614230 260855 614282 260861
rect 620962 260845 620990 275784
rect 622498 270169 622526 275650
rect 623650 272727 623678 275650
rect 623636 272718 623692 272727
rect 623636 272653 623692 272662
rect 624898 272315 624926 275650
rect 624886 272309 624938 272315
rect 624886 272251 624938 272257
rect 626050 270687 626078 275650
rect 627298 272579 627326 275650
rect 627284 272570 627340 272579
rect 627284 272505 627340 272514
rect 626038 270681 626090 270687
rect 626038 270623 626090 270629
rect 622486 270163 622538 270169
rect 622486 270105 622538 270111
rect 628450 261923 628478 275650
rect 629698 269503 629726 275650
rect 630850 272431 630878 275650
rect 630836 272422 630892 272431
rect 630836 272357 630892 272366
rect 632098 270243 632126 275650
rect 632086 270237 632138 270243
rect 632086 270179 632138 270185
rect 633154 269725 633182 275650
rect 633142 269719 633194 269725
rect 633142 269661 633194 269667
rect 629686 269497 629738 269503
rect 629686 269439 629738 269445
rect 628436 261914 628492 261923
rect 628436 261849 628492 261858
rect 588020 260813 588076 260822
rect 620950 260839 621002 260845
rect 620950 260781 621002 260787
rect 634402 260739 634430 275650
rect 635554 261627 635582 275650
rect 636514 269429 636542 275784
rect 636502 269423 636554 269429
rect 636502 269365 636554 269371
rect 635540 261618 635596 261627
rect 635540 261553 635596 261562
rect 634388 260730 634444 260739
rect 634388 260665 634444 260674
rect 637954 260591 637982 275650
rect 639106 269207 639134 275650
rect 640354 269355 640382 275650
rect 641506 272283 641534 275650
rect 641492 272274 641548 272283
rect 641492 272209 641548 272218
rect 640342 269349 640394 269355
rect 640342 269291 640394 269297
rect 639094 269201 639146 269207
rect 639094 269143 639146 269149
rect 642754 260697 642782 275650
rect 643906 269281 643934 275650
rect 645154 272135 645182 275650
rect 645140 272126 645196 272135
rect 645140 272061 645196 272070
rect 646306 270317 646334 275650
rect 646294 270311 646346 270317
rect 646294 270253 646346 270259
rect 643894 269275 643946 269281
rect 643894 269217 643946 269223
rect 647554 269027 647582 275650
rect 647540 269018 647596 269027
rect 647540 268953 647596 268962
rect 648706 263551 648734 275650
rect 649378 275053 649406 987757
rect 649462 984929 649514 984935
rect 649462 984871 649514 984877
rect 649474 275645 649502 984871
rect 649570 951857 649598 993857
rect 649654 983819 649706 983825
rect 649654 983761 649706 983767
rect 649558 951851 649610 951857
rect 649558 951793 649610 951799
rect 649558 927431 649610 927437
rect 649558 927373 649610 927379
rect 649462 275639 649514 275645
rect 649462 275581 649514 275587
rect 649366 275047 649418 275053
rect 649366 274989 649418 274995
rect 648692 263542 648748 263551
rect 648692 263477 648748 263486
rect 642742 260691 642794 260697
rect 642742 260633 642794 260639
rect 637940 260582 637996 260591
rect 637940 260517 637996 260526
rect 563060 260434 563116 260443
rect 563060 260369 563116 260378
rect 559124 260286 559180 260295
rect 559124 260221 559180 260230
rect 639286 256399 639338 256405
rect 639286 256341 639338 256347
rect 494516 243414 494572 243423
rect 494516 243349 494572 243358
rect 521300 243414 521356 243423
rect 521300 243349 521356 243358
rect 421844 242230 421900 242239
rect 421844 242165 421900 242174
rect 415316 240454 415372 240463
rect 415316 240389 415372 240398
rect 421858 239089 421886 242165
rect 494530 242091 494558 243349
rect 494516 242082 494572 242091
rect 494516 242017 494572 242026
rect 494530 239385 494558 242017
rect 549046 240489 549098 240495
rect 549046 240431 549098 240437
rect 494518 239379 494570 239385
rect 494518 239321 494570 239327
rect 497206 239379 497258 239385
rect 497206 239321 497258 239327
rect 420598 239083 420650 239089
rect 420598 239025 420650 239031
rect 421846 239083 421898 239089
rect 421846 239025 421898 239031
rect 420610 233780 420638 239025
rect 420562 233752 420638 233780
rect 420562 233618 420590 233752
rect 497218 233632 497246 239321
rect 505556 239270 505612 239279
rect 505556 239205 505558 239214
rect 505610 239205 505612 239214
rect 505558 239173 505610 239179
rect 414838 233607 414890 233613
rect 306932 233581 306988 233590
rect 497218 233604 497472 233632
rect 505570 233618 505598 239173
rect 510370 239163 510398 239191
rect 510358 239157 510410 239163
rect 510356 239122 510358 239131
rect 510410 239122 510412 239131
rect 549058 239089 549086 240431
rect 637558 239601 637610 239607
rect 637558 239543 637610 239549
rect 510356 239057 510412 239066
rect 541462 239083 541514 239089
rect 510370 233618 510398 239057
rect 541462 239025 541514 239031
rect 549046 239083 549098 239089
rect 549046 239025 549098 239031
rect 541474 234691 541502 239025
rect 541460 234682 541516 234691
rect 541460 234617 541516 234626
rect 549058 233928 549086 239025
rect 549010 233900 549086 233928
rect 549010 233618 549038 233900
rect 637172 233794 637228 233803
rect 637172 233729 637228 233738
rect 637186 233632 637214 233729
rect 637570 233632 637598 239543
rect 638038 239527 638090 239533
rect 638038 239469 638090 239475
rect 637654 239453 637706 239459
rect 637654 239395 637706 239401
rect 637666 233951 637694 239395
rect 638050 234099 638078 239469
rect 638806 239379 638858 239385
rect 638806 239321 638858 239327
rect 638420 239122 638476 239131
rect 638420 239057 638476 239066
rect 638036 234090 638092 234099
rect 638036 234025 638092 234034
rect 637652 233942 637708 233951
rect 637652 233877 637708 233886
rect 637186 233604 637598 233632
rect 637666 233618 637694 233877
rect 638050 233618 638078 234025
rect 638132 233646 638188 233655
rect 638434 233632 638462 239057
rect 638188 233618 638462 233632
rect 638516 233646 638572 233655
rect 638188 233604 638448 233618
rect 638132 233581 638188 233590
rect 638818 233632 638846 239321
rect 639298 239131 639326 256341
rect 649570 239385 649598 927373
rect 649666 752395 649694 983761
rect 649846 981821 649898 981827
rect 649846 981763 649898 981769
rect 649652 752386 649708 752395
rect 649652 752321 649708 752330
rect 649654 748869 649706 748875
rect 649654 748811 649706 748817
rect 649558 239379 649610 239385
rect 649558 239321 649610 239327
rect 639382 239305 639434 239311
rect 639382 239247 639434 239253
rect 639284 239122 639340 239131
rect 639284 239057 639340 239066
rect 639284 233794 639340 233803
rect 639284 233729 639340 233738
rect 639298 233632 639326 233729
rect 639394 233632 639422 239247
rect 639766 239083 639818 239089
rect 639766 239025 639818 239031
rect 639778 233632 639806 239025
rect 638572 233604 638846 233632
rect 639168 233604 639422 233632
rect 639552 233604 639806 233632
rect 638516 233581 638572 233590
rect 414838 233549 414890 233555
rect 305376 233456 305438 233484
rect 210178 208592 210302 208620
rect 210178 169973 210206 208592
rect 210262 208521 210314 208527
rect 210262 208463 210314 208469
rect 210166 169967 210218 169973
rect 210166 169909 210218 169915
rect 210164 161274 210220 161283
rect 210164 161209 210220 161218
rect 210178 153291 210206 161209
rect 210164 153282 210220 153291
rect 210164 153217 210220 153226
rect 210166 148285 210218 148291
rect 210166 148227 210218 148233
rect 210070 147027 210122 147033
rect 210070 146969 210122 146975
rect 209974 146805 210026 146811
rect 209974 146747 210026 146753
rect 210178 146756 210206 148227
rect 210274 146885 210302 208463
rect 210262 146879 210314 146885
rect 210262 146821 210314 146827
rect 209986 127053 210014 146747
rect 210070 146731 210122 146737
rect 210178 146728 210302 146756
rect 210070 146673 210122 146679
rect 209974 127047 210026 127053
rect 209974 126989 210026 126995
rect 209974 126751 210026 126757
rect 209974 126693 210026 126699
rect 209986 71891 210014 126693
rect 209972 71882 210028 71891
rect 209972 71817 210028 71826
rect 209974 71769 210026 71775
rect 209974 71711 210026 71717
rect 209986 71225 210014 71711
rect 209972 71216 210028 71225
rect 209972 71151 210028 71160
rect 209972 60856 210028 60865
rect 209972 60791 210028 60800
rect 209986 60675 210014 60791
rect 209974 60669 210026 60675
rect 209974 60611 210026 60617
rect 209974 60373 210026 60379
rect 209974 60315 210026 60321
rect 209986 59237 210014 60315
rect 209972 59228 210028 59237
rect 209972 59163 210028 59172
rect 209972 58118 210028 58127
rect 209972 58053 210028 58062
rect 209986 53127 210014 58053
rect 210082 54385 210110 146673
rect 210274 126924 210302 146728
rect 210178 126896 210302 126924
rect 210178 126757 210206 126896
rect 210166 126751 210218 126757
rect 210166 126693 210218 126699
rect 210262 126751 210314 126757
rect 210262 126693 210314 126699
rect 210166 103515 210218 103521
rect 210166 103457 210218 103463
rect 210178 101121 210206 103457
rect 210164 101112 210220 101121
rect 210164 101047 210220 101056
rect 210166 100555 210218 100561
rect 210166 100497 210218 100503
rect 210178 99493 210206 100497
rect 210164 99484 210220 99493
rect 210164 99419 210220 99428
rect 210164 97856 210220 97865
rect 210164 97791 210166 97800
rect 210218 97791 210220 97800
rect 210166 97759 210218 97765
rect 210166 97521 210218 97527
rect 210166 97463 210218 97469
rect 210178 96237 210206 97463
rect 210164 96228 210220 96237
rect 210164 96163 210220 96172
rect 210166 94857 210218 94863
rect 210166 94799 210218 94805
rect 210178 94609 210206 94799
rect 210164 94600 210220 94609
rect 210164 94535 210220 94544
rect 210164 87718 210220 87727
rect 210164 87653 210220 87662
rect 210178 62895 210206 87653
rect 210274 83435 210302 126693
rect 210260 83426 210316 83435
rect 210260 83361 210316 83370
rect 210260 77728 210316 77737
rect 210260 77663 210316 77672
rect 210274 77399 210302 77663
rect 210262 77393 210314 77399
rect 210262 77335 210314 77341
rect 210262 74507 210314 74513
rect 210260 74472 210262 74481
rect 210314 74472 210316 74481
rect 210260 74407 210316 74416
rect 210166 62889 210218 62895
rect 210166 62831 210218 62837
rect 210164 57082 210220 57091
rect 210164 57017 210220 57026
rect 210070 54379 210122 54385
rect 210070 54321 210122 54327
rect 210068 54122 210124 54131
rect 210068 54057 210124 54066
rect 209974 53121 210026 53127
rect 209974 53063 210026 53069
rect 210082 52905 210110 54057
rect 210178 53201 210206 57017
rect 210260 56490 210316 56499
rect 210260 56425 210316 56434
rect 210274 53645 210302 56425
rect 210356 54418 210412 54427
rect 210356 54353 210412 54362
rect 210644 54418 210700 54427
rect 220628 54418 220684 54427
rect 213744 54385 213854 54404
rect 215952 54385 216062 54404
rect 213744 54379 213866 54385
rect 213744 54376 213814 54379
rect 210644 54353 210700 54362
rect 210262 53639 210314 53645
rect 210262 53581 210314 53587
rect 210370 53571 210398 54353
rect 210658 53867 210686 54353
rect 213814 54321 213866 54327
rect 214198 54379 214250 54385
rect 215952 54379 216074 54385
rect 215952 54376 216022 54379
rect 214198 54321 214250 54327
rect 216022 54321 216074 54327
rect 218818 54376 218928 54404
rect 214210 54131 214238 54321
rect 216406 54305 216458 54311
rect 218612 54270 218668 54279
rect 216458 54253 216528 54256
rect 216406 54247 216528 54253
rect 216418 54228 216528 54247
rect 218160 54237 218270 54256
rect 218160 54231 218282 54237
rect 218160 54228 218230 54231
rect 218612 54205 218668 54214
rect 218230 54173 218282 54179
rect 214196 54122 214252 54131
rect 218626 54108 218654 54205
rect 218242 54089 218352 54108
rect 214196 54057 214252 54066
rect 218230 54083 218352 54089
rect 218282 54080 218352 54083
rect 218626 54080 218736 54108
rect 218230 54025 218282 54031
rect 218422 54009 218474 54015
rect 214848 53932 214910 53960
rect 216226 53941 216336 53960
rect 210646 53861 210698 53867
rect 210646 53803 210698 53809
rect 210754 53784 211008 53812
rect 211138 53784 211200 53812
rect 210358 53565 210410 53571
rect 210358 53507 210410 53513
rect 210166 53195 210218 53201
rect 210166 53137 210218 53143
rect 210070 52899 210122 52905
rect 210070 52841 210122 52847
rect 209878 51863 209930 51869
rect 209878 51805 209930 51811
rect 209302 48829 209354 48835
rect 209302 48771 209354 48777
rect 209014 48681 209066 48687
rect 209014 48623 209066 48629
rect 208726 48607 208778 48613
rect 208726 48549 208778 48555
rect 208822 48607 208874 48613
rect 208822 48549 208874 48555
rect 208738 48243 208766 48549
rect 208630 48237 208682 48243
rect 208630 48179 208682 48185
rect 208726 48237 208778 48243
rect 208726 48179 208778 48185
rect 208438 48163 208490 48169
rect 208438 48105 208490 48111
rect 208534 48163 208586 48169
rect 208534 48105 208586 48111
rect 208246 48089 208298 48095
rect 208246 48031 208298 48037
rect 208150 48015 208202 48021
rect 208150 47957 208202 47963
rect 208054 47571 208106 47577
rect 208054 47513 208106 47519
rect 208450 47503 208478 48105
rect 208438 47497 208490 47503
rect 208438 47439 208490 47445
rect 207286 42169 207338 42175
rect 207286 42111 207338 42117
rect 187604 41838 187660 41847
rect 187344 41796 187604 41824
rect 194324 41838 194380 41847
rect 194064 41796 194324 41824
rect 187604 41773 187660 41782
rect 194324 41773 194380 41782
rect 210754 40811 210782 53784
rect 211138 51573 211166 53784
rect 211126 51567 211178 51573
rect 211126 51509 211178 51515
rect 210838 50309 210890 50315
rect 210838 50251 210890 50257
rect 210850 49723 210878 50251
rect 210838 49717 210890 49723
rect 210838 49659 210890 49665
rect 211330 45251 211358 53798
rect 211522 51499 211550 53798
rect 211510 51493 211562 51499
rect 211510 51435 211562 51441
rect 211316 45242 211372 45251
rect 211316 45177 211372 45186
rect 211714 45103 211742 53798
rect 211796 53530 211852 53539
rect 211796 53465 211852 53474
rect 211810 53053 211838 53465
rect 211798 53047 211850 53053
rect 211798 52989 211850 52995
rect 211906 51911 211934 53798
rect 211892 51902 211948 51911
rect 211892 51837 211948 51846
rect 212098 45399 212126 53798
rect 212290 52239 212318 53798
rect 212278 52233 212330 52239
rect 212278 52175 212330 52181
rect 212084 45390 212140 45399
rect 212084 45325 212140 45334
rect 211700 45094 211756 45103
rect 211700 45029 211756 45038
rect 212482 42397 212510 53798
rect 212640 53784 212702 53812
rect 212832 53784 212894 53812
rect 212674 52059 212702 53784
rect 212660 52050 212716 52059
rect 212660 51985 212716 51994
rect 212866 44839 212894 53784
rect 213010 53664 213038 53798
rect 212962 53636 213038 53664
rect 213154 53784 213216 53812
rect 213346 53784 213408 53812
rect 212962 53391 212990 53636
rect 212948 53382 213004 53391
rect 212948 53317 213004 53326
rect 213154 44955 213182 53784
rect 213346 51795 213374 53784
rect 213334 51789 213386 51795
rect 213334 51731 213386 51737
rect 213140 44946 213196 44955
rect 213140 44881 213196 44890
rect 212854 44833 212906 44839
rect 212854 44775 212906 44781
rect 212470 42391 212522 42397
rect 212470 42333 212522 42339
rect 213538 42101 213566 53798
rect 213922 44765 213950 53798
rect 214114 51721 214142 53798
rect 214102 51715 214154 51721
rect 214102 51657 214154 51663
rect 213910 44759 213962 44765
rect 213910 44701 213962 44707
rect 213526 42095 213578 42101
rect 213526 42037 213578 42043
rect 214306 41731 214334 53798
rect 214498 51869 214526 53798
rect 214486 51863 214538 51869
rect 214486 51805 214538 51811
rect 214690 44691 214718 53798
rect 214882 53539 214910 53932
rect 216214 53935 216336 53941
rect 216266 53932 216336 53935
rect 217248 53932 217310 53960
rect 218422 53951 218474 53957
rect 216214 53877 216266 53883
rect 215040 53784 215102 53812
rect 214868 53530 214924 53539
rect 214868 53465 214924 53474
rect 215074 44807 215102 53784
rect 215218 53650 215246 53798
rect 215362 53784 215424 53812
rect 215554 53784 215616 53812
rect 215204 53641 215260 53650
rect 215204 53576 215260 53585
rect 215060 44798 215116 44807
rect 215060 44733 215116 44742
rect 214678 44685 214730 44691
rect 215362 44659 215390 53784
rect 215554 53275 215582 53784
rect 215542 53269 215594 53275
rect 215542 53211 215594 53217
rect 215746 52165 215774 53798
rect 216130 52609 216158 53798
rect 216706 53095 216734 53798
rect 216692 53086 216748 53095
rect 216692 53021 216748 53030
rect 216118 52603 216170 52609
rect 216118 52545 216170 52551
rect 215734 52159 215786 52165
rect 215734 52101 215786 52107
rect 216898 52017 216926 53798
rect 217042 53650 217070 53798
rect 217028 53641 217084 53650
rect 217028 53576 217084 53585
rect 217282 53497 217310 53932
rect 217426 53664 217454 53798
rect 217378 53636 217454 53664
rect 217570 53784 217632 53812
rect 217270 53491 217322 53497
rect 217270 53433 217322 53439
rect 217378 53349 217406 53636
rect 217570 53423 217598 53784
rect 217810 53571 217838 53798
rect 217798 53565 217850 53571
rect 217798 53507 217850 53513
rect 217558 53417 217610 53423
rect 217558 53359 217610 53365
rect 217366 53343 217418 53349
rect 217366 53285 217418 53291
rect 217954 52461 217982 53798
rect 218434 53497 218462 53951
rect 218544 53784 218654 53812
rect 218422 53491 218474 53497
rect 218422 53433 218474 53439
rect 217942 52455 217994 52461
rect 217942 52397 217994 52403
rect 216886 52011 216938 52017
rect 216886 51953 216938 51959
rect 218626 49131 218654 53784
rect 218818 52905 218846 54376
rect 220628 54353 220684 54362
rect 220438 54157 220490 54163
rect 220368 54105 220438 54108
rect 220368 54099 220490 54105
rect 220368 54080 220478 54099
rect 218806 52899 218858 52905
rect 218806 52841 218858 52847
rect 218614 49125 218666 49131
rect 218614 49067 218666 49073
rect 219106 48835 219134 53798
rect 219264 53784 219326 53812
rect 219298 52979 219326 53784
rect 219442 53645 219470 53798
rect 219430 53639 219482 53645
rect 219430 53581 219482 53587
rect 219634 53516 219662 53798
rect 219586 53497 219662 53516
rect 219574 53491 219662 53497
rect 219626 53488 219662 53491
rect 219778 53784 219840 53812
rect 219970 53784 220032 53812
rect 219574 53433 219626 53439
rect 219286 52973 219338 52979
rect 219286 52915 219338 52921
rect 219478 51789 219530 51795
rect 219478 51731 219530 51737
rect 219490 51499 219518 51731
rect 219478 51493 219530 51499
rect 219478 51435 219530 51441
rect 219094 48829 219146 48835
rect 219094 48771 219146 48777
rect 219778 48687 219806 53784
rect 219970 48803 219998 53784
rect 219956 48794 220012 48803
rect 219956 48729 220012 48738
rect 219766 48681 219818 48687
rect 219766 48623 219818 48629
rect 220162 48243 220190 53798
rect 220438 52233 220490 52239
rect 220438 52175 220490 52181
rect 220450 51869 220478 52175
rect 220438 51863 220490 51869
rect 220438 51805 220490 51811
rect 220546 48613 220574 53798
rect 220642 53497 220670 54353
rect 229652 53974 229708 53983
rect 229652 53909 229708 53918
rect 220630 53491 220682 53497
rect 220630 53433 220682 53439
rect 220534 48607 220586 48613
rect 220534 48549 220586 48555
rect 220150 48237 220202 48243
rect 220150 48179 220202 48185
rect 220738 47767 220766 53798
rect 220930 52091 220958 53798
rect 221122 53243 221150 53798
rect 221108 53234 221164 53243
rect 221108 53169 221164 53178
rect 220918 52085 220970 52091
rect 220918 52027 220970 52033
rect 220724 47758 220780 47767
rect 221314 47725 221342 53798
rect 221458 53645 221486 53798
rect 221664 53784 221726 53812
rect 221446 53639 221498 53645
rect 221446 53581 221498 53587
rect 221698 47799 221726 53784
rect 221842 53516 221870 53798
rect 221986 53784 222048 53812
rect 222178 53784 222240 53812
rect 221842 53488 221918 53516
rect 221782 53121 221834 53127
rect 221782 53063 221834 53069
rect 221794 52979 221822 53063
rect 221782 52973 221834 52979
rect 221782 52915 221834 52921
rect 221890 52651 221918 53488
rect 221876 52642 221932 52651
rect 221876 52577 221932 52586
rect 221986 48169 222014 53784
rect 222178 48761 222206 53784
rect 222166 48755 222218 48761
rect 222166 48697 222218 48703
rect 221974 48163 222026 48169
rect 221974 48105 222026 48111
rect 222370 48095 222398 53798
rect 222562 52503 222590 53798
rect 222548 52494 222604 52503
rect 222548 52429 222604 52438
rect 222358 48089 222410 48095
rect 222358 48031 222410 48037
rect 222754 48021 222782 53798
rect 222946 48835 222974 53798
rect 223138 50167 223166 53798
rect 223330 52207 223358 53798
rect 223316 52198 223372 52207
rect 223316 52133 223372 52142
rect 223126 50161 223178 50167
rect 223126 50103 223178 50109
rect 223522 50093 223550 53798
rect 223680 53784 223742 53812
rect 223872 53784 223934 53812
rect 223714 52355 223742 53784
rect 223700 52346 223756 52355
rect 223700 52281 223756 52290
rect 223606 52011 223658 52017
rect 223606 51953 223658 51959
rect 223618 51647 223646 51953
rect 223606 51641 223658 51647
rect 223606 51583 223658 51589
rect 223510 50087 223562 50093
rect 223510 50029 223562 50035
rect 222934 48829 222986 48835
rect 222934 48771 222986 48777
rect 222742 48015 222794 48021
rect 222742 47957 222794 47963
rect 223906 47947 223934 53784
rect 224050 53516 224078 53798
rect 224194 53784 224256 53812
rect 224050 53488 224126 53516
rect 224098 48909 224126 53488
rect 224194 50019 224222 53784
rect 224182 50013 224234 50019
rect 224182 49955 224234 49961
rect 224086 48903 224138 48909
rect 224086 48845 224138 48851
rect 223894 47941 223946 47947
rect 223894 47883 223946 47889
rect 221686 47793 221738 47799
rect 221686 47735 221738 47741
rect 220724 47693 220780 47702
rect 221302 47719 221354 47725
rect 221302 47661 221354 47667
rect 224578 47577 224606 53798
rect 224962 50463 224990 53798
rect 224950 50457 225002 50463
rect 224950 50399 225002 50405
rect 224566 47571 224618 47577
rect 224566 47513 224618 47519
rect 225346 47503 225374 53798
rect 225730 50241 225758 53798
rect 226080 53784 226142 53812
rect 226114 50389 226142 53784
rect 226402 53784 226464 53812
rect 226102 50383 226154 50389
rect 226102 50325 226154 50331
rect 225718 50235 225770 50241
rect 225718 50177 225770 50183
rect 226402 48687 226430 53784
rect 226786 49723 226814 53798
rect 227170 50315 227198 53798
rect 227554 51943 227582 53798
rect 227542 51937 227594 51943
rect 227542 51879 227594 51885
rect 227158 50309 227210 50315
rect 227158 50251 227210 50257
rect 226774 49717 226826 49723
rect 226774 49659 226826 49665
rect 226390 48681 226442 48687
rect 226390 48623 226442 48629
rect 227938 48391 227966 53798
rect 228034 53784 228288 53812
rect 228418 53784 228672 53812
rect 227926 48385 227978 48391
rect 227926 48327 227978 48333
rect 225334 47497 225386 47503
rect 225334 47439 225386 47445
rect 228034 46541 228062 53784
rect 228418 50759 228446 53784
rect 228994 50907 229022 53798
rect 228982 50901 229034 50907
rect 228982 50843 229034 50849
rect 228406 50753 228458 50759
rect 228406 50695 228458 50701
rect 229378 50611 229406 53798
rect 229666 53391 229694 53909
rect 229652 53382 229708 53391
rect 229652 53317 229708 53326
rect 229762 50685 229790 53798
rect 229750 50679 229802 50685
rect 229750 50621 229802 50627
rect 229366 50605 229418 50611
rect 229366 50547 229418 50553
rect 230146 48317 230174 53798
rect 230496 53784 230558 53812
rect 230530 50981 230558 53784
rect 230626 53784 230880 53812
rect 230518 50975 230570 50981
rect 230518 50917 230570 50923
rect 230134 48311 230186 48317
rect 230134 48253 230186 48259
rect 230626 46763 230654 53784
rect 231202 51129 231230 53798
rect 231190 51123 231242 51129
rect 231190 51065 231242 51071
rect 231586 51055 231614 53798
rect 231766 53639 231818 53645
rect 231766 53581 231818 53587
rect 231778 52979 231806 53581
rect 231766 52973 231818 52979
rect 231766 52915 231818 52921
rect 231970 51203 231998 53798
rect 231958 51197 232010 51203
rect 231958 51139 232010 51145
rect 231574 51049 231626 51055
rect 231574 50991 231626 50997
rect 230614 46757 230666 46763
rect 230614 46699 230666 46705
rect 232354 46615 232382 53798
rect 232450 53784 232704 53812
rect 232834 53784 233088 53812
rect 232450 49797 232478 53784
rect 232438 49791 232490 49797
rect 232438 49733 232490 49739
rect 232834 46689 232862 53784
rect 233410 47429 233438 53798
rect 233794 51425 233822 53798
rect 233782 51419 233834 51425
rect 233782 51361 233834 51367
rect 233398 47423 233450 47429
rect 233398 47365 233450 47371
rect 234178 46837 234206 53798
rect 234562 49649 234590 53798
rect 234658 53784 234912 53812
rect 235042 53784 235296 53812
rect 234658 49871 234686 53784
rect 235042 51277 235070 53784
rect 235030 51271 235082 51277
rect 235030 51213 235082 51219
rect 235618 49945 235646 53798
rect 236002 51351 236030 53798
rect 235990 51345 236042 51351
rect 235990 51287 236042 51293
rect 235606 49939 235658 49945
rect 235606 49881 235658 49887
rect 234646 49865 234698 49871
rect 234646 49807 234698 49813
rect 234550 49643 234602 49649
rect 234550 49585 234602 49591
rect 234166 46831 234218 46837
rect 234166 46773 234218 46779
rect 232822 46683 232874 46689
rect 232822 46625 232874 46631
rect 232342 46609 232394 46615
rect 232342 46551 232394 46557
rect 228022 46535 228074 46541
rect 228022 46477 228074 46483
rect 236386 46171 236414 53798
rect 236770 49575 236798 53798
rect 236866 53784 237120 53812
rect 237250 53784 237504 53812
rect 236758 49569 236810 49575
rect 236758 49511 236810 49517
rect 236866 46393 236894 53784
rect 237250 51319 237278 53784
rect 237236 51310 237292 51319
rect 237236 51245 237292 51254
rect 237826 51171 237854 53798
rect 237812 51162 237868 51171
rect 237812 51097 237868 51106
rect 238210 50875 238238 53798
rect 238196 50866 238252 50875
rect 238196 50801 238252 50810
rect 238594 47651 238622 53798
rect 238582 47645 238634 47651
rect 238582 47587 238634 47593
rect 238978 46467 239006 53798
rect 239074 53784 239328 53812
rect 239458 53784 239712 53812
rect 239074 46911 239102 53784
rect 239458 48211 239486 53784
rect 239444 48202 239500 48211
rect 239444 48137 239500 48146
rect 240034 48063 240062 53798
rect 240020 48054 240076 48063
rect 240020 47989 240076 47998
rect 240418 47873 240446 53798
rect 240802 48539 240830 53798
rect 241186 52017 241214 53798
rect 241282 53784 241536 53812
rect 241666 53784 241920 53812
rect 241174 52011 241226 52017
rect 241174 51953 241226 51959
rect 240790 48533 240842 48539
rect 240790 48475 240842 48481
rect 241282 48465 241310 53784
rect 241270 48459 241322 48465
rect 241270 48401 241322 48407
rect 241666 47915 241694 53784
rect 241846 53565 241898 53571
rect 241942 53565 241994 53571
rect 241898 53513 241942 53516
rect 241846 53507 241994 53513
rect 241858 53488 241982 53507
rect 242242 48507 242270 53798
rect 242228 48498 242284 48507
rect 242228 48433 242284 48442
rect 241652 47906 241708 47915
rect 240406 47867 240458 47873
rect 241652 47841 241708 47850
rect 240406 47809 240458 47815
rect 242626 47619 242654 53798
rect 243010 48655 243038 53798
rect 242996 48646 243052 48655
rect 242996 48581 243052 48590
rect 243394 48359 243422 53798
rect 243490 53784 243744 53812
rect 243874 53784 244128 53812
rect 282262 53787 282314 53793
rect 243490 51023 243518 53784
rect 243476 51014 243532 51023
rect 243476 50949 243532 50958
rect 243874 50833 243902 53784
rect 282262 53729 282314 53735
rect 246742 53713 246794 53719
rect 246742 53655 246794 53661
rect 282070 53713 282122 53719
rect 282274 53664 282302 53729
rect 282122 53661 282302 53664
rect 282070 53655 282302 53661
rect 345622 53713 345674 53719
rect 345622 53655 345674 53661
rect 246754 53349 246782 53655
rect 282082 53636 282302 53655
rect 289174 53491 289226 53497
rect 289174 53433 289226 53439
rect 262102 53417 262154 53423
rect 262198 53417 262250 53423
rect 262154 53365 262198 53368
rect 262102 53359 262250 53365
rect 246742 53343 246794 53349
rect 262114 53340 262238 53359
rect 246742 53285 246794 53291
rect 262390 53269 262442 53275
rect 262114 53229 262390 53257
rect 262114 53220 262142 53229
rect 261922 53192 262142 53220
rect 262390 53211 262442 53217
rect 282358 53269 282410 53275
rect 282358 53211 282410 53217
rect 283606 53269 283658 53275
rect 283606 53211 283658 53217
rect 261922 53053 261950 53192
rect 273622 53121 273674 53127
rect 273622 53063 273674 53069
rect 261910 53047 261962 53053
rect 261910 52989 261962 52995
rect 273634 52905 273662 53063
rect 282370 52979 282398 53211
rect 282358 52973 282410 52979
rect 282358 52915 282410 52921
rect 283618 52905 283646 53211
rect 273622 52899 273674 52905
rect 273622 52841 273674 52847
rect 283606 52899 283658 52905
rect 283606 52841 283658 52847
rect 289186 50907 289214 53433
rect 316918 53343 316970 53349
rect 316918 53285 316970 53291
rect 293782 53269 293834 53275
rect 316930 53220 316958 53285
rect 293782 53211 293834 53217
rect 293686 53195 293738 53201
rect 293686 53137 293738 53143
rect 293698 52979 293726 53137
rect 293794 52979 293822 53211
rect 296566 53195 296618 53201
rect 296758 53195 296810 53201
rect 296618 53155 296758 53183
rect 296566 53137 296618 53143
rect 296758 53137 296810 53143
rect 316738 53192 316958 53220
rect 328546 53201 328670 53220
rect 328534 53195 328670 53201
rect 316738 53127 316766 53192
rect 328586 53192 328670 53195
rect 328534 53137 328586 53143
rect 328642 53127 328670 53192
rect 313846 53121 313898 53127
rect 313846 53063 313898 53069
rect 316726 53121 316778 53127
rect 316726 53063 316778 53069
rect 328630 53121 328682 53127
rect 328630 53063 328682 53069
rect 313858 52979 313886 53063
rect 293686 52973 293738 52979
rect 293686 52915 293738 52921
rect 293782 52973 293834 52979
rect 293782 52915 293834 52921
rect 313846 52973 313898 52979
rect 313846 52915 313898 52921
rect 289174 50901 289226 50907
rect 289174 50843 289226 50849
rect 302422 50901 302474 50907
rect 302422 50843 302474 50849
rect 243862 50827 243914 50833
rect 243862 50769 243914 50775
rect 302434 48951 302462 50843
rect 345634 49057 345662 53655
rect 380182 53565 380234 53571
rect 380182 53507 380234 53513
rect 354260 53234 354316 53243
rect 354260 53169 354262 53178
rect 354314 53169 354316 53178
rect 354262 53137 354314 53143
rect 374326 53121 374378 53127
rect 374326 53063 374378 53069
rect 374338 52947 374366 53063
rect 374324 52938 374380 52947
rect 374324 52873 374380 52882
rect 362902 51715 362954 51721
rect 362902 51657 362954 51663
rect 348406 51641 348458 51647
rect 348502 51641 348554 51647
rect 348458 51589 348502 51592
rect 362914 51615 362942 51657
rect 348406 51583 348554 51589
rect 362900 51606 362956 51615
rect 348418 51564 348542 51583
rect 362900 51541 362956 51550
rect 345622 49051 345674 49057
rect 345622 48993 345674 48999
rect 353590 49051 353642 49057
rect 353590 48993 353642 48999
rect 302420 48942 302476 48951
rect 302420 48877 302476 48886
rect 243380 48350 243436 48359
rect 243380 48285 243436 48294
rect 242612 47610 242668 47619
rect 242612 47545 242668 47554
rect 239062 46905 239114 46911
rect 239062 46847 239114 46853
rect 238966 46461 239018 46467
rect 238966 46403 239018 46409
rect 236854 46387 236906 46393
rect 236854 46329 236906 46335
rect 236374 46165 236426 46171
rect 353602 46139 353630 48993
rect 380194 48317 380222 53507
rect 417622 53491 417674 53497
rect 417622 53433 417674 53439
rect 440566 53491 440618 53497
rect 440566 53433 440618 53439
rect 383170 53349 383294 53368
rect 383158 53343 383306 53349
rect 383210 53340 383254 53343
rect 383158 53285 383210 53291
rect 383254 53285 383306 53291
rect 417634 53275 417662 53433
rect 423284 53382 423340 53391
rect 423284 53317 423286 53326
rect 423338 53317 423340 53326
rect 423286 53285 423338 53291
rect 440578 53275 440606 53433
rect 463702 53417 463754 53423
rect 443444 53382 443500 53391
rect 463702 53359 463754 53365
rect 443444 53317 443500 53326
rect 463606 53343 463658 53349
rect 417622 53269 417674 53275
rect 417622 53211 417674 53217
rect 440566 53269 440618 53275
rect 440566 53211 440618 53217
rect 443458 53220 443486 53317
rect 463606 53285 463658 53291
rect 443458 53192 443582 53220
rect 443554 53127 443582 53192
rect 463618 53127 463646 53285
rect 443542 53121 443594 53127
rect 443542 53063 443594 53069
rect 463606 53121 463658 53127
rect 463606 53063 463658 53069
rect 434900 51754 434956 51763
rect 403222 51715 403274 51721
rect 434900 51689 434902 51698
rect 403222 51657 403274 51663
rect 434954 51689 434956 51698
rect 459284 51754 459340 51763
rect 459284 51689 459340 51698
rect 434902 51657 434954 51663
rect 403234 51615 403262 51657
rect 459298 51647 459326 51689
rect 459286 51641 459338 51647
rect 382964 51606 383020 51615
rect 403220 51606 403276 51615
rect 383020 51573 383102 51592
rect 383020 51567 383114 51573
rect 383020 51564 383062 51567
rect 382964 51541 383020 51550
rect 403220 51541 403276 51550
rect 423284 51606 423340 51615
rect 423340 51573 423422 51592
rect 459286 51583 459338 51589
rect 423340 51567 423434 51573
rect 423340 51564 423382 51567
rect 423284 51541 423340 51550
rect 383062 51509 383114 51515
rect 423382 51509 423434 51515
rect 463714 49057 463742 53359
rect 498742 53343 498794 53349
rect 498742 53285 498794 53291
rect 489622 51641 489674 51647
rect 489620 51606 489622 51615
rect 489674 51606 489676 51615
rect 489620 51541 489676 51550
rect 498754 50981 498782 53285
rect 509878 53269 509930 53275
rect 509698 53217 509878 53220
rect 509698 53211 509930 53217
rect 525910 53269 525962 53275
rect 525910 53211 525962 53217
rect 509698 53201 509918 53211
rect 509686 53195 509918 53201
rect 509738 53192 509918 53195
rect 509686 53137 509738 53143
rect 509602 51721 509726 51740
rect 509602 51715 509738 51721
rect 509602 51712 509686 51715
rect 509602 51615 509630 51712
rect 509686 51657 509738 51663
rect 520246 51715 520298 51721
rect 520246 51657 520298 51663
rect 509588 51606 509644 51615
rect 520258 51573 520286 51657
rect 509588 51541 509644 51550
rect 520246 51567 520298 51573
rect 520246 51509 520298 51515
rect 498742 50975 498794 50981
rect 498742 50917 498794 50923
rect 504022 50975 504074 50981
rect 504022 50917 504074 50923
rect 463702 49051 463754 49057
rect 463702 48993 463754 48999
rect 471382 49051 471434 49057
rect 471382 48993 471434 48999
rect 380182 48311 380234 48317
rect 380182 48253 380234 48259
rect 394582 48311 394634 48317
rect 394582 48253 394634 48259
rect 236374 46107 236426 46113
rect 353588 46130 353644 46139
rect 353588 46065 353644 46074
rect 214678 44627 214730 44633
rect 215348 44650 215404 44659
rect 215348 44585 215404 44594
rect 302516 43318 302572 43327
rect 302516 43253 302572 43262
rect 361748 43318 361804 43327
rect 361748 43253 361804 43262
rect 364916 43318 364972 43327
rect 364916 43253 364972 43262
rect 302530 42120 302558 43253
rect 310102 42391 310154 42397
rect 310102 42333 310154 42339
rect 306740 42134 306796 42143
rect 302530 42092 302688 42120
rect 306796 42092 307008 42120
rect 310114 42106 310142 42333
rect 357140 42134 357196 42143
rect 306740 42069 306796 42078
rect 357196 42092 357456 42120
rect 361762 42106 361790 43253
rect 364930 42106 364958 43253
rect 394594 43211 394622 48253
rect 408886 44833 408938 44839
rect 408886 44775 408938 44781
rect 394582 43205 394634 43211
rect 394582 43147 394634 43153
rect 405238 42169 405290 42175
rect 408898 42143 408926 44775
rect 457750 44759 457802 44765
rect 457750 44701 457802 44707
rect 410804 43318 410860 43327
rect 410804 43253 410860 43262
rect 408982 43205 409034 43211
rect 408982 43147 409034 43153
rect 408884 42134 408940 42143
rect 405290 42117 405552 42120
rect 405238 42111 405552 42117
rect 405250 42092 405552 42111
rect 357140 42069 357196 42078
rect 408884 42069 408940 42078
rect 408994 41824 409022 43147
rect 410818 41824 410846 43253
rect 416276 42134 416332 42143
rect 416332 42092 416592 42120
rect 416276 42069 416332 42078
rect 408994 41796 409296 41824
rect 410818 41796 411120 41824
rect 214294 41725 214346 41731
rect 214294 41667 214346 41673
rect 210740 40802 210796 40811
rect 210740 40737 210796 40746
rect 457762 40367 457790 44701
rect 460066 42101 460368 42120
rect 471394 42106 471422 48993
rect 504034 48687 504062 50917
rect 504022 48681 504074 48687
rect 504022 48623 504074 48629
rect 512566 48681 512618 48687
rect 512566 48623 512618 48629
rect 509782 44685 509834 44691
rect 509782 44627 509834 44633
rect 509794 43285 509822 44627
rect 509782 43279 509834 43285
rect 509782 43221 509834 43227
rect 512578 42175 512606 48623
rect 518804 44798 518860 44807
rect 518804 44733 518860 44742
rect 512566 42169 512618 42175
rect 512566 42111 512618 42117
rect 518818 42106 518846 44733
rect 521590 43205 521642 43211
rect 521590 43147 521642 43153
rect 520342 42169 520394 42175
rect 521602 42120 521630 43147
rect 525922 42120 525950 53211
rect 639682 51943 639710 233604
rect 649666 233243 649694 748811
rect 649750 702767 649802 702773
rect 649750 702709 649802 702715
rect 649762 239311 649790 702709
rect 649858 668141 649886 981763
rect 649954 846227 649982 995157
rect 650230 989517 650282 989523
rect 650230 989459 650282 989465
rect 650038 988555 650090 988561
rect 650038 988497 650090 988503
rect 650050 892847 650078 988497
rect 650134 981377 650186 981383
rect 650134 981319 650186 981325
rect 650036 892838 650092 892847
rect 650036 892773 650092 892782
rect 649940 846218 649996 846227
rect 649940 846153 649996 846162
rect 650146 809259 650174 981319
rect 650134 809253 650186 809259
rect 650134 809195 650186 809201
rect 650242 705479 650270 989459
rect 652246 983745 652298 983751
rect 652246 983687 652298 983693
rect 650902 983523 650954 983529
rect 650902 983465 650954 983471
rect 650228 705470 650284 705479
rect 650228 705405 650284 705414
rect 649846 668135 649898 668141
rect 649846 668077 649898 668083
rect 649846 656739 649898 656745
rect 649846 656681 649898 656687
rect 649750 239305 649802 239311
rect 649750 239247 649802 239253
rect 645526 233237 645578 233243
rect 645526 233179 645578 233185
rect 649654 233237 649706 233243
rect 649654 233179 649706 233185
rect 645334 233089 645386 233095
rect 645334 233031 645386 233037
rect 645142 233015 645194 233021
rect 645142 232957 645194 232963
rect 645154 231139 645182 232957
rect 645238 232941 645290 232947
rect 645238 232883 645290 232889
rect 645250 231731 645278 232883
rect 645236 231722 645292 231731
rect 645236 231657 645292 231666
rect 645140 231130 645196 231139
rect 645140 231065 645196 231074
rect 640726 79243 640778 79249
rect 640726 79185 640778 79191
rect 625750 51937 625802 51943
rect 625750 51879 625802 51885
rect 639670 51937 639722 51943
rect 639670 51879 639722 51885
rect 601940 51754 601996 51763
rect 558838 51715 558890 51721
rect 601940 51689 601942 51698
rect 558838 51657 558890 51663
rect 601994 51689 601996 51698
rect 622004 51754 622060 51763
rect 622004 51689 622060 51698
rect 601942 51657 601994 51663
rect 550006 51641 550058 51647
rect 550102 51641 550154 51647
rect 550058 51589 550102 51592
rect 550006 51583 550154 51589
rect 550018 51564 550142 51583
rect 558850 51573 558878 51657
rect 622018 51647 622046 51689
rect 625762 51647 625790 51879
rect 622006 51641 622058 51647
rect 622006 51583 622058 51589
rect 625750 51641 625802 51647
rect 625750 51583 625802 51589
rect 558838 51567 558890 51573
rect 558838 51509 558890 51515
rect 640738 49057 640766 79185
rect 625078 49051 625130 49057
rect 625078 48993 625130 48999
rect 640726 49051 640778 49057
rect 640726 48993 640778 48999
rect 529268 44650 529324 44659
rect 529268 44585 529324 44594
rect 520394 42117 520656 42120
rect 520342 42111 520656 42117
rect 460054 42095 460368 42101
rect 460106 42092 460368 42095
rect 520354 42092 520656 42111
rect 521602 42092 521856 42120
rect 525922 42092 526176 42120
rect 529282 42106 529310 44585
rect 460054 42037 460106 42043
rect 463700 41838 463756 41847
rect 465716 41838 465772 41847
rect 463756 41796 464016 41824
rect 463700 41773 463756 41782
rect 465772 41796 465936 41824
rect 514882 41805 515136 41824
rect 514870 41799 515136 41805
rect 465716 41773 465772 41782
rect 514922 41796 515136 41799
rect 514870 41741 514922 41747
rect 625090 40663 625118 48993
rect 645154 48835 645182 231065
rect 645142 48829 645194 48835
rect 645142 48771 645194 48777
rect 645250 48761 645278 231657
rect 645346 230547 645374 233031
rect 645538 232323 645566 233179
rect 649858 233169 649886 656681
rect 649942 613523 649994 613529
rect 649942 613465 649994 613471
rect 649954 239089 649982 613465
rect 650038 567421 650090 567427
rect 650038 567363 650090 567369
rect 649942 239083 649994 239089
rect 649942 239025 649994 239031
rect 645718 233163 645770 233169
rect 645718 233105 645770 233111
rect 649846 233163 649898 233169
rect 649846 233105 649898 233111
rect 645730 232767 645758 233105
rect 650050 233095 650078 567363
rect 650134 521319 650186 521325
rect 650134 521261 650186 521267
rect 650146 239607 650174 521261
rect 650230 478177 650282 478183
rect 650230 478119 650282 478125
rect 650134 239601 650186 239607
rect 650134 239543 650186 239549
rect 650242 239459 650270 478119
rect 650326 391745 650378 391751
rect 650326 391687 650378 391693
rect 650230 239453 650282 239459
rect 650230 239395 650282 239401
rect 650038 233089 650090 233095
rect 650038 233031 650090 233037
rect 650338 233021 650366 391687
rect 650422 345643 650474 345649
rect 650422 345585 650474 345591
rect 650434 239533 650462 345585
rect 650518 299615 650570 299621
rect 650518 299557 650570 299563
rect 650422 239527 650474 239533
rect 650422 239469 650474 239475
rect 650326 233015 650378 233021
rect 650326 232957 650378 232963
rect 650530 232947 650558 299557
rect 650914 240495 650942 983465
rect 652258 941941 652286 983687
rect 658006 983671 658058 983677
rect 658006 983613 658058 983619
rect 655124 974682 655180 974691
rect 655124 974617 655180 974626
rect 653782 951851 653834 951857
rect 653782 951793 653834 951799
rect 652246 941935 652298 941941
rect 652246 941877 652298 941883
rect 653794 939467 653822 951793
rect 654356 951150 654412 951159
rect 654356 951085 654412 951094
rect 654370 942089 654398 951085
rect 655138 944679 655166 974617
rect 655220 962842 655276 962851
rect 655220 962777 655276 962786
rect 655234 944901 655262 962777
rect 655222 944895 655274 944901
rect 655222 944837 655274 944843
rect 655126 944673 655178 944679
rect 655126 944615 655178 944621
rect 654358 942083 654410 942089
rect 654358 942025 654410 942031
rect 653780 939458 653836 939467
rect 653780 939393 653836 939402
rect 658018 939129 658046 983613
rect 658102 983597 658154 983603
rect 658102 983539 658154 983545
rect 658114 942237 658142 983539
rect 675094 980785 675146 980791
rect 675094 980727 675146 980733
rect 675106 960573 675134 980727
rect 675286 980711 675338 980717
rect 675286 980653 675338 980659
rect 675298 961348 675326 980653
rect 675394 966403 675422 966736
rect 675380 966394 675436 966403
rect 675380 966329 675436 966338
rect 675778 965811 675806 966070
rect 675764 965802 675820 965811
rect 675764 965737 675820 965746
rect 675778 965071 675806 965435
rect 675764 965062 675820 965071
rect 675764 964997 675820 965006
rect 675394 963295 675422 963595
rect 675380 963286 675436 963295
rect 675380 963221 675436 963230
rect 675490 962703 675518 963036
rect 675476 962694 675532 962703
rect 675476 962629 675532 962638
rect 675394 962259 675422 962399
rect 675380 962250 675436 962259
rect 675380 962185 675436 962194
rect 675778 961371 675806 961778
rect 675764 961362 675820 961371
rect 675298 961320 675422 961348
rect 675394 961200 675422 961320
rect 675764 961297 675820 961306
rect 675394 961186 675696 961200
rect 675408 961172 675710 961186
rect 675682 960779 675710 961172
rect 675668 960770 675724 960779
rect 675668 960705 675724 960714
rect 675106 960559 675504 960573
rect 675106 960545 675518 960559
rect 675490 960187 675518 960545
rect 675476 960178 675532 960187
rect 675476 960113 675532 960122
rect 675490 959035 675518 959262
rect 673942 959029 673994 959035
rect 673942 958971 673994 958977
rect 675478 959029 675530 959035
rect 675478 958971 675530 958977
rect 669526 954737 669578 954743
rect 669526 954679 669578 954685
rect 658102 942231 658154 942237
rect 658102 942173 658154 942179
rect 658006 939123 658058 939129
rect 658006 939065 658058 939071
rect 654452 927618 654508 927627
rect 654452 927553 654508 927562
rect 654466 927511 654494 927553
rect 654454 927505 654506 927511
rect 654454 927447 654506 927453
rect 666742 927505 666794 927511
rect 666742 927447 666794 927453
rect 654452 915926 654508 915935
rect 654452 915861 654454 915870
rect 654506 915861 654508 915870
rect 660982 915887 661034 915893
rect 654454 915829 654506 915835
rect 660982 915829 661034 915835
rect 654452 904234 654508 904243
rect 654452 904169 654508 904178
rect 654466 901537 654494 904169
rect 654454 901531 654506 901537
rect 654454 901473 654506 901479
rect 654452 880702 654508 880711
rect 654452 880637 654508 880646
rect 654466 878449 654494 880637
rect 654454 878443 654506 878449
rect 654454 878385 654506 878391
rect 660886 878443 660938 878449
rect 660886 878385 660938 878391
rect 654452 869010 654508 869019
rect 654452 868945 654508 868954
rect 654466 866979 654494 868945
rect 654454 866973 654506 866979
rect 654454 866915 654506 866921
rect 654452 857318 654508 857327
rect 654452 857253 654508 857262
rect 654466 855435 654494 857253
rect 654454 855429 654506 855435
rect 654454 855371 654506 855377
rect 654452 833786 654508 833795
rect 654452 833721 654508 833730
rect 654466 832421 654494 833721
rect 654454 832415 654506 832421
rect 654454 832357 654506 832363
rect 654452 822094 654508 822103
rect 654452 822029 654508 822038
rect 654466 820877 654494 822029
rect 654454 820871 654506 820877
rect 654454 820813 654506 820819
rect 654452 810402 654508 810411
rect 654452 810337 654508 810346
rect 654466 809333 654494 810337
rect 654454 809327 654506 809333
rect 654454 809269 654506 809275
rect 653782 809253 653834 809259
rect 653782 809195 653834 809201
rect 653794 798719 653822 809195
rect 653780 798710 653836 798719
rect 653780 798645 653836 798654
rect 654452 786870 654508 786879
rect 654452 786805 654508 786814
rect 654466 786319 654494 786805
rect 654454 786313 654506 786319
rect 654454 786255 654506 786261
rect 654452 775178 654508 775187
rect 654452 775113 654508 775122
rect 654466 774775 654494 775113
rect 654454 774769 654506 774775
rect 654454 774711 654506 774717
rect 654452 763338 654508 763347
rect 654452 763273 654454 763282
rect 654506 763273 654508 763282
rect 654454 763241 654506 763247
rect 654452 739954 654508 739963
rect 654452 739889 654508 739898
rect 654466 737331 654494 739889
rect 654454 737325 654506 737331
rect 654454 737267 654506 737273
rect 655220 728262 655276 728271
rect 655220 728197 655276 728206
rect 654452 716422 654508 716431
rect 654452 716357 654508 716366
rect 654466 714317 654494 716357
rect 654454 714311 654506 714317
rect 654454 714253 654506 714259
rect 654452 693038 654508 693047
rect 654452 692973 654508 692982
rect 654466 691303 654494 692973
rect 654454 691297 654506 691303
rect 654454 691239 654506 691245
rect 654452 669506 654508 669515
rect 654452 669441 654508 669450
rect 654466 668215 654494 669441
rect 654454 668209 654506 668215
rect 654454 668151 654506 668157
rect 652246 668135 652298 668141
rect 652246 668077 652298 668083
rect 652258 658563 652286 668077
rect 652244 658554 652300 658563
rect 652244 658489 652300 658498
rect 654452 646122 654508 646131
rect 654452 646057 654508 646066
rect 654466 645275 654494 646057
rect 654454 645269 654506 645275
rect 654454 645211 654506 645217
rect 654454 613449 654506 613455
rect 654454 613391 654506 613397
rect 654466 611055 654494 613391
rect 654452 611046 654508 611055
rect 654452 610981 654508 610990
rect 654452 599206 654508 599215
rect 654452 599141 654508 599150
rect 654466 599099 654494 599141
rect 654454 599093 654506 599099
rect 654454 599035 654506 599041
rect 655124 587366 655180 587375
rect 655124 587301 655180 587310
rect 654452 575674 654508 575683
rect 654452 575609 654508 575618
rect 654466 573199 654494 575609
rect 654454 573193 654506 573199
rect 654454 573135 654506 573141
rect 654454 564461 654506 564467
rect 654454 564403 654506 564409
rect 654466 564139 654494 564403
rect 654452 564130 654508 564139
rect 654452 564065 654508 564074
rect 654452 552290 654508 552299
rect 654452 552225 654508 552234
rect 654466 550185 654494 552225
rect 654454 550179 654506 550185
rect 654454 550121 654506 550127
rect 654452 540450 654508 540459
rect 654452 540385 654508 540394
rect 654466 538641 654494 540385
rect 654454 538635 654506 538641
rect 654454 538577 654506 538583
rect 654452 528758 654508 528767
rect 654452 528693 654508 528702
rect 654466 527097 654494 528693
rect 654454 527091 654506 527097
rect 654454 527033 654506 527039
rect 654070 517323 654122 517329
rect 654070 517265 654122 517271
rect 654082 517223 654110 517265
rect 654068 517214 654124 517223
rect 654068 517149 654124 517158
rect 654932 505374 654988 505383
rect 654932 505309 654988 505318
rect 654946 504083 654974 505309
rect 654934 504077 654986 504083
rect 654934 504019 654986 504025
rect 654452 481842 654508 481851
rect 654452 481777 654508 481786
rect 654466 480995 654494 481777
rect 654454 480989 654506 480995
rect 654454 480931 654506 480937
rect 654454 470629 654506 470635
rect 654454 470571 654506 470577
rect 654466 470307 654494 470571
rect 654452 470298 654508 470307
rect 654452 470233 654508 470242
rect 654452 446618 654508 446627
rect 654452 446553 654508 446562
rect 654466 446437 654494 446553
rect 654454 446431 654506 446437
rect 654454 446373 654506 446379
rect 654454 434961 654506 434967
rect 654452 434926 654454 434935
rect 654506 434926 654508 434935
rect 654452 434861 654508 434870
rect 654452 423382 654508 423391
rect 654452 423317 654454 423326
rect 654506 423317 654508 423326
rect 654454 423285 654506 423291
rect 654452 411394 654508 411403
rect 654452 411329 654508 411338
rect 654466 408993 654494 411329
rect 655138 409141 655166 587301
rect 655234 584817 655262 728197
rect 660898 721791 660926 878385
rect 660994 767523 661022 915829
rect 663958 901531 664010 901537
rect 663958 901473 664010 901479
rect 661174 855429 661226 855435
rect 661174 855371 661226 855377
rect 660982 767517 661034 767523
rect 660982 767459 661034 767465
rect 661078 763299 661130 763305
rect 661078 763241 661130 763247
rect 660982 737399 661034 737405
rect 660982 737341 661034 737347
rect 660886 721785 660938 721791
rect 660886 721727 660938 721733
rect 655412 681346 655468 681355
rect 655412 681281 655468 681290
rect 655316 634430 655372 634439
rect 655316 634365 655372 634374
rect 655222 584811 655274 584817
rect 655222 584753 655274 584759
rect 655330 495573 655358 634365
rect 655426 541527 655454 681281
rect 656372 622590 656428 622599
rect 656372 622525 656428 622534
rect 656386 622113 656414 622525
rect 656374 622107 656426 622113
rect 656374 622049 656426 622055
rect 660886 555877 660938 555883
rect 660886 555819 660938 555825
rect 655414 541521 655466 541527
rect 655414 541463 655466 541469
rect 655318 495567 655370 495573
rect 655318 495509 655370 495515
rect 655220 493534 655276 493543
rect 655220 493469 655276 493478
rect 655126 409135 655178 409141
rect 655126 409077 655178 409083
rect 654454 408987 654506 408993
rect 654454 408929 654506 408935
rect 654644 399702 654700 399711
rect 654644 399637 654700 399646
rect 654658 397523 654686 399637
rect 654646 397517 654698 397523
rect 654646 397459 654698 397465
rect 654452 388010 654508 388019
rect 654452 387945 654508 387954
rect 654466 385979 654494 387945
rect 654454 385973 654506 385979
rect 654454 385915 654506 385921
rect 654454 377241 654506 377247
rect 654454 377183 654506 377189
rect 654466 376475 654494 377183
rect 654452 376466 654508 376475
rect 654452 376401 654508 376410
rect 654452 364478 654508 364487
rect 654452 364413 654508 364422
rect 654466 363557 654494 364413
rect 654454 363551 654506 363557
rect 654454 363493 654506 363499
rect 654452 341094 654508 341103
rect 654452 341029 654508 341038
rect 654466 339877 654494 341029
rect 654454 339871 654506 339877
rect 654454 339813 654506 339819
rect 654070 329659 654122 329665
rect 654070 329601 654122 329607
rect 654082 329559 654110 329601
rect 654068 329550 654124 329559
rect 654068 329485 654124 329494
rect 655234 319749 655262 493469
rect 656372 458458 656428 458467
rect 656372 458393 656428 458402
rect 656386 457981 656414 458393
rect 656374 457975 656426 457981
rect 656374 457917 656426 457923
rect 655316 352786 655372 352795
rect 655316 352721 655372 352730
rect 655222 319743 655274 319749
rect 655222 319685 655274 319691
rect 655124 317562 655180 317571
rect 655124 317497 655180 317506
rect 654454 283039 654506 283045
rect 654454 282981 654506 282987
rect 654466 282643 654494 282981
rect 654452 282634 654508 282643
rect 654452 282569 654508 282578
rect 650902 240489 650954 240495
rect 650902 240431 650954 240437
rect 650518 232941 650570 232947
rect 650518 232883 650570 232889
rect 645716 232758 645772 232767
rect 645716 232693 645772 232702
rect 645524 232314 645580 232323
rect 645524 232249 645580 232258
rect 645332 230538 645388 230547
rect 645332 230473 645388 230482
rect 645346 48909 645374 230473
rect 645538 51869 645566 232249
rect 645622 210297 645674 210303
rect 645622 210239 645674 210245
rect 645526 51863 645578 51869
rect 645526 51805 645578 51811
rect 645634 48983 645662 210239
rect 645730 51795 645758 232693
rect 646100 211002 646156 211011
rect 646100 210937 646156 210946
rect 646114 210303 646142 210937
rect 646102 210297 646154 210303
rect 646102 210239 646154 210245
rect 647926 167229 647978 167235
rect 647926 167171 647978 167177
rect 646196 166898 646252 166907
rect 646196 166833 646252 166842
rect 645908 166454 645964 166463
rect 645908 166389 645964 166398
rect 645922 164201 645950 166389
rect 646210 164275 646238 166833
rect 647938 165871 647966 167171
rect 647924 165862 647980 165871
rect 647924 165797 647980 165806
rect 646198 164269 646250 164275
rect 646198 164211 646250 164217
rect 645910 164195 645962 164201
rect 645910 164137 645962 164143
rect 655138 138449 655166 317497
rect 655220 305870 655276 305879
rect 655220 305805 655276 305814
rect 655234 138597 655262 305805
rect 655330 184403 655358 352721
rect 655412 294178 655468 294187
rect 655412 294113 655468 294122
rect 655318 184397 655370 184403
rect 655318 184339 655370 184345
rect 655222 138591 655274 138597
rect 655222 138533 655274 138539
rect 655126 138443 655178 138449
rect 655126 138385 655178 138391
rect 655426 135637 655454 294113
rect 660898 283045 660926 555819
rect 660994 470635 661022 737341
rect 661090 630623 661118 763241
rect 661186 720903 661214 855371
rect 663766 820871 663818 820877
rect 663766 820813 663818 820819
rect 661174 720897 661226 720903
rect 661174 720839 661226 720845
rect 661270 691297 661322 691303
rect 661270 691239 661322 691245
rect 661078 630617 661130 630623
rect 661078 630559 661130 630565
rect 661174 573193 661226 573199
rect 661174 573135 661226 573141
rect 661078 538635 661130 538641
rect 661078 538577 661130 538583
rect 660982 470629 661034 470635
rect 660982 470571 661034 470577
rect 661090 364963 661118 538577
rect 661186 408475 661214 573135
rect 661282 541379 661310 691239
rect 663778 677391 663806 820813
rect 663862 780615 663914 780621
rect 663862 780557 663914 780563
rect 663766 677385 663818 677391
rect 663766 677327 663818 677333
rect 663766 602053 663818 602059
rect 663766 601995 663818 602001
rect 661270 541373 661322 541379
rect 661270 541315 661322 541321
rect 661174 408469 661226 408475
rect 661174 408411 661226 408417
rect 661174 397517 661226 397523
rect 661174 397459 661226 397465
rect 661078 364957 661130 364963
rect 661078 364899 661130 364905
rect 660982 363551 661034 363557
rect 660982 363493 661034 363499
rect 660886 283039 660938 283045
rect 660886 282981 660938 282987
rect 660994 183959 661022 363493
rect 661186 229543 661214 397459
rect 663778 329665 663806 601995
rect 663874 517329 663902 780557
rect 663970 765895 663998 901473
rect 666646 865345 666698 865351
rect 666646 865287 666698 865293
rect 664054 809327 664106 809333
rect 664054 809269 664106 809275
rect 663958 765889 664010 765895
rect 663958 765831 664010 765837
rect 663958 737325 664010 737331
rect 663958 737267 664010 737273
rect 663970 586371 663998 737267
rect 664066 675763 664094 809269
rect 664054 675757 664106 675763
rect 664054 675699 664106 675705
rect 664054 668209 664106 668215
rect 664054 668151 664106 668157
rect 663958 586365 664010 586371
rect 663958 586307 664010 586313
rect 663958 550179 664010 550185
rect 663958 550121 664010 550127
rect 663862 517323 663914 517329
rect 663862 517265 663914 517271
rect 663862 457975 663914 457981
rect 663862 457917 663914 457923
rect 663766 329659 663818 329665
rect 663766 329601 663818 329607
rect 663874 274091 663902 457917
rect 663970 363927 663998 550121
rect 664066 540491 664094 668151
rect 666658 564467 666686 865287
rect 666754 766931 666782 927447
rect 666838 832415 666890 832421
rect 666838 832357 666890 832363
rect 666742 766925 666794 766931
rect 666742 766867 666794 766873
rect 666850 676503 666878 832357
rect 666934 714311 666986 714317
rect 666934 714253 666986 714259
rect 666838 676497 666890 676503
rect 666838 676439 666890 676445
rect 666838 645269 666890 645275
rect 666838 645211 666890 645217
rect 666742 645195 666794 645201
rect 666742 645137 666794 645143
rect 666646 564461 666698 564467
rect 666646 564403 666698 564409
rect 664054 540485 664106 540491
rect 664054 540427 664106 540433
rect 666646 504077 666698 504083
rect 666646 504019 666698 504025
rect 664054 434961 664106 434967
rect 664054 434903 664106 434909
rect 663958 363921 664010 363927
rect 663958 363863 664010 363869
rect 663862 274085 663914 274091
rect 663862 274027 663914 274033
rect 664066 273351 664094 434903
rect 666658 318935 666686 504019
rect 666754 377247 666782 645137
rect 666850 497571 666878 645211
rect 666946 585483 666974 714253
rect 669538 613455 669566 954679
rect 672310 942379 672362 942385
rect 672310 942321 672362 942327
rect 669622 866973 669674 866979
rect 669622 866915 669674 866921
rect 669634 722531 669662 866915
rect 669718 786313 669770 786319
rect 669718 786255 669770 786261
rect 669622 722525 669674 722531
rect 669622 722467 669674 722473
rect 669622 686265 669674 686271
rect 669622 686207 669674 686213
rect 669526 613449 669578 613455
rect 669526 613391 669578 613397
rect 669526 599093 669578 599099
rect 669526 599035 669578 599041
rect 666934 585477 666986 585483
rect 666934 585419 666986 585425
rect 666838 497565 666890 497571
rect 666838 497507 666890 497513
rect 666838 480989 666890 480995
rect 666838 480931 666890 480937
rect 666742 377241 666794 377247
rect 666742 377183 666794 377189
rect 666742 339871 666794 339877
rect 666742 339813 666794 339819
rect 666646 318929 666698 318935
rect 666646 318871 666698 318877
rect 664054 273345 664106 273351
rect 664054 273287 664106 273293
rect 661174 229537 661226 229543
rect 661174 229479 661226 229485
rect 660982 183953 661034 183959
rect 660982 183895 661034 183901
rect 666754 182923 666782 339813
rect 666850 318343 666878 480931
rect 669538 409215 669566 599035
rect 669634 423349 669662 686207
rect 669730 631807 669758 786255
rect 672214 779357 672266 779363
rect 672214 779299 672266 779305
rect 672022 777655 672074 777661
rect 672022 777597 672074 777603
rect 669814 774769 669866 774775
rect 669814 774711 669866 774717
rect 669826 632547 669854 774711
rect 671926 719195 671978 719201
rect 671926 719137 671978 719143
rect 671938 674875 671966 719137
rect 672034 709951 672062 777597
rect 672118 733625 672170 733631
rect 672118 733567 672170 733573
rect 672022 709945 672074 709951
rect 672022 709887 672074 709893
rect 672022 688633 672074 688639
rect 672022 688575 672074 688581
rect 671926 674869 671978 674875
rect 671926 674811 671978 674817
rect 671926 648303 671978 648309
rect 671926 648245 671978 648251
rect 671638 644825 671690 644831
rect 671638 644767 671690 644773
rect 671446 642309 671498 642315
rect 671446 642251 671498 642257
rect 669814 632541 669866 632547
rect 669814 632483 669866 632489
rect 669718 631801 669770 631807
rect 669718 631743 669770 631749
rect 670966 628175 671018 628181
rect 670966 628117 671018 628123
rect 670870 627805 670922 627811
rect 670870 627747 670922 627753
rect 669718 622107 669770 622113
rect 669718 622049 669770 622055
rect 669730 496683 669758 622049
rect 670882 587555 670910 627747
rect 670870 587549 670922 587555
rect 670870 587491 670922 587497
rect 670978 583231 671006 628117
rect 670964 583222 671020 583231
rect 670964 583157 671020 583166
rect 671458 574531 671486 642251
rect 671542 599315 671594 599321
rect 671542 599257 671594 599263
rect 671446 574525 671498 574531
rect 671446 574467 671498 574473
rect 671554 529243 671582 599257
rect 671650 572015 671678 644767
rect 671734 628471 671786 628477
rect 671734 628413 671786 628419
rect 671746 584891 671774 628413
rect 671830 603903 671882 603909
rect 671830 603845 671882 603851
rect 671734 584885 671786 584891
rect 671734 584827 671786 584833
rect 671638 572009 671690 572015
rect 671638 571951 671690 571957
rect 671842 532721 671870 603845
rect 671938 575419 671966 648245
rect 672034 617895 672062 688575
rect 672130 661407 672158 733567
rect 672226 709063 672254 779299
rect 672322 765303 672350 942321
rect 673954 937247 673982 958971
rect 675394 958443 675422 958744
rect 675094 958437 675146 958443
rect 675094 958379 675146 958385
rect 675382 958437 675434 958443
rect 675382 958379 675434 958385
rect 674134 953923 674186 953929
rect 674134 953865 674186 953871
rect 674038 952073 674090 952079
rect 674038 952015 674090 952021
rect 673940 937238 673996 937247
rect 673940 937173 673996 937182
rect 674050 936359 674078 952015
rect 674146 939615 674174 953865
rect 675106 953527 675134 958379
rect 675394 957671 675422 958078
rect 675380 957662 675436 957671
rect 675380 957597 675436 957606
rect 675490 957037 675518 957412
rect 675190 957031 675242 957037
rect 675190 956973 675242 956979
rect 675478 957031 675530 957037
rect 675478 956973 675530 956979
rect 675092 953518 675148 953527
rect 675092 953453 675148 953462
rect 675202 953379 675230 956973
rect 675490 956043 675518 956228
rect 675476 956034 675532 956043
rect 675476 955969 675532 955978
rect 675394 954743 675422 955044
rect 675382 954737 675434 954743
rect 675382 954679 675434 954685
rect 675490 953929 675518 954378
rect 675478 953923 675530 953929
rect 675478 953865 675530 953871
rect 675188 953370 675244 953379
rect 675188 953305 675244 953314
rect 675490 952079 675518 952528
rect 675478 952073 675530 952079
rect 675478 952015 675530 952021
rect 674708 945378 674764 945387
rect 674708 945313 674764 945322
rect 674722 944901 674750 945313
rect 674710 944895 674762 944901
rect 674710 944837 674762 944843
rect 674708 944786 674764 944795
rect 674708 944721 674764 944730
rect 674722 944679 674750 944721
rect 674710 944673 674762 944679
rect 674710 944615 674762 944621
rect 674612 944046 674668 944055
rect 674612 943981 674668 943990
rect 674626 942089 674654 943981
rect 674804 943306 674860 943315
rect 674804 943241 674860 943250
rect 674708 942418 674764 942427
rect 674708 942353 674710 942362
rect 674762 942353 674764 942362
rect 674710 942321 674762 942327
rect 674710 942231 674762 942237
rect 674710 942173 674762 942179
rect 674722 942131 674750 942173
rect 674708 942122 674764 942131
rect 674614 942083 674666 942089
rect 674708 942057 674764 942066
rect 674614 942025 674666 942031
rect 674818 941941 674846 943241
rect 674806 941935 674858 941941
rect 674806 941877 674858 941883
rect 674708 940790 674764 940799
rect 674708 940725 674764 940734
rect 674132 939606 674188 939615
rect 674132 939541 674188 939550
rect 674722 939129 674750 940725
rect 674710 939123 674762 939129
rect 674710 939065 674762 939071
rect 674036 936350 674092 936359
rect 674036 936285 674092 936294
rect 679796 928654 679852 928663
rect 679796 928589 679852 928598
rect 679810 928071 679838 928589
rect 679796 928062 679852 928071
rect 679796 927997 679852 928006
rect 679810 927437 679838 927997
rect 679798 927431 679850 927437
rect 679798 927373 679850 927379
rect 675106 877509 675408 877537
rect 675106 876419 675134 877509
rect 675778 876419 675806 876900
rect 675092 876410 675148 876419
rect 675092 876345 675148 876354
rect 675764 876410 675820 876419
rect 675764 876345 675820 876354
rect 675092 876262 675148 876271
rect 675148 876220 675408 876248
rect 675092 876197 675148 876206
rect 675284 875818 675340 875827
rect 675284 875753 675340 875762
rect 675188 875670 675244 875679
rect 675188 875605 675244 875614
rect 674998 872153 675050 872159
rect 674998 872095 675050 872101
rect 674518 871709 674570 871715
rect 674518 871651 674570 871657
rect 674326 869045 674378 869051
rect 674326 868987 674378 868993
rect 674230 868379 674282 868385
rect 674230 868321 674282 868327
rect 673654 867861 673706 867867
rect 673654 867803 673706 867809
rect 672886 783501 672938 783507
rect 672886 783443 672938 783449
rect 672790 782243 672842 782249
rect 672790 782185 672842 782191
rect 672502 779801 672554 779807
rect 672502 779743 672554 779749
rect 672310 765297 672362 765303
rect 672310 765239 672362 765245
rect 672406 762559 672458 762565
rect 672406 762501 672458 762507
rect 672310 738139 672362 738145
rect 672310 738081 672362 738087
rect 672214 709057 672266 709063
rect 672214 708999 672266 709005
rect 672322 699887 672350 738081
rect 672418 717721 672446 762501
rect 672406 717715 672458 717721
rect 672406 717657 672458 717663
rect 672310 699881 672362 699887
rect 672310 699823 672362 699829
rect 672214 692925 672266 692931
rect 672214 692867 672266 692873
rect 672118 661401 672170 661407
rect 672118 661343 672170 661349
rect 672226 619227 672254 692867
rect 672418 671027 672446 717657
rect 672514 707435 672542 779743
rect 672598 778617 672650 778623
rect 672598 778559 672650 778565
rect 672502 707429 672554 707435
rect 672502 707371 672554 707377
rect 672610 706843 672638 778559
rect 672694 763299 672746 763305
rect 672694 763241 672746 763247
rect 672706 718503 672734 763241
rect 672802 745989 672830 782185
rect 672790 745983 672842 745989
rect 672790 745925 672842 745931
rect 672692 718494 672748 718503
rect 672692 718429 672748 718438
rect 672694 715347 672746 715353
rect 672694 715289 672746 715295
rect 672598 706837 672650 706843
rect 672598 706779 672650 706785
rect 672598 699881 672650 699887
rect 672598 699823 672650 699829
rect 672610 692709 672638 699823
rect 672598 692703 672650 692709
rect 672598 692645 672650 692651
rect 672502 674055 672554 674061
rect 672502 673997 672554 674003
rect 672406 671021 672458 671027
rect 672406 670963 672458 670969
rect 672310 644085 672362 644091
rect 672310 644027 672362 644033
rect 672214 619221 672266 619227
rect 672214 619163 672266 619169
rect 672022 617889 672074 617895
rect 672022 617831 672074 617837
rect 672214 603681 672266 603687
rect 672214 603623 672266 603629
rect 672022 599611 672074 599617
rect 672022 599553 672074 599559
rect 671926 575413 671978 575419
rect 671926 575355 671978 575361
rect 671830 532715 671882 532721
rect 671830 532657 671882 532663
rect 671542 529237 671594 529243
rect 671542 529179 671594 529185
rect 669814 527091 669866 527097
rect 669814 527033 669866 527039
rect 669718 496677 669770 496683
rect 669718 496619 669770 496625
rect 669718 446431 669770 446437
rect 669718 446373 669770 446379
rect 669622 423343 669674 423349
rect 669622 423285 669674 423291
rect 669526 409209 669578 409215
rect 669526 409151 669578 409157
rect 669622 408987 669674 408993
rect 669622 408929 669674 408935
rect 669526 385973 669578 385979
rect 669526 385915 669578 385921
rect 666838 318337 666890 318343
rect 666838 318279 666890 318285
rect 669538 227915 669566 385915
rect 669634 228951 669662 408929
rect 669730 274979 669758 446373
rect 669826 363335 669854 527033
rect 672034 526949 672062 599553
rect 672118 598427 672170 598433
rect 672118 598369 672170 598375
rect 672022 526943 672074 526949
rect 672022 526885 672074 526891
rect 672130 526801 672158 598369
rect 672226 564467 672254 603623
rect 672322 573643 672350 644027
rect 672514 630327 672542 673997
rect 672610 653785 672638 692645
rect 672706 673363 672734 715289
rect 672898 710543 672926 783443
rect 673666 751655 673694 867803
rect 674242 780515 674270 868321
rect 674338 781972 674366 868987
rect 674530 785080 674558 871651
rect 675010 864019 675038 872095
rect 675202 871715 675230 875605
rect 675190 871709 675242 871715
rect 675190 871651 675242 871657
rect 675298 871364 675326 875753
rect 675490 874051 675518 874384
rect 675476 874042 675532 874051
rect 675476 873977 675532 873986
rect 675394 873459 675422 873866
rect 675380 873450 675436 873459
rect 675380 873385 675436 873394
rect 675394 872867 675422 873200
rect 675380 872858 675436 872867
rect 675380 872793 675436 872802
rect 675490 872159 675518 872534
rect 675478 872153 675530 872159
rect 675478 872095 675530 872101
rect 675394 871715 675422 872016
rect 675382 871709 675434 871715
rect 675382 871651 675434 871657
rect 675202 871336 675408 871364
rect 675202 871216 675230 871336
rect 675106 871188 675230 871216
rect 674902 864013 674954 864019
rect 674902 863955 674954 863961
rect 674998 864013 675050 864019
rect 674998 863955 675050 863961
rect 674914 843891 674942 863955
rect 675106 862632 675134 871188
rect 675394 869907 675422 870092
rect 675380 869898 675436 869907
rect 675380 869833 675436 869842
rect 675490 869051 675518 869500
rect 675478 869045 675530 869051
rect 675478 868987 675530 868993
rect 675394 868385 675422 868875
rect 675382 868379 675434 868385
rect 675382 868321 675434 868327
rect 675394 867867 675422 868242
rect 675382 867861 675434 867867
rect 675382 867803 675434 867809
rect 675394 866947 675422 867058
rect 675380 866938 675436 866947
rect 675380 866873 675436 866882
rect 675394 865351 675422 865839
rect 675382 865345 675434 865351
rect 675382 865287 675434 865293
rect 675682 864727 675710 865208
rect 675668 864718 675724 864727
rect 675668 864653 675724 864662
rect 675490 862951 675518 863358
rect 675476 862942 675532 862951
rect 675476 862877 675532 862886
rect 675106 862604 675230 862632
rect 675202 846703 675230 862604
rect 675190 846697 675242 846703
rect 675190 846639 675242 846645
rect 675382 846697 675434 846703
rect 675382 846639 675434 846645
rect 674806 843885 674858 843891
rect 674806 843827 674858 843833
rect 674902 843885 674954 843891
rect 674902 843827 674954 843833
rect 674818 826691 674846 843827
rect 674804 826682 674860 826691
rect 675394 826649 675422 846639
rect 674804 826617 674860 826626
rect 675382 826643 675434 826649
rect 675382 826585 675434 826591
rect 675574 826643 675626 826649
rect 675574 826585 675626 826591
rect 674900 826534 674956 826543
rect 674900 826469 674956 826478
rect 674914 792017 674942 826469
rect 675586 816456 675614 826585
rect 675298 816428 675614 816456
rect 674710 792011 674762 792017
rect 674710 791953 674762 791959
rect 674902 792011 674954 792017
rect 674902 791953 674954 791959
rect 674530 785052 674654 785080
rect 674518 784981 674570 784987
rect 674518 784923 674570 784929
rect 674338 781944 674462 781972
rect 674228 780506 674284 780515
rect 674228 780441 674284 780450
rect 674230 775509 674282 775515
rect 674230 775451 674282 775457
rect 673748 764226 673804 764235
rect 673748 764161 673804 764170
rect 673652 751646 673708 751655
rect 673652 751581 673708 751590
rect 673762 720575 673790 764161
rect 674038 741617 674090 741623
rect 674038 741559 674090 741565
rect 673748 720566 673804 720575
rect 673748 720501 673804 720510
rect 673652 718494 673708 718503
rect 673652 718429 673708 718438
rect 673666 715353 673694 718429
rect 673654 715347 673706 715353
rect 673654 715289 673706 715295
rect 674050 714507 674078 741559
rect 674134 732367 674186 732373
rect 674134 732309 674186 732315
rect 674036 714498 674092 714507
rect 674036 714433 674092 714442
rect 672886 710537 672938 710543
rect 672886 710479 672938 710485
rect 674036 679570 674092 679579
rect 674036 679505 674092 679514
rect 672692 673354 672748 673363
rect 672692 673289 672748 673298
rect 672598 653779 672650 653785
rect 672598 653721 672650 653727
rect 672598 643419 672650 643425
rect 672598 643361 672650 643367
rect 672502 630321 672554 630327
rect 672502 630263 672554 630269
rect 672502 597169 672554 597175
rect 672502 597111 672554 597117
rect 672406 583627 672458 583633
rect 672406 583569 672458 583575
rect 672418 578897 672446 583569
rect 672406 578891 672458 578897
rect 672406 578833 672458 578839
rect 672310 573637 672362 573643
rect 672310 573579 672362 573585
rect 672214 564461 672266 564467
rect 672214 564403 672266 564409
rect 672214 564313 672266 564319
rect 672214 564255 672266 564261
rect 672226 541453 672254 564255
rect 672214 541447 672266 541453
rect 672214 541389 672266 541395
rect 672514 529909 672542 597111
rect 672610 571423 672638 643361
rect 672706 628181 672734 673289
rect 674050 670403 674078 679505
rect 674036 670394 674092 670403
rect 674036 670329 674092 670338
rect 674146 664483 674174 732309
rect 674242 716135 674270 775451
rect 674326 773659 674378 773665
rect 674326 773601 674378 773607
rect 674228 716126 674284 716135
rect 674228 716061 674284 716070
rect 674338 713027 674366 773601
rect 674434 772671 674462 781944
rect 674420 772662 674476 772671
rect 674420 772597 674476 772606
rect 674422 767517 674474 767523
rect 674420 767482 674422 767491
rect 674474 767482 674476 767491
rect 674420 767417 674476 767426
rect 674422 765889 674474 765895
rect 674420 765854 674422 765863
rect 674474 765854 674476 765863
rect 674420 765789 674476 765798
rect 674530 761844 674558 784923
rect 674626 782249 674654 785052
rect 674614 782243 674666 782249
rect 674614 782185 674666 782191
rect 674722 777407 674750 791953
rect 675298 784192 675326 816428
rect 675778 787915 675806 788322
rect 675764 787906 675820 787915
rect 675764 787841 675820 787850
rect 675490 787471 675518 787656
rect 675476 787462 675532 787471
rect 675476 787397 675532 787406
rect 675778 786731 675806 787035
rect 675764 786722 675820 786731
rect 675764 786657 675820 786666
rect 675394 784987 675422 785214
rect 675382 784981 675434 784987
rect 675382 784923 675434 784929
rect 675778 784215 675806 784622
rect 675106 784164 675326 784192
rect 675764 784206 675820 784215
rect 674998 782909 675050 782915
rect 674998 782851 675050 782857
rect 674902 780467 674954 780473
rect 674902 780409 674954 780415
rect 674708 777398 674764 777407
rect 674708 777333 674764 777342
rect 674710 766925 674762 766931
rect 674708 766890 674710 766899
rect 674762 766890 674764 766899
rect 674708 766825 674764 766834
rect 674710 765297 674762 765303
rect 674708 765262 674710 765271
rect 674762 765262 674764 765271
rect 674708 765197 674764 765206
rect 674708 763338 674764 763347
rect 674708 763273 674710 763282
rect 674762 763273 674764 763282
rect 674710 763241 674762 763247
rect 674708 762598 674764 762607
rect 674708 762533 674710 762542
rect 674762 762533 674764 762542
rect 674710 762501 674762 762507
rect 674434 761816 674558 761844
rect 674434 741623 674462 761816
rect 674914 751780 674942 780409
rect 675010 777555 675038 782851
rect 675106 782120 675134 784164
rect 675764 784141 675820 784150
rect 675298 783985 675408 784013
rect 675298 783507 675326 783985
rect 675286 783501 675338 783507
rect 675286 783443 675338 783449
rect 675298 783350 675408 783378
rect 675298 782915 675326 783350
rect 675286 782909 675338 782915
rect 675286 782851 675338 782857
rect 675298 782789 675408 782817
rect 675298 782249 675326 782789
rect 675286 782243 675338 782249
rect 675286 782185 675338 782191
rect 675408 782180 675792 782194
rect 675394 782166 675806 782180
rect 675394 782120 675422 782166
rect 675106 782092 675422 782120
rect 675778 781995 675806 782166
rect 675764 781986 675820 781995
rect 675764 781921 675820 781930
rect 675094 780615 675146 780621
rect 675094 780557 675146 780563
rect 674996 777546 675052 777555
rect 674996 777481 675052 777490
rect 675106 777069 675134 780557
rect 675490 780473 675518 780848
rect 675478 780467 675530 780473
rect 675478 780409 675530 780415
rect 675394 779807 675422 780330
rect 675382 779801 675434 779807
rect 675382 779743 675434 779749
rect 675490 779363 675518 779664
rect 675478 779357 675530 779363
rect 675478 779299 675530 779305
rect 675394 778623 675422 779031
rect 675382 778617 675434 778623
rect 675382 778559 675434 778565
rect 675490 777661 675518 777814
rect 675478 777655 675530 777661
rect 675478 777597 675530 777603
rect 675094 777063 675146 777069
rect 675094 777005 675146 777011
rect 675382 777063 675434 777069
rect 675382 777005 675434 777011
rect 675394 776630 675422 777005
rect 675394 775515 675422 775995
rect 675382 775509 675434 775515
rect 675382 775451 675434 775457
rect 675394 773665 675422 774155
rect 675382 773659 675434 773665
rect 675382 773601 675434 773607
rect 674722 751752 674942 751780
rect 674722 745915 674750 751752
rect 679700 750166 679756 750175
rect 679700 750101 679756 750110
rect 679714 749583 679742 750101
rect 679700 749574 679756 749583
rect 679700 749509 679756 749518
rect 679714 748875 679742 749509
rect 679702 748869 679754 748875
rect 679702 748811 679754 748817
rect 674998 745983 675050 745989
rect 674998 745925 675050 745931
rect 674710 745909 674762 745915
rect 674710 745851 674762 745857
rect 674902 745909 674954 745915
rect 674902 745851 674954 745857
rect 674422 741617 674474 741623
rect 674422 741559 674474 741565
rect 674914 738071 674942 745851
rect 675010 738145 675038 745925
rect 675092 743358 675148 743367
rect 675148 743316 675408 743344
rect 675092 743293 675148 743302
rect 675298 742724 675422 742752
rect 675298 742678 675326 742724
rect 675106 742650 675326 742678
rect 675394 742664 675422 742724
rect 675106 742183 675134 742650
rect 675092 742174 675148 742183
rect 675092 742109 675148 742118
rect 675106 742021 675408 742049
rect 675106 740259 675134 742021
rect 675092 740250 675148 740259
rect 675092 740185 675148 740194
rect 675394 740111 675422 740222
rect 675380 740102 675436 740111
rect 675380 740037 675436 740046
rect 675490 739223 675518 739630
rect 675476 739214 675532 739223
rect 675476 739149 675532 739158
rect 675778 738779 675806 738999
rect 675764 738770 675820 738779
rect 675764 738705 675820 738714
rect 674998 738139 675050 738145
rect 674998 738081 675050 738087
rect 674902 738065 674954 738071
rect 674902 738007 674954 738013
rect 674998 737991 675050 737997
rect 674998 737933 675050 737939
rect 674902 737917 674954 737923
rect 674902 737859 674954 737865
rect 674518 735697 674570 735703
rect 674518 735639 674570 735645
rect 674422 722525 674474 722531
rect 674420 722490 674422 722499
rect 674474 722490 674476 722499
rect 674420 722425 674476 722434
rect 674422 721785 674474 721791
rect 674420 721750 674422 721759
rect 674474 721750 674476 721759
rect 674420 721685 674476 721694
rect 674422 720897 674474 720903
rect 674420 720862 674422 720871
rect 674474 720862 674476 720871
rect 674420 720797 674476 720806
rect 674420 719234 674476 719243
rect 674420 719169 674422 719178
rect 674474 719169 674476 719178
rect 674422 719137 674474 719143
rect 674420 717754 674476 717763
rect 674420 717689 674422 717698
rect 674474 717689 674476 717698
rect 674422 717657 674474 717663
rect 674324 713018 674380 713027
rect 674324 712953 674380 712962
rect 674422 710537 674474 710543
rect 674420 710502 674422 710511
rect 674474 710502 674476 710511
rect 674420 710437 674476 710446
rect 674422 709057 674474 709063
rect 674420 709022 674422 709031
rect 674474 709022 674476 709031
rect 674420 708957 674476 708966
rect 674422 707429 674474 707435
rect 674420 707394 674422 707403
rect 674474 707394 674476 707403
rect 674420 707329 674476 707338
rect 674326 690705 674378 690711
rect 674326 690647 674378 690653
rect 674230 687375 674282 687381
rect 674230 687317 674282 687323
rect 674132 664474 674188 664483
rect 674132 664409 674188 664418
rect 672886 648081 672938 648087
rect 672886 648023 672938 648029
rect 672694 628175 672746 628181
rect 672694 628117 672746 628123
rect 672694 601979 672746 601985
rect 672694 601921 672746 601927
rect 672598 571417 672650 571423
rect 672598 571359 672650 571365
rect 672706 532795 672734 601921
rect 672790 578891 672842 578897
rect 672790 578833 672842 578839
rect 672802 564319 672830 578833
rect 672898 573051 672926 648023
rect 674132 630730 674188 630739
rect 674132 630665 674188 630674
rect 674146 630623 674174 630665
rect 674134 630617 674186 630623
rect 674134 630559 674186 630565
rect 673846 630321 673898 630327
rect 673846 630263 673898 630269
rect 673858 629851 673886 630263
rect 673844 629842 673900 629851
rect 673844 629777 673900 629786
rect 673844 629102 673900 629111
rect 673844 629037 673900 629046
rect 673858 628477 673886 629037
rect 673846 628471 673898 628477
rect 673846 628413 673898 628419
rect 673844 628362 673900 628371
rect 673844 628297 673900 628306
rect 673858 628181 673886 628297
rect 673846 628175 673898 628181
rect 673846 628117 673898 628123
rect 674242 619491 674270 687317
rect 674338 623635 674366 690647
rect 674422 689373 674474 689379
rect 674422 689315 674474 689321
rect 674434 679727 674462 689315
rect 674420 679718 674476 679727
rect 674420 679653 674476 679662
rect 674422 677385 674474 677391
rect 674420 677350 674422 677359
rect 674474 677350 674476 677359
rect 674420 677285 674476 677294
rect 674422 676497 674474 676503
rect 674420 676462 674422 676471
rect 674474 676462 674476 676471
rect 674420 676397 674476 676406
rect 674422 675757 674474 675763
rect 674420 675722 674422 675731
rect 674474 675722 674476 675731
rect 674420 675657 674476 675666
rect 674422 674869 674474 674875
rect 674420 674834 674422 674843
rect 674474 674834 674476 674843
rect 674420 674769 674476 674778
rect 674420 674094 674476 674103
rect 674420 674029 674422 674038
rect 674474 674029 674476 674038
rect 674422 673997 674474 674003
rect 674530 668775 674558 735639
rect 674710 730517 674762 730523
rect 674710 730459 674762 730465
rect 674614 728667 674666 728673
rect 674614 728609 674666 728615
rect 674516 668766 674572 668775
rect 674516 668701 674572 668710
rect 674626 668035 674654 728609
rect 674722 671143 674750 730459
rect 674806 709945 674858 709951
rect 674804 709910 674806 709919
rect 674858 709910 674860 709919
rect 674804 709845 674860 709854
rect 674806 706837 674858 706843
rect 674804 706802 674806 706811
rect 674858 706802 674860 706811
rect 674804 706737 674860 706746
rect 674914 688311 674942 737859
rect 675010 714063 675038 737933
rect 675394 737923 675422 738372
rect 675478 738139 675530 738145
rect 675478 738081 675530 738087
rect 675382 737917 675434 737923
rect 675382 737859 675434 737865
rect 675490 737780 675518 738081
rect 675764 737734 675820 737743
rect 675764 737669 675820 737678
rect 675190 737399 675242 737405
rect 675190 737341 675242 737347
rect 675202 732077 675230 737341
rect 675778 737159 675806 737669
rect 675490 735703 675518 735856
rect 675478 735697 675530 735703
rect 675478 735639 675530 735645
rect 675778 734931 675806 735338
rect 675764 734922 675820 734931
rect 675764 734857 675820 734866
rect 675394 734191 675422 734672
rect 675380 734182 675436 734191
rect 675380 734117 675436 734126
rect 675490 733631 675518 734006
rect 675478 733625 675530 733631
rect 675478 733567 675530 733573
rect 675490 732373 675518 732822
rect 675478 732367 675530 732373
rect 675478 732309 675530 732315
rect 675190 732071 675242 732077
rect 675190 732013 675242 732019
rect 675382 732071 675434 732077
rect 675382 732013 675434 732019
rect 675394 731638 675422 732013
rect 675490 730523 675518 730972
rect 675478 730517 675530 730523
rect 675478 730459 675530 730465
rect 675490 728673 675518 729155
rect 675478 728667 675530 728673
rect 675478 728609 675530 728615
rect 674996 714054 675052 714063
rect 674996 713989 675052 713998
rect 679700 705174 679756 705183
rect 679700 705109 679756 705118
rect 679714 704591 679742 705109
rect 679700 704582 679756 704591
rect 679700 704517 679756 704526
rect 679714 702773 679742 704517
rect 679702 702767 679754 702773
rect 679702 702709 679754 702715
rect 674996 702510 675052 702519
rect 674996 702445 675052 702454
rect 674900 688302 674956 688311
rect 674900 688237 674956 688246
rect 674806 685525 674858 685531
rect 674806 685467 674858 685473
rect 674708 671134 674764 671143
rect 674708 671069 674764 671078
rect 674612 668026 674668 668035
rect 674612 667961 674668 667970
rect 674422 661401 674474 661407
rect 674420 661366 674422 661375
rect 674474 661366 674476 661375
rect 674420 661301 674476 661310
rect 674422 656147 674474 656153
rect 674422 656089 674474 656095
rect 674324 623626 674380 623635
rect 674324 623561 674380 623570
rect 674434 622747 674462 656089
rect 674518 646453 674570 646459
rect 674518 646395 674570 646401
rect 674420 622738 674476 622747
rect 674420 622673 674476 622682
rect 674228 619482 674284 619491
rect 674228 619417 674284 619426
rect 673846 619221 673898 619227
rect 673846 619163 673898 619169
rect 673858 618011 673886 619163
rect 673844 618002 673900 618011
rect 673844 617937 673900 617946
rect 673846 617889 673898 617895
rect 673846 617831 673898 617837
rect 673858 616383 673886 617831
rect 673844 616374 673900 616383
rect 673844 616309 673900 616318
rect 674530 603687 674558 646395
rect 674614 645343 674666 645349
rect 674614 645285 674666 645291
rect 674626 624925 674654 645285
rect 674710 632541 674762 632547
rect 674708 632506 674710 632515
rect 674762 632506 674764 632515
rect 674708 632441 674764 632450
rect 674710 631801 674762 631807
rect 674708 631766 674710 631775
rect 674762 631766 674764 631775
rect 674708 631701 674764 631710
rect 674818 626151 674846 685467
rect 674902 683675 674954 683681
rect 674902 683617 674954 683623
rect 674914 656153 674942 683617
rect 675010 679727 675038 702445
rect 675394 697931 675422 698338
rect 675380 697922 675436 697931
rect 675380 697857 675436 697866
rect 675490 697339 675518 697672
rect 675476 697330 675532 697339
rect 675476 697265 675532 697274
rect 675764 697182 675820 697191
rect 675764 697117 675820 697126
rect 675778 697035 675806 697117
rect 675490 694823 675518 695195
rect 675476 694814 675532 694823
rect 675476 694749 675532 694758
rect 675778 694379 675806 694638
rect 675284 694370 675340 694379
rect 675284 694305 675340 694314
rect 675764 694370 675820 694379
rect 675764 694305 675820 694314
rect 675298 692173 675326 694305
rect 675490 693491 675518 693972
rect 675476 693482 675532 693491
rect 675476 693417 675532 693426
rect 675394 692931 675422 693380
rect 675382 692925 675434 692931
rect 675382 692867 675434 692873
rect 675490 692709 675518 692788
rect 675478 692703 675530 692709
rect 675478 692645 675530 692651
rect 675298 692159 675408 692173
rect 675298 692145 675422 692159
rect 675394 692011 675422 692145
rect 675380 692002 675436 692011
rect 675380 691937 675436 691946
rect 675490 690711 675518 690864
rect 675478 690705 675530 690711
rect 675478 690647 675530 690653
rect 675394 689823 675422 690346
rect 675094 689817 675146 689823
rect 675094 689759 675146 689765
rect 675382 689817 675434 689823
rect 675382 689759 675434 689765
rect 675106 685647 675134 689759
rect 675394 689379 675422 689680
rect 675382 689373 675434 689379
rect 675382 689315 675434 689321
rect 675490 688639 675518 689014
rect 675478 688633 675530 688639
rect 675478 688575 675530 688581
rect 675490 687381 675518 687830
rect 675478 687375 675530 687381
rect 675478 687317 675530 687323
rect 675394 686271 675422 686646
rect 675382 686265 675434 686271
rect 675382 686207 675434 686213
rect 675092 685638 675148 685647
rect 675092 685573 675148 685582
rect 675490 685531 675518 685980
rect 675478 685525 675530 685531
rect 675478 685467 675530 685473
rect 675490 683681 675518 684130
rect 675478 683675 675530 683681
rect 675478 683617 675530 683623
rect 674996 679718 675052 679727
rect 674996 679653 675052 679662
rect 674996 679570 675052 679579
rect 674996 679505 675052 679514
rect 675860 679570 675916 679579
rect 675860 679505 675916 679514
rect 675010 671587 675038 679505
rect 675188 672318 675244 672327
rect 675188 672253 675244 672262
rect 674996 671578 675052 671587
rect 674996 671513 675052 671522
rect 675092 671282 675148 671291
rect 675092 671217 675148 671226
rect 675106 670699 675134 671217
rect 675202 671027 675230 672253
rect 675190 671021 675242 671027
rect 675190 670963 675242 670969
rect 675092 670690 675148 670699
rect 675092 670625 675148 670634
rect 675202 664460 675230 670963
rect 675874 670699 675902 679505
rect 675860 670690 675916 670699
rect 675860 670625 675916 670634
rect 675106 664432 675230 664460
rect 674902 656147 674954 656153
rect 674902 656089 674954 656095
rect 674998 653779 675050 653785
rect 674998 653721 675050 653727
rect 674902 649561 674954 649567
rect 674902 649503 674954 649509
rect 674914 646459 674942 649503
rect 675010 647736 675038 653721
rect 675106 647865 675134 664432
rect 679700 660034 679756 660043
rect 679700 659969 679756 659978
rect 679714 659303 679742 659969
rect 679700 659294 679756 659303
rect 679700 659229 679756 659238
rect 679714 656745 679742 659229
rect 679702 656739 679754 656745
rect 679702 656681 679754 656687
rect 675778 652643 675806 653124
rect 675764 652634 675820 652643
rect 675764 652569 675820 652578
rect 675490 652199 675518 652458
rect 675476 652190 675532 652199
rect 675476 652125 675532 652134
rect 675490 651459 675518 651835
rect 675476 651450 675532 651459
rect 675476 651385 675532 651394
rect 675188 651006 675244 651015
rect 675188 650941 675244 650950
rect 675202 649567 675230 650941
rect 675778 649683 675806 650016
rect 675764 649674 675820 649683
rect 675764 649609 675820 649618
rect 675190 649561 675242 649567
rect 675190 649503 675242 649509
rect 675298 649484 675422 649512
rect 675298 649438 675326 649484
rect 675202 649410 675326 649438
rect 675394 649424 675422 649484
rect 675202 648055 675230 649410
rect 675298 648785 675408 648813
rect 675298 648309 675326 648785
rect 675286 648303 675338 648309
rect 675286 648245 675338 648251
rect 675298 648152 675408 648180
rect 675298 648087 675326 648152
rect 675286 648081 675338 648087
rect 675188 648046 675244 648055
rect 675286 648023 675338 648029
rect 675188 647981 675244 647990
rect 675094 647859 675146 647865
rect 675094 647801 675146 647807
rect 675010 647708 675230 647736
rect 675202 647617 675230 647708
rect 675202 647589 675408 647617
rect 675094 647563 675146 647569
rect 675094 647505 675146 647511
rect 674902 646453 674954 646459
rect 674902 646395 674954 646401
rect 675106 640809 675134 647505
rect 675202 645349 675230 647589
rect 675394 646459 675422 646982
rect 675382 646453 675434 646459
rect 675382 646395 675434 646401
rect 675490 645391 675518 645650
rect 675476 645382 675532 645391
rect 675190 645343 675242 645349
rect 675476 645317 675532 645326
rect 675190 645285 675242 645291
rect 675190 645195 675242 645201
rect 675190 645137 675242 645143
rect 675202 641871 675230 645137
rect 675394 644831 675422 645132
rect 675382 644825 675434 644831
rect 675382 644767 675434 644773
rect 675490 644091 675518 644466
rect 675478 644085 675530 644091
rect 675478 644027 675530 644033
rect 675394 643425 675422 643831
rect 675382 643419 675434 643425
rect 675382 643361 675434 643367
rect 675490 642315 675518 642616
rect 675478 642309 675530 642315
rect 675478 642251 675530 642257
rect 675190 641865 675242 641871
rect 675190 641807 675242 641813
rect 675382 641865 675434 641871
rect 675382 641807 675434 641813
rect 675394 641432 675422 641807
rect 675106 640781 675230 640809
rect 675202 628075 675230 640781
rect 675778 640359 675806 640795
rect 675764 640350 675820 640359
rect 675764 640285 675820 640294
rect 675394 638583 675422 638955
rect 675380 638574 675436 638583
rect 675380 638509 675436 638518
rect 675188 628066 675244 628075
rect 675188 628001 675244 628010
rect 675202 627811 675230 628001
rect 675190 627805 675242 627811
rect 675190 627747 675242 627753
rect 674804 626142 674860 626151
rect 674804 626077 674860 626086
rect 674614 624919 674666 624925
rect 674614 624861 674666 624867
rect 674902 624919 674954 624925
rect 674902 624861 674954 624867
rect 674914 604987 674942 624861
rect 679700 615042 679756 615051
rect 679700 614977 679756 614986
rect 679714 614459 679742 614977
rect 679700 614450 679756 614459
rect 679700 614385 679756 614394
rect 679714 613529 679742 614385
rect 679702 613523 679754 613529
rect 679702 613465 679754 613471
rect 675106 608118 675408 608146
rect 675106 607799 675134 608118
rect 675092 607790 675148 607799
rect 675092 607725 675148 607734
rect 675092 607494 675148 607503
rect 675148 607452 675408 607480
rect 675092 607429 675148 607438
rect 675490 606467 675518 606835
rect 675476 606458 675532 606467
rect 675476 606393 675532 606402
rect 674900 604978 674956 604987
rect 674900 604913 674956 604922
rect 675106 604981 675408 605009
rect 675106 604839 675134 604981
rect 674708 604830 674764 604839
rect 674708 604765 674764 604774
rect 675092 604830 675148 604839
rect 675092 604765 675148 604774
rect 674518 603681 674570 603687
rect 674518 603623 674570 603629
rect 674722 602873 674750 604765
rect 675106 604418 675408 604446
rect 675106 603909 675134 604418
rect 675094 603903 675146 603909
rect 675094 603845 675146 603851
rect 675106 603785 675408 603813
rect 673750 602867 673802 602873
rect 673750 602809 673802 602815
rect 674710 602867 674762 602873
rect 674710 602809 674762 602815
rect 673174 602719 673226 602725
rect 673174 602661 673226 602667
rect 672886 573045 672938 573051
rect 672886 572987 672938 572993
rect 672790 564313 672842 564319
rect 672790 564255 672842 564261
rect 672694 532789 672746 532795
rect 672694 532731 672746 532737
rect 672502 529903 672554 529909
rect 672502 529845 672554 529851
rect 673186 527879 673214 602661
rect 673762 561655 673790 602809
rect 675106 601985 675134 603785
rect 675286 603681 675338 603687
rect 675286 603623 675338 603629
rect 675190 602053 675242 602059
rect 675190 601995 675242 602001
rect 675094 601979 675146 601985
rect 675094 601921 675146 601927
rect 675202 596879 675230 601995
rect 675298 601973 675326 603623
rect 675394 602725 675422 603174
rect 675478 602867 675530 602873
rect 675478 602809 675530 602815
rect 675382 602719 675434 602725
rect 675382 602661 675434 602667
rect 675490 602582 675518 602809
rect 675298 601945 675408 601973
rect 675778 600251 675806 600658
rect 675764 600242 675820 600251
rect 675764 600177 675820 600186
rect 675394 599617 675422 600140
rect 675382 599611 675434 599617
rect 675382 599553 675434 599559
rect 675394 599321 675422 599474
rect 675382 599315 675434 599321
rect 675382 599257 675434 599263
rect 675490 598433 675518 598808
rect 675478 598427 675530 598433
rect 675478 598369 675530 598375
rect 675490 597175 675518 597624
rect 675478 597169 675530 597175
rect 675478 597111 675530 597117
rect 675190 596873 675242 596879
rect 675190 596815 675242 596821
rect 675382 596873 675434 596879
rect 675382 596815 675434 596821
rect 675394 596440 675422 596815
rect 675778 595367 675806 595774
rect 675764 595358 675820 595367
rect 675764 595293 675820 595302
rect 675778 593443 675806 593955
rect 675764 593434 675820 593443
rect 675764 593369 675820 593378
rect 676822 587549 676874 587555
rect 676822 587491 676874 587497
rect 674708 586478 674764 586487
rect 674708 586413 674764 586422
rect 674422 586365 674474 586371
rect 674420 586330 674422 586339
rect 674474 586330 674476 586339
rect 674420 586265 674476 586274
rect 674422 585477 674474 585483
rect 674420 585442 674422 585451
rect 674474 585442 674476 585451
rect 674420 585377 674476 585386
rect 674614 584885 674666 584891
rect 674612 584850 674614 584859
rect 674666 584850 674668 584859
rect 674722 584817 674750 586413
rect 674612 584785 674668 584794
rect 674710 584811 674762 584817
rect 674710 584753 674762 584759
rect 674708 583666 674764 583675
rect 674708 583601 674710 583610
rect 674762 583601 674764 583610
rect 674710 583569 674762 583575
rect 674420 583222 674476 583231
rect 674420 583157 674476 583166
rect 674434 578939 674462 583157
rect 676834 582639 676862 587491
rect 676820 582630 676876 582639
rect 675190 582591 675242 582597
rect 676820 582565 676822 582574
rect 675190 582533 675242 582539
rect 676874 582565 676876 582574
rect 676822 582533 676874 582539
rect 674420 578930 674476 578939
rect 674420 578865 674476 578874
rect 674710 575413 674762 575419
rect 674708 575378 674710 575387
rect 674762 575378 674764 575387
rect 674708 575313 674764 575322
rect 674710 574525 674762 574531
rect 674708 574490 674710 574499
rect 674762 574490 674764 574499
rect 674708 574425 674764 574434
rect 674422 573637 674474 573643
rect 674420 573602 674422 573611
rect 674474 573602 674476 573611
rect 674420 573537 674476 573546
rect 674710 573045 674762 573051
rect 674708 573010 674710 573019
rect 674762 573010 674764 573019
rect 674708 572945 674764 572954
rect 674422 572009 674474 572015
rect 674420 571974 674422 571983
rect 674474 571974 674476 571983
rect 674420 571909 674476 571918
rect 674710 571417 674762 571423
rect 674708 571382 674710 571391
rect 674762 571382 674764 571391
rect 674708 571317 674764 571326
rect 675202 564560 675230 582533
rect 676834 582505 676862 582533
rect 679796 569754 679852 569763
rect 679796 569689 679852 569698
rect 679810 569171 679838 569689
rect 679796 569162 679852 569171
rect 679796 569097 679852 569106
rect 679810 567427 679838 569097
rect 679798 567421 679850 567427
rect 679798 567363 679850 567369
rect 674818 564532 675230 564560
rect 673750 561649 673802 561655
rect 673750 561591 673802 561597
rect 674326 559577 674378 559583
rect 674326 559519 674378 559525
rect 673942 558097 673994 558103
rect 673942 558039 673994 558045
rect 673846 541447 673898 541453
rect 673846 541389 673898 541395
rect 673858 539719 673886 541389
rect 673954 540140 673982 558039
rect 674134 553953 674186 553959
rect 674134 553895 674186 553901
rect 674146 540288 674174 553895
rect 674230 541373 674282 541379
rect 674228 541338 674230 541347
rect 674282 541338 674284 541347
rect 674228 541273 674284 541282
rect 674230 540485 674282 540491
rect 674228 540450 674230 540459
rect 674282 540450 674284 540459
rect 674228 540385 674284 540394
rect 674146 540260 674270 540288
rect 673954 540112 674174 540140
rect 673844 539710 673900 539719
rect 673844 539645 673900 539654
rect 674038 538635 674090 538641
rect 674038 538577 674090 538583
rect 673846 532789 673898 532795
rect 673846 532731 673898 532737
rect 673750 532715 673802 532721
rect 673750 532657 673802 532663
rect 673762 530987 673790 532657
rect 673748 530978 673804 530987
rect 673748 530913 673804 530922
rect 673858 530099 673886 532731
rect 673844 530090 673900 530099
rect 673844 530025 673900 530034
rect 673846 529903 673898 529909
rect 673846 529845 673898 529851
rect 673858 529359 673886 529845
rect 673844 529350 673900 529359
rect 673844 529285 673900 529294
rect 673846 529237 673898 529243
rect 673846 529179 673898 529185
rect 673858 528619 673886 529179
rect 673844 528610 673900 528619
rect 673844 528545 673900 528554
rect 673172 527870 673228 527879
rect 673172 527805 673228 527814
rect 673844 526982 673900 526991
rect 673844 526917 673846 526926
rect 673898 526917 673900 526926
rect 673846 526885 673898 526891
rect 672118 526795 672170 526801
rect 672118 526737 672170 526743
rect 673846 526795 673898 526801
rect 673846 526737 673898 526743
rect 673858 526251 673886 526737
rect 673844 526242 673900 526251
rect 673844 526177 673900 526186
rect 673942 508369 673994 508375
rect 673942 508311 673994 508317
rect 673954 486143 673982 508311
rect 673940 486134 673996 486143
rect 673940 486069 673996 486078
rect 674050 483035 674078 538577
rect 674146 508375 674174 540112
rect 674134 508369 674186 508375
rect 674134 508311 674186 508317
rect 674242 508172 674270 540260
rect 674146 508144 674270 508172
rect 674338 508153 674366 559519
rect 674518 555063 674570 555069
rect 674518 555005 674570 555011
rect 674422 551955 674474 551961
rect 674422 551897 674474 551903
rect 674326 508147 674378 508153
rect 674146 484663 674174 508144
rect 674326 508089 674378 508095
rect 674434 508024 674462 551897
rect 674530 518365 674558 555005
rect 674818 553312 674846 564532
rect 674998 564461 675050 564467
rect 674998 564403 675050 564409
rect 675010 557456 675038 564403
rect 675284 562946 675340 562955
rect 675340 562904 675408 562932
rect 675284 562881 675340 562890
rect 675298 562312 675422 562340
rect 675298 562266 675326 562312
rect 675106 562238 675326 562266
rect 675394 562252 675422 562312
rect 675106 561771 675134 562238
rect 675092 561762 675148 561771
rect 675092 561697 675148 561706
rect 675094 561649 675146 561655
rect 675094 561591 675146 561597
rect 675284 561614 675340 561623
rect 675106 557604 675134 561591
rect 675394 561600 675422 561660
rect 675340 561572 675422 561600
rect 675284 561549 675340 561558
rect 675394 559583 675422 559810
rect 675382 559577 675434 559583
rect 675382 559519 675434 559525
rect 675490 558959 675518 559218
rect 675476 558950 675532 558959
rect 675476 558885 675532 558894
rect 675394 558103 675422 558626
rect 675382 558097 675434 558103
rect 675382 558039 675434 558045
rect 675394 557775 675422 557960
rect 675380 557766 675436 557775
rect 675380 557701 675436 557710
rect 675106 557576 675422 557604
rect 675010 557428 675230 557456
rect 675202 556790 675230 557428
rect 675394 557403 675422 557576
rect 675202 556762 675326 556790
rect 675298 556716 675326 556762
rect 675394 556716 675422 556776
rect 675298 556688 675422 556716
rect 675190 555877 675242 555883
rect 675190 555819 675242 555825
rect 675094 554545 675146 554551
rect 675094 554487 675146 554493
rect 674818 553284 675038 553312
rect 674806 553213 674858 553219
rect 674806 553155 674858 553161
rect 674614 548255 674666 548261
rect 674614 548197 674666 548203
rect 674518 518359 674570 518365
rect 674518 518301 674570 518307
rect 674242 507996 674462 508024
rect 674242 485329 674270 507996
rect 674326 507925 674378 507931
rect 674326 507867 674378 507873
rect 674422 507925 674474 507931
rect 674422 507867 674474 507873
rect 674338 490139 674366 507867
rect 674324 490130 674380 490139
rect 674324 490065 674380 490074
rect 674434 489399 674462 507867
rect 674518 497565 674570 497571
rect 674516 497530 674518 497539
rect 674570 497530 674572 497539
rect 674516 497465 674572 497474
rect 674518 496677 674570 496683
rect 674516 496642 674518 496651
rect 674570 496642 674572 496651
rect 674516 496577 674572 496586
rect 674420 489390 674476 489399
rect 674420 489325 674476 489334
rect 674626 488807 674654 548197
rect 674708 541634 674764 541643
rect 674708 541569 674764 541578
rect 674722 541527 674750 541569
rect 674710 541521 674762 541527
rect 674710 541463 674762 541469
rect 674710 541373 674762 541379
rect 674710 541315 674762 541321
rect 674722 497960 674750 541315
rect 674818 498108 674846 553155
rect 675010 550227 675038 553284
rect 674996 550218 675052 550227
rect 674996 550153 675052 550162
rect 675106 538641 675134 554487
rect 675202 551665 675230 555819
rect 675490 555069 675518 555444
rect 675478 555063 675530 555069
rect 675478 555005 675530 555011
rect 675394 554551 675422 554926
rect 675382 554545 675434 554551
rect 675382 554487 675434 554493
rect 675490 553959 675518 554260
rect 675478 553953 675530 553959
rect 675478 553895 675530 553901
rect 675394 553219 675422 553631
rect 675382 553213 675434 553219
rect 675382 553155 675434 553161
rect 675490 551961 675518 552410
rect 675478 551955 675530 551961
rect 675478 551897 675530 551903
rect 675190 551659 675242 551665
rect 675190 551601 675242 551607
rect 675382 551659 675434 551665
rect 675382 551601 675434 551607
rect 675394 551226 675422 551601
rect 675490 550111 675518 550595
rect 675190 550105 675242 550111
rect 675190 550047 675242 550053
rect 675478 550105 675530 550111
rect 675478 550047 675530 550053
rect 675202 541379 675230 550047
rect 675394 548261 675422 548755
rect 675382 548255 675434 548261
rect 675382 548197 675434 548203
rect 676532 547110 676588 547119
rect 676532 547045 676588 547054
rect 675190 541373 675242 541379
rect 675190 541315 675242 541321
rect 675094 538635 675146 538641
rect 675094 538577 675146 538583
rect 676546 537943 676574 547045
rect 676628 546962 676684 546971
rect 676628 546897 676684 546906
rect 676532 537934 676588 537943
rect 676532 537869 676588 537878
rect 674902 518359 674954 518365
rect 674902 518301 674954 518307
rect 674914 507931 674942 518301
rect 674902 507925 674954 507931
rect 674902 507867 674954 507873
rect 674818 498080 674942 498108
rect 674722 497932 674846 497960
rect 674708 497826 674764 497835
rect 674708 497761 674764 497770
rect 674722 495573 674750 497761
rect 674710 495567 674762 495573
rect 674710 495509 674762 495515
rect 674818 491915 674846 497932
rect 674804 491906 674860 491915
rect 674804 491841 674860 491850
rect 674612 488798 674668 488807
rect 674612 488733 674668 488742
rect 674228 485320 674284 485329
rect 674228 485255 674284 485264
rect 674132 484654 674188 484663
rect 674132 484589 674188 484598
rect 674036 483026 674092 483035
rect 674036 482961 674092 482970
rect 674914 482443 674942 498080
rect 676546 493987 676574 537869
rect 676642 537203 676670 546897
rect 676724 538674 676780 538683
rect 676724 538609 676780 538618
rect 676628 537194 676684 537203
rect 676628 537129 676684 537138
rect 676532 493978 676588 493987
rect 676532 493913 676588 493922
rect 674900 482434 674956 482443
rect 674900 482369 674956 482378
rect 676546 412143 676574 493913
rect 676642 493099 676670 537129
rect 676738 495911 676766 538609
rect 679796 524762 679852 524771
rect 679796 524697 679852 524706
rect 679810 524179 679838 524697
rect 679796 524170 679852 524179
rect 679796 524105 679852 524114
rect 679810 521325 679838 524105
rect 679798 521319 679850 521325
rect 679798 521261 679850 521267
rect 676724 495902 676780 495911
rect 676724 495837 676780 495846
rect 676724 494570 676780 494579
rect 676724 494505 676780 494514
rect 676628 493090 676684 493099
rect 676628 493025 676684 493034
rect 676532 412134 676588 412143
rect 676532 412069 676588 412078
rect 676642 411995 676670 493025
rect 676628 411986 676684 411995
rect 676628 411921 676684 411930
rect 674708 409322 674764 409331
rect 674708 409257 674764 409266
rect 674422 409209 674474 409215
rect 674422 409151 674474 409157
rect 674434 409109 674462 409151
rect 674722 409141 674750 409257
rect 674710 409135 674762 409141
rect 674420 409100 674476 409109
rect 674710 409077 674762 409083
rect 674420 409035 674476 409044
rect 674710 408469 674762 408475
rect 674708 408434 674710 408443
rect 674762 408434 674764 408443
rect 674708 408369 674764 408378
rect 676738 407703 676766 494505
rect 679796 480806 679852 480815
rect 679796 480741 679852 480750
rect 679810 480075 679838 480741
rect 679796 480066 679852 480075
rect 679796 480001 679852 480010
rect 679810 478183 679838 480001
rect 679798 478177 679850 478183
rect 679798 478119 679850 478125
rect 676724 407694 676780 407703
rect 676724 407629 676780 407638
rect 673844 406658 673900 406667
rect 673844 406593 673900 406602
rect 669814 363329 669866 363335
rect 669814 363271 669866 363277
rect 673858 362267 673886 406593
rect 674900 404142 674956 404151
rect 674900 404077 674956 404086
rect 674036 401922 674092 401931
rect 674036 401857 674092 401866
rect 673940 397186 673996 397195
rect 673940 397121 673996 397130
rect 673954 375767 673982 397121
rect 674050 383167 674078 401857
rect 674516 397778 674572 397787
rect 674516 397713 674572 397722
rect 674420 396446 674476 396455
rect 674420 396381 674476 396390
rect 674324 394004 674380 394013
rect 674324 393939 674380 393948
rect 674038 383161 674090 383167
rect 674038 383103 674090 383109
rect 674338 376877 674366 393939
rect 674434 377617 674462 396381
rect 674530 384351 674558 397713
rect 674804 395410 674860 395419
rect 674804 395345 674860 395354
rect 674708 394522 674764 394531
rect 674708 394457 674764 394466
rect 674518 384345 674570 384351
rect 674518 384287 674570 384293
rect 674722 378209 674750 394457
rect 674818 381336 674846 395345
rect 674914 384943 674942 404077
rect 675284 402514 675340 402523
rect 675284 402449 675340 402458
rect 675188 399406 675244 399415
rect 675188 399341 675244 399350
rect 674996 398518 675052 398527
rect 674996 398453 675052 398462
rect 675010 385036 675038 398453
rect 675202 385110 675230 399341
rect 675298 385737 675326 402449
rect 679700 392598 679756 392607
rect 679700 392533 679756 392542
rect 679714 392163 679742 392533
rect 679700 392154 679756 392163
rect 679700 392089 679756 392098
rect 679714 391751 679742 392089
rect 679702 391745 679754 391751
rect 679702 391687 679754 391693
rect 675298 385709 675408 385737
rect 675202 385082 675326 385110
rect 675298 385036 675326 385082
rect 675394 385036 675422 385096
rect 675010 385008 675230 385036
rect 675298 385008 675422 385036
rect 674902 384937 674954 384943
rect 674902 384879 674954 384885
rect 675094 384345 675146 384351
rect 675094 384287 675146 384293
rect 675106 381410 675134 384287
rect 675202 382076 675230 385008
rect 675286 384937 675338 384943
rect 675286 384879 675338 384885
rect 675298 384444 675326 384879
rect 675298 384416 675408 384444
rect 675382 383161 675434 383167
rect 675382 383103 675434 383109
rect 675394 382580 675422 383103
rect 675202 382048 675326 382076
rect 675298 381928 675326 382048
rect 675394 381928 675422 382062
rect 675298 381900 675422 381928
rect 675106 381382 675408 381410
rect 674818 381308 675422 381336
rect 675394 380730 675422 381308
rect 675106 380198 675408 380226
rect 674710 378203 674762 378209
rect 674710 378145 674762 378151
rect 674422 377611 674474 377617
rect 674422 377553 674474 377559
rect 674326 376871 674378 376877
rect 674326 376813 674378 376819
rect 673942 375761 673994 375767
rect 673942 375703 673994 375709
rect 675106 374551 675134 380198
rect 675202 379532 675408 379560
rect 675092 374542 675148 374551
rect 675092 374477 675148 374486
rect 675202 371739 675230 379532
rect 675476 378834 675532 378843
rect 675476 378769 675532 378778
rect 675490 378288 675518 378769
rect 675382 378203 675434 378209
rect 675382 378145 675434 378151
rect 675394 377696 675422 378145
rect 675382 377611 675434 377617
rect 675382 377553 675434 377559
rect 675394 377075 675422 377553
rect 675478 376871 675530 376877
rect 675478 376813 675530 376819
rect 675490 376438 675518 376813
rect 675478 375761 675530 375767
rect 675478 375703 675530 375709
rect 675490 375254 675518 375703
rect 675476 373950 675532 373959
rect 675476 373885 675532 373894
rect 675490 373404 675518 373885
rect 675380 372026 675436 372035
rect 675380 371961 675436 371970
rect 675188 371730 675244 371739
rect 675188 371665 675244 371674
rect 675394 371554 675422 371961
rect 674710 364957 674762 364963
rect 674708 364922 674710 364931
rect 674762 364922 674764 364931
rect 674708 364857 674764 364866
rect 674422 363921 674474 363927
rect 674420 363886 674422 363895
rect 674474 363886 674476 363895
rect 674420 363821 674476 363830
rect 674710 363329 674762 363335
rect 674708 363294 674710 363303
rect 674762 363294 674764 363303
rect 674708 363229 674764 363238
rect 673844 362258 673900 362267
rect 673844 362193 673900 362202
rect 674036 359150 674092 359159
rect 674036 359085 674092 359094
rect 674050 339581 674078 359085
rect 677108 358114 677164 358123
rect 677108 358049 677164 358058
rect 674612 357226 674668 357235
rect 674612 357161 674668 357170
rect 674516 352490 674572 352499
rect 674516 352425 674572 352434
rect 674228 351306 674284 351315
rect 674228 351241 674284 351250
rect 674132 348790 674188 348799
rect 674132 348725 674188 348734
rect 674038 339575 674090 339581
rect 674038 339517 674090 339523
rect 674146 331589 674174 348725
rect 674242 332255 674270 351241
rect 674324 349604 674380 349613
rect 674324 349539 674380 349548
rect 674338 332773 674366 349539
rect 674530 336621 674558 352425
rect 674626 340987 674654 357161
rect 675188 356486 675244 356495
rect 675188 356421 675244 356430
rect 675092 353378 675148 353387
rect 675092 353313 675148 353322
rect 674804 350270 674860 350279
rect 674804 350205 674860 350214
rect 674614 340981 674666 340987
rect 674614 340923 674666 340929
rect 674518 336615 674570 336621
rect 674518 336557 674570 336563
rect 674818 335569 674846 350205
rect 675106 336862 675134 353313
rect 675202 337409 675230 356421
rect 676916 355746 676972 355755
rect 676916 355681 676972 355690
rect 675284 354118 675340 354127
rect 675284 354053 675340 354062
rect 675298 339896 675326 354053
rect 676820 351750 676876 351759
rect 676820 351685 676876 351694
rect 676834 344507 676862 351685
rect 676930 345395 676958 355681
rect 677012 355006 677068 355015
rect 677012 354941 677068 354950
rect 676916 345386 676972 345395
rect 676916 345321 676972 345330
rect 677026 345247 677054 354941
rect 677122 345543 677150 358049
rect 679796 347458 679852 347467
rect 679796 347393 679852 347402
rect 679810 346727 679838 347393
rect 679796 346718 679852 346727
rect 679796 346653 679852 346662
rect 679810 345649 679838 346653
rect 679798 345643 679850 345649
rect 679798 345585 679850 345591
rect 677108 345534 677164 345543
rect 677108 345469 677164 345478
rect 677012 345238 677068 345247
rect 677012 345173 677068 345182
rect 676820 344498 676876 344507
rect 676820 344433 676876 344442
rect 675478 340981 675530 340987
rect 675478 340923 675530 340929
rect 675490 340548 675518 340923
rect 675298 339868 675408 339896
rect 675382 339575 675434 339581
rect 675382 339517 675434 339523
rect 675394 339216 675422 339517
rect 675202 337381 675408 337409
rect 675106 336834 675408 336862
rect 675382 336615 675434 336621
rect 675382 336557 675434 336563
rect 675394 336182 675422 336557
rect 674818 335541 675408 335569
rect 675284 335026 675340 335035
rect 675202 334984 675284 335012
rect 674326 332767 674378 332773
rect 674326 332709 674378 332715
rect 674230 332249 674282 332255
rect 674230 332191 674282 332197
rect 674134 331583 674186 331589
rect 674134 331525 674186 331531
rect 675202 329559 675230 334984
rect 675340 334984 675408 335012
rect 675284 334961 675340 334970
rect 675298 334901 675326 334961
rect 675586 333851 675614 334332
rect 675572 333842 675628 333851
rect 675572 333777 675628 333786
rect 675764 333546 675820 333555
rect 675764 333481 675820 333490
rect 675778 333074 675806 333481
rect 675382 332767 675434 332773
rect 675382 332709 675434 332715
rect 675394 332519 675422 332709
rect 675478 332249 675530 332255
rect 675478 332191 675530 332197
rect 675490 331890 675518 332191
rect 675382 331583 675434 331589
rect 675382 331525 675434 331531
rect 675394 331224 675422 331525
rect 675764 330586 675820 330595
rect 675764 330521 675820 330530
rect 675778 330040 675806 330521
rect 675188 329550 675244 329559
rect 675188 329485 675244 329494
rect 675778 328079 675806 328190
rect 675764 328070 675820 328079
rect 675764 328005 675820 328014
rect 675764 326886 675820 326895
rect 675764 326821 675820 326830
rect 675778 326340 675806 326821
rect 674422 319743 674474 319749
rect 674420 319708 674422 319717
rect 674474 319708 674476 319717
rect 674420 319643 674476 319652
rect 674422 318929 674474 318935
rect 674420 318894 674422 318903
rect 674474 318894 674476 318903
rect 674420 318829 674476 318838
rect 674710 318337 674762 318343
rect 674708 318302 674710 318311
rect 674762 318302 674764 318311
rect 674708 318237 674764 318246
rect 673940 314158 673996 314167
rect 673940 314093 673996 314102
rect 673954 294589 673982 314093
rect 674324 312530 674380 312539
rect 674324 312465 674380 312474
rect 674228 304612 674284 304621
rect 674228 304547 674284 304556
rect 674132 303798 674188 303807
rect 674132 303733 674188 303742
rect 673942 294583 673994 294589
rect 673942 294525 673994 294531
rect 674146 286597 674174 303733
rect 674242 287781 674270 304547
rect 674338 295995 674366 312465
rect 677108 311494 677164 311503
rect 677108 311429 677164 311438
rect 676916 310754 676972 310763
rect 676916 310689 676972 310698
rect 674516 309126 674572 309135
rect 674516 309061 674572 309070
rect 674420 305426 674476 305435
rect 674420 305361 674476 305370
rect 674326 295989 674378 295995
rect 674326 295931 674378 295937
rect 674434 291111 674462 305361
rect 674530 295403 674558 309061
rect 675092 308386 675148 308395
rect 675092 308321 675148 308330
rect 674996 307498 675052 307507
rect 674996 307433 675052 307442
rect 674806 299541 674858 299547
rect 674806 299483 674858 299489
rect 674518 295397 674570 295403
rect 674518 295339 674570 295345
rect 674422 291105 674474 291111
rect 674422 291047 674474 291053
rect 674230 287775 674282 287781
rect 674230 287717 674282 287723
rect 674818 287411 674846 299483
rect 674902 299467 674954 299473
rect 674902 299409 674954 299415
rect 674914 288595 674942 299409
rect 675010 291204 675038 307433
rect 675106 291870 675134 308321
rect 676820 306018 676876 306027
rect 676820 305953 676876 305962
rect 676834 299547 676862 305953
rect 676822 299541 676874 299547
rect 676822 299483 676874 299489
rect 676930 299473 676958 310689
rect 677012 306758 677068 306767
rect 677012 306693 677068 306702
rect 677026 299515 677054 306693
rect 677012 299506 677068 299515
rect 676918 299467 676970 299473
rect 677012 299441 677068 299450
rect 676918 299409 676970 299415
rect 677122 299399 677150 311429
rect 677204 310014 677260 310023
rect 677204 309949 677260 309958
rect 675286 299393 675338 299399
rect 675286 299335 675338 299341
rect 677110 299393 677162 299399
rect 677218 299367 677246 309949
rect 679796 302466 679852 302475
rect 679796 302401 679852 302410
rect 679810 301735 679838 302401
rect 679796 301726 679852 301735
rect 679796 301661 679852 301670
rect 679810 299621 679838 301661
rect 679798 299615 679850 299621
rect 679798 299557 679850 299563
rect 677110 299335 677162 299341
rect 677204 299358 677260 299367
rect 675298 292832 675326 299335
rect 677204 299293 677260 299302
rect 675382 295989 675434 295995
rect 675382 295931 675434 295937
rect 675394 295523 675422 295931
rect 675478 295397 675530 295403
rect 675478 295339 675530 295345
rect 675490 294890 675518 295339
rect 675382 294583 675434 294589
rect 675382 294525 675434 294531
rect 675394 294224 675422 294525
rect 675298 292804 675422 292832
rect 675394 292374 675422 292804
rect 675106 291842 675408 291870
rect 675010 291176 675408 291204
rect 675094 291105 675146 291111
rect 675094 291047 675146 291053
rect 675106 290569 675134 291047
rect 675106 290541 675408 290569
rect 675284 290034 675340 290043
rect 675010 289992 675284 290020
rect 674902 288589 674954 288595
rect 674902 288531 674954 288537
rect 674806 287405 674858 287411
rect 674806 287347 674858 287353
rect 674134 286591 674186 286597
rect 674134 286533 674186 286539
rect 675010 285011 675038 289992
rect 675340 289992 675408 290020
rect 675284 289969 675340 289978
rect 675298 289909 675326 289969
rect 675476 289590 675532 289599
rect 675476 289525 675532 289534
rect 675298 289400 675422 289428
rect 675298 289354 675326 289400
rect 675106 289326 675326 289354
rect 675394 289354 675422 289400
rect 675490 289354 675518 289525
rect 675394 289340 675518 289354
rect 675408 289326 675504 289340
rect 674996 285002 675052 285011
rect 674996 284937 675052 284946
rect 675106 284863 675134 289326
rect 675478 288589 675530 288595
rect 675478 288531 675530 288537
rect 675490 288082 675518 288531
rect 675382 287775 675434 287781
rect 675382 287717 675434 287723
rect 675394 287519 675422 287717
rect 675478 287405 675530 287411
rect 675478 287347 675530 287353
rect 675490 286898 675518 287347
rect 675382 286591 675434 286597
rect 675382 286533 675434 286539
rect 675394 286232 675422 286533
rect 675668 285298 675724 285307
rect 675668 285233 675724 285242
rect 675682 285048 675710 285233
rect 674132 284854 674188 284863
rect 674132 284789 674188 284798
rect 675092 284854 675148 284863
rect 675092 284789 675148 284798
rect 674146 275391 674174 284789
rect 675380 283670 675436 283679
rect 675380 283605 675436 283614
rect 675394 283198 675422 283605
rect 675764 281894 675820 281903
rect 675764 281829 675820 281838
rect 675778 281348 675806 281829
rect 674132 275382 674188 275391
rect 674132 275317 674188 275326
rect 669718 274973 669770 274979
rect 669718 274915 669770 274921
rect 674146 274059 674174 275317
rect 674710 274973 674762 274979
rect 674708 274938 674710 274947
rect 674762 274938 674764 274947
rect 674708 274873 674764 274882
rect 674710 274085 674762 274091
rect 674132 274050 674188 274059
rect 674132 273985 674188 273994
rect 674708 274050 674710 274059
rect 674762 274050 674764 274059
rect 674708 273985 674764 273994
rect 674710 273345 674762 273351
rect 674708 273310 674710 273319
rect 674762 273310 674764 273319
rect 674708 273245 674764 273254
rect 673940 267538 673996 267547
rect 673940 267473 673996 267482
rect 673954 251003 673982 267473
rect 678260 266502 678316 266511
rect 678260 266437 678316 266446
rect 678164 265762 678220 265771
rect 678164 265697 678220 265706
rect 674612 264134 674668 264143
rect 674612 264069 674668 264078
rect 674324 263542 674380 263551
rect 674324 263477 674380 263486
rect 674132 258806 674188 258815
rect 674132 258741 674188 258750
rect 673942 250997 673994 251003
rect 673942 250939 673994 250945
rect 674146 241605 674174 258741
rect 674338 247081 674366 263477
rect 674420 262802 674476 262811
rect 674420 262737 674476 262746
rect 674326 247075 674378 247081
rect 674326 247017 674378 247023
rect 674434 247007 674462 262737
rect 674626 250411 674654 264069
rect 676916 261766 676972 261775
rect 676916 261701 676972 261710
rect 676820 261026 676876 261035
rect 676820 260961 676876 260970
rect 674708 259842 674764 259851
rect 674708 259777 674764 259786
rect 674614 250405 674666 250411
rect 674614 250347 674666 250353
rect 674422 247001 674474 247007
rect 674422 246943 674474 246949
rect 674722 246119 674750 259777
rect 675092 259398 675148 259407
rect 675092 259333 675148 259342
rect 675106 253612 675134 259333
rect 674914 253584 675134 253612
rect 674806 251663 674858 251669
rect 674806 251605 674858 251611
rect 674710 246113 674762 246119
rect 674710 246055 674762 246061
rect 674134 241599 674186 241605
rect 674134 241541 674186 241547
rect 674818 240569 674846 251605
rect 674914 242789 674942 253584
rect 675094 253513 675146 253519
rect 675094 253455 675146 253461
rect 674998 251589 675050 251595
rect 674998 251531 675050 251537
rect 674902 242783 674954 242789
rect 674902 242725 674954 242731
rect 675010 242419 675038 251531
rect 675106 247396 675134 253455
rect 676834 251595 676862 260961
rect 676930 251669 676958 261701
rect 678178 253487 678206 265697
rect 678274 253519 678302 266437
rect 678356 265022 678412 265031
rect 678356 264957 678412 264966
rect 678370 253635 678398 264957
rect 679796 257474 679852 257483
rect 679796 257409 679852 257418
rect 679810 256891 679838 257409
rect 679796 256882 679852 256891
rect 679796 256817 679852 256826
rect 679810 256405 679838 256817
rect 679798 256399 679850 256405
rect 679798 256341 679850 256347
rect 678356 253626 678412 253635
rect 678356 253561 678412 253570
rect 678262 253513 678314 253519
rect 678164 253478 678220 253487
rect 678262 253455 678314 253461
rect 678164 253413 678220 253422
rect 676918 251663 676970 251669
rect 676918 251605 676970 251611
rect 676822 251589 676874 251595
rect 676822 251531 676874 251537
rect 675382 250997 675434 251003
rect 675382 250939 675434 250945
rect 675284 250518 675340 250527
rect 675394 250523 675422 250939
rect 675284 250453 675340 250462
rect 675298 249246 675326 250453
rect 675478 250405 675530 250411
rect 675478 250347 675530 250353
rect 675490 249898 675518 250347
rect 675298 249218 675408 249246
rect 675106 247368 675408 247396
rect 675478 247075 675530 247081
rect 675478 247017 675530 247023
rect 675286 247001 675338 247007
rect 675286 246943 675338 246949
rect 675298 246212 675326 246943
rect 675490 246864 675518 247017
rect 675298 246184 675408 246212
rect 675382 246113 675434 246119
rect 675382 246055 675434 246061
rect 675394 245532 675422 246055
rect 675764 245190 675820 245199
rect 675764 245125 675820 245134
rect 675092 245042 675148 245051
rect 675778 245028 675806 245125
rect 675148 245014 675806 245028
rect 675148 245000 675792 245014
rect 675092 244977 675148 244986
rect 674998 242413 675050 242419
rect 674998 242355 675050 242361
rect 675106 241351 675134 244977
rect 675298 244334 675408 244362
rect 675188 244302 675244 244311
rect 675298 244288 675326 244334
rect 675244 244260 675326 244288
rect 675188 244237 675244 244246
rect 675092 241342 675148 241351
rect 675092 241277 675148 241286
rect 674806 240563 674858 240569
rect 674806 240505 674858 240511
rect 674612 239270 674668 239279
rect 674612 239205 674614 239214
rect 674666 239205 674668 239214
rect 674996 239270 675052 239279
rect 674996 239205 675052 239214
rect 675094 239231 675146 239237
rect 674614 239173 674666 239179
rect 675010 239163 675038 239205
rect 675094 239173 675146 239179
rect 674998 239157 675050 239163
rect 674998 239099 675050 239105
rect 675010 235241 675038 239099
rect 675106 235315 675134 239173
rect 675202 238983 675230 244237
rect 675764 243562 675820 243571
rect 675764 243497 675820 243506
rect 675778 243090 675806 243497
rect 675382 242783 675434 242789
rect 675382 242725 675434 242731
rect 675394 242498 675422 242725
rect 675382 242413 675434 242419
rect 675382 242355 675434 242361
rect 675394 241875 675422 242355
rect 675478 241599 675530 241605
rect 675478 241541 675530 241547
rect 675490 241240 675518 241541
rect 675478 240563 675530 240569
rect 675478 240505 675530 240511
rect 675490 240056 675518 240505
rect 675188 238974 675244 238983
rect 675188 238909 675244 238918
rect 675476 238678 675532 238687
rect 675476 238613 675532 238622
rect 675490 238206 675518 238613
rect 675764 236902 675820 236911
rect 675764 236837 675820 236846
rect 675778 236356 675806 236837
rect 675094 235309 675146 235315
rect 675094 235251 675146 235257
rect 679798 235309 679850 235315
rect 679798 235251 679850 235257
rect 674998 235235 675050 235241
rect 674998 235177 675050 235183
rect 674422 229537 674474 229543
rect 674420 229502 674422 229511
rect 674474 229502 674476 229511
rect 674420 229437 674476 229446
rect 669622 228945 669674 228951
rect 674710 228945 674762 228951
rect 669622 228887 669674 228893
rect 674708 228910 674710 228919
rect 674762 228910 674764 228919
rect 674708 228845 674764 228854
rect 669526 227909 669578 227915
rect 674422 227909 674474 227915
rect 669526 227851 669578 227857
rect 674420 227874 674422 227883
rect 674474 227874 674476 227883
rect 674420 227809 674476 227818
rect 679810 225811 679838 235251
rect 679990 235235 680042 235241
rect 679990 235177 680042 235183
rect 679796 225802 679852 225811
rect 679796 225737 679852 225746
rect 677204 223730 677260 223739
rect 677204 223665 677260 223674
rect 674420 222250 674476 222259
rect 674420 222185 674476 222194
rect 674324 217514 674380 217523
rect 674324 217449 674380 217458
rect 674338 201349 674366 217449
rect 674434 205789 674462 222185
rect 674996 221214 675052 221223
rect 674996 221149 675052 221158
rect 674900 214998 674956 215007
rect 674900 214933 674956 214942
rect 674804 214258 674860 214267
rect 674804 214193 674860 214202
rect 674708 213370 674764 213379
rect 674708 213305 674764 213314
rect 674614 210223 674666 210229
rect 674614 210165 674666 210171
rect 674422 205783 674474 205789
rect 674422 205725 674474 205731
rect 674326 201343 674378 201349
rect 674326 201285 674378 201291
rect 674626 197057 674654 210165
rect 674614 197051 674666 197057
rect 674614 196993 674666 196999
rect 674722 196613 674750 213305
rect 674818 197649 674846 214193
rect 674914 200369 674942 214933
rect 675010 204772 675038 221149
rect 677012 220622 677068 220631
rect 677012 220557 677068 220566
rect 675188 218550 675244 218559
rect 675188 218485 675244 218494
rect 675092 218106 675148 218115
rect 675092 218041 675148 218050
rect 675106 204901 675134 218041
rect 675202 205197 675230 218485
rect 675284 217810 675340 217819
rect 675284 217745 675340 217754
rect 675298 211751 675326 217745
rect 676916 216478 676972 216487
rect 676916 216413 676972 216422
rect 676820 215886 676876 215895
rect 676820 215821 676876 215830
rect 675284 211742 675340 211751
rect 675284 211677 675340 211686
rect 676834 210229 676862 215821
rect 676930 210271 676958 216413
rect 676916 210262 676972 210271
rect 676822 210223 676874 210229
rect 676916 210197 676972 210206
rect 676822 210165 676874 210171
rect 677026 210123 677054 220557
rect 677108 219734 677164 219743
rect 677108 219669 677164 219678
rect 677012 210114 677068 210123
rect 677012 210049 677068 210058
rect 677122 209975 677150 219669
rect 677108 209966 677164 209975
rect 677108 209901 677164 209910
rect 677218 209827 677246 223665
rect 679700 212186 679756 212195
rect 679700 212121 679756 212130
rect 679714 211455 679742 212121
rect 679700 211446 679756 211455
rect 679700 211381 679756 211390
rect 679714 210303 679742 211381
rect 679702 210297 679754 210303
rect 679702 210239 679754 210245
rect 677204 209818 677260 209827
rect 677204 209753 677260 209762
rect 679810 209679 679838 225737
rect 680002 224923 680030 235177
rect 679988 224914 680044 224923
rect 679988 224849 680044 224858
rect 679796 209670 679852 209679
rect 679796 209605 679852 209614
rect 680002 209531 680030 224849
rect 679988 209522 680044 209531
rect 679988 209457 680044 209466
rect 675478 205783 675530 205789
rect 675478 205725 675530 205731
rect 675490 205350 675518 205725
rect 675190 205191 675242 205197
rect 675190 205133 675242 205139
rect 675478 205191 675530 205197
rect 675478 205133 675530 205139
rect 675094 204895 675146 204901
rect 675094 204837 675146 204843
rect 675010 204744 675134 204772
rect 675106 204698 675134 204744
rect 674998 204673 675050 204679
rect 675106 204670 675230 204698
rect 675490 204684 675518 205133
rect 674998 204615 675050 204621
rect 675010 201664 675038 204615
rect 675202 202182 675230 204670
rect 675764 204342 675820 204351
rect 675764 204277 675820 204286
rect 675778 204018 675806 204277
rect 675298 202228 675422 202256
rect 675298 202182 675326 202228
rect 675202 202154 675326 202182
rect 675394 202168 675422 202228
rect 675010 201636 675408 201664
rect 675382 201343 675434 201349
rect 675382 201285 675434 201291
rect 675394 200984 675422 201285
rect 674914 200341 675408 200369
rect 675202 199786 675408 199814
rect 675092 199754 675148 199763
rect 675202 199740 675230 199786
rect 675148 199712 675230 199740
rect 675092 199689 675148 199698
rect 674806 197643 674858 197649
rect 674806 197585 674858 197591
rect 674710 196607 674762 196613
rect 674710 196549 674762 196555
rect 675106 195619 675134 199689
rect 675298 199268 675422 199296
rect 675188 199162 675244 199171
rect 675298 199148 675326 199268
rect 675244 199120 675326 199148
rect 675394 199134 675422 199268
rect 675188 199097 675244 199106
rect 675202 195767 675230 199097
rect 675476 198422 675532 198431
rect 675476 198357 675532 198366
rect 675490 197876 675518 198357
rect 675382 197643 675434 197649
rect 675382 197585 675434 197591
rect 675394 197319 675422 197585
rect 675478 197051 675530 197057
rect 675478 196993 675530 196999
rect 675490 196692 675518 196993
rect 675382 196607 675434 196613
rect 675382 196549 675434 196555
rect 675394 196026 675422 196549
rect 675188 195758 675244 195767
rect 675188 195693 675244 195702
rect 675092 195610 675148 195619
rect 675092 195545 675148 195554
rect 675764 195314 675820 195323
rect 675764 195249 675820 195258
rect 675778 194842 675806 195249
rect 675380 193538 675436 193547
rect 675380 193473 675436 193482
rect 675394 192992 675422 193473
rect 675764 191614 675820 191623
rect 675764 191549 675820 191558
rect 675778 191142 675806 191549
rect 674420 184510 674476 184519
rect 674420 184445 674476 184454
rect 674434 184403 674462 184445
rect 674422 184397 674474 184403
rect 674422 184339 674474 184345
rect 674710 183953 674762 183959
rect 674708 183918 674710 183927
rect 674762 183918 674764 183927
rect 674708 183853 674764 183862
rect 666742 182917 666794 182923
rect 674422 182917 674474 182923
rect 666742 182859 666794 182865
rect 674420 182882 674422 182891
rect 674474 182882 674476 182891
rect 674420 182817 674476 182826
rect 679700 179922 679756 179931
rect 679700 179857 679756 179866
rect 674036 178886 674092 178895
rect 674036 178821 674092 178830
rect 674050 159465 674078 178821
rect 674420 177258 674476 177267
rect 674420 177193 674476 177202
rect 674324 169414 674380 169423
rect 674324 169349 674380 169358
rect 674038 159459 674090 159465
rect 674038 159401 674090 159407
rect 674338 152657 674366 169349
rect 674434 160797 674462 177193
rect 677012 176222 677068 176231
rect 677012 176157 677068 176166
rect 676916 175630 676972 175639
rect 676916 175565 676972 175574
rect 675188 174002 675244 174011
rect 675188 173937 675244 173946
rect 674900 173114 674956 173123
rect 674900 173049 674956 173058
rect 674516 168378 674572 168387
rect 674516 168313 674572 168322
rect 674422 160791 674474 160797
rect 674422 160733 674474 160739
rect 674326 152651 674378 152657
rect 674326 152593 674378 152599
rect 674530 151473 674558 168313
rect 674708 167342 674764 167351
rect 674708 167277 674764 167286
rect 674722 167235 674750 167277
rect 674710 167229 674762 167235
rect 674710 167171 674762 167177
rect 674612 166602 674668 166611
rect 674612 166537 674668 166546
rect 674626 164275 674654 166537
rect 674708 165714 674764 165723
rect 674708 165649 674764 165658
rect 674614 164269 674666 164275
rect 674614 164211 674666 164217
rect 674722 164201 674750 165649
rect 674710 164195 674762 164201
rect 674710 164137 674762 164143
rect 674806 163307 674858 163313
rect 674806 163249 674858 163255
rect 674818 152213 674846 163249
rect 674914 156949 674942 173049
rect 674996 172374 675052 172383
rect 674996 172309 675052 172318
rect 675010 157097 675038 172309
rect 675092 170006 675148 170015
rect 675092 169941 675148 169950
rect 674998 157091 675050 157097
rect 674998 157033 675050 157039
rect 674902 156943 674954 156949
rect 674902 156885 674954 156891
rect 675106 156080 675134 169941
rect 675202 160057 675230 173937
rect 676820 170894 676876 170903
rect 676820 170829 676876 170838
rect 675284 166454 675340 166463
rect 675284 166389 675340 166398
rect 675298 165575 675326 166389
rect 675284 165566 675340 165575
rect 675284 165501 675340 165510
rect 675286 164121 675338 164127
rect 675286 164063 675338 164069
rect 675190 160051 675242 160057
rect 675190 159993 675242 159999
rect 675298 159780 675326 164063
rect 676834 163313 676862 170829
rect 676930 164095 676958 175565
rect 677026 164127 677054 176157
rect 677204 174742 677260 174751
rect 677204 174677 677260 174686
rect 677108 171486 677164 171495
rect 677108 171421 677164 171430
rect 677014 164121 677066 164127
rect 676916 164086 676972 164095
rect 677014 164063 677066 164069
rect 676916 164021 676972 164030
rect 677122 163651 677150 171421
rect 677218 163947 677246 174677
rect 679714 166611 679742 179857
rect 679796 179478 679852 179487
rect 679796 179413 679852 179422
rect 679700 166602 679756 166611
rect 679700 166537 679756 166546
rect 679810 166463 679838 179413
rect 679796 166454 679852 166463
rect 679796 166389 679852 166398
rect 677204 163938 677260 163947
rect 677204 163873 677260 163882
rect 677108 163642 677164 163651
rect 677108 163577 677164 163586
rect 676822 163307 676874 163313
rect 676822 163249 676874 163255
rect 675382 160791 675434 160797
rect 675382 160733 675434 160739
rect 675394 160323 675422 160733
rect 675478 160051 675530 160057
rect 675478 159993 675530 159999
rect 675202 159752 675326 159780
rect 675202 157190 675230 159752
rect 675490 159692 675518 159993
rect 675382 159459 675434 159465
rect 675382 159401 675434 159407
rect 675394 159026 675422 159401
rect 675202 157162 675326 157190
rect 675298 157116 675326 157162
rect 675490 157116 675518 157176
rect 675190 157091 675242 157097
rect 675298 157088 675518 157116
rect 675190 157033 675242 157039
rect 675010 156052 675134 156080
rect 675010 155369 675038 156052
rect 675202 156006 675230 157033
rect 675478 156943 675530 156949
rect 675478 156885 675530 156891
rect 675490 156658 675518 156885
rect 675202 155978 675408 156006
rect 675010 155341 675408 155369
rect 675490 154623 675518 154808
rect 675476 154614 675532 154623
rect 675476 154549 675532 154558
rect 675380 154318 675436 154327
rect 675380 154253 675436 154262
rect 675394 154142 675422 154253
rect 675764 153430 675820 153439
rect 675764 153365 675820 153374
rect 675778 152884 675806 153365
rect 675382 152651 675434 152657
rect 675382 152593 675434 152599
rect 675394 152292 675422 152593
rect 674806 152207 674858 152213
rect 674806 152149 674858 152155
rect 675478 152207 675530 152213
rect 675478 152149 675530 152155
rect 675490 151700 675518 152149
rect 674518 151467 674570 151473
rect 674518 151409 674570 151415
rect 675382 151467 675434 151473
rect 675382 151409 675434 151415
rect 675394 151034 675422 151409
rect 675764 150322 675820 150331
rect 675764 150257 675820 150266
rect 675778 149850 675806 150257
rect 675476 148546 675532 148555
rect 675476 148481 675532 148490
rect 675490 148000 675518 148481
rect 675764 146622 675820 146631
rect 675764 146557 675820 146566
rect 675778 146150 675806 146557
rect 674708 139074 674764 139083
rect 674708 139009 674764 139018
rect 674722 138597 674750 139009
rect 674710 138591 674762 138597
rect 674710 138533 674762 138539
rect 674420 138482 674476 138491
rect 674420 138417 674422 138426
rect 674474 138417 674476 138426
rect 674422 138385 674474 138391
rect 674612 137298 674668 137307
rect 674612 137233 674668 137242
rect 674626 135637 674654 137233
rect 674708 135670 674764 135679
rect 655414 135631 655466 135637
rect 655414 135573 655466 135579
rect 674614 135631 674666 135637
rect 674708 135605 674764 135614
rect 674614 135573 674666 135579
rect 674722 135415 674750 135605
rect 646486 135409 646538 135415
rect 646486 135351 646538 135357
rect 674710 135409 674762 135415
rect 674710 135351 674762 135357
rect 646498 120139 646526 135351
rect 673364 134930 673420 134939
rect 673420 134888 673486 134916
rect 673364 134865 673420 134874
rect 674420 133746 674476 133755
rect 674420 133681 674476 133690
rect 674132 131230 674188 131239
rect 674132 131165 674188 131174
rect 674036 123386 674092 123395
rect 674036 123321 674092 123330
rect 647828 121758 647884 121767
rect 647828 121693 647884 121702
rect 647842 121281 647870 121693
rect 647830 121275 647882 121281
rect 647830 121217 647882 121223
rect 647926 121201 647978 121207
rect 647924 121166 647926 121175
rect 647978 121166 647980 121175
rect 647830 121127 647882 121133
rect 647924 121101 647980 121110
rect 647830 121069 647882 121075
rect 647842 120731 647870 121069
rect 647828 120722 647884 120731
rect 647828 120657 647884 120666
rect 646484 120130 646540 120139
rect 646484 120065 646540 120074
rect 674050 119228 674078 123321
rect 673954 119200 674078 119228
rect 647926 112913 647978 112919
rect 665206 112913 665258 112919
rect 647926 112855 647978 112861
rect 665204 112878 665206 112887
rect 665258 112878 665260 112887
rect 647938 104451 647966 112855
rect 665204 112813 665260 112822
rect 665204 111546 665260 111555
rect 665204 111481 665260 111490
rect 647924 104442 647980 104451
rect 647924 104377 647980 104386
rect 665218 96491 665246 111481
rect 673954 106185 673982 119200
rect 674146 119080 674174 131165
rect 674228 128122 674284 128131
rect 674228 128057 674284 128066
rect 674050 119052 674174 119080
rect 674050 113659 674078 119052
rect 674134 118981 674186 118987
rect 674134 118923 674186 118929
rect 674146 114177 674174 118923
rect 674134 114171 674186 114177
rect 674134 114113 674186 114119
rect 674038 113653 674090 113659
rect 674038 113595 674090 113601
rect 674242 113363 674270 128057
rect 674324 127382 674380 127391
rect 674324 127317 674380 127326
rect 674230 113357 674282 113363
rect 674230 113299 674282 113305
rect 674338 111217 674366 127317
rect 674434 118987 674462 133681
rect 675092 131822 675148 131831
rect 675092 131757 675148 131766
rect 674900 124866 674956 124875
rect 674900 124801 674956 124810
rect 674516 123978 674572 123987
rect 674516 123913 674572 123922
rect 674422 118981 674474 118987
rect 674422 118923 674474 118929
rect 674422 118019 674474 118025
rect 674422 117961 674474 117967
rect 674326 111211 674378 111217
rect 674326 111153 674378 111159
rect 673942 106179 673994 106185
rect 673942 106121 673994 106127
rect 674434 105223 674462 117961
rect 674530 107369 674558 123913
rect 674804 122202 674860 122211
rect 674804 122137 674860 122146
rect 674612 121610 674668 121619
rect 674612 121545 674668 121554
rect 674626 121133 674654 121545
rect 674708 121314 674764 121323
rect 674708 121249 674710 121258
rect 674762 121249 674764 121258
rect 674710 121217 674762 121223
rect 674818 121207 674846 122137
rect 674806 121201 674858 121207
rect 674806 121143 674858 121149
rect 674614 121127 674666 121133
rect 674614 121069 674666 121075
rect 674914 120116 674942 124801
rect 674722 120088 674942 120116
rect 674614 118093 674666 118099
rect 674614 118035 674666 118041
rect 674518 107363 674570 107369
rect 674518 107305 674570 107311
rect 674626 106999 674654 118035
rect 674722 110169 674750 120088
rect 674806 120017 674858 120023
rect 674806 119959 674858 119965
rect 674818 114492 674846 119959
rect 675106 115158 675134 131757
rect 677012 130342 677068 130351
rect 677012 130277 677068 130286
rect 675188 128714 675244 128723
rect 675188 128649 675244 128658
rect 675202 120023 675230 128649
rect 676916 126346 676972 126355
rect 676916 126281 676972 126290
rect 676820 125606 676876 125615
rect 676820 125541 676876 125550
rect 675190 120017 675242 120023
rect 675190 119959 675242 119965
rect 676834 118099 676862 125541
rect 676822 118093 676874 118099
rect 676822 118035 676874 118041
rect 676930 118025 676958 126281
rect 677026 120435 677054 130277
rect 677108 129602 677164 129611
rect 677108 129537 677164 129546
rect 677012 120426 677068 120435
rect 677012 120361 677068 120370
rect 677122 118067 677150 129537
rect 677108 118058 677164 118067
rect 676918 118019 676970 118025
rect 677108 117993 677164 118002
rect 676918 117961 676970 117967
rect 675106 115130 675326 115158
rect 675298 115084 675326 115130
rect 675394 115084 675422 115144
rect 675298 115056 675422 115084
rect 674818 114464 675408 114492
rect 675382 114171 675434 114177
rect 675382 114113 675434 114119
rect 675394 113812 675422 114113
rect 675190 113653 675242 113659
rect 675190 113595 675242 113601
rect 675094 113357 675146 113363
rect 675094 113299 675146 113305
rect 675106 111458 675134 113299
rect 675202 112009 675230 113595
rect 675202 111981 675408 112009
rect 675106 111430 675408 111458
rect 675382 111211 675434 111217
rect 675382 111153 675434 111159
rect 675394 110778 675422 111153
rect 674722 110141 675408 110169
rect 675476 110066 675532 110075
rect 675476 110001 675532 110010
rect 675490 109594 675518 110001
rect 675380 109474 675436 109483
rect 675380 109409 675436 109418
rect 675394 108959 675422 109409
rect 675668 108142 675724 108151
rect 675668 108077 675724 108086
rect 675682 107670 675710 108077
rect 675382 107363 675434 107369
rect 675382 107305 675434 107311
rect 675394 107119 675422 107305
rect 674614 106993 674666 106999
rect 674614 106935 674666 106941
rect 675478 106993 675530 106999
rect 675478 106935 675530 106941
rect 675490 106486 675518 106935
rect 675382 106179 675434 106185
rect 675382 106121 675434 106127
rect 675394 105820 675422 106121
rect 674422 105217 674474 105223
rect 674422 105159 674474 105165
rect 675382 105217 675434 105223
rect 675382 105159 675434 105165
rect 675394 104636 675422 105159
rect 675380 103258 675436 103267
rect 675380 103193 675436 103202
rect 675394 102786 675422 103193
rect 675764 101482 675820 101491
rect 675764 101417 675820 101426
rect 675778 100936 675806 101417
rect 663190 96485 663242 96491
rect 663190 96427 663242 96433
rect 665206 96485 665258 96491
rect 665206 96427 665258 96433
rect 646486 92711 646538 92717
rect 646486 92653 646538 92659
rect 659830 92711 659882 92717
rect 659830 92653 659882 92659
rect 646102 92489 646154 92495
rect 646102 92431 646154 92437
rect 646114 86395 646142 92431
rect 646292 88606 646348 88615
rect 646292 88541 646348 88550
rect 646306 87611 646334 88541
rect 646294 87605 646346 87611
rect 646294 87547 646346 87553
rect 646388 86978 646444 86987
rect 646388 86913 646444 86922
rect 646402 86797 646430 86913
rect 646390 86791 646442 86797
rect 646390 86733 646442 86739
rect 646100 86386 646156 86395
rect 646100 86321 646156 86330
rect 646498 85040 646526 92653
rect 647542 92637 647594 92643
rect 647542 92579 647594 92585
rect 647350 92563 647402 92569
rect 647350 92505 647402 92511
rect 647254 92267 647306 92273
rect 647254 92209 647306 92215
rect 646582 92193 646634 92199
rect 646582 92135 646634 92141
rect 646402 85012 646526 85040
rect 646004 84314 646060 84323
rect 646004 84249 646060 84258
rect 646018 81839 646046 84249
rect 646294 83165 646346 83171
rect 646292 83130 646294 83139
rect 646346 83130 646348 83139
rect 646292 83065 646348 83074
rect 646100 82686 646156 82695
rect 646100 82621 646156 82630
rect 646114 81913 646142 82621
rect 646102 81907 646154 81913
rect 646102 81849 646154 81855
rect 646006 81833 646058 81839
rect 646006 81775 646058 81781
rect 646294 77615 646346 77621
rect 646294 77557 646346 77563
rect 646306 76479 646334 77557
rect 646292 76470 646348 76479
rect 646292 76405 646348 76414
rect 646100 74102 646156 74111
rect 646100 74037 646156 74046
rect 646114 72441 646142 74037
rect 646292 73362 646348 73371
rect 646292 73297 646348 73306
rect 646306 72589 646334 73297
rect 646402 73223 646430 85012
rect 646486 84941 646538 84947
rect 646486 84883 646538 84889
rect 646498 84767 646526 84883
rect 646484 84758 646540 84767
rect 646484 84693 646540 84702
rect 646484 78986 646540 78995
rect 646484 78921 646540 78930
rect 646498 78287 646526 78921
rect 646486 78281 646538 78287
rect 646486 78223 646538 78229
rect 646594 76456 646622 92135
rect 647266 85951 647294 92209
rect 647252 85942 647308 85951
rect 647252 85877 647308 85886
rect 647362 81363 647390 92505
rect 647444 87570 647500 87579
rect 647444 87505 647500 87514
rect 647348 81354 647404 81363
rect 647348 81289 647404 81298
rect 646870 80279 646922 80285
rect 646870 80221 646922 80227
rect 646882 79883 646910 80221
rect 646868 79874 646924 79883
rect 646868 79809 646924 79818
rect 646870 78947 646922 78953
rect 646870 78889 646922 78895
rect 646882 78847 646910 78889
rect 646868 78838 646924 78847
rect 646868 78773 646924 78782
rect 646870 78355 646922 78361
rect 646870 78297 646922 78303
rect 646882 78255 646910 78297
rect 646868 78246 646924 78255
rect 646868 78181 646924 78190
rect 646678 77689 646730 77695
rect 646678 77631 646730 77637
rect 646690 76627 646718 77631
rect 647458 77473 647486 87505
rect 647554 82103 647582 92579
rect 647830 92341 647882 92347
rect 647830 92283 647882 92289
rect 647636 89198 647692 89207
rect 647636 89133 647692 89142
rect 647540 82094 647596 82103
rect 647540 82029 647596 82038
rect 647650 81691 647678 89133
rect 647842 85359 647870 92283
rect 658870 92193 658922 92199
rect 658870 92135 658922 92141
rect 647924 88014 647980 88023
rect 658882 87986 658910 92135
rect 659842 88000 659870 92653
rect 661750 92637 661802 92643
rect 661750 92579 661802 92585
rect 660694 92563 660746 92569
rect 660694 92505 660746 92511
rect 659842 87972 660144 88000
rect 660706 87986 660734 92505
rect 661174 92267 661226 92273
rect 661174 92209 661226 92215
rect 661186 88000 661214 92209
rect 661762 88000 661790 92579
rect 663094 92489 663146 92495
rect 663094 92431 663146 92437
rect 662518 92341 662570 92347
rect 662518 92283 662570 92289
rect 661186 87972 661440 88000
rect 661762 87972 662016 88000
rect 662530 87986 662558 92283
rect 663106 87986 663134 92431
rect 647924 87949 647980 87958
rect 647938 87093 647966 87949
rect 650998 87605 651050 87611
rect 650998 87547 651050 87553
rect 647926 87087 647978 87093
rect 647926 87029 647978 87035
rect 650900 86978 650956 86987
rect 650900 86913 650956 86922
rect 647828 85350 647884 85359
rect 647828 85285 647884 85294
rect 650914 84947 650942 86913
rect 651010 85359 651038 87547
rect 659362 87389 659616 87408
rect 652342 87383 652394 87389
rect 652342 87325 652394 87331
rect 659350 87383 659616 87389
rect 659402 87380 659616 87383
rect 659350 87325 659402 87331
rect 651094 86791 651146 86797
rect 651094 86733 651146 86739
rect 650996 85350 651052 85359
rect 650996 85285 651052 85294
rect 650902 84941 650954 84947
rect 650902 84883 650954 84889
rect 650996 84314 651052 84323
rect 650996 84249 651052 84258
rect 650900 82686 650956 82695
rect 650900 82621 650956 82630
rect 647638 81685 647690 81691
rect 647638 81627 647690 81633
rect 647924 81502 647980 81511
rect 647924 81437 647926 81446
rect 647978 81437 647980 81446
rect 647926 81405 647978 81411
rect 647924 80466 647980 80475
rect 647924 80401 647980 80410
rect 647938 79397 647966 80401
rect 647926 79391 647978 79397
rect 647926 79333 647978 79339
rect 647926 77763 647978 77769
rect 647926 77705 647978 77711
rect 647828 77654 647884 77663
rect 647828 77589 647884 77598
rect 647842 77547 647870 77589
rect 647830 77541 647882 77547
rect 647830 77483 647882 77489
rect 647446 77467 647498 77473
rect 647446 77409 647498 77415
rect 647938 77219 647966 77705
rect 650914 77621 650942 82621
rect 650902 77615 650954 77621
rect 650902 77557 650954 77563
rect 651010 77547 651038 84249
rect 651106 83435 651134 86733
rect 651188 86238 651244 86247
rect 651188 86173 651244 86182
rect 651092 83426 651148 83435
rect 651092 83361 651148 83370
rect 651202 78361 651230 86173
rect 652354 83731 652382 87325
rect 658006 87309 658058 87315
rect 656866 87232 657792 87260
rect 658058 87257 658320 87260
rect 658006 87251 658320 87257
rect 658018 87232 658320 87251
rect 652340 83722 652396 83731
rect 652340 83657 652396 83666
rect 651190 78355 651242 78361
rect 651190 78297 651242 78303
rect 650998 77541 651050 77547
rect 650998 77483 651050 77489
rect 647924 77210 647980 77219
rect 647924 77145 647980 77154
rect 646676 76618 646732 76627
rect 646676 76553 646732 76562
rect 646594 76428 646718 76456
rect 646486 75691 646538 75697
rect 646486 75633 646538 75639
rect 646498 75591 646526 75633
rect 646484 75582 646540 75591
rect 646484 75517 646540 75526
rect 646388 73214 646444 73223
rect 646388 73149 646444 73158
rect 646294 72583 646346 72589
rect 646294 72525 646346 72531
rect 646102 72435 646154 72441
rect 646102 72377 646154 72383
rect 646690 72335 646718 76428
rect 647926 76135 647978 76141
rect 647926 76077 647978 76083
rect 647938 74999 647966 76077
rect 656866 75697 656894 87232
rect 657046 87161 657098 87167
rect 657046 87103 657098 87109
rect 657058 83171 657086 87103
rect 657046 83165 657098 83171
rect 657046 83107 657098 83113
rect 661078 81685 661130 81691
rect 661130 81633 661440 81636
rect 661078 81627 661440 81633
rect 661090 81608 661440 81627
rect 657538 81469 657792 81488
rect 657526 81463 657792 81469
rect 657578 81460 657792 81463
rect 657526 81405 657578 81411
rect 662900 81206 662956 81215
rect 662900 81141 662956 81150
rect 656962 81016 657216 81044
rect 656962 80285 656990 81016
rect 656950 80279 657002 80285
rect 656950 80221 657002 80227
rect 658306 77695 658334 81030
rect 658882 78953 658910 81030
rect 659602 80748 659630 81030
rect 659554 80729 659630 80748
rect 659446 80723 659498 80729
rect 659446 80665 659498 80671
rect 659542 80723 659630 80729
rect 659594 80720 659630 80723
rect 659542 80665 659594 80671
rect 658870 78947 658922 78953
rect 658870 78889 658922 78895
rect 658294 77689 658346 77695
rect 658294 77631 658346 77637
rect 659458 77473 659486 80665
rect 659446 77467 659498 77473
rect 659446 77409 659498 77415
rect 656854 75691 656906 75697
rect 656854 75633 656906 75639
rect 647924 74990 647980 74999
rect 647924 74925 647980 74934
rect 647156 73954 647212 73963
rect 647156 73889 647212 73898
rect 646676 72326 646732 72335
rect 646676 72261 646732 72270
rect 647170 72219 647198 73889
rect 660130 72219 660158 81030
rect 660706 79397 660734 81030
rect 661762 81016 662016 81044
rect 660694 79391 660746 79397
rect 660694 79333 660746 79339
rect 661762 76141 661790 81016
rect 662530 78287 662558 81030
rect 662518 78281 662570 78287
rect 662518 78223 662570 78229
rect 662914 77769 662942 81141
rect 663202 79249 663230 96427
rect 663286 87087 663338 87093
rect 663286 87029 663338 87035
rect 663298 85211 663326 87029
rect 663572 85646 663628 85655
rect 663572 85581 663628 85590
rect 663284 85202 663340 85211
rect 663284 85137 663340 85146
rect 663476 84758 663532 84767
rect 663476 84693 663532 84702
rect 663380 82834 663436 82843
rect 663380 82769 663436 82778
rect 663284 82094 663340 82103
rect 663284 82029 663340 82038
rect 663298 81913 663326 82029
rect 663286 81907 663338 81913
rect 663286 81849 663338 81855
rect 663394 81839 663422 82769
rect 663382 81833 663434 81839
rect 663382 81775 663434 81781
rect 663490 80156 663518 84693
rect 663298 80128 663518 80156
rect 663190 79243 663242 79249
rect 663190 79185 663242 79191
rect 662902 77763 662954 77769
rect 662902 77705 662954 77711
rect 661750 76135 661802 76141
rect 661750 76077 661802 76083
rect 663298 72589 663326 80128
rect 663586 80008 663614 85581
rect 663490 79980 663614 80008
rect 663286 72583 663338 72589
rect 663286 72525 663338 72531
rect 663490 72441 663518 79980
rect 663478 72435 663530 72441
rect 663478 72377 663530 72383
rect 647158 72213 647210 72219
rect 647158 72155 647210 72161
rect 660118 72213 660170 72219
rect 660118 72155 660170 72161
rect 645718 51789 645770 51795
rect 645718 51731 645770 51737
rect 645622 48977 645674 48983
rect 645622 48919 645674 48925
rect 645334 48903 645386 48909
rect 645334 48845 645386 48851
rect 645238 48755 645290 48761
rect 645238 48697 645290 48703
rect 625076 40654 625132 40663
rect 625076 40589 625132 40598
rect 141812 40358 141868 40367
rect 141812 40293 141868 40302
rect 457748 40358 457804 40367
rect 457748 40293 457804 40302
<< via2 >>
rect 108596 1005449 108598 1005466
rect 108598 1005449 108650 1005466
rect 108650 1005449 108652 1005466
rect 108596 1005410 108652 1005449
rect 114164 1005427 114220 1005466
rect 114164 1005410 114166 1005427
rect 114166 1005410 114218 1005427
rect 114218 1005410 114220 1005427
rect 308756 1005427 308812 1005466
rect 308756 1005410 308758 1005427
rect 308758 1005410 308810 1005427
rect 308810 1005410 308812 1005427
rect 321044 1005410 321100 1005466
rect 321428 1005410 321484 1005466
rect 325460 1005410 325516 1005466
rect 357908 1005449 357910 1005466
rect 357910 1005449 357962 1005466
rect 357962 1005449 357964 1005466
rect 357908 1005410 357964 1005449
rect 364148 1005427 364204 1005466
rect 364148 1005410 364150 1005427
rect 364150 1005410 364202 1005427
rect 364202 1005410 364204 1005427
rect 81044 995790 81100 995846
rect 85940 995642 85996 995698
rect 61844 993866 61900 993922
rect 42068 968706 42124 968762
rect 41780 967078 41836 967134
rect 41780 965006 41836 965062
rect 42164 963970 42220 964026
rect 41780 963378 41836 963434
rect 42164 962786 42220 962842
rect 42548 962490 42604 962546
rect 41876 962046 41932 962102
rect 42356 962046 42412 962102
rect 41780 959678 41836 959734
rect 41780 959086 41836 959142
rect 41972 958346 42028 958402
rect 41780 957754 41836 957810
rect 41780 956126 41836 956182
rect 42164 949318 42220 949374
rect 42548 953166 42604 953222
rect 42356 948430 42412 948486
rect 42644 947542 42700 947598
rect 40340 946506 40396 946562
rect 40052 945026 40108 945082
rect 42836 942214 42892 942270
rect 43124 947838 43180 947894
rect 43028 946950 43084 947006
rect 42932 939106 42988 939162
rect 44756 945618 44812 945674
rect 44564 944730 44620 944786
rect 43028 933038 43084 933094
rect 42356 932594 42412 932650
rect 42356 930983 42412 931022
rect 42356 930966 42358 930983
rect 42358 930966 42410 930983
rect 42410 930966 42412 930983
rect 43124 907138 43180 907194
rect 43124 887158 43180 887214
rect 42356 823853 42358 823870
rect 42358 823853 42410 823870
rect 42410 823853 42412 823870
rect 42356 823814 42412 823853
rect 42452 822630 42508 822686
rect 42356 822225 42358 822242
rect 42358 822225 42410 822242
rect 42410 822225 42412 822242
rect 42356 822186 42412 822225
rect 43220 821150 43276 821206
rect 40340 820706 40396 820762
rect 40052 820114 40108 820170
rect 37460 819078 37516 819134
rect 41684 817894 41740 817950
rect 40148 816710 40204 816766
rect 37364 812714 37420 812770
rect 40244 815822 40300 815878
rect 37364 802206 37420 802262
rect 37268 802058 37324 802114
rect 41588 815230 41644 815286
rect 40244 801910 40300 801966
rect 41972 814342 42028 814398
rect 41876 813602 41932 813658
rect 41780 809606 41836 809662
rect 41780 800282 41836 800338
rect 42356 812270 42412 812326
rect 42068 811086 42124 811142
rect 42164 808274 42220 808330
rect 42068 800282 42124 800338
rect 42260 805183 42316 805222
rect 42260 805166 42262 805183
rect 42262 805166 42314 805183
rect 42314 805166 42316 805183
rect 43124 810346 43180 810402
rect 43028 809310 43084 809366
rect 42452 807534 42508 807590
rect 42452 803538 42508 803594
rect 42260 799986 42316 800042
rect 42452 797914 42508 797970
rect 41780 794214 41836 794270
rect 41780 791254 41836 791310
rect 42164 790958 42220 791014
rect 42740 794806 42796 794862
rect 42452 791846 42508 791902
rect 42740 791698 42796 791754
rect 42740 780467 42796 780506
rect 42740 780450 42742 780467
rect 42742 780450 42794 780467
rect 42794 780450 42796 780467
rect 42452 779897 42454 779914
rect 42454 779897 42506 779914
rect 42506 779897 42508 779914
rect 42452 779858 42508 779897
rect 42740 778861 42742 778878
rect 42742 778861 42794 778878
rect 42794 778861 42796 778878
rect 42740 778822 42796 778861
rect 43316 777934 43372 777990
rect 43220 777194 43276 777250
rect 42836 774826 42892 774882
rect 38996 773494 39052 773550
rect 38804 772606 38860 772662
rect 37364 769498 37420 769554
rect 42452 771126 42508 771182
rect 41780 770386 41836 770442
rect 38804 760174 38860 760230
rect 37364 758546 37420 758602
rect 41876 769054 41932 769110
rect 41972 767870 42028 767926
rect 42068 765206 42124 765262
rect 42740 763726 42796 763782
rect 42740 762263 42796 762302
rect 42740 762246 42742 762263
rect 42742 762246 42794 762263
rect 42794 762246 42796 762263
rect 41780 751738 41836 751794
rect 41780 748630 41836 748686
rect 42164 747446 42220 747502
rect 41972 747298 42028 747354
rect 42932 772458 42988 772514
rect 43124 767722 43180 767778
rect 43028 766982 43084 767038
rect 42836 751886 42892 751942
rect 42836 751590 42892 751646
rect 42740 746854 42796 746910
rect 42932 747150 42988 747206
rect 42644 737251 42700 737290
rect 42644 737234 42646 737251
rect 42646 737234 42698 737251
rect 42698 737234 42700 737251
rect 42356 736681 42358 736698
rect 42358 736681 42410 736698
rect 42410 736681 42412 736698
rect 42356 736642 42412 736681
rect 42068 735902 42124 735958
rect 40148 730278 40204 730334
rect 37364 726282 37420 726338
rect 37364 716958 37420 717014
rect 40244 729538 40300 729594
rect 41684 728798 41740 728854
rect 41588 727170 41644 727226
rect 40244 716662 40300 716718
rect 41972 727910 42028 727966
rect 41780 725838 41836 725894
rect 42356 735475 42412 735514
rect 42356 735458 42358 735475
rect 42358 735458 42410 735475
rect 42410 735458 42412 735475
rect 43220 734866 43276 734922
rect 42932 731610 42988 731666
rect 42068 725838 42124 725894
rect 42068 724654 42124 724710
rect 41972 716070 42028 716126
rect 42164 724062 42220 724118
rect 41876 713850 41932 713906
rect 42068 713850 42124 713906
rect 41876 711630 41932 711686
rect 43028 722138 43084 722194
rect 42836 710742 42892 710798
rect 41780 708522 41836 708578
rect 42164 707782 42220 707838
rect 41780 706746 41836 706802
rect 42164 706154 42220 706210
rect 41780 704674 41836 704730
rect 41780 704082 41836 704138
rect 42260 703638 42316 703694
rect 43316 733978 43372 734034
rect 43316 720510 43372 720566
rect 43316 719030 43372 719086
rect 42836 703490 42892 703546
rect 42260 700826 42316 700882
rect 42260 700530 42316 700586
rect 42644 694035 42700 694074
rect 42644 694018 42646 694035
rect 42646 694018 42698 694035
rect 42698 694018 42700 694035
rect 42356 693426 42412 693482
rect 41396 692686 41452 692742
rect 40244 687062 40300 687118
rect 41300 679958 41356 680014
rect 42644 692429 42646 692446
rect 42646 692429 42698 692446
rect 42698 692429 42700 692446
rect 42644 692390 42700 692429
rect 43508 691650 43564 691706
rect 43220 690762 43276 690818
rect 41876 688246 41932 688302
rect 41780 683954 41836 684010
rect 41396 670930 41452 670986
rect 42740 686026 42796 686082
rect 42068 684842 42124 684898
rect 41972 679514 42028 679570
rect 42164 682622 42220 682678
rect 42260 681438 42316 681494
rect 42356 677146 42412 677202
rect 43124 678182 43180 678238
rect 42356 675683 42412 675722
rect 42356 675666 42358 675683
rect 42358 675666 42410 675683
rect 42410 675666 42412 675683
rect 42164 670634 42220 670690
rect 42644 670930 42700 670986
rect 42452 669302 42508 669358
rect 42548 668858 42604 668914
rect 42548 668710 42604 668766
rect 41780 666638 41836 666694
rect 42836 666490 42892 666546
rect 42164 661458 42220 661514
rect 41876 660718 41932 660774
rect 43028 664714 43084 664770
rect 41780 656722 41836 656778
rect 41780 656130 41836 656186
rect 42836 650802 42892 650858
rect 42452 649783 42508 649822
rect 42452 649766 42454 649783
rect 42454 649766 42506 649783
rect 42506 649766 42508 649783
rect 42452 649509 42454 649526
rect 42454 649509 42506 649526
rect 42506 649509 42508 649526
rect 42452 649470 42508 649509
rect 43220 648434 43276 648490
rect 43124 645326 43180 645382
rect 40052 643846 40108 643902
rect 41876 642366 41932 642422
rect 41780 640738 41836 640794
rect 41492 638370 41548 638426
rect 42164 641626 42220 641682
rect 41972 639406 42028 639462
rect 41876 627418 41932 627474
rect 42068 636742 42124 636798
rect 43028 636594 43084 636650
rect 42644 635706 42700 635762
rect 42452 632467 42508 632506
rect 42452 632450 42454 632467
rect 42454 632450 42506 632467
rect 42506 632450 42508 632467
rect 42164 627418 42220 627474
rect 42932 634966 42988 635022
rect 43124 627862 43180 627918
rect 42164 623422 42220 623478
rect 42068 620166 42124 620222
rect 42452 623866 42508 623922
rect 42452 623274 42508 623330
rect 41972 618390 42028 618446
rect 41780 617798 41836 617854
rect 42932 620758 42988 620814
rect 42740 618242 42796 618298
rect 42836 618094 42892 618150
rect 42740 607699 42742 607716
rect 42742 607699 42794 607716
rect 42794 607699 42796 607716
rect 42740 607660 42796 607699
rect 42740 606863 42796 606902
rect 42740 606846 42742 606863
rect 42742 606846 42794 606863
rect 42794 606846 42796 606863
rect 42452 606254 42508 606310
rect 43508 647546 43564 647602
rect 43796 646954 43852 647010
rect 43604 646066 43660 646122
rect 43508 605218 43564 605274
rect 43220 604626 43276 604682
rect 43412 603738 43468 603794
rect 43124 602110 43180 602166
rect 40052 600630 40108 600686
rect 43028 599594 43084 599650
rect 41876 598410 41932 598466
rect 41780 597522 41836 597578
rect 42068 596190 42124 596246
rect 41972 595154 42028 595210
rect 41876 584202 41932 584258
rect 42836 594858 42892 594914
rect 42164 593674 42220 593730
rect 42068 584202 42124 584258
rect 42548 593526 42604 593582
rect 42548 592342 42604 592398
rect 42452 590566 42508 590622
rect 42452 589251 42508 589290
rect 42452 589234 42454 589251
rect 42454 589234 42506 589251
rect 42506 589234 42508 589251
rect 42548 584646 42604 584702
rect 42932 591750 42988 591806
rect 43028 585386 43084 585442
rect 42452 584498 42508 584554
rect 42452 584202 42508 584258
rect 41780 577098 41836 577154
rect 42260 575914 42316 575970
rect 41972 575174 42028 575230
rect 41780 574582 41836 574638
rect 43028 580058 43084 580114
rect 42932 578282 42988 578338
rect 42452 573990 42508 574046
rect 42836 573842 42892 573898
rect 34484 564666 34540 564722
rect 42452 563499 42508 563538
rect 42452 563482 42454 563499
rect 42454 563482 42506 563499
rect 42506 563482 42508 563499
rect 42356 563038 42412 563094
rect 43220 562002 43276 562058
rect 41972 558598 42028 558654
rect 40052 557414 40108 557470
rect 37364 553566 37420 553622
rect 40148 556674 40204 556730
rect 41876 555934 41932 555990
rect 41684 555194 41740 555250
rect 40148 544242 40204 544298
rect 37364 542910 37420 542966
rect 41780 554306 41836 554362
rect 41684 541282 41740 541338
rect 41876 541134 41932 541190
rect 42068 552974 42124 553030
rect 42356 551938 42412 551994
rect 42164 550014 42220 550070
rect 42068 540986 42124 541042
rect 43028 551642 43084 551698
rect 42932 551050 42988 551106
rect 42836 548534 42892 548590
rect 42644 546257 42700 546296
rect 42644 546240 42646 546257
rect 42646 546240 42698 546257
rect 42698 546240 42700 546257
rect 43124 549274 43180 549330
rect 43028 538766 43084 538822
rect 42932 536842 42988 536898
rect 42836 535658 42892 535714
rect 41876 531958 41932 532014
rect 41780 531218 41836 531274
rect 42740 532550 42796 532606
rect 42644 532254 42700 532310
rect 43796 603738 43852 603794
rect 43604 602850 43660 602906
rect 43508 561558 43564 561614
rect 43412 560522 43468 560578
rect 42644 436907 42646 436924
rect 42646 436907 42698 436924
rect 42698 436907 42700 436924
rect 42644 436868 42700 436907
rect 42644 436093 42646 436110
rect 42646 436093 42698 436110
rect 42698 436093 42700 436110
rect 42644 436054 42700 436093
rect 42356 435462 42412 435518
rect 43220 433538 43276 433594
rect 43604 559782 43660 559838
rect 43508 434426 43564 434482
rect 43412 432946 43468 433002
rect 42164 429838 42220 429894
rect 41780 426730 41836 426786
rect 37364 424362 37420 424418
rect 37268 421994 37324 422050
rect 40148 423178 40204 423234
rect 40244 420514 40300 420570
rect 43604 432058 43660 432114
rect 42740 424066 42796 424122
rect 42644 420070 42700 420126
rect 42644 418607 42700 418646
rect 42644 418590 42646 418607
rect 42646 418590 42698 418607
rect 42698 418590 42700 418607
rect 43028 421254 43084 421310
rect 41780 406010 41836 406066
rect 41972 404826 42028 404882
rect 41780 403790 41836 403846
rect 42164 402606 42220 402662
rect 41780 401866 41836 401922
rect 41780 400090 41836 400146
rect 42260 399942 42316 399998
rect 41780 399498 41836 399554
rect 41780 398758 41836 398814
rect 42356 393913 42358 393930
rect 42358 393913 42410 393930
rect 42410 393913 42412 393930
rect 42356 393874 42412 393913
rect 42356 393173 42358 393190
rect 42358 393173 42410 393190
rect 42410 393173 42412 393190
rect 42356 393134 42412 393173
rect 42356 392285 42358 392302
rect 42358 392285 42410 392302
rect 42410 392285 42412 392302
rect 42356 392246 42412 392285
rect 43220 391210 43276 391266
rect 43124 390914 43180 390970
rect 43028 387214 43084 387270
rect 35924 384402 35980 384458
rect 41780 383514 41836 383570
rect 37172 381146 37228 381202
rect 40052 380406 40108 380462
rect 37268 378778 37324 378834
rect 37364 378038 37420 378094
rect 40148 377446 40204 377502
rect 35924 371526 35980 371582
rect 42932 380258 42988 380314
rect 42356 376706 42412 376762
rect 42356 375243 42412 375282
rect 42356 375226 42358 375243
rect 42358 375226 42410 375243
rect 42410 375226 42412 375243
rect 42068 362794 42124 362850
rect 41876 361906 41932 361962
rect 41780 361314 41836 361370
rect 41780 359390 41836 359446
rect 41780 358650 41836 358706
rect 41876 356874 41932 356930
rect 41780 356430 41836 356486
rect 41780 355542 41836 355598
rect 42356 350697 42358 350714
rect 42358 350697 42410 350714
rect 42410 350697 42412 350714
rect 42356 350658 42412 350697
rect 42644 349661 42646 349678
rect 42646 349661 42698 349678
rect 42698 349661 42700 349678
rect 42644 349622 42700 349661
rect 42356 349069 42358 349086
rect 42358 349069 42410 349086
rect 42410 349069 42412 349086
rect 42356 349030 42412 349069
rect 43220 347698 43276 347754
rect 43220 347550 43276 347606
rect 42740 344072 42796 344128
rect 39956 340298 40012 340354
rect 37172 337338 37228 337394
rect 42356 337930 42412 337986
rect 40052 337190 40108 337246
rect 40244 334082 40300 334138
rect 42164 333490 42220 333546
rect 42164 332027 42220 332066
rect 42164 332010 42166 332027
rect 42166 332010 42218 332027
rect 42218 332010 42220 332027
rect 42356 327422 42412 327478
rect 43124 335414 43180 335470
rect 42356 322982 42412 323038
rect 41780 319726 41836 319782
rect 41876 318690 41932 318746
rect 41780 317950 41836 318006
rect 42164 317358 42220 317414
rect 41780 316174 41836 316230
rect 41780 315434 41836 315490
rect 41780 313658 41836 313714
rect 41780 313214 41836 313270
rect 41780 312326 41836 312382
rect 42260 307481 42262 307498
rect 42262 307481 42314 307498
rect 42314 307481 42316 307498
rect 42260 307442 42316 307481
rect 42260 306741 42262 306758
rect 42262 306741 42314 306758
rect 42314 306741 42316 306758
rect 42260 306702 42316 306741
rect 42836 305666 42892 305722
rect 43220 304038 43276 304094
rect 43220 303890 43276 303946
rect 41972 300338 42028 300394
rect 39956 297230 40012 297286
rect 37364 293974 37420 294030
rect 40148 293974 40204 294030
rect 40244 290866 40300 290922
rect 42164 294714 42220 294770
rect 42260 292642 42316 292698
rect 42836 292198 42892 292254
rect 42548 290274 42604 290330
rect 42644 289107 42700 289146
rect 42644 289090 42646 289107
rect 42646 289090 42698 289107
rect 42698 289090 42700 289107
rect 42260 283614 42316 283670
rect 42548 281542 42604 281598
rect 41780 276510 41836 276566
rect 41972 275178 42028 275234
rect 41780 274586 41836 274642
rect 41780 272810 41836 272866
rect 41780 272366 41836 272422
rect 41780 270590 41836 270646
rect 42260 270442 42316 270498
rect 41780 269998 41836 270054
rect 41780 269110 41836 269166
rect 42260 264265 42262 264282
rect 42262 264265 42314 264282
rect 42314 264265 42316 264282
rect 42260 264226 42316 264265
rect 42260 263525 42262 263542
rect 42262 263525 42314 263542
rect 42314 263525 42316 263542
rect 42260 263486 42316 263525
rect 42260 262637 42262 262654
rect 42262 262637 42314 262654
rect 42314 262637 42316 262654
rect 42260 262598 42316 262637
rect 41780 259490 41836 259546
rect 40244 254014 40300 254070
rect 37364 250758 37420 250814
rect 40052 250758 40108 250814
rect 37268 249130 37324 249186
rect 40148 247946 40204 248002
rect 43028 259342 43084 259398
rect 41972 257122 42028 257178
rect 42068 251498 42124 251554
rect 42260 248390 42316 248446
rect 42068 240694 42124 240750
rect 42356 245430 42412 245486
rect 42356 240694 42412 240750
rect 43412 261562 43468 261618
rect 43220 260822 43276 260878
rect 43124 245282 43180 245338
rect 43124 243358 43180 243414
rect 42452 237882 42508 237938
rect 47444 946210 47500 946266
rect 41780 233294 41836 233350
rect 41876 231666 41932 231722
rect 41780 231074 41836 231130
rect 42068 230482 42124 230538
rect 41780 229594 41836 229650
rect 41780 229002 41836 229058
rect 41780 227226 41836 227282
rect 41780 226782 41836 226838
rect 41780 225894 41836 225950
rect 42356 221049 42358 221066
rect 42358 221049 42410 221066
rect 42410 221049 42412 221066
rect 42356 221010 42412 221049
rect 42356 220309 42358 220326
rect 42358 220309 42410 220326
rect 42410 220309 42412 220326
rect 42356 220270 42412 220309
rect 42356 219421 42358 219438
rect 42358 219421 42410 219438
rect 42410 219421 42412 219438
rect 42356 219382 42412 219421
rect 43220 217606 43276 217662
rect 43508 216866 43564 216922
rect 43316 216126 43372 216182
rect 41972 213906 42028 213962
rect 41876 210798 41932 210854
rect 37268 207690 37324 207746
rect 40148 207098 40204 207154
rect 37364 206062 37420 206118
rect 40244 204582 40300 204638
rect 43124 209762 43180 209818
rect 42068 208282 42124 208338
rect 42356 205470 42412 205526
rect 42164 204325 42166 204342
rect 42166 204325 42218 204342
rect 42218 204325 42220 204342
rect 42164 204286 42220 204325
rect 42164 202954 42220 203010
rect 42164 197626 42220 197682
rect 42356 197330 42412 197386
rect 42356 195110 42412 195166
rect 42068 190966 42124 191022
rect 41780 190078 41836 190134
rect 41876 189042 41932 189098
rect 41780 188302 41836 188358
rect 59540 973146 59596 973202
rect 62036 992090 62092 992146
rect 78356 993718 78412 993774
rect 82580 995050 82636 995106
rect 82580 993866 82636 993922
rect 85364 995346 85420 995402
rect 86420 995198 86476 995254
rect 84500 994606 84556 994662
rect 83444 993570 83500 993626
rect 93044 993570 93100 993626
rect 83444 992090 83500 992146
rect 62036 962490 62092 962546
rect 61844 962046 61900 962102
rect 59540 958790 59596 958846
rect 59540 944599 59596 944638
rect 59540 944582 59542 944599
rect 59542 944582 59594 944599
rect 59594 944582 59596 944599
rect 59540 930078 59596 930134
rect 59540 915722 59596 915778
rect 58196 901531 58252 901570
rect 58196 901514 58198 901531
rect 58198 901514 58250 901531
rect 58250 901514 58252 901531
rect 59540 887010 59596 887066
rect 58964 872506 59020 872562
rect 59540 858315 59596 858354
rect 59540 858298 59542 858315
rect 59542 858298 59594 858315
rect 59594 858298 59596 858315
rect 59540 843942 59596 843998
rect 59540 829586 59596 829642
rect 59540 815230 59596 815286
rect 59540 800726 59596 800782
rect 58964 786518 59020 786574
rect 59540 772014 59596 772070
rect 59540 757658 59596 757714
rect 59540 743302 59596 743358
rect 58388 728946 58444 729002
rect 58388 714590 58444 714646
rect 57812 700234 57868 700290
rect 59540 685878 59596 685934
rect 59444 671522 59500 671578
rect 59540 657166 59596 657222
rect 59252 642810 59308 642866
rect 58004 628454 58060 628510
rect 59444 613950 59500 614006
rect 59540 599742 59596 599798
rect 59540 585386 59596 585442
rect 59540 570882 59596 570938
rect 59540 556674 59596 556730
rect 59540 542318 59596 542374
rect 59540 527814 59596 527870
rect 59348 513458 59404 513514
rect 57812 499102 57868 499158
rect 59540 484746 59596 484802
rect 59540 470390 59596 470446
rect 59540 456034 59596 456090
rect 57812 441530 57868 441586
rect 59540 427322 59596 427378
rect 59540 412818 59596 412874
rect 58964 398610 59020 398666
rect 59540 384106 59596 384162
rect 59540 369750 59596 369806
rect 59540 355542 59596 355598
rect 59540 341038 59596 341094
rect 59540 326682 59596 326738
rect 59540 312326 59596 312382
rect 59540 297970 59596 298026
rect 59540 283614 59596 283670
rect 217268 1005279 217324 1005318
rect 217268 1005262 217270 1005279
rect 217270 1005262 217322 1005279
rect 217322 1005262 217324 1005279
rect 218900 1005279 218956 1005318
rect 218900 1005262 218902 1005279
rect 218902 1005262 218954 1005279
rect 218954 1005262 218956 1005279
rect 223124 1005262 223180 1005318
rect 115220 1005153 115222 1005170
rect 115222 1005153 115274 1005170
rect 115274 1005153 115276 1005170
rect 115220 1005114 115276 1005153
rect 221876 1005114 221932 1005170
rect 150356 1002489 150358 1002506
rect 150358 1002489 150410 1002506
rect 150410 1002489 150412 1002506
rect 100628 995955 100684 995994
rect 100628 995938 100630 995955
rect 100630 995938 100682 995955
rect 100682 995938 100684 995955
rect 107252 995938 107308 995994
rect 94868 995790 94924 995846
rect 99956 995829 99958 995846
rect 99958 995829 100010 995846
rect 100010 995829 100012 995846
rect 99956 995790 100012 995829
rect 102164 995807 102220 995846
rect 102164 995790 102166 995807
rect 102166 995790 102218 995807
rect 102218 995790 102220 995807
rect 105332 995790 105388 995846
rect 94964 995642 95020 995698
rect 98996 995642 99052 995698
rect 94676 995346 94732 995402
rect 94868 995346 94924 995402
rect 102164 995511 102220 995550
rect 102164 995494 102166 995511
rect 102166 995494 102218 995511
rect 102218 995494 102220 995511
rect 98996 995198 99052 995254
rect 100724 995198 100780 995254
rect 100820 985469 100822 985486
rect 100822 985469 100874 985486
rect 100874 985469 100876 985486
rect 100820 985430 100876 985469
rect 106580 995198 106636 995254
rect 106580 994606 106636 994662
rect 113300 995807 113356 995846
rect 113300 995790 113302 995807
rect 113302 995790 113354 995807
rect 113354 995790 113356 995807
rect 113492 995829 113494 995846
rect 113494 995829 113546 995846
rect 113546 995829 113548 995846
rect 113492 995790 113548 995829
rect 115220 995494 115276 995550
rect 108212 995198 108268 995254
rect 108404 995198 108460 995254
rect 108404 993718 108460 993774
rect 115316 995346 115372 995402
rect 120980 995642 121036 995698
rect 131732 995790 131788 995846
rect 133076 995346 133132 995402
rect 134228 995050 134284 995106
rect 136724 995642 136780 995698
rect 134612 994754 134668 994810
rect 137396 995494 137452 995550
rect 136148 994014 136204 994070
rect 150356 1002450 150412 1002489
rect 153620 1002341 153622 1002358
rect 153622 1002341 153674 1002358
rect 153674 1002341 153676 1002358
rect 153620 1002302 153676 1002341
rect 160244 1000839 160300 1000878
rect 160244 1000822 160246 1000839
rect 160246 1000822 160298 1000839
rect 160298 1000822 160300 1000839
rect 155156 999507 155212 999546
rect 155156 999490 155158 999507
rect 155158 999490 155210 999507
rect 155210 999490 155212 999507
rect 158612 999529 158614 999546
rect 158614 999529 158666 999546
rect 158666 999529 158668 999546
rect 158612 999490 158668 999529
rect 156884 999381 156886 999398
rect 156886 999381 156938 999398
rect 156938 999381 156940 999398
rect 156884 999342 156940 999381
rect 162260 996273 162262 996290
rect 162262 996273 162314 996290
rect 162314 996273 162316 996290
rect 144212 995790 144268 995846
rect 162260 996234 162316 996273
rect 163124 996103 163180 996142
rect 163124 996086 163126 996103
rect 163126 996086 163178 996103
rect 163178 996086 163180 996103
rect 145268 995938 145324 995994
rect 149108 995938 149164 995994
rect 149492 995938 149548 995994
rect 152084 995955 152140 995994
rect 152084 995938 152086 995955
rect 152086 995938 152138 995955
rect 152138 995938 152140 995955
rect 143636 995050 143692 995106
rect 141236 994497 141238 994514
rect 141238 994497 141290 994514
rect 141290 994497 141292 994514
rect 141236 994458 141292 994497
rect 140372 993718 140428 993774
rect 120884 985469 120886 985486
rect 120886 985469 120938 985486
rect 120938 985469 120940 985486
rect 120884 985430 120940 985469
rect 164180 995955 164236 995994
rect 164180 995938 164182 995955
rect 164182 995938 164234 995955
rect 164234 995938 164236 995955
rect 164564 995977 164566 995994
rect 164566 995977 164618 995994
rect 164618 995977 164620 995994
rect 164564 995938 164620 995977
rect 165620 995807 165676 995846
rect 165620 995790 165622 995807
rect 165622 995790 165674 995807
rect 165674 995790 165676 995807
rect 166292 995790 166348 995846
rect 208436 1000839 208492 1000878
rect 208436 1000822 208438 1000839
rect 208438 1000822 208490 1000839
rect 208490 1000822 208492 1000839
rect 152564 995198 152620 995254
rect 156692 995198 156748 995254
rect 159572 995198 159628 995254
rect 161204 995198 161260 995254
rect 146996 994606 147052 994662
rect 158420 994623 158476 994662
rect 158420 994606 158422 994623
rect 158422 994606 158474 994623
rect 158474 994606 158476 994623
rect 156692 994014 156748 994070
rect 185108 995790 185164 995846
rect 170228 995642 170284 995698
rect 178484 994623 178540 994662
rect 178484 994606 178486 994623
rect 178486 994606 178538 994623
rect 178538 994606 178540 994623
rect 183764 995346 183820 995402
rect 188084 995790 188140 995846
rect 195380 995642 195436 995698
rect 198548 995938 198604 995994
rect 198644 995790 198700 995846
rect 185780 994606 185836 994662
rect 189428 995494 189484 995550
rect 188852 995346 188908 995402
rect 187316 994162 187372 994218
rect 185780 994014 185836 994070
rect 192404 995198 192460 995254
rect 191540 993866 191596 993922
rect 205652 996547 205708 996586
rect 205652 996530 205654 996547
rect 205654 996530 205706 996547
rect 205706 996530 205708 996547
rect 211700 996547 211756 996586
rect 211700 996530 211702 996547
rect 211702 996530 211754 996547
rect 211754 996530 211756 996547
rect 203636 996125 203638 996142
rect 203638 996125 203690 996142
rect 203690 996125 203692 996142
rect 203636 996086 203692 996125
rect 213332 996103 213388 996142
rect 213332 996086 213334 996103
rect 213334 996086 213386 996103
rect 213386 996086 213388 996103
rect 202964 995977 202966 995994
rect 202966 995977 203018 995994
rect 203018 995977 203020 995994
rect 202964 995938 203020 995977
rect 206612 995938 206668 995994
rect 201812 995790 201868 995846
rect 204980 995807 205036 995846
rect 204980 995790 204982 995807
rect 204982 995790 205034 995807
rect 205034 995790 205036 995807
rect 201620 995198 201676 995254
rect 198644 994902 198700 994958
rect 206996 995659 207052 995698
rect 206996 995642 206998 995659
rect 206998 995642 207050 995659
rect 207050 995642 207052 995659
rect 201812 995494 201868 995550
rect 212660 995494 212716 995550
rect 207380 995198 207436 995254
rect 211028 995198 211084 995254
rect 207284 995050 207340 995106
rect 207380 994162 207436 994218
rect 215636 995955 215692 995994
rect 215636 995938 215638 995955
rect 215638 995938 215690 995955
rect 215690 995938 215692 995955
rect 216884 995977 216886 995994
rect 216886 995977 216938 995994
rect 216938 995977 216940 995994
rect 216884 995938 216940 995977
rect 214100 995829 214102 995846
rect 214102 995829 214154 995846
rect 214154 995829 214156 995846
rect 214100 995790 214156 995829
rect 218900 995642 218956 995698
rect 246836 1005114 246892 1005170
rect 239540 995790 239596 995846
rect 246452 995790 246508 995846
rect 241844 995642 241900 995698
rect 231476 994162 231532 994218
rect 237428 995050 237484 995106
rect 240212 995494 240268 995550
rect 254036 1002467 254092 1002506
rect 254036 1002450 254038 1002467
rect 254038 1002450 254090 1002467
rect 254090 1002450 254092 1002467
rect 253172 1002319 253228 1002358
rect 253172 1002302 253174 1002319
rect 253174 1002302 253226 1002319
rect 253226 1002302 253228 1002319
rect 243572 995198 243628 995254
rect 238676 994606 238732 994662
rect 237428 994014 237484 994070
rect 247604 995385 247606 995402
rect 247606 995385 247658 995402
rect 247658 995385 247660 995402
rect 247604 995346 247660 995385
rect 259604 999381 259606 999398
rect 259606 999381 259658 999398
rect 259658 999381 259660 999398
rect 259604 999342 259660 999381
rect 259124 995938 259180 995994
rect 261428 995938 261484 995994
rect 261812 995938 261868 995994
rect 250484 995198 250540 995254
rect 250676 995198 250732 995254
rect 254804 995790 254860 995846
rect 255956 995790 256012 995846
rect 260468 995790 260524 995846
rect 255956 995494 256012 995550
rect 260468 994606 260524 994662
rect 263060 999507 263116 999546
rect 263060 999490 263062 999507
rect 263062 999490 263114 999507
rect 263114 999490 263116 999507
rect 265940 996103 265996 996142
rect 265940 996086 265942 996103
rect 265942 996086 265994 996103
rect 265994 996086 265996 996103
rect 266804 996125 266806 996142
rect 266806 996125 266858 996142
rect 266858 996125 266860 996142
rect 266804 996086 266860 996125
rect 265076 995977 265078 995994
rect 265078 995977 265130 995994
rect 265130 995977 265132 995994
rect 265076 995938 265132 995977
rect 266996 995955 267052 995994
rect 266996 995938 266998 995955
rect 266998 995938 267050 995955
rect 267050 995938 267052 995955
rect 268628 995790 268684 995846
rect 273620 995790 273676 995846
rect 264020 995346 264076 995402
rect 261812 994162 261868 994218
rect 161300 981007 161356 981046
rect 161300 980990 161302 981007
rect 161302 980990 161354 981007
rect 161354 980990 161356 981007
rect 171284 980990 171340 981046
rect 239060 985282 239116 985338
rect 239540 985282 239596 985338
rect 239156 985151 239212 985190
rect 239156 985134 239158 985151
rect 239158 985134 239210 985151
rect 239210 985134 239212 985151
rect 239732 985151 239788 985190
rect 239732 985134 239734 985151
rect 239734 985134 239786 985151
rect 239786 985134 239788 985151
rect 292436 995790 292492 995846
rect 293588 995790 293644 995846
rect 298292 995790 298348 995846
rect 273716 995642 273772 995698
rect 291092 995642 291148 995698
rect 307988 1005279 308044 1005318
rect 307988 1005262 307990 1005279
rect 307990 1005262 308042 1005279
rect 308042 1005262 308044 1005279
rect 309620 1005301 309622 1005318
rect 309622 1005301 309674 1005318
rect 309674 1005301 309676 1005318
rect 309620 1005262 309676 1005301
rect 318644 1005279 318700 1005318
rect 318644 1005262 318646 1005279
rect 318646 1005262 318698 1005279
rect 318698 1005262 318700 1005279
rect 365012 1005449 365014 1005466
rect 365014 1005449 365066 1005466
rect 365066 1005449 365068 1005466
rect 365012 1005410 365068 1005449
rect 365780 1005279 365836 1005318
rect 365780 1005262 365782 1005279
rect 365782 1005262 365834 1005279
rect 365834 1005262 365836 1005279
rect 366740 1005301 366742 1005318
rect 366742 1005301 366794 1005318
rect 366794 1005301 366796 1005318
rect 366740 1005262 366796 1005301
rect 315188 1005153 315190 1005170
rect 315190 1005153 315242 1005170
rect 315242 1005153 315244 1005170
rect 298580 1002302 298636 1002358
rect 286004 994162 286060 994218
rect 279284 993609 279286 993626
rect 279286 993609 279338 993626
rect 279338 993609 279340 993626
rect 279284 993570 279340 993609
rect 288788 995050 288844 995106
rect 291764 995494 291820 995550
rect 290324 994458 290380 994514
rect 295412 994310 295468 994366
rect 288788 994014 288844 994070
rect 288404 993570 288460 993626
rect 288404 992090 288460 992146
rect 299540 995642 299596 995698
rect 299732 995938 299788 995994
rect 299636 995494 299692 995550
rect 315188 1005114 315244 1005153
rect 305588 1002467 305644 1002506
rect 305588 1002450 305590 1002467
rect 305590 1002450 305642 1002467
rect 305642 1002450 305644 1002467
rect 307604 1002489 307606 1002506
rect 307606 1002489 307658 1002506
rect 307658 1002489 307660 1002506
rect 307604 1002450 307660 1002489
rect 304724 1002319 304780 1002358
rect 304724 1002302 304726 1002319
rect 304726 1002302 304778 1002319
rect 304778 1002302 304780 1002319
rect 306548 1002341 306550 1002358
rect 306550 1002341 306602 1002358
rect 306602 1002341 306604 1002358
rect 306548 1002302 306604 1002341
rect 311156 999507 311212 999546
rect 311156 999490 311158 999507
rect 311158 999490 311210 999507
rect 311210 999490 311212 999507
rect 310292 999381 310294 999398
rect 310294 999381 310346 999398
rect 310346 999381 310348 999398
rect 310292 999342 310348 999381
rect 317108 996103 317164 996142
rect 317108 996086 317110 996103
rect 317110 996086 317162 996103
rect 317162 996086 317164 996103
rect 318644 996125 318646 996142
rect 318646 996125 318698 996142
rect 318698 996125 318700 996142
rect 318644 996086 318700 996125
rect 363476 1005153 363478 1005170
rect 363478 1005153 363530 1005170
rect 363530 1005153 363532 1005170
rect 313844 995938 313900 995994
rect 316340 995977 316342 995994
rect 316342 995977 316394 995994
rect 316394 995977 316396 995994
rect 316340 995938 316396 995977
rect 326804 995938 326860 995994
rect 310292 995642 310348 995698
rect 311060 995198 311116 995254
rect 310292 994458 310348 994514
rect 311060 994162 311116 994218
rect 323924 995642 323980 995698
rect 363476 1005114 363532 1005153
rect 359924 1003969 359926 1003986
rect 359926 1003969 359978 1003986
rect 359978 1003969 359980 1003986
rect 359924 1003930 359980 1003969
rect 358388 1003799 358444 1003838
rect 358388 1003782 358390 1003799
rect 358390 1003782 358442 1003799
rect 358442 1003782 358444 1003799
rect 359060 1003821 359062 1003838
rect 359062 1003821 359114 1003838
rect 359114 1003821 359116 1003838
rect 359060 1003782 359116 1003821
rect 360692 1003673 360694 1003690
rect 360694 1003673 360746 1003690
rect 360746 1003673 360748 1003690
rect 360692 1003634 360748 1003673
rect 361556 1000839 361612 1000878
rect 361556 1000822 361558 1000839
rect 361558 1000822 361610 1000839
rect 361610 1000822 361612 1000839
rect 356276 998049 356278 998066
rect 356278 998049 356330 998066
rect 356330 998049 356332 998066
rect 356276 998010 356332 998049
rect 357044 998027 357100 998066
rect 357044 998010 357046 998027
rect 357046 998010 357098 998027
rect 357098 998010 357100 998027
rect 367892 997901 367894 997918
rect 367894 997901 367946 997918
rect 367946 997901 367948 997918
rect 367892 997862 367948 997901
rect 362324 995938 362380 995994
rect 367124 995977 367126 995994
rect 367126 995977 367178 995994
rect 367178 995977 367180 995994
rect 367124 995938 367180 995977
rect 343892 995642 343948 995698
rect 369044 997879 369100 997918
rect 369044 997862 369046 997879
rect 369046 997862 369098 997879
rect 369098 997862 369100 997879
rect 370580 995955 370636 995994
rect 370580 995938 370582 995955
rect 370582 995938 370634 995955
rect 370634 995938 370636 995955
rect 371348 995807 371404 995846
rect 371348 995790 371350 995807
rect 371350 995790 371402 995807
rect 371402 995790 371404 995807
rect 371540 995642 371596 995698
rect 377300 995938 377356 995994
rect 380180 995790 380236 995846
rect 380276 995642 380332 995698
rect 430868 1005449 430870 1005466
rect 430870 1005449 430922 1005466
rect 430922 1005449 430924 1005466
rect 430868 1005410 430924 1005449
rect 424532 1005301 424534 1005318
rect 424534 1005301 424586 1005318
rect 424586 1005301 424588 1005318
rect 424532 1005262 424588 1005301
rect 425300 1005279 425356 1005318
rect 425300 1005262 425302 1005279
rect 425302 1005262 425354 1005279
rect 425354 1005262 425356 1005279
rect 430772 1005262 430828 1005318
rect 426068 1005153 426070 1005170
rect 426070 1005153 426122 1005170
rect 426122 1005153 426124 1005170
rect 426068 1005114 426124 1005153
rect 433172 1005131 433228 1005170
rect 433172 1005114 433174 1005131
rect 433174 1005114 433226 1005131
rect 433226 1005114 433228 1005131
rect 435572 1005114 435628 1005170
rect 423380 1003947 423436 1003986
rect 423380 1003930 423382 1003947
rect 423382 1003930 423434 1003947
rect 423434 1003930 423436 1003947
rect 426452 1003821 426454 1003838
rect 426454 1003821 426506 1003838
rect 426506 1003821 426508 1003838
rect 426452 1003782 426508 1003821
rect 388820 995790 388876 995846
rect 428084 1003673 428086 1003690
rect 428086 1003673 428138 1003690
rect 428138 1003673 428140 1003690
rect 428084 1003634 428140 1003673
rect 434132 1001135 434188 1001174
rect 434132 1001118 434134 1001135
rect 434134 1001118 434186 1001135
rect 434186 1001118 434188 1001135
rect 432500 1000987 432556 1001026
rect 432500 1000970 432502 1000987
rect 432502 1000970 432554 1000987
rect 432554 1000970 432556 1000987
rect 427316 1000839 427372 1000878
rect 427316 1000822 427318 1000839
rect 427318 1000822 427370 1000839
rect 427370 1000822 427372 1000839
rect 428948 1000861 428950 1000878
rect 428950 1000861 429002 1000878
rect 429002 1000861 429004 1000878
rect 428948 1000822 429004 1000861
rect 436340 996234 436396 996290
rect 436436 996125 436438 996142
rect 436438 996125 436490 996142
rect 436490 996125 436492 996142
rect 436436 996086 436492 996125
rect 429716 995938 429772 995994
rect 434132 995977 434134 995994
rect 434134 995977 434186 995994
rect 434186 995977 434188 995994
rect 434132 995938 434188 995977
rect 445076 995938 445132 995994
rect 422516 995790 422572 995846
rect 396692 995642 396748 995698
rect 390836 994014 390892 994070
rect 438740 995807 438796 995846
rect 438740 995790 438742 995807
rect 438742 995790 438794 995807
rect 438794 995790 438796 995807
rect 440660 995642 440716 995698
rect 390164 993570 390220 993626
rect 390164 992090 390220 992146
rect 471476 995494 471532 995550
rect 466484 995346 466540 995402
rect 501140 1005427 501196 1005466
rect 501140 1005410 501142 1005427
rect 501142 1005410 501194 1005427
rect 501194 1005410 501196 1005427
rect 504596 1005279 504652 1005318
rect 504596 1005262 504598 1005279
rect 504598 1005262 504650 1005279
rect 504650 1005262 504652 1005279
rect 554516 1005301 554518 1005318
rect 554518 1005301 554570 1005318
rect 554570 1005301 554572 1005318
rect 554516 1005262 554572 1005301
rect 555764 1005279 555820 1005318
rect 555764 1005262 555766 1005279
rect 555766 1005262 555818 1005279
rect 555818 1005262 555820 1005279
rect 500756 1005153 500758 1005170
rect 500758 1005153 500810 1005170
rect 500810 1005153 500812 1005170
rect 500756 1005114 500812 1005153
rect 471956 995938 472012 995994
rect 472052 995642 472108 995698
rect 472244 995790 472300 995846
rect 488852 999490 488908 999546
rect 480980 995790 481036 995846
rect 485684 995790 485740 995846
rect 477044 995642 477100 995698
rect 476468 995346 476524 995402
rect 469460 993587 469516 993626
rect 479924 995642 479980 995698
rect 488852 995642 488908 995698
rect 482036 995494 482092 995550
rect 479828 994014 479884 994070
rect 485588 994014 485644 994070
rect 497588 999529 497590 999546
rect 497590 999529 497642 999546
rect 497642 999529 497644 999546
rect 497588 999490 497644 999529
rect 502772 1002467 502828 1002506
rect 502772 1002450 502774 1002467
rect 502774 1002450 502826 1002467
rect 502826 1002450 502828 1002467
rect 503444 1002489 503446 1002506
rect 503446 1002489 503498 1002506
rect 503498 1002489 503500 1002506
rect 503444 1002450 503500 1002489
rect 505076 1002341 505078 1002358
rect 505078 1002341 505130 1002358
rect 505130 1002341 505132 1002358
rect 505076 1002302 505132 1002341
rect 511028 1001283 511084 1001322
rect 511028 1001266 511030 1001283
rect 511030 1001266 511082 1001283
rect 511082 1001266 511084 1001283
rect 509396 1001009 509398 1001026
rect 509398 1001009 509450 1001026
rect 509450 1001009 509452 1001026
rect 509396 1000970 509452 1001009
rect 507764 1000713 507766 1000730
rect 507766 1000713 507818 1000730
rect 507818 1000713 507820 1000730
rect 507764 1000674 507820 1000713
rect 506324 999507 506380 999546
rect 506324 999490 506326 999507
rect 506326 999490 506378 999507
rect 506378 999490 506380 999507
rect 502388 999359 502444 999398
rect 502388 999342 502390 999359
rect 502390 999342 502442 999359
rect 502442 999342 502444 999359
rect 508628 996547 508684 996586
rect 508628 996530 508630 996547
rect 508630 996530 508682 996547
rect 508682 996530 508684 996547
rect 510260 996569 510262 996586
rect 510262 996569 510314 996586
rect 510314 996569 510316 996586
rect 510260 996530 510316 996569
rect 511124 995955 511180 995994
rect 511124 995938 511126 995955
rect 511126 995938 511178 995955
rect 511178 995938 511180 995955
rect 499988 995790 500044 995846
rect 511892 995829 511894 995846
rect 511894 995829 511946 995846
rect 511946 995829 511948 995846
rect 511892 995790 511948 995829
rect 506612 995198 506668 995254
rect 516692 1001283 516748 1001322
rect 516692 1001266 516694 1001283
rect 516694 1001266 516746 1001283
rect 516746 1001266 516748 1001283
rect 516692 1001009 516694 1001026
rect 516694 1001009 516746 1001026
rect 516746 1001009 516748 1001026
rect 516692 1000970 516748 1001009
rect 516692 1000713 516694 1000730
rect 516694 1000713 516746 1000730
rect 516746 1000713 516748 1000730
rect 516692 1000674 516748 1000713
rect 516692 999786 516748 999842
rect 516788 999507 516844 999546
rect 516788 999490 516790 999507
rect 516790 999490 516842 999507
rect 516842 999490 516844 999507
rect 516692 999359 516748 999398
rect 516692 999342 516694 999359
rect 516694 999342 516746 999359
rect 516746 999342 516748 999359
rect 513428 996125 513430 996142
rect 513430 996125 513482 996142
rect 513482 996125 513484 996142
rect 513428 996086 513484 996125
rect 513428 995977 513430 995994
rect 513430 995977 513482 995994
rect 513482 995977 513484 995994
rect 513428 995938 513484 995977
rect 518420 995642 518476 995698
rect 469460 993570 469462 993587
rect 469462 993570 469514 993587
rect 469514 993570 469516 993587
rect 518612 995494 518668 995550
rect 553748 1005153 553750 1005170
rect 553750 1005153 553802 1005170
rect 553802 1005153 553804 1005170
rect 521396 999638 521452 999694
rect 553748 1005114 553804 1005153
rect 552596 1003821 552598 1003838
rect 552598 1003821 552650 1003838
rect 552650 1003821 552652 1003838
rect 552596 1003782 552652 1003821
rect 556532 1003799 556588 1003838
rect 556532 1003782 556534 1003799
rect 556534 1003782 556586 1003799
rect 556586 1003782 556588 1003799
rect 551732 1003673 551734 1003690
rect 551734 1003673 551786 1003690
rect 551786 1003673 551788 1003690
rect 551732 1003634 551788 1003673
rect 559220 1002637 559222 1002654
rect 559222 1002637 559274 1002654
rect 559274 1002637 559276 1002654
rect 559220 1002598 559276 1002637
rect 559988 1002615 560044 1002654
rect 559988 1002598 559990 1002615
rect 559990 1002598 560042 1002615
rect 560042 1002598 560044 1002615
rect 562196 1002489 562198 1002506
rect 562198 1002489 562250 1002506
rect 562250 1002489 562252 1002506
rect 562196 1002450 562252 1002489
rect 564596 1002467 564652 1002506
rect 564596 1002450 564598 1002467
rect 564598 1002450 564650 1002467
rect 564650 1002450 564652 1002467
rect 544244 1002302 544300 1002358
rect 560468 1002341 560470 1002358
rect 560470 1002341 560522 1002358
rect 560522 1002341 560524 1002358
rect 560468 1002302 560524 1002341
rect 561524 1002319 561580 1002358
rect 561524 1002302 561526 1002319
rect 561526 1002302 561578 1002319
rect 561578 1002302 561580 1002319
rect 523604 1001266 523660 1001322
rect 523508 1000674 523564 1000730
rect 521588 999934 521644 999990
rect 523316 999786 523372 999842
rect 521492 999490 521548 999546
rect 521108 999342 521164 999398
rect 520916 995494 520972 995550
rect 521300 995938 521356 995994
rect 521204 995790 521260 995846
rect 523316 995346 523372 995402
rect 523508 995938 523564 995994
rect 523700 1000970 523756 1001026
rect 523604 995642 523660 995698
rect 523892 999934 523948 999990
rect 523796 999342 523852 999398
rect 523988 999638 524044 999694
rect 524084 999490 524140 999546
rect 527924 995790 527980 995846
rect 532244 995790 532300 995846
rect 526100 995642 526156 995698
rect 530900 995346 530956 995402
rect 531188 994162 531244 994218
rect 535316 995494 535372 995550
rect 555284 998027 555340 998066
rect 555284 998010 555286 998027
rect 555286 998010 555338 998027
rect 555338 998010 555340 998027
rect 557300 997879 557356 997918
rect 557300 997862 557302 997879
rect 557302 997862 557354 997879
rect 557354 997862 557356 997879
rect 564788 995977 564790 995994
rect 564790 995977 564842 995994
rect 564842 995977 564844 995994
rect 564788 995938 564844 995977
rect 562772 995642 562828 995698
rect 563540 995659 563596 995698
rect 563540 995642 563542 995659
rect 563542 995642 563594 995659
rect 563594 995642 563596 995659
rect 557972 995346 558028 995402
rect 567572 994458 567628 994514
rect 570356 995642 570412 995698
rect 570548 995494 570604 995550
rect 570452 994310 570508 994366
rect 573140 995790 573196 995846
rect 573236 994606 573292 994662
rect 628148 994458 628204 994514
rect 604724 994014 604780 994070
rect 622004 993718 622060 993774
rect 631796 994606 631852 994662
rect 631028 994162 631084 994218
rect 218900 980733 218902 980750
rect 218902 980733 218954 980750
rect 218954 980733 218956 980750
rect 218900 980694 218956 980733
rect 238964 980694 239020 980750
rect 634292 994310 634348 994366
rect 632756 994162 632812 994218
rect 649556 993866 649612 993922
rect 70580 262746 70636 262802
rect 77780 269258 77836 269314
rect 83636 264078 83692 264134
rect 88436 269406 88492 269462
rect 86036 263930 86092 263986
rect 82868 263782 82924 263838
rect 95636 269702 95692 269758
rect 96788 269554 96844 269610
rect 99188 264522 99244 264578
rect 102644 269998 102700 270054
rect 103892 269850 103948 269906
rect 106292 264670 106348 264726
rect 100244 264374 100300 264430
rect 93236 264226 93292 264282
rect 111092 270294 111148 270350
rect 109844 270146 109900 270202
rect 121748 270442 121804 270498
rect 118100 264818 118156 264874
rect 129236 270590 129292 270646
rect 135956 269110 136012 269166
rect 125300 263338 125356 263394
rect 65204 246318 65260 246374
rect 65012 246170 65068 246226
rect 80660 245321 80662 245338
rect 80662 245321 80714 245338
rect 80714 245321 80716 245338
rect 80660 245282 80716 245321
rect 100724 245134 100780 245190
rect 126548 245134 126604 245190
rect 126740 245134 126796 245190
rect 139220 263190 139276 263246
rect 140660 239214 140716 239270
rect 140756 239066 140812 239122
rect 143156 268814 143212 268870
rect 146036 240546 146092 240602
rect 144020 239806 144076 239862
rect 144116 238622 144172 238678
rect 144020 236271 144076 236310
rect 144020 236254 144022 236271
rect 144022 236254 144074 236271
rect 144074 236254 144076 236271
rect 144020 233590 144076 233646
rect 144116 232110 144172 232166
rect 144020 231370 144076 231426
rect 144212 230186 144268 230242
rect 144020 228410 144076 228466
rect 144116 227670 144172 227726
rect 144020 226634 144076 226690
rect 144020 225006 144076 225062
rect 144116 223674 144172 223730
rect 144020 222934 144076 222990
rect 144020 220122 144076 220178
rect 144020 218198 144076 218254
rect 144116 215238 144172 215294
rect 144020 213314 144076 213370
rect 145364 214498 145420 214554
rect 144020 211686 144076 211742
rect 144116 209762 144172 209818
rect 144020 207433 144022 207450
rect 144022 207433 144074 207450
rect 144074 207433 144076 207450
rect 144020 207394 144076 207433
rect 144212 203250 144268 203306
rect 144788 196590 144844 196646
rect 144596 194814 144652 194870
rect 41780 185934 41836 185990
rect 41780 184158 41836 184214
rect 41780 183566 41836 183622
rect 41780 182826 41836 182882
rect 144020 184454 144076 184510
rect 144020 181790 144076 181846
rect 144116 180458 144172 180514
rect 144020 178573 144022 178590
rect 144022 178573 144074 178590
rect 144074 178573 144076 178590
rect 144020 178534 144076 178573
rect 42740 177054 42796 177110
rect 144020 176758 144076 176814
rect 144020 173354 144076 173410
rect 144020 171282 144076 171338
rect 144116 168322 144172 168378
rect 144020 167582 144076 167638
rect 144020 166546 144076 166602
rect 144116 163586 144172 163642
rect 144020 162846 144076 162902
rect 144500 159886 144556 159942
rect 144020 159294 144076 159350
rect 144308 158110 144364 158166
rect 144212 156334 144268 156390
rect 144020 155611 144076 155650
rect 144020 155594 144022 155611
rect 144022 155594 144074 155611
rect 144074 155594 144076 155611
rect 144116 154410 144172 154466
rect 144020 152930 144076 152986
rect 144116 151598 144172 151654
rect 144020 150858 144076 150914
rect 144020 147158 144076 147214
rect 141524 137538 141580 137594
rect 141524 120962 141580 121018
rect 141044 118594 141100 118650
rect 141044 118298 141100 118354
rect 144212 147898 144268 147954
rect 144212 145974 144268 146030
rect 144212 142422 144268 142478
rect 144212 138426 144268 138482
rect 144212 132802 144268 132858
rect 144212 131026 144268 131082
rect 144212 129990 144268 130046
rect 144116 105866 144172 105922
rect 144020 104830 144076 104886
rect 144020 103942 144076 103998
rect 144116 102758 144172 102814
rect 144020 101278 144076 101334
rect 144020 99798 144076 99854
rect 144116 99058 144172 99114
rect 144020 98039 144076 98078
rect 144020 98022 144022 98039
rect 144022 98022 144074 98039
rect 144074 98022 144076 98039
rect 144020 96246 144076 96302
rect 144116 94322 144172 94378
rect 144020 92694 144076 92750
rect 144500 149082 144556 149138
rect 144404 143162 144460 143218
rect 144404 139462 144460 139518
rect 144692 141238 144748 141294
rect 144500 135022 144556 135078
rect 144404 133986 144460 134042
rect 144404 120962 144460 121018
rect 144308 106458 144364 106514
rect 144116 90770 144172 90826
rect 144020 89586 144076 89642
rect 144020 87810 144076 87866
rect 144020 85886 144076 85942
rect 144020 82334 144076 82390
rect 144020 81150 144076 81206
rect 144116 79374 144172 79430
rect 144020 78634 144076 78690
rect 144116 75674 144172 75730
rect 144020 75082 144076 75138
rect 144020 73898 144076 73954
rect 144116 72714 144172 72770
rect 144020 70938 144076 70994
rect 144020 69754 144076 69810
rect 144020 67534 144076 67590
rect 144020 66350 144076 66406
rect 144020 64761 144022 64778
rect 144022 64761 144074 64778
rect 144074 64761 144076 64778
rect 144020 64722 144076 64761
rect 144020 62650 144076 62706
rect 144020 58654 144076 58710
rect 144212 69014 144268 69070
rect 144020 57322 144076 57378
rect 144116 56434 144172 56490
rect 144020 54675 144076 54714
rect 144020 54658 144022 54675
rect 144022 54658 144074 54675
rect 144074 54658 144076 54675
rect 144020 53770 144076 53826
rect 144692 135910 144748 135966
rect 144596 124366 144652 124422
rect 144596 121554 144652 121610
rect 144596 120814 144652 120870
rect 144596 118315 144652 118354
rect 144596 118298 144598 118315
rect 144598 118298 144650 118315
rect 144650 118298 144652 118315
rect 144596 116670 144652 116726
rect 144596 114154 144652 114210
rect 144596 112395 144652 112434
rect 144596 112378 144598 112395
rect 144598 112378 144650 112395
rect 144650 112378 144652 112395
rect 144596 109714 144652 109770
rect 144596 107511 144652 107550
rect 144596 107494 144598 107511
rect 144598 107494 144650 107511
rect 144650 107494 144652 107511
rect 144884 174390 144940 174446
rect 145076 172022 145132 172078
rect 144980 161366 145036 161422
rect 144884 144198 144940 144254
rect 144788 125106 144844 125162
rect 144788 122590 144844 122646
rect 144788 119038 144844 119094
rect 144788 113118 144844 113174
rect 144788 111194 144844 111250
rect 144692 106606 144748 106662
rect 144596 106310 144652 106366
rect 144692 100834 144748 100890
rect 144788 87070 144844 87126
rect 145268 170098 145324 170154
rect 145172 164770 145228 164826
rect 145460 210502 145516 210558
rect 145556 207986 145612 208042
rect 145652 205618 145708 205674
rect 145844 205026 145900 205082
rect 145748 201326 145804 201382
rect 145940 190078 145996 190134
rect 149588 240398 149644 240454
rect 146228 236846 146284 236902
rect 146132 186378 146188 186434
rect 146036 108234 146092 108290
rect 145940 83518 145996 83574
rect 146420 235070 146476 235126
rect 146900 230077 146902 230094
rect 146902 230077 146954 230094
rect 146954 230077 146956 230094
rect 146900 230038 146956 230077
rect 146804 202066 146860 202122
rect 146324 185194 146380 185250
rect 146228 91362 146284 91418
rect 146228 65462 146284 65518
rect 146420 183270 146476 183326
rect 146708 199550 146764 199606
rect 146804 198975 146860 199014
rect 146804 198958 146806 198975
rect 146806 198958 146858 198975
rect 146858 198958 146860 198975
rect 146804 197774 146860 197830
rect 146804 193630 146860 193686
rect 146804 192890 146860 192946
rect 146708 191706 146764 191762
rect 146708 189338 146764 189394
rect 146804 188154 146860 188210
rect 146804 179718 146860 179774
rect 146612 176018 146668 176074
rect 146804 157222 146860 157278
rect 146612 156778 146668 156834
rect 146516 129250 146572 129306
rect 146708 115355 146764 115394
rect 146708 115338 146710 115355
rect 146710 115338 146762 115355
rect 146762 115338 146764 115355
rect 146708 115190 146764 115246
rect 146516 95506 146572 95562
rect 146516 84110 146572 84166
rect 146900 127474 146956 127530
rect 146900 126882 146956 126938
rect 147092 115190 147148 115246
rect 146900 77450 146956 77506
rect 146516 59542 146572 59598
rect 146900 62354 146956 62410
rect 146900 60726 146956 60782
rect 158420 245025 158422 245042
rect 158422 245025 158474 245042
rect 158474 245025 158476 245042
rect 158420 244986 158476 245025
rect 162644 47850 162700 47906
rect 166868 230055 166924 230094
rect 166868 230038 166870 230055
rect 166870 230038 166922 230055
rect 166922 230038 166924 230055
rect 168500 244838 168556 244894
rect 168404 48590 168460 48646
rect 171284 48442 171340 48498
rect 174164 48294 174220 48350
rect 165524 47554 165580 47610
rect 216596 263486 216652 263542
rect 252020 266907 252076 266946
rect 252020 266890 252022 266907
rect 252022 266890 252074 266907
rect 252074 266890 252076 266907
rect 255668 266002 255724 266058
rect 256148 267778 256204 267834
rect 256916 267334 256972 267390
rect 256532 266907 256588 266946
rect 256532 266890 256534 266907
rect 256534 266890 256586 266907
rect 256586 266890 256588 266907
rect 256724 266150 256780 266206
rect 257300 267186 257356 267242
rect 257780 267038 257836 267094
rect 258452 266890 258508 266946
rect 258932 266742 258988 266798
rect 259028 266594 259084 266650
rect 259508 266446 259564 266502
rect 259988 266298 260044 266354
rect 263444 262006 263500 262062
rect 263252 260378 263308 260434
rect 262772 260230 262828 260286
rect 263924 261710 263980 261766
rect 264308 261414 264364 261470
rect 264884 261266 264940 261322
rect 265460 261118 265516 261174
rect 265844 260970 265900 261026
rect 266036 260822 266092 260878
rect 268244 273550 268300 273606
rect 267764 273402 267820 273458
rect 267572 271922 267628 271978
rect 268724 273254 268780 273310
rect 269108 273106 269164 273162
rect 269780 272958 269836 273014
rect 270260 272810 270316 272866
rect 270452 272662 270508 272718
rect 270836 272514 270892 272570
rect 271316 272366 271372 272422
rect 272564 272218 272620 272274
rect 271988 260674 272044 260730
rect 272372 260526 272428 260582
rect 273044 272070 273100 272126
rect 279284 263042 279340 263098
rect 319220 267630 319276 267686
rect 320276 267482 320332 267538
rect 319604 265854 319660 265910
rect 321908 265854 321964 265910
rect 326804 268666 326860 268722
rect 326900 261858 326956 261914
rect 327476 261562 327532 261618
rect 367988 262894 368044 262950
rect 380084 265262 380140 265318
rect 382388 265301 382390 265318
rect 382390 265301 382442 265318
rect 382442 265301 382444 265318
rect 382388 265262 382444 265301
rect 382580 262154 382636 262210
rect 383636 268518 383692 268574
rect 384788 268962 384844 269018
rect 385460 262746 385516 262802
rect 386132 269406 386188 269462
rect 386516 262894 386572 262950
rect 387668 269258 387724 269314
rect 386708 262154 386764 262210
rect 389012 269998 389068 270054
rect 388532 269258 388588 269314
rect 388820 263782 388876 263838
rect 389396 264078 389452 264134
rect 389780 263930 389836 263986
rect 392180 270590 392236 270646
rect 390644 270294 390700 270350
rect 391604 269702 391660 269758
rect 391796 269275 391852 269314
rect 391796 269258 391798 269275
rect 391798 269258 391850 269275
rect 391850 269258 391852 269275
rect 391988 264226 392044 264282
rect 392564 269554 392620 269610
rect 392180 264078 392236 264134
rect 393044 264522 393100 264578
rect 393716 264374 393772 264430
rect 394484 262302 394540 262358
rect 394772 264670 394828 264726
rect 395060 269850 395116 269906
rect 395924 270146 395980 270202
rect 395348 268518 395404 268574
rect 397076 262319 397132 262358
rect 397076 262302 397078 262319
rect 397078 262302 397130 262319
rect 397130 262302 397132 262319
rect 397844 264818 397900 264874
rect 398996 270442 399052 270498
rect 398612 268814 398668 268870
rect 399572 263338 399628 263394
rect 400724 264078 400780 264134
rect 401108 263042 401164 263098
rect 402260 269110 402316 269166
rect 403316 263190 403372 263246
rect 210164 256382 210220 256438
rect 204788 230482 204844 230538
rect 201716 229446 201772 229502
rect 201620 228410 201676 228466
rect 204884 230038 204940 230094
rect 201812 227818 201868 227874
rect 193748 64130 193804 64186
rect 194132 62502 194188 62558
rect 188564 48146 188620 48202
rect 194420 90770 194476 90826
rect 194612 81298 194668 81354
rect 194516 79670 194572 79726
rect 195572 76414 195628 76470
rect 194708 69014 194764 69070
rect 194324 47998 194380 48054
rect 197588 225598 197644 225654
rect 201716 227226 201772 227282
rect 201812 226782 201868 226838
rect 201620 226190 201676 226246
rect 201524 225154 201580 225210
rect 201716 224579 201772 224618
rect 201716 224562 201718 224579
rect 201718 224562 201770 224579
rect 201770 224562 201772 224579
rect 201620 223970 201676 224026
rect 201716 223526 201772 223582
rect 201812 222934 201868 222990
rect 201524 222342 201580 222398
rect 198644 221306 198700 221362
rect 201716 220714 201772 220770
rect 201620 219678 201676 219734
rect 201812 219086 201868 219142
rect 201716 218050 201772 218106
rect 198164 217458 198220 217514
rect 197588 216422 197644 216478
rect 201716 215830 201772 215886
rect 201620 214794 201676 214850
rect 201236 214202 201292 214258
rect 201812 213166 201868 213222
rect 201716 212574 201772 212630
rect 201620 211538 201676 211594
rect 197300 93286 197356 93342
rect 199988 102166 200044 102222
rect 197684 91658 197740 91714
rect 198740 88550 198796 88606
rect 197780 82077 197782 82094
rect 197782 82077 197834 82094
rect 197834 82077 197836 82094
rect 197780 82038 197836 82077
rect 197396 79818 197452 79874
rect 198356 73306 198412 73362
rect 199316 61318 199372 61374
rect 200180 93434 200236 93490
rect 201716 101574 201772 101630
rect 201716 100577 201718 100594
rect 201718 100577 201770 100594
rect 201770 100577 201772 100594
rect 201716 100538 201772 100577
rect 201716 99946 201772 100002
rect 201620 98910 201676 98966
rect 201812 98318 201868 98374
rect 201716 96690 201772 96746
rect 201620 95654 201676 95710
rect 202964 97282 203020 97338
rect 201812 95062 201868 95118
rect 201716 94026 201772 94082
rect 201620 92398 201676 92454
rect 201716 91806 201772 91862
rect 201620 90178 201676 90234
rect 201812 89586 201868 89642
rect 201716 89142 201772 89198
rect 201524 87958 201580 88014
rect 201620 87514 201676 87570
rect 201812 86922 201868 86978
rect 201716 86330 201772 86386
rect 201716 85886 201772 85942
rect 201620 85294 201676 85350
rect 201812 84702 201868 84758
rect 201524 84258 201580 84314
rect 201908 83666 201964 83722
rect 201044 83074 201100 83130
rect 201716 82630 201772 82686
rect 201620 81446 201676 81502
rect 200276 80410 200332 80466
rect 200372 78782 200428 78838
rect 201716 78190 201772 78246
rect 201716 77154 201772 77210
rect 201620 76562 201676 76618
rect 201812 75526 201868 75582
rect 201524 74934 201580 74990
rect 201044 73898 201100 73954
rect 200948 73158 201004 73214
rect 201716 72270 201772 72326
rect 201716 71695 201772 71734
rect 201716 71678 201718 71695
rect 201718 71678 201770 71695
rect 201770 71678 201772 71695
rect 201620 70642 201676 70698
rect 201812 70050 201868 70106
rect 200468 69458 200524 69514
rect 201716 68422 201772 68478
rect 201620 67830 201676 67886
rect 201812 67386 201868 67442
rect 201524 66794 201580 66850
rect 201620 66202 201676 66258
rect 201716 65758 201772 65814
rect 200180 65166 200236 65222
rect 201716 64574 201772 64630
rect 201716 63538 201772 63594
rect 201716 62946 201772 63002
rect 201620 61910 201676 61966
rect 201620 60282 201676 60338
rect 201716 59690 201772 59746
rect 203156 54214 203212 54270
rect 206804 232702 206860 232758
rect 206708 231666 206764 231722
rect 206612 231074 206668 231130
rect 206516 230038 206572 230094
rect 206420 202806 206476 202862
rect 206900 232110 206956 232166
rect 206996 230482 207052 230538
rect 215540 252090 215596 252146
rect 209972 242174 210028 242230
rect 208340 242026 208396 242082
rect 207284 241878 207340 241934
rect 207284 55546 207340 55602
rect 207188 48738 207244 48794
rect 205172 47702 205228 47758
rect 208724 241878 208780 241934
rect 208916 240398 208972 240454
rect 208724 239806 208780 239862
rect 208916 239658 208972 239714
rect 209876 239658 209932 239714
rect 211508 237142 211564 237198
rect 211892 234034 211948 234090
rect 211508 233738 211564 233794
rect 210068 228854 210124 228910
rect 209972 221824 210028 221880
rect 209972 220196 210028 220252
rect 209972 218568 210028 218624
rect 209972 215312 210028 215368
rect 209972 212056 210028 212112
rect 209684 53326 209740 53382
rect 211316 233590 211372 233646
rect 212276 233886 212332 233942
rect 214196 233590 214252 233646
rect 215636 248538 215692 248594
rect 215540 243358 215596 243414
rect 215060 241730 215116 241786
rect 215444 239658 215500 239714
rect 216020 244098 216076 244154
rect 215828 240546 215884 240602
rect 215924 240398 215980 240454
rect 217076 237882 217132 237938
rect 216692 233738 216748 233794
rect 217652 243506 217708 243562
rect 218804 237734 218860 237790
rect 218996 237586 219052 237642
rect 221588 243654 221644 243710
rect 221012 238326 221068 238382
rect 223604 243950 223660 244006
rect 222740 238474 222796 238530
rect 224468 245282 224524 245338
rect 224468 244690 224524 244746
rect 224660 244690 224716 244746
rect 224180 238030 224236 238086
rect 226388 243802 226444 243858
rect 225812 238178 225868 238234
rect 228116 244542 228172 244598
rect 227444 238622 227500 238678
rect 229652 244394 229708 244450
rect 231188 243062 231244 243118
rect 230228 238770 230284 238826
rect 232052 238918 232108 238974
rect 232916 244246 232972 244302
rect 234356 242914 234412 242970
rect 235988 243210 236044 243266
rect 235124 237438 235180 237494
rect 238196 237290 238252 237346
rect 240596 241878 240652 241934
rect 241556 240842 241612 240898
rect 240980 240694 241036 240750
rect 242420 241286 242476 241342
rect 242324 241138 242380 241194
rect 241844 240102 241900 240158
rect 242804 241434 242860 241490
rect 243380 241582 243436 241638
rect 259220 245134 259276 245190
rect 259220 244986 259276 245042
rect 272372 233738 272428 233794
rect 279284 245134 279340 245190
rect 279284 244838 279340 244894
rect 280340 233738 280396 233794
rect 285428 241007 285484 241046
rect 285428 240990 285430 241007
rect 285430 240990 285482 241007
rect 285482 240990 285484 241007
rect 285716 240250 285772 240306
rect 285428 239806 285484 239862
rect 286676 240990 286732 241046
rect 289844 240990 289900 241046
rect 293300 239806 293356 239862
rect 294452 240990 294508 241046
rect 296660 244986 296716 245042
rect 296660 244838 296716 244894
rect 299156 240250 299212 240306
rect 210164 216940 210220 216996
rect 210164 213684 210220 213740
rect 306548 233738 306604 233794
rect 306932 233590 306988 233646
rect 325460 241730 325516 241786
rect 325460 239658 325516 239714
rect 331220 241878 331276 241934
rect 335156 244098 335212 244154
rect 338996 238326 339052 238382
rect 339860 245134 339916 245190
rect 339764 244986 339820 245042
rect 340820 243654 340876 243710
rect 341780 243950 341836 244006
rect 341204 238474 341260 238530
rect 342548 244690 342604 244746
rect 342164 238030 342220 238086
rect 343028 243802 343084 243858
rect 342836 240267 342892 240306
rect 342836 240250 342838 240267
rect 342838 240250 342890 240267
rect 342890 240250 342892 240267
rect 342740 239993 342742 240010
rect 342742 239993 342794 240010
rect 342794 239993 342796 240010
rect 342740 239954 342796 239993
rect 342740 238178 342796 238234
rect 343988 244542 344044 244598
rect 343412 238622 343468 238678
rect 344756 244394 344812 244450
rect 344372 237882 344428 237938
rect 345236 243062 345292 243118
rect 344852 238770 344908 238826
rect 346196 244246 346252 244302
rect 345620 238918 345676 238974
rect 347444 243210 347500 243266
rect 346964 242914 347020 242970
rect 347060 237438 347116 237494
rect 348404 243506 348460 243562
rect 348788 237290 348844 237346
rect 351380 240250 351436 240306
rect 350612 239954 350668 240010
rect 352244 237734 352300 237790
rect 354452 237586 354508 237642
rect 358868 239510 358924 239566
rect 359444 239362 359500 239418
rect 365684 241878 365740 241934
rect 365588 241730 365644 241786
rect 365396 241582 365452 241638
rect 365204 240250 365260 240306
rect 365780 241582 365836 241638
rect 365780 241138 365836 241194
rect 366068 241434 366124 241490
rect 366452 241434 366508 241490
rect 366452 241286 366508 241342
rect 366068 241138 366124 241194
rect 367604 241582 367660 241638
rect 367796 241582 367852 241638
rect 367412 240990 367468 241046
rect 369140 240842 369196 240898
rect 370196 240694 370252 240750
rect 368468 240102 368524 240158
rect 377108 240694 377164 240750
rect 377012 239806 377068 239862
rect 377492 239954 377548 240010
rect 378452 240102 378508 240158
rect 379220 241434 379276 241490
rect 377876 239658 377932 239714
rect 379316 240842 379372 240898
rect 383060 239510 383116 239566
rect 385076 243358 385132 243414
rect 394772 240546 394828 240602
rect 395252 239510 395308 239566
rect 403028 244986 403084 245042
rect 403220 244986 403276 245042
rect 408116 240250 408172 240306
rect 408980 241730 409036 241786
rect 409844 241878 409900 241934
rect 409364 240694 409420 240750
rect 410516 241138 410572 241194
rect 410324 239954 410380 240010
rect 408308 239806 408364 239862
rect 411572 241286 411628 241342
rect 413108 241582 413164 241638
rect 412628 241434 412684 241490
rect 412532 240990 412588 241046
rect 413780 240842 413836 240898
rect 412052 240102 412108 240158
rect 410900 239658 410956 239714
rect 420500 244838 420556 244894
rect 502292 266002 502348 266058
rect 505940 267778 505996 267834
rect 512756 267334 512812 267390
rect 516596 267186 516652 267242
rect 509492 266150 509548 266206
rect 520148 267038 520204 267094
rect 463604 245578 463660 245634
rect 440564 245282 440620 245338
rect 463604 245134 463660 245190
rect 523796 266890 523852 266946
rect 527348 266742 527404 266798
rect 530900 266594 530956 266650
rect 534452 266446 534508 266502
rect 538004 266298 538060 266354
rect 548756 268666 548812 268722
rect 567764 267630 567820 267686
rect 566516 262006 566572 262062
rect 570164 261710 570220 261766
rect 574580 267482 574636 267538
rect 573716 261414 573772 261470
rect 577268 261266 577324 261322
rect 580916 261118 580972 261174
rect 584372 260970 584428 261026
rect 598772 271922 598828 271978
rect 602228 273402 602284 273458
rect 605492 273550 605548 273606
rect 609428 273254 609484 273310
rect 612980 273106 613036 273162
rect 616532 272958 616588 273014
rect 620084 272810 620140 272866
rect 588020 260822 588076 260878
rect 623636 272662 623692 272718
rect 627284 272514 627340 272570
rect 630836 272366 630892 272422
rect 628436 261858 628492 261914
rect 635540 261562 635596 261618
rect 634388 260674 634444 260730
rect 641492 272218 641548 272274
rect 645140 272070 645196 272126
rect 647540 268962 647596 269018
rect 648692 263486 648748 263542
rect 637940 260526 637996 260582
rect 563060 260378 563116 260434
rect 559124 260230 559180 260286
rect 494516 243358 494572 243414
rect 521300 243358 521356 243414
rect 421844 242174 421900 242230
rect 415316 240398 415372 240454
rect 494516 242026 494572 242082
rect 505556 239231 505612 239270
rect 505556 239214 505558 239231
rect 505558 239214 505610 239231
rect 505610 239214 505612 239231
rect 510356 239105 510358 239122
rect 510358 239105 510410 239122
rect 510410 239105 510412 239122
rect 510356 239066 510412 239105
rect 541460 234626 541516 234682
rect 637172 233738 637228 233794
rect 638420 239066 638476 239122
rect 638036 234034 638092 234090
rect 637652 233886 637708 233942
rect 638132 233590 638188 233646
rect 638516 233590 638572 233646
rect 649652 752330 649708 752386
rect 639284 239066 639340 239122
rect 639284 233738 639340 233794
rect 210164 161218 210220 161274
rect 210164 153226 210220 153282
rect 209972 71826 210028 71882
rect 209972 71160 210028 71216
rect 209972 60800 210028 60856
rect 209972 59172 210028 59228
rect 209972 58062 210028 58118
rect 210164 101056 210220 101112
rect 210164 99428 210220 99484
rect 210164 97817 210220 97856
rect 210164 97800 210166 97817
rect 210166 97800 210218 97817
rect 210218 97800 210220 97817
rect 210164 96172 210220 96228
rect 210164 94544 210220 94600
rect 210164 87662 210220 87718
rect 210260 83370 210316 83426
rect 210260 77672 210316 77728
rect 210260 74455 210262 74472
rect 210262 74455 210314 74472
rect 210314 74455 210316 74472
rect 210260 74416 210316 74455
rect 210164 57026 210220 57082
rect 210068 54066 210124 54122
rect 210260 56434 210316 56490
rect 210356 54362 210412 54418
rect 210644 54362 210700 54418
rect 218612 54214 218668 54270
rect 214196 54066 214252 54122
rect 187604 41782 187660 41838
rect 194324 41782 194380 41838
rect 211316 45186 211372 45242
rect 211796 53474 211852 53530
rect 211892 51846 211948 51902
rect 212084 45334 212140 45390
rect 211700 45038 211756 45094
rect 212660 51994 212716 52050
rect 212948 53326 213004 53382
rect 213140 44890 213196 44946
rect 214868 53474 214924 53530
rect 215204 53585 215260 53641
rect 215060 44742 215116 44798
rect 216692 53030 216748 53086
rect 217028 53585 217084 53641
rect 220628 54362 220684 54418
rect 219956 48738 220012 48794
rect 229652 53918 229708 53974
rect 221108 53178 221164 53234
rect 220724 47702 220780 47758
rect 221876 52586 221932 52642
rect 222548 52438 222604 52494
rect 223316 52142 223372 52198
rect 223700 52290 223756 52346
rect 229652 53326 229708 53382
rect 237236 51254 237292 51310
rect 237812 51106 237868 51162
rect 238196 50810 238252 50866
rect 239444 48146 239500 48202
rect 240020 47998 240076 48054
rect 242228 48442 242284 48498
rect 241652 47850 241708 47906
rect 242996 48590 243052 48646
rect 243476 50958 243532 51014
rect 354260 53195 354316 53234
rect 354260 53178 354262 53195
rect 354262 53178 354314 53195
rect 354314 53178 354316 53195
rect 374324 52882 374380 52938
rect 362900 51550 362956 51606
rect 302420 48886 302476 48942
rect 243380 48294 243436 48350
rect 242612 47554 242668 47610
rect 423284 53343 423340 53382
rect 423284 53326 423286 53343
rect 423286 53326 423338 53343
rect 423338 53326 423340 53343
rect 443444 53326 443500 53382
rect 434900 51715 434956 51754
rect 434900 51698 434902 51715
rect 434902 51698 434954 51715
rect 434954 51698 434956 51715
rect 459284 51698 459340 51754
rect 382964 51550 383020 51606
rect 403220 51550 403276 51606
rect 423284 51550 423340 51606
rect 489620 51589 489622 51606
rect 489622 51589 489674 51606
rect 489674 51589 489676 51606
rect 489620 51550 489676 51589
rect 509588 51550 509644 51606
rect 353588 46074 353644 46130
rect 215348 44594 215404 44650
rect 302516 43262 302572 43318
rect 361748 43262 361804 43318
rect 364916 43262 364972 43318
rect 306740 42078 306796 42134
rect 357140 42078 357196 42134
rect 410804 43262 410860 43318
rect 408884 42078 408940 42134
rect 416276 42078 416332 42134
rect 210740 40746 210796 40802
rect 518804 44742 518860 44798
rect 650036 892782 650092 892838
rect 649940 846162 649996 846218
rect 650228 705414 650284 705470
rect 645236 231666 645292 231722
rect 645140 231074 645196 231130
rect 601940 51715 601996 51754
rect 601940 51698 601942 51715
rect 601942 51698 601994 51715
rect 601994 51698 601996 51715
rect 622004 51698 622060 51754
rect 529268 44594 529324 44650
rect 463700 41782 463756 41838
rect 465716 41782 465772 41838
rect 655124 974626 655180 974682
rect 654356 951094 654412 951150
rect 655220 962786 655276 962842
rect 653780 939402 653836 939458
rect 675380 966338 675436 966394
rect 675764 965746 675820 965802
rect 675764 965006 675820 965062
rect 675380 963230 675436 963286
rect 675476 962638 675532 962694
rect 675380 962194 675436 962250
rect 675764 961306 675820 961362
rect 675668 960714 675724 960770
rect 675476 960122 675532 960178
rect 654452 927562 654508 927618
rect 654452 915887 654508 915926
rect 654452 915870 654454 915887
rect 654454 915870 654506 915887
rect 654506 915870 654508 915887
rect 654452 904178 654508 904234
rect 654452 880646 654508 880702
rect 654452 868954 654508 869010
rect 654452 857262 654508 857318
rect 654452 833730 654508 833786
rect 654452 822038 654508 822094
rect 654452 810346 654508 810402
rect 653780 798654 653836 798710
rect 654452 786814 654508 786870
rect 654452 775122 654508 775178
rect 654452 763299 654508 763338
rect 654452 763282 654454 763299
rect 654454 763282 654506 763299
rect 654506 763282 654508 763299
rect 654452 739898 654508 739954
rect 655220 728206 655276 728262
rect 654452 716366 654508 716422
rect 654452 692982 654508 693038
rect 654452 669450 654508 669506
rect 652244 658498 652300 658554
rect 654452 646066 654508 646122
rect 654452 610990 654508 611046
rect 654452 599150 654508 599206
rect 655124 587310 655180 587366
rect 654452 575618 654508 575674
rect 654452 564074 654508 564130
rect 654452 552234 654508 552290
rect 654452 540394 654508 540450
rect 654452 528702 654508 528758
rect 654068 517158 654124 517214
rect 654932 505318 654988 505374
rect 654452 481786 654508 481842
rect 654452 470242 654508 470298
rect 654452 446562 654508 446618
rect 654452 434909 654454 434926
rect 654454 434909 654506 434926
rect 654506 434909 654508 434926
rect 654452 434870 654508 434909
rect 654452 423343 654508 423382
rect 654452 423326 654454 423343
rect 654454 423326 654506 423343
rect 654506 423326 654508 423343
rect 654452 411338 654508 411394
rect 655412 681290 655468 681346
rect 655316 634374 655372 634430
rect 656372 622534 656428 622590
rect 655220 493478 655276 493534
rect 654644 399646 654700 399702
rect 654452 387954 654508 388010
rect 654452 376410 654508 376466
rect 654452 364422 654508 364478
rect 654452 341038 654508 341094
rect 654068 329494 654124 329550
rect 656372 458402 656428 458458
rect 655316 352730 655372 352786
rect 655124 317506 655180 317562
rect 654452 282578 654508 282634
rect 645716 232702 645772 232758
rect 645524 232258 645580 232314
rect 645332 230482 645388 230538
rect 646100 210946 646156 211002
rect 646196 166842 646252 166898
rect 645908 166398 645964 166454
rect 647924 165806 647980 165862
rect 655220 305814 655276 305870
rect 655412 294122 655468 294178
rect 670964 583166 671020 583222
rect 673940 937182 673996 937238
rect 675380 957606 675436 957662
rect 675092 953462 675148 953518
rect 675476 955978 675532 956034
rect 675188 953314 675244 953370
rect 674708 945322 674764 945378
rect 674708 944730 674764 944786
rect 674612 943990 674668 944046
rect 674804 943250 674860 943306
rect 674708 942379 674764 942418
rect 674708 942362 674710 942379
rect 674710 942362 674762 942379
rect 674762 942362 674764 942379
rect 674708 942066 674764 942122
rect 674708 940734 674764 940790
rect 674132 939550 674188 939606
rect 674036 936294 674092 936350
rect 679796 928598 679852 928654
rect 679796 928006 679852 928062
rect 675092 876354 675148 876410
rect 675764 876354 675820 876410
rect 675092 876206 675148 876262
rect 675284 875762 675340 875818
rect 675188 875614 675244 875670
rect 672692 718438 672748 718494
rect 675476 873986 675532 874042
rect 675380 873394 675436 873450
rect 675380 872802 675436 872858
rect 675380 869842 675436 869898
rect 675380 866882 675436 866938
rect 675668 864662 675724 864718
rect 675476 862886 675532 862942
rect 674804 826626 674860 826682
rect 674900 826478 674956 826534
rect 674228 780450 674284 780506
rect 673748 764170 673804 764226
rect 673652 751590 673708 751646
rect 673748 720510 673804 720566
rect 673652 718438 673708 718494
rect 674036 714442 674092 714498
rect 674036 679514 674092 679570
rect 672692 673298 672748 673354
rect 674036 670338 674092 670394
rect 674228 716070 674284 716126
rect 674420 772606 674476 772662
rect 674420 767465 674422 767482
rect 674422 767465 674474 767482
rect 674474 767465 674476 767482
rect 674420 767426 674476 767465
rect 674420 765837 674422 765854
rect 674422 765837 674474 765854
rect 674474 765837 674476 765854
rect 674420 765798 674476 765837
rect 675764 787850 675820 787906
rect 675476 787406 675532 787462
rect 675764 786666 675820 786722
rect 674708 777342 674764 777398
rect 674708 766873 674710 766890
rect 674710 766873 674762 766890
rect 674762 766873 674764 766890
rect 674708 766834 674764 766873
rect 674708 765245 674710 765262
rect 674710 765245 674762 765262
rect 674762 765245 674764 765262
rect 674708 765206 674764 765245
rect 674708 763299 674764 763338
rect 674708 763282 674710 763299
rect 674710 763282 674762 763299
rect 674762 763282 674764 763299
rect 674708 762559 674764 762598
rect 674708 762542 674710 762559
rect 674710 762542 674762 762559
rect 674762 762542 674764 762559
rect 675764 784150 675820 784206
rect 675764 781930 675820 781986
rect 674996 777490 675052 777546
rect 679700 750110 679756 750166
rect 679700 749518 679756 749574
rect 675092 743302 675148 743358
rect 675092 742118 675148 742174
rect 675092 740194 675148 740250
rect 675380 740046 675436 740102
rect 675476 739158 675532 739214
rect 675764 738714 675820 738770
rect 674420 722473 674422 722490
rect 674422 722473 674474 722490
rect 674474 722473 674476 722490
rect 674420 722434 674476 722473
rect 674420 721733 674422 721750
rect 674422 721733 674474 721750
rect 674474 721733 674476 721750
rect 674420 721694 674476 721733
rect 674420 720845 674422 720862
rect 674422 720845 674474 720862
rect 674474 720845 674476 720862
rect 674420 720806 674476 720845
rect 674420 719195 674476 719234
rect 674420 719178 674422 719195
rect 674422 719178 674474 719195
rect 674474 719178 674476 719195
rect 674420 717715 674476 717754
rect 674420 717698 674422 717715
rect 674422 717698 674474 717715
rect 674474 717698 674476 717715
rect 674324 712962 674380 713018
rect 674420 710485 674422 710502
rect 674422 710485 674474 710502
rect 674474 710485 674476 710502
rect 674420 710446 674476 710485
rect 674420 709005 674422 709022
rect 674422 709005 674474 709022
rect 674474 709005 674476 709022
rect 674420 708966 674476 709005
rect 674420 707377 674422 707394
rect 674422 707377 674474 707394
rect 674474 707377 674476 707394
rect 674420 707338 674476 707377
rect 674132 664418 674188 664474
rect 674132 630674 674188 630730
rect 673844 629786 673900 629842
rect 673844 629046 673900 629102
rect 673844 628306 673900 628362
rect 674420 679662 674476 679718
rect 674420 677333 674422 677350
rect 674422 677333 674474 677350
rect 674474 677333 674476 677350
rect 674420 677294 674476 677333
rect 674420 676445 674422 676462
rect 674422 676445 674474 676462
rect 674474 676445 674476 676462
rect 674420 676406 674476 676445
rect 674420 675705 674422 675722
rect 674422 675705 674474 675722
rect 674474 675705 674476 675722
rect 674420 675666 674476 675705
rect 674420 674817 674422 674834
rect 674422 674817 674474 674834
rect 674474 674817 674476 674834
rect 674420 674778 674476 674817
rect 674420 674055 674476 674094
rect 674420 674038 674422 674055
rect 674422 674038 674474 674055
rect 674474 674038 674476 674055
rect 674516 668710 674572 668766
rect 674804 709893 674806 709910
rect 674806 709893 674858 709910
rect 674858 709893 674860 709910
rect 674804 709854 674860 709893
rect 674804 706785 674806 706802
rect 674806 706785 674858 706802
rect 674858 706785 674860 706802
rect 674804 706746 674860 706785
rect 675764 737678 675820 737734
rect 675764 734866 675820 734922
rect 675380 734126 675436 734182
rect 674996 713998 675052 714054
rect 679700 705118 679756 705174
rect 679700 704526 679756 704582
rect 674996 702454 675052 702510
rect 674900 688246 674956 688302
rect 674708 671078 674764 671134
rect 674612 667970 674668 668026
rect 674420 661349 674422 661366
rect 674422 661349 674474 661366
rect 674474 661349 674476 661366
rect 674420 661310 674476 661349
rect 674324 623570 674380 623626
rect 674420 622682 674476 622738
rect 674228 619426 674284 619482
rect 673844 617946 673900 618002
rect 673844 616318 673900 616374
rect 674708 632489 674710 632506
rect 674710 632489 674762 632506
rect 674762 632489 674764 632506
rect 674708 632450 674764 632489
rect 674708 631749 674710 631766
rect 674710 631749 674762 631766
rect 674762 631749 674764 631766
rect 674708 631710 674764 631749
rect 675380 697866 675436 697922
rect 675476 697274 675532 697330
rect 675764 697126 675820 697182
rect 675476 694758 675532 694814
rect 675284 694314 675340 694370
rect 675764 694314 675820 694370
rect 675476 693426 675532 693482
rect 675380 691946 675436 692002
rect 675092 685582 675148 685638
rect 674996 679662 675052 679718
rect 674996 679514 675052 679570
rect 675860 679514 675916 679570
rect 675188 672262 675244 672318
rect 674996 671522 675052 671578
rect 675092 671226 675148 671282
rect 675092 670634 675148 670690
rect 675860 670634 675916 670690
rect 679700 659978 679756 660034
rect 679700 659238 679756 659294
rect 675764 652578 675820 652634
rect 675476 652134 675532 652190
rect 675476 651394 675532 651450
rect 675188 650950 675244 651006
rect 675764 649618 675820 649674
rect 675188 647990 675244 648046
rect 675476 645326 675532 645382
rect 675764 640294 675820 640350
rect 675380 638518 675436 638574
rect 675188 628010 675244 628066
rect 674804 626086 674860 626142
rect 679700 614986 679756 615042
rect 679700 614394 679756 614450
rect 675092 607734 675148 607790
rect 675092 607438 675148 607494
rect 675476 606402 675532 606458
rect 674900 604922 674956 604978
rect 674708 604774 674764 604830
rect 675092 604774 675148 604830
rect 675764 600186 675820 600242
rect 675764 595302 675820 595358
rect 675764 593378 675820 593434
rect 674708 586422 674764 586478
rect 674420 586313 674422 586330
rect 674422 586313 674474 586330
rect 674474 586313 674476 586330
rect 674420 586274 674476 586313
rect 674420 585425 674422 585442
rect 674422 585425 674474 585442
rect 674474 585425 674476 585442
rect 674420 585386 674476 585425
rect 674612 584833 674614 584850
rect 674614 584833 674666 584850
rect 674666 584833 674668 584850
rect 674612 584794 674668 584833
rect 674708 583627 674764 583666
rect 674708 583610 674710 583627
rect 674710 583610 674762 583627
rect 674762 583610 674764 583627
rect 674420 583166 674476 583222
rect 676820 582591 676876 582630
rect 676820 582574 676822 582591
rect 676822 582574 676874 582591
rect 676874 582574 676876 582591
rect 674420 578874 674476 578930
rect 674708 575361 674710 575378
rect 674710 575361 674762 575378
rect 674762 575361 674764 575378
rect 674708 575322 674764 575361
rect 674708 574473 674710 574490
rect 674710 574473 674762 574490
rect 674762 574473 674764 574490
rect 674708 574434 674764 574473
rect 674420 573585 674422 573602
rect 674422 573585 674474 573602
rect 674474 573585 674476 573602
rect 674420 573546 674476 573585
rect 674708 572993 674710 573010
rect 674710 572993 674762 573010
rect 674762 572993 674764 573010
rect 674708 572954 674764 572993
rect 674420 571957 674422 571974
rect 674422 571957 674474 571974
rect 674474 571957 674476 571974
rect 674420 571918 674476 571957
rect 674708 571365 674710 571382
rect 674710 571365 674762 571382
rect 674762 571365 674764 571382
rect 674708 571326 674764 571365
rect 679796 569698 679852 569754
rect 679796 569106 679852 569162
rect 674228 541321 674230 541338
rect 674230 541321 674282 541338
rect 674282 541321 674284 541338
rect 674228 541282 674284 541321
rect 674228 540433 674230 540450
rect 674230 540433 674282 540450
rect 674282 540433 674284 540450
rect 674228 540394 674284 540433
rect 673844 539654 673900 539710
rect 673748 530922 673804 530978
rect 673844 530034 673900 530090
rect 673844 529294 673900 529350
rect 673844 528554 673900 528610
rect 673172 527814 673228 527870
rect 673844 526943 673900 526982
rect 673844 526926 673846 526943
rect 673846 526926 673898 526943
rect 673898 526926 673900 526943
rect 673844 526186 673900 526242
rect 673940 486078 673996 486134
rect 675284 562890 675340 562946
rect 675092 561706 675148 561762
rect 675284 561558 675340 561614
rect 675476 558894 675532 558950
rect 675380 557710 675436 557766
rect 674324 490074 674380 490130
rect 674516 497513 674518 497530
rect 674518 497513 674570 497530
rect 674570 497513 674572 497530
rect 674516 497474 674572 497513
rect 674516 496625 674518 496642
rect 674518 496625 674570 496642
rect 674570 496625 674572 496642
rect 674516 496586 674572 496625
rect 674420 489334 674476 489390
rect 674708 541578 674764 541634
rect 674996 550162 675052 550218
rect 676532 547054 676588 547110
rect 676628 546906 676684 546962
rect 676532 537878 676588 537934
rect 674708 497770 674764 497826
rect 674804 491850 674860 491906
rect 674612 488742 674668 488798
rect 674228 485264 674284 485320
rect 674132 484598 674188 484654
rect 674036 482970 674092 483026
rect 676724 538618 676780 538674
rect 676628 537138 676684 537194
rect 676532 493922 676588 493978
rect 674900 482378 674956 482434
rect 679796 524706 679852 524762
rect 679796 524114 679852 524170
rect 676724 495846 676780 495902
rect 676724 494514 676780 494570
rect 676628 493034 676684 493090
rect 676532 412078 676588 412134
rect 676628 411930 676684 411986
rect 674708 409266 674764 409322
rect 674420 409044 674476 409100
rect 674708 408417 674710 408434
rect 674710 408417 674762 408434
rect 674762 408417 674764 408434
rect 674708 408378 674764 408417
rect 679796 480750 679852 480806
rect 679796 480010 679852 480066
rect 676724 407638 676780 407694
rect 673844 406602 673900 406658
rect 674900 404086 674956 404142
rect 674036 401866 674092 401922
rect 673940 397130 673996 397186
rect 674516 397722 674572 397778
rect 674420 396390 674476 396446
rect 674324 393948 674380 394004
rect 674804 395354 674860 395410
rect 674708 394466 674764 394522
rect 675284 402458 675340 402514
rect 675188 399350 675244 399406
rect 674996 398462 675052 398518
rect 679700 392542 679756 392598
rect 679700 392098 679756 392154
rect 675092 374486 675148 374542
rect 675476 378778 675532 378834
rect 675476 373894 675532 373950
rect 675380 371970 675436 372026
rect 675188 371674 675244 371730
rect 674708 364905 674710 364922
rect 674710 364905 674762 364922
rect 674762 364905 674764 364922
rect 674708 364866 674764 364905
rect 674420 363869 674422 363886
rect 674422 363869 674474 363886
rect 674474 363869 674476 363886
rect 674420 363830 674476 363869
rect 674708 363277 674710 363294
rect 674710 363277 674762 363294
rect 674762 363277 674764 363294
rect 674708 363238 674764 363277
rect 673844 362202 673900 362258
rect 674036 359094 674092 359150
rect 677108 358058 677164 358114
rect 674612 357170 674668 357226
rect 674516 352434 674572 352490
rect 674228 351250 674284 351306
rect 674132 348734 674188 348790
rect 674324 349548 674380 349604
rect 675188 356430 675244 356486
rect 675092 353322 675148 353378
rect 674804 350214 674860 350270
rect 676916 355690 676972 355746
rect 675284 354062 675340 354118
rect 676820 351694 676876 351750
rect 677012 354950 677068 355006
rect 676916 345330 676972 345386
rect 679796 347402 679852 347458
rect 679796 346662 679852 346718
rect 677108 345478 677164 345534
rect 677012 345182 677068 345238
rect 676820 344442 676876 344498
rect 675284 334970 675340 335026
rect 675572 333786 675628 333842
rect 675764 333490 675820 333546
rect 675764 330530 675820 330586
rect 675188 329494 675244 329550
rect 675764 328014 675820 328070
rect 675764 326830 675820 326886
rect 674420 319691 674422 319708
rect 674422 319691 674474 319708
rect 674474 319691 674476 319708
rect 674420 319652 674476 319691
rect 674420 318877 674422 318894
rect 674422 318877 674474 318894
rect 674474 318877 674476 318894
rect 674420 318838 674476 318877
rect 674708 318285 674710 318302
rect 674710 318285 674762 318302
rect 674762 318285 674764 318302
rect 674708 318246 674764 318285
rect 673940 314102 673996 314158
rect 674324 312474 674380 312530
rect 674228 304556 674284 304612
rect 674132 303742 674188 303798
rect 677108 311438 677164 311494
rect 676916 310698 676972 310754
rect 674516 309070 674572 309126
rect 674420 305370 674476 305426
rect 675092 308330 675148 308386
rect 674996 307442 675052 307498
rect 676820 305962 676876 306018
rect 677012 306702 677068 306758
rect 677012 299450 677068 299506
rect 677204 309958 677260 310014
rect 679796 302410 679852 302466
rect 679796 301670 679852 301726
rect 677204 299302 677260 299358
rect 675284 289978 675340 290034
rect 675476 289534 675532 289590
rect 674996 284946 675052 285002
rect 675668 285242 675724 285298
rect 674132 284798 674188 284854
rect 675092 284798 675148 284854
rect 675380 283614 675436 283670
rect 675764 281838 675820 281894
rect 674132 275326 674188 275382
rect 674708 274921 674710 274938
rect 674710 274921 674762 274938
rect 674762 274921 674764 274938
rect 674708 274882 674764 274921
rect 674132 273994 674188 274050
rect 674708 274033 674710 274050
rect 674710 274033 674762 274050
rect 674762 274033 674764 274050
rect 674708 273994 674764 274033
rect 674708 273293 674710 273310
rect 674710 273293 674762 273310
rect 674762 273293 674764 273310
rect 674708 273254 674764 273293
rect 673940 267482 673996 267538
rect 678260 266446 678316 266502
rect 678164 265706 678220 265762
rect 674612 264078 674668 264134
rect 674324 263486 674380 263542
rect 674132 258750 674188 258806
rect 674420 262746 674476 262802
rect 676916 261710 676972 261766
rect 676820 260970 676876 261026
rect 674708 259786 674764 259842
rect 675092 259342 675148 259398
rect 678356 264966 678412 265022
rect 679796 257418 679852 257474
rect 679796 256826 679852 256882
rect 678356 253570 678412 253626
rect 678164 253422 678220 253478
rect 675284 250462 675340 250518
rect 675764 245134 675820 245190
rect 675092 244986 675148 245042
rect 675188 244246 675244 244302
rect 675092 241286 675148 241342
rect 674612 239231 674668 239270
rect 674612 239214 674614 239231
rect 674614 239214 674666 239231
rect 674666 239214 674668 239231
rect 674996 239214 675052 239270
rect 675764 243506 675820 243562
rect 675188 238918 675244 238974
rect 675476 238622 675532 238678
rect 675764 236846 675820 236902
rect 674420 229485 674422 229502
rect 674422 229485 674474 229502
rect 674474 229485 674476 229502
rect 674420 229446 674476 229485
rect 674708 228893 674710 228910
rect 674710 228893 674762 228910
rect 674762 228893 674764 228910
rect 674708 228854 674764 228893
rect 674420 227857 674422 227874
rect 674422 227857 674474 227874
rect 674474 227857 674476 227874
rect 674420 227818 674476 227857
rect 679796 225746 679852 225802
rect 677204 223674 677260 223730
rect 674420 222194 674476 222250
rect 674324 217458 674380 217514
rect 674996 221158 675052 221214
rect 674900 214942 674956 214998
rect 674804 214202 674860 214258
rect 674708 213314 674764 213370
rect 677012 220566 677068 220622
rect 675188 218494 675244 218550
rect 675092 218050 675148 218106
rect 675284 217754 675340 217810
rect 676916 216422 676972 216478
rect 676820 215830 676876 215886
rect 675284 211686 675340 211742
rect 676916 210206 676972 210262
rect 677108 219678 677164 219734
rect 677012 210058 677068 210114
rect 677108 209910 677164 209966
rect 679700 212130 679756 212186
rect 679700 211390 679756 211446
rect 677204 209762 677260 209818
rect 679988 224858 680044 224914
rect 679796 209614 679852 209670
rect 679988 209466 680044 209522
rect 675764 204286 675820 204342
rect 675092 199698 675148 199754
rect 675188 199106 675244 199162
rect 675476 198366 675532 198422
rect 675188 195702 675244 195758
rect 675092 195554 675148 195610
rect 675764 195258 675820 195314
rect 675380 193482 675436 193538
rect 675764 191558 675820 191614
rect 674420 184454 674476 184510
rect 674708 183901 674710 183918
rect 674710 183901 674762 183918
rect 674762 183901 674764 183918
rect 674708 183862 674764 183901
rect 674420 182865 674422 182882
rect 674422 182865 674474 182882
rect 674474 182865 674476 182882
rect 674420 182826 674476 182865
rect 679700 179866 679756 179922
rect 674036 178830 674092 178886
rect 674420 177202 674476 177258
rect 674324 169358 674380 169414
rect 677012 176166 677068 176222
rect 676916 175574 676972 175630
rect 675188 173946 675244 174002
rect 674900 173058 674956 173114
rect 674516 168322 674572 168378
rect 674708 167286 674764 167342
rect 674612 166546 674668 166602
rect 674708 165658 674764 165714
rect 674996 172318 675052 172374
rect 675092 169950 675148 170006
rect 676820 170838 676876 170894
rect 675284 166398 675340 166454
rect 675284 165510 675340 165566
rect 677204 174686 677260 174742
rect 677108 171430 677164 171486
rect 676916 164030 676972 164086
rect 679796 179422 679852 179478
rect 679700 166546 679756 166602
rect 679796 166398 679852 166454
rect 677204 163882 677260 163938
rect 677108 163586 677164 163642
rect 675476 154558 675532 154614
rect 675380 154262 675436 154318
rect 675764 153374 675820 153430
rect 675764 150266 675820 150322
rect 675476 148490 675532 148546
rect 675764 146566 675820 146622
rect 674708 139018 674764 139074
rect 674420 138443 674476 138482
rect 674420 138426 674422 138443
rect 674422 138426 674474 138443
rect 674474 138426 674476 138443
rect 674612 137242 674668 137298
rect 674708 135614 674764 135670
rect 673364 134874 673420 134930
rect 674420 133690 674476 133746
rect 674132 131174 674188 131230
rect 674036 123330 674092 123386
rect 647828 121702 647884 121758
rect 647924 121149 647926 121166
rect 647926 121149 647978 121166
rect 647978 121149 647980 121166
rect 647924 121110 647980 121149
rect 647828 120666 647884 120722
rect 646484 120074 646540 120130
rect 665204 112861 665206 112878
rect 665206 112861 665258 112878
rect 665258 112861 665260 112878
rect 665204 112822 665260 112861
rect 665204 111490 665260 111546
rect 647924 104386 647980 104442
rect 674228 128066 674284 128122
rect 674324 127326 674380 127382
rect 675092 131766 675148 131822
rect 674900 124810 674956 124866
rect 674516 123922 674572 123978
rect 674804 122146 674860 122202
rect 674612 121554 674668 121610
rect 674708 121275 674764 121314
rect 674708 121258 674710 121275
rect 674710 121258 674762 121275
rect 674762 121258 674764 121275
rect 677012 130286 677068 130342
rect 675188 128658 675244 128714
rect 676916 126290 676972 126346
rect 676820 125550 676876 125606
rect 677108 129546 677164 129602
rect 677012 120370 677068 120426
rect 677108 118002 677164 118058
rect 675476 110010 675532 110066
rect 675380 109418 675436 109474
rect 675668 108086 675724 108142
rect 675380 103202 675436 103258
rect 675764 101426 675820 101482
rect 646292 88550 646348 88606
rect 646388 86922 646444 86978
rect 646100 86330 646156 86386
rect 646004 84258 646060 84314
rect 646292 83113 646294 83130
rect 646294 83113 646346 83130
rect 646346 83113 646348 83130
rect 646292 83074 646348 83113
rect 646100 82630 646156 82686
rect 646292 76414 646348 76470
rect 646100 74046 646156 74102
rect 646292 73306 646348 73362
rect 646484 84702 646540 84758
rect 646484 78930 646540 78986
rect 647252 85886 647308 85942
rect 647444 87514 647500 87570
rect 647348 81298 647404 81354
rect 646868 79818 646924 79874
rect 646868 78782 646924 78838
rect 646868 78190 646924 78246
rect 647636 89142 647692 89198
rect 647540 82038 647596 82094
rect 647924 87958 647980 88014
rect 650900 86922 650956 86978
rect 647828 85294 647884 85350
rect 650996 85294 651052 85350
rect 650996 84258 651052 84314
rect 650900 82630 650956 82686
rect 647924 81463 647980 81502
rect 647924 81446 647926 81463
rect 647926 81446 647978 81463
rect 647978 81446 647980 81463
rect 647924 80410 647980 80466
rect 647828 77598 647884 77654
rect 651188 86182 651244 86238
rect 651092 83370 651148 83426
rect 652340 83666 652396 83722
rect 647924 77154 647980 77210
rect 646676 76562 646732 76618
rect 646484 75526 646540 75582
rect 646388 73158 646444 73214
rect 662900 81150 662956 81206
rect 647924 74934 647980 74990
rect 647156 73898 647212 73954
rect 646676 72270 646732 72326
rect 663572 85590 663628 85646
rect 663284 85146 663340 85202
rect 663476 84702 663532 84758
rect 663380 82778 663436 82834
rect 663284 82038 663340 82094
rect 625076 40598 625132 40654
rect 141812 40302 141868 40358
rect 457748 40302 457804 40358
<< metal3 >>
rect 251778 1019912 252990 1019972
rect 251778 1019824 251838 1019912
rect 251424 1019794 251838 1019824
rect 252930 1019794 252990 1019912
rect 251394 1019764 251838 1019794
rect 108591 1005468 108657 1005471
rect 114159 1005468 114225 1005471
rect 108591 1005466 109152 1005468
rect 108591 1005410 108596 1005466
rect 108652 1005410 109152 1005466
rect 108591 1005408 109152 1005410
rect 114159 1005466 114720 1005468
rect 114159 1005410 114164 1005466
rect 114220 1005410 114720 1005466
rect 114159 1005408 114720 1005410
rect 108591 1005405 108657 1005408
rect 114159 1005405 114225 1005408
rect 217263 1005320 217329 1005323
rect 216672 1005318 217329 1005320
rect 216672 1005262 217268 1005318
rect 217324 1005262 217329 1005318
rect 216672 1005260 217329 1005262
rect 217263 1005257 217329 1005260
rect 218895 1005320 218961 1005323
rect 223119 1005320 223185 1005323
rect 218895 1005318 223185 1005320
rect 218895 1005262 218900 1005318
rect 218956 1005262 223124 1005318
rect 223180 1005262 223185 1005318
rect 218895 1005260 223185 1005262
rect 218895 1005257 218961 1005260
rect 223119 1005257 223185 1005260
rect 115215 1005172 115281 1005175
rect 221871 1005172 221937 1005175
rect 115215 1005170 115488 1005172
rect 115215 1005114 115220 1005170
rect 115276 1005114 115488 1005170
rect 115215 1005112 115488 1005114
rect 218304 1005170 221937 1005172
rect 218304 1005114 221876 1005170
rect 221932 1005114 221937 1005170
rect 218304 1005112 221937 1005114
rect 115215 1005109 115281 1005112
rect 221871 1005109 221937 1005112
rect 246831 1005172 246897 1005175
rect 251394 1005172 251454 1019764
rect 308751 1005468 308817 1005471
rect 321039 1005468 321105 1005471
rect 308751 1005466 309312 1005468
rect 308751 1005410 308756 1005466
rect 308812 1005410 309312 1005466
rect 308751 1005408 309312 1005410
rect 320448 1005466 321105 1005468
rect 320448 1005410 321044 1005466
rect 321100 1005410 321105 1005466
rect 320448 1005408 321105 1005410
rect 308751 1005405 308817 1005408
rect 321039 1005405 321105 1005408
rect 321423 1005468 321489 1005471
rect 325455 1005468 325521 1005471
rect 357903 1005468 357969 1005471
rect 364143 1005468 364209 1005471
rect 365007 1005468 365073 1005471
rect 430863 1005468 430929 1005471
rect 501135 1005468 501201 1005471
rect 321423 1005466 325521 1005468
rect 321423 1005410 321428 1005466
rect 321484 1005410 325460 1005466
rect 325516 1005410 325521 1005466
rect 321423 1005408 325521 1005410
rect 357408 1005466 357969 1005468
rect 357408 1005410 357908 1005466
rect 357964 1005410 357969 1005466
rect 357408 1005408 357969 1005410
rect 363648 1005466 364209 1005468
rect 363648 1005410 364148 1005466
rect 364204 1005410 364209 1005466
rect 363648 1005408 364209 1005410
rect 364512 1005466 365073 1005468
rect 364512 1005410 365012 1005466
rect 365068 1005410 365073 1005466
rect 364512 1005408 365073 1005410
rect 430368 1005466 430929 1005468
rect 430368 1005410 430868 1005466
rect 430924 1005410 430929 1005466
rect 430368 1005408 430929 1005410
rect 501024 1005466 501201 1005468
rect 501024 1005410 501140 1005466
rect 501196 1005410 501201 1005466
rect 501024 1005408 501201 1005410
rect 321423 1005405 321489 1005408
rect 325455 1005405 325521 1005408
rect 357903 1005405 357969 1005408
rect 364143 1005405 364209 1005408
rect 365007 1005405 365073 1005408
rect 430863 1005405 430929 1005408
rect 501135 1005405 501201 1005408
rect 307983 1005320 308049 1005323
rect 309615 1005320 309681 1005323
rect 318639 1005320 318705 1005323
rect 365775 1005320 365841 1005323
rect 366735 1005320 366801 1005323
rect 424527 1005320 424593 1005323
rect 425295 1005320 425361 1005323
rect 307983 1005318 308448 1005320
rect 307983 1005262 307988 1005318
rect 308044 1005262 308448 1005318
rect 307983 1005260 308448 1005262
rect 309615 1005318 310176 1005320
rect 309615 1005262 309620 1005318
rect 309676 1005262 310176 1005318
rect 309615 1005260 310176 1005262
rect 318048 1005318 318705 1005320
rect 318048 1005262 318644 1005318
rect 318700 1005262 318705 1005318
rect 318048 1005260 318705 1005262
rect 365280 1005318 365841 1005320
rect 365280 1005262 365780 1005318
rect 365836 1005262 365841 1005318
rect 365280 1005260 365841 1005262
rect 366048 1005318 366801 1005320
rect 366048 1005262 366740 1005318
rect 366796 1005262 366801 1005318
rect 366048 1005260 366801 1005262
rect 424032 1005318 424593 1005320
rect 424032 1005262 424532 1005318
rect 424588 1005262 424593 1005318
rect 424032 1005260 424593 1005262
rect 424800 1005318 425361 1005320
rect 424800 1005262 425300 1005318
rect 425356 1005262 425361 1005318
rect 424800 1005260 425361 1005262
rect 307983 1005257 308049 1005260
rect 309615 1005257 309681 1005260
rect 318639 1005257 318705 1005260
rect 365775 1005257 365841 1005260
rect 366735 1005257 366801 1005260
rect 424527 1005257 424593 1005260
rect 425295 1005257 425361 1005260
rect 430767 1005320 430833 1005323
rect 504591 1005320 504657 1005323
rect 554511 1005320 554577 1005323
rect 555759 1005320 555825 1005323
rect 430767 1005318 431040 1005320
rect 430767 1005262 430772 1005318
rect 430828 1005262 431040 1005318
rect 430767 1005260 431040 1005262
rect 504096 1005318 504657 1005320
rect 504096 1005262 504596 1005318
rect 504652 1005262 504657 1005318
rect 504096 1005260 504657 1005262
rect 554016 1005318 554577 1005320
rect 554016 1005262 554516 1005318
rect 554572 1005262 554577 1005318
rect 554016 1005260 554577 1005262
rect 555552 1005318 555825 1005320
rect 555552 1005262 555764 1005318
rect 555820 1005262 555825 1005318
rect 555552 1005260 555825 1005262
rect 430767 1005257 430833 1005260
rect 504591 1005257 504657 1005260
rect 554511 1005257 554577 1005260
rect 555759 1005257 555825 1005260
rect 246831 1005170 251454 1005172
rect 246831 1005114 246836 1005170
rect 246892 1005142 251454 1005170
rect 315183 1005172 315249 1005175
rect 363471 1005172 363537 1005175
rect 426063 1005172 426129 1005175
rect 433167 1005172 433233 1005175
rect 435567 1005172 435633 1005175
rect 500751 1005172 500817 1005175
rect 553743 1005172 553809 1005175
rect 315183 1005170 315744 1005172
rect 246892 1005114 251424 1005142
rect 246831 1005112 251424 1005114
rect 315183 1005114 315188 1005170
rect 315244 1005114 315744 1005170
rect 315183 1005112 315744 1005114
rect 362976 1005170 363537 1005172
rect 362976 1005114 363476 1005170
rect 363532 1005114 363537 1005170
rect 362976 1005112 363537 1005114
rect 425568 1005170 426129 1005172
rect 425568 1005114 426068 1005170
rect 426124 1005114 426129 1005170
rect 425568 1005112 426129 1005114
rect 432672 1005170 433233 1005172
rect 432672 1005114 433172 1005170
rect 433228 1005114 433233 1005170
rect 432672 1005112 433233 1005114
rect 435168 1005170 435633 1005172
rect 435168 1005114 435572 1005170
rect 435628 1005114 435633 1005170
rect 435168 1005112 435633 1005114
rect 500160 1005170 500817 1005172
rect 500160 1005114 500756 1005170
rect 500812 1005114 500817 1005170
rect 500160 1005112 500817 1005114
rect 553248 1005170 553809 1005172
rect 553248 1005114 553748 1005170
rect 553804 1005114 553809 1005170
rect 553248 1005112 553809 1005114
rect 246831 1005109 246897 1005112
rect 315183 1005109 315249 1005112
rect 363471 1005109 363537 1005112
rect 426063 1005109 426129 1005112
rect 433167 1005109 433233 1005112
rect 435567 1005109 435633 1005112
rect 500751 1005109 500817 1005112
rect 553743 1005109 553809 1005112
rect 359919 1003988 359985 1003991
rect 423375 1003988 423441 1003991
rect 359712 1003986 359985 1003988
rect 359712 1003930 359924 1003986
rect 359980 1003930 359985 1003986
rect 359712 1003928 359985 1003930
rect 423168 1003986 423441 1003988
rect 423168 1003930 423380 1003986
rect 423436 1003930 423441 1003986
rect 423168 1003928 423441 1003930
rect 359919 1003925 359985 1003928
rect 423375 1003925 423441 1003928
rect 358383 1003840 358449 1003843
rect 359055 1003840 359121 1003843
rect 426447 1003840 426513 1003843
rect 552591 1003840 552657 1003843
rect 556527 1003840 556593 1003843
rect 358176 1003838 358449 1003840
rect 358176 1003782 358388 1003838
rect 358444 1003782 358449 1003838
rect 358176 1003780 358449 1003782
rect 358944 1003838 359121 1003840
rect 358944 1003782 359060 1003838
rect 359116 1003782 359121 1003838
rect 358944 1003780 359121 1003782
rect 426336 1003838 426513 1003840
rect 426336 1003782 426452 1003838
rect 426508 1003782 426513 1003838
rect 426336 1003780 426513 1003782
rect 552384 1003838 552657 1003840
rect 552384 1003782 552596 1003838
rect 552652 1003782 552657 1003838
rect 552384 1003780 552657 1003782
rect 556320 1003838 556593 1003840
rect 556320 1003782 556532 1003838
rect 556588 1003782 556593 1003838
rect 556320 1003780 556593 1003782
rect 358383 1003777 358449 1003780
rect 359055 1003777 359121 1003780
rect 426447 1003777 426513 1003780
rect 552591 1003777 552657 1003780
rect 556527 1003777 556593 1003780
rect 360687 1003692 360753 1003695
rect 428079 1003692 428145 1003695
rect 551727 1003692 551793 1003695
rect 360480 1003690 360753 1003692
rect 360480 1003634 360692 1003690
rect 360748 1003634 360753 1003690
rect 360480 1003632 360753 1003634
rect 427872 1003690 428145 1003692
rect 427872 1003634 428084 1003690
rect 428140 1003634 428145 1003690
rect 427872 1003632 428145 1003634
rect 551520 1003690 551793 1003692
rect 551520 1003634 551732 1003690
rect 551788 1003634 551793 1003690
rect 551520 1003632 551793 1003634
rect 360687 1003629 360753 1003632
rect 428079 1003629 428145 1003632
rect 551727 1003629 551793 1003632
rect 559215 1002656 559281 1002659
rect 559983 1002656 560049 1002659
rect 558816 1002654 559281 1002656
rect 558816 1002598 559220 1002654
rect 559276 1002598 559281 1002654
rect 558816 1002596 559281 1002598
rect 559488 1002654 560049 1002656
rect 559488 1002598 559988 1002654
rect 560044 1002598 560049 1002654
rect 559488 1002596 560049 1002598
rect 559215 1002593 559281 1002596
rect 559983 1002593 560049 1002596
rect 150351 1002508 150417 1002511
rect 254031 1002508 254097 1002511
rect 305583 1002508 305649 1002511
rect 307599 1002508 307665 1002511
rect 502767 1002508 502833 1002511
rect 503439 1002508 503505 1002511
rect 562191 1002508 562257 1002511
rect 564591 1002508 564657 1002511
rect 150351 1002506 151008 1002508
rect 150351 1002450 150356 1002506
rect 150412 1002450 151008 1002506
rect 150351 1002448 151008 1002450
rect 254031 1002506 254592 1002508
rect 254031 1002450 254036 1002506
rect 254092 1002450 254592 1002506
rect 254031 1002448 254592 1002450
rect 305583 1002506 306144 1002508
rect 305583 1002450 305588 1002506
rect 305644 1002450 306144 1002506
rect 305583 1002448 306144 1002450
rect 307599 1002506 307872 1002508
rect 307599 1002450 307604 1002506
rect 307660 1002450 307872 1002506
rect 307599 1002448 307872 1002450
rect 502560 1002506 502833 1002508
rect 502560 1002450 502772 1002506
rect 502828 1002450 502833 1002506
rect 502560 1002448 502833 1002450
rect 503328 1002506 503505 1002508
rect 503328 1002450 503444 1002506
rect 503500 1002450 503505 1002506
rect 503328 1002448 503505 1002450
rect 561888 1002506 562257 1002508
rect 561888 1002450 562196 1002506
rect 562252 1002450 562257 1002506
rect 561888 1002448 562257 1002450
rect 564192 1002506 564657 1002508
rect 564192 1002450 564596 1002506
rect 564652 1002450 564657 1002506
rect 564192 1002448 564657 1002450
rect 150351 1002445 150417 1002448
rect 254031 1002445 254097 1002448
rect 305583 1002445 305649 1002448
rect 307599 1002445 307665 1002448
rect 502767 1002445 502833 1002448
rect 503439 1002445 503505 1002448
rect 562191 1002445 562257 1002448
rect 564591 1002445 564657 1002448
rect 153615 1002360 153681 1002363
rect 253167 1002360 253233 1002363
rect 298575 1002360 298641 1002363
rect 304719 1002360 304785 1002363
rect 306543 1002360 306609 1002363
rect 505071 1002360 505137 1002363
rect 153615 1002358 154080 1002360
rect 153615 1002302 153620 1002358
rect 153676 1002302 154080 1002358
rect 153615 1002300 154080 1002302
rect 253167 1002358 253728 1002360
rect 253167 1002302 253172 1002358
rect 253228 1002302 253728 1002358
rect 253167 1002300 253728 1002302
rect 298575 1002358 303072 1002360
rect 298575 1002302 298580 1002358
rect 298636 1002330 303072 1002358
rect 304719 1002358 305376 1002360
rect 298636 1002302 303102 1002330
rect 298575 1002300 303102 1002302
rect 153615 1002297 153681 1002300
rect 253167 1002297 253233 1002300
rect 298575 1002297 298641 1002300
rect 160239 1000880 160305 1000883
rect 208431 1000880 208497 1000883
rect 160239 1000878 160512 1000880
rect 160239 1000822 160244 1000878
rect 160300 1000822 160512 1000878
rect 160239 1000820 160512 1000822
rect 208431 1000878 208800 1000880
rect 208431 1000822 208436 1000878
rect 208492 1000822 208800 1000878
rect 208431 1000820 208800 1000822
rect 160239 1000817 160305 1000820
rect 208431 1000817 208497 1000820
rect 155151 999548 155217 999551
rect 158607 999548 158673 999551
rect 263055 999548 263121 999551
rect 155151 999546 155712 999548
rect 155151 999490 155156 999546
rect 155212 999490 155712 999546
rect 155151 999488 155712 999490
rect 158607 999546 158880 999548
rect 158607 999490 158612 999546
rect 158668 999490 158880 999546
rect 158607 999488 158880 999490
rect 263055 999546 263328 999548
rect 263055 999490 263060 999546
rect 263116 999490 263328 999546
rect 263055 999488 263328 999490
rect 155151 999485 155217 999488
rect 158607 999485 158673 999488
rect 263055 999485 263121 999488
rect 156879 999400 156945 999403
rect 259599 999400 259665 999403
rect 156879 999398 157344 999400
rect 156879 999342 156884 999398
rect 156940 999342 157344 999398
rect 156879 999340 157344 999342
rect 259599 999398 260160 999400
rect 259599 999342 259604 999398
rect 259660 999342 260160 999398
rect 259599 999340 260160 999342
rect 156879 999337 156945 999340
rect 259599 999337 259665 999340
rect 205647 996588 205713 996591
rect 211695 996588 211761 996591
rect 205647 996586 206304 996588
rect 205647 996530 205652 996586
rect 205708 996530 206304 996586
rect 205647 996528 206304 996530
rect 211695 996586 211872 996588
rect 211695 996530 211700 996586
rect 211756 996530 211872 996586
rect 211695 996528 211872 996530
rect 205647 996525 205713 996528
rect 211695 996525 211761 996528
rect 162255 996292 162321 996295
rect 162144 996290 162321 996292
rect 162144 996234 162260 996290
rect 162316 996234 162321 996290
rect 162144 996232 162321 996234
rect 162255 996229 162321 996232
rect 163119 996144 163185 996147
rect 162912 996142 163185 996144
rect 162912 996086 163124 996142
rect 163180 996086 163185 996142
rect 162912 996084 163185 996086
rect 163119 996081 163185 996084
rect 203631 996144 203697 996147
rect 213327 996144 213393 996147
rect 265935 996144 266001 996147
rect 266799 996144 266865 996147
rect 203631 996142 204000 996144
rect 203631 996086 203636 996142
rect 203692 996086 204000 996142
rect 203631 996084 204000 996086
rect 213327 996142 213504 996144
rect 213327 996086 213332 996142
rect 213388 996086 213504 996142
rect 213327 996084 213504 996086
rect 265728 996142 266001 996144
rect 265728 996086 265940 996142
rect 265996 996086 266001 996142
rect 265728 996084 266001 996086
rect 266400 996142 266865 996144
rect 266400 996086 266804 996142
rect 266860 996086 266865 996142
rect 266400 996084 266865 996086
rect 203631 996081 203697 996084
rect 213327 996081 213393 996084
rect 265935 996081 266001 996084
rect 266799 996081 266865 996084
rect 100623 995996 100689 995999
rect 107247 995996 107313 995999
rect 145263 995996 145329 995999
rect 149103 995996 149169 995999
rect 100623 995994 101184 995996
rect 100623 995938 100628 995994
rect 100684 995938 101184 995994
rect 100623 995936 101184 995938
rect 107247 995994 107424 995996
rect 107247 995938 107252 995994
rect 107308 995938 107424 995994
rect 107247 995936 107424 995938
rect 145263 995994 149169 995996
rect 145263 995938 145268 995994
rect 145324 995938 149108 995994
rect 149164 995938 149169 995994
rect 145263 995936 149169 995938
rect 100623 995933 100689 995936
rect 107247 995933 107313 995936
rect 145263 995933 145329 995936
rect 149103 995933 149169 995936
rect 149487 995996 149553 995999
rect 152079 995996 152145 995999
rect 164175 995996 164241 995999
rect 164559 995996 164625 995999
rect 198543 995996 198609 995999
rect 202959 995996 203025 995999
rect 206607 995996 206673 995999
rect 215631 995996 215697 995999
rect 216879 995996 216945 995999
rect 259119 995996 259185 995999
rect 261423 995996 261489 995999
rect 261807 995996 261873 995999
rect 265071 995996 265137 995999
rect 149487 995994 150144 995996
rect 149487 995938 149492 995994
rect 149548 995938 150144 995994
rect 149487 995936 150144 995938
rect 152079 995994 152544 995996
rect 152079 995938 152084 995994
rect 152140 995938 152544 995994
rect 152079 995936 152544 995938
rect 163680 995994 164241 995996
rect 163680 995938 164180 995994
rect 164236 995938 164241 995994
rect 163680 995936 164241 995938
rect 164448 995994 164625 995996
rect 164448 995938 164564 995994
rect 164620 995938 164625 995994
rect 164448 995936 164625 995938
rect 149487 995933 149553 995936
rect 152079 995933 152145 995936
rect 164175 995933 164241 995936
rect 164559 995933 164625 995936
rect 185922 995994 198609 995996
rect 185922 995938 198548 995994
rect 198604 995938 198609 995994
rect 185922 995936 198609 995938
rect 81039 995848 81105 995851
rect 94863 995848 94929 995851
rect 81039 995846 94929 995848
rect 81039 995790 81044 995846
rect 81100 995790 94868 995846
rect 94924 995790 94929 995846
rect 99951 995848 100017 995851
rect 102159 995848 102225 995851
rect 105327 995848 105393 995851
rect 113295 995848 113361 995851
rect 99951 995846 100416 995848
rect 81039 995788 94929 995790
rect 81039 995785 81105 995788
rect 94863 995785 94929 995788
rect 85935 995700 86001 995703
rect 94959 995700 95025 995703
rect 97218 995700 97278 995818
rect 98754 995700 98814 995818
rect 85935 995698 94206 995700
rect 85935 995642 85940 995698
rect 85996 995642 94206 995698
rect 85935 995640 94206 995642
rect 85935 995637 86001 995640
rect 94146 995552 94206 995640
rect 94959 995698 98814 995700
rect 94959 995642 94964 995698
rect 95020 995642 98814 995698
rect 94959 995640 98814 995642
rect 98991 995700 99057 995703
rect 99522 995700 99582 995818
rect 99951 995790 99956 995846
rect 100012 995790 100416 995846
rect 102159 995846 102720 995848
rect 99951 995788 100416 995790
rect 99951 995785 100017 995788
rect 98991 995698 99582 995700
rect 98991 995642 98996 995698
rect 99052 995642 99582 995698
rect 98991 995640 99582 995642
rect 94959 995637 95025 995640
rect 98991 995637 99057 995640
rect 102018 995552 102078 995818
rect 102159 995790 102164 995846
rect 102220 995790 102720 995846
rect 105327 995846 105984 995848
rect 102159 995788 102720 995790
rect 102159 995785 102225 995788
rect 94146 995492 102078 995552
rect 102159 995552 102225 995555
rect 103458 995552 103518 995818
rect 102159 995550 103518 995552
rect 102159 995494 102164 995550
rect 102220 995494 103518 995550
rect 102159 995492 103518 995494
rect 102159 995489 102225 995492
rect 85359 995404 85425 995407
rect 94671 995404 94737 995407
rect 85359 995402 94737 995404
rect 85359 995346 85364 995402
rect 85420 995346 94676 995402
rect 94732 995346 94737 995402
rect 85359 995344 94737 995346
rect 85359 995341 85425 995344
rect 94671 995341 94737 995344
rect 94863 995404 94929 995407
rect 104322 995404 104382 995818
rect 94863 995402 104382 995404
rect 94863 995346 94868 995402
rect 94924 995346 104382 995402
rect 94863 995344 104382 995346
rect 94863 995341 94929 995344
rect 86415 995256 86481 995259
rect 98991 995256 99057 995259
rect 86415 995254 99057 995256
rect 86415 995198 86420 995254
rect 86476 995198 98996 995254
rect 99052 995198 99057 995254
rect 86415 995196 99057 995198
rect 86415 995193 86481 995196
rect 98991 995193 99057 995196
rect 100719 995256 100785 995259
rect 105090 995256 105150 995818
rect 105327 995790 105332 995846
rect 105388 995790 105984 995846
rect 105327 995788 105984 995790
rect 105327 995785 105393 995788
rect 100719 995254 105150 995256
rect 100719 995198 100724 995254
rect 100780 995198 105150 995254
rect 100719 995196 105150 995198
rect 106575 995256 106641 995259
rect 106722 995256 106782 995818
rect 108258 995259 108318 995818
rect 106575 995254 106782 995256
rect 106575 995198 106580 995254
rect 106636 995198 106782 995254
rect 106575 995196 106782 995198
rect 108207 995254 108318 995259
rect 108207 995198 108212 995254
rect 108268 995198 108318 995254
rect 108207 995196 108318 995198
rect 108399 995256 108465 995259
rect 109890 995256 109950 995818
rect 110688 995788 110910 995848
rect 112992 995846 113361 995848
rect 110850 995404 110910 995788
rect 111522 995552 111582 995818
rect 112194 995700 112254 995818
rect 112992 995790 113300 995846
rect 113356 995790 113361 995846
rect 112992 995788 113361 995790
rect 113295 995785 113361 995788
rect 113487 995848 113553 995851
rect 131727 995848 131793 995851
rect 144207 995848 144273 995851
rect 165615 995848 165681 995851
rect 166287 995848 166353 995851
rect 185103 995848 185169 995851
rect 185922 995848 185982 995936
rect 198543 995933 198609 995936
rect 200898 995936 201504 995996
rect 202959 995994 203232 995996
rect 202959 995938 202964 995994
rect 203020 995938 203232 995994
rect 202959 995936 203232 995938
rect 204546 995936 204768 995996
rect 206607 995994 207072 995996
rect 206607 995938 206612 995994
rect 206668 995938 207072 995994
rect 206607 995936 207072 995938
rect 215631 995994 215808 995996
rect 215631 995938 215636 995994
rect 215692 995938 215808 995994
rect 215631 995936 215808 995938
rect 216879 995994 217440 995996
rect 216879 995938 216884 995994
rect 216940 995938 217440 995994
rect 216879 995936 217440 995938
rect 259119 995994 259296 995996
rect 259119 995938 259124 995994
rect 259180 995938 259296 995994
rect 259119 995936 259296 995938
rect 261423 995994 261600 995996
rect 261423 995938 261428 995994
rect 261484 995938 261600 995994
rect 261423 995936 261600 995938
rect 261807 995994 262464 995996
rect 261807 995938 261812 995994
rect 261868 995938 262464 995994
rect 261807 995936 262464 995938
rect 264864 995994 265137 995996
rect 264864 995938 265076 995994
rect 265132 995938 265137 995994
rect 264864 995936 265137 995938
rect 113487 995846 113856 995848
rect 113487 995790 113492 995846
rect 113548 995790 113856 995846
rect 113487 995788 113856 995790
rect 131727 995846 144273 995848
rect 131727 995790 131732 995846
rect 131788 995790 144212 995846
rect 144268 995790 144273 995846
rect 131727 995788 144273 995790
rect 113487 995785 113553 995788
rect 131727 995785 131793 995788
rect 144207 995785 144273 995788
rect 120975 995700 121041 995703
rect 112194 995698 121041 995700
rect 112194 995642 120980 995698
rect 121036 995642 121041 995698
rect 112194 995640 121041 995642
rect 120975 995637 121041 995640
rect 136719 995700 136785 995703
rect 151746 995700 151806 995818
rect 136719 995698 151806 995700
rect 136719 995642 136724 995698
rect 136780 995642 151806 995698
rect 136719 995640 151806 995642
rect 136719 995637 136785 995640
rect 115215 995552 115281 995555
rect 111522 995550 115281 995552
rect 111522 995494 115220 995550
rect 115276 995494 115281 995550
rect 111522 995492 115281 995494
rect 115215 995489 115281 995492
rect 137391 995552 137457 995555
rect 153378 995552 153438 995818
rect 137391 995550 153438 995552
rect 137391 995494 137396 995550
rect 137452 995494 153438 995550
rect 137391 995492 153438 995494
rect 137391 995489 137457 995492
rect 115311 995404 115377 995407
rect 110850 995402 115377 995404
rect 110850 995346 115316 995402
rect 115372 995346 115377 995402
rect 110850 995344 115377 995346
rect 115311 995341 115377 995344
rect 133071 995404 133137 995407
rect 154914 995404 154974 995818
rect 133071 995402 154974 995404
rect 133071 995346 133076 995402
rect 133132 995346 154974 995402
rect 133071 995344 154974 995346
rect 133071 995341 133137 995344
rect 108399 995254 109950 995256
rect 108399 995198 108404 995254
rect 108460 995198 109950 995254
rect 108399 995196 109950 995198
rect 152559 995256 152625 995259
rect 156546 995256 156606 995818
rect 152559 995254 156606 995256
rect 152559 995198 152564 995254
rect 152620 995198 156606 995254
rect 152559 995196 156606 995198
rect 156687 995256 156753 995259
rect 158178 995256 158238 995818
rect 159618 995259 159678 995818
rect 161250 995259 161310 995818
rect 165216 995788 165438 995848
rect 165378 995700 165438 995788
rect 165615 995846 166080 995848
rect 165615 995790 165620 995846
rect 165676 995790 166080 995846
rect 165615 995788 166080 995790
rect 166287 995846 166944 995848
rect 166287 995790 166292 995846
rect 166348 995790 166944 995846
rect 166287 995788 166944 995790
rect 185103 995846 185982 995848
rect 185103 995790 185108 995846
rect 185164 995790 185982 995846
rect 185103 995788 185982 995790
rect 188079 995848 188145 995851
rect 198639 995848 198705 995851
rect 188079 995846 198705 995848
rect 188079 995790 188084 995846
rect 188140 995790 198644 995846
rect 198700 995790 198705 995846
rect 188079 995788 198705 995790
rect 165615 995785 165681 995788
rect 166287 995785 166353 995788
rect 185103 995785 185169 995788
rect 188079 995785 188145 995788
rect 198639 995785 198705 995788
rect 170223 995700 170289 995703
rect 165378 995698 170289 995700
rect 165378 995642 170228 995698
rect 170284 995642 170289 995698
rect 165378 995640 170289 995642
rect 170223 995637 170289 995640
rect 195375 995700 195441 995703
rect 200034 995700 200094 995818
rect 200898 995700 200958 995936
rect 202959 995933 203025 995936
rect 201807 995848 201873 995851
rect 201807 995846 202368 995848
rect 201807 995790 201812 995846
rect 201868 995790 202368 995846
rect 201807 995788 202368 995790
rect 201807 995785 201873 995788
rect 195375 995698 200958 995700
rect 195375 995642 195380 995698
rect 195436 995642 200958 995698
rect 195375 995640 200958 995642
rect 195375 995637 195441 995640
rect 189423 995552 189489 995555
rect 201807 995552 201873 995555
rect 189423 995550 201873 995552
rect 189423 995494 189428 995550
rect 189484 995494 201812 995550
rect 201868 995494 201873 995550
rect 189423 995492 201873 995494
rect 189423 995489 189489 995492
rect 201807 995489 201873 995492
rect 183759 995404 183825 995407
rect 188847 995404 188913 995407
rect 204546 995404 204606 995936
rect 206607 995933 206673 995936
rect 215631 995933 215697 995936
rect 216879 995933 216945 995936
rect 259119 995933 259185 995936
rect 261423 995933 261489 995936
rect 261807 995933 261873 995936
rect 265071 995933 265137 995936
rect 266991 995996 267057 995999
rect 299727 995996 299793 995999
rect 266991 995994 267264 995996
rect 266991 995938 266996 995994
rect 267052 995938 267264 995994
rect 266991 995936 267264 995938
rect 293442 995994 299793 995996
rect 293442 995938 299732 995994
rect 299788 995938 299793 995994
rect 293442 995936 299793 995938
rect 266991 995933 267057 995936
rect 204975 995848 205041 995851
rect 214095 995848 214161 995851
rect 239535 995848 239601 995851
rect 246447 995848 246513 995851
rect 204975 995846 205536 995848
rect 204975 995790 204980 995846
rect 205036 995790 205536 995846
rect 214095 995846 214368 995848
rect 204975 995788 205536 995790
rect 204975 995785 205041 995788
rect 206991 995700 207057 995703
rect 207906 995700 207966 995818
rect 206991 995698 207966 995700
rect 206991 995642 206996 995698
rect 207052 995642 207966 995698
rect 206991 995640 207966 995642
rect 206991 995637 207057 995640
rect 183759 995402 188670 995404
rect 183759 995346 183764 995402
rect 183820 995346 188670 995402
rect 183759 995344 188670 995346
rect 183759 995341 183825 995344
rect 156687 995254 158238 995256
rect 156687 995198 156692 995254
rect 156748 995198 158238 995254
rect 156687 995196 158238 995198
rect 159567 995254 159678 995259
rect 159567 995198 159572 995254
rect 159628 995198 159678 995254
rect 159567 995196 159678 995198
rect 161199 995254 161310 995259
rect 161199 995198 161204 995254
rect 161260 995198 161310 995254
rect 161199 995196 161310 995198
rect 100719 995193 100785 995196
rect 106575 995193 106641 995196
rect 108207 995193 108273 995196
rect 108399 995193 108465 995196
rect 152559 995193 152625 995196
rect 156687 995193 156753 995196
rect 159567 995193 159633 995196
rect 161199 995193 161265 995196
rect 82575 995108 82641 995111
rect 134223 995108 134289 995111
rect 143631 995108 143697 995111
rect 82575 995106 143697 995108
rect 82575 995050 82580 995106
rect 82636 995050 134228 995106
rect 134284 995050 143636 995106
rect 143692 995050 143697 995106
rect 82575 995048 143697 995050
rect 82575 995045 82641 995048
rect 134223 995045 134289 995048
rect 143631 995045 143697 995048
rect 188610 994960 188670 995344
rect 188847 995402 204606 995404
rect 188847 995346 188852 995402
rect 188908 995346 204606 995402
rect 188847 995344 204606 995346
rect 188847 995341 188913 995344
rect 192399 995256 192465 995259
rect 201615 995256 201681 995259
rect 192399 995254 201681 995256
rect 192399 995198 192404 995254
rect 192460 995198 201620 995254
rect 201676 995198 201681 995254
rect 192399 995196 201681 995198
rect 192399 995193 192465 995196
rect 201615 995193 201681 995196
rect 207375 995256 207441 995259
rect 209538 995256 209598 995818
rect 207375 995254 209598 995256
rect 207375 995198 207380 995254
rect 207436 995198 209598 995254
rect 207375 995196 209598 995198
rect 207375 995193 207441 995196
rect 207279 995108 207345 995111
rect 210210 995108 210270 995818
rect 211074 995259 211134 995818
rect 212706 995555 212766 995818
rect 214095 995790 214100 995846
rect 214156 995790 214368 995846
rect 239535 995846 246513 995848
rect 214095 995788 214368 995790
rect 214095 995785 214161 995788
rect 215010 995700 215070 995818
rect 239535 995790 239540 995846
rect 239596 995790 246452 995846
rect 246508 995790 246513 995846
rect 239535 995788 246513 995790
rect 239535 995785 239601 995788
rect 246447 995785 246513 995788
rect 254799 995848 254865 995851
rect 255951 995848 256017 995851
rect 260463 995848 260529 995851
rect 268623 995848 268689 995851
rect 273615 995848 273681 995851
rect 254799 995846 255456 995848
rect 254799 995790 254804 995846
rect 254860 995790 255456 995846
rect 254799 995788 255456 995790
rect 255951 995846 256224 995848
rect 255951 995790 255956 995846
rect 256012 995790 256224 995846
rect 255951 995788 256224 995790
rect 254799 995785 254865 995788
rect 255951 995785 256017 995788
rect 218895 995700 218961 995703
rect 215010 995698 218961 995700
rect 215010 995642 218900 995698
rect 218956 995642 218961 995698
rect 215010 995640 218961 995642
rect 218895 995637 218961 995640
rect 241839 995700 241905 995703
rect 256866 995700 256926 995818
rect 241839 995698 256926 995700
rect 241839 995642 241844 995698
rect 241900 995642 256926 995698
rect 241839 995640 256926 995642
rect 257538 995788 257760 995848
rect 260463 995846 261024 995848
rect 241839 995637 241905 995640
rect 212655 995550 212766 995555
rect 212655 995494 212660 995550
rect 212716 995494 212766 995550
rect 212655 995492 212766 995494
rect 240207 995552 240273 995555
rect 255951 995552 256017 995555
rect 240207 995550 256017 995552
rect 240207 995494 240212 995550
rect 240268 995494 255956 995550
rect 256012 995494 256017 995550
rect 240207 995492 256017 995494
rect 212655 995489 212721 995492
rect 240207 995489 240273 995492
rect 255951 995489 256017 995492
rect 247599 995404 247665 995407
rect 257538 995404 257598 995788
rect 247599 995402 257598 995404
rect 247599 995346 247604 995402
rect 247660 995346 257598 995402
rect 247599 995344 257598 995346
rect 247599 995341 247665 995344
rect 211023 995254 211134 995259
rect 211023 995198 211028 995254
rect 211084 995198 211134 995254
rect 211023 995196 211134 995198
rect 243567 995256 243633 995259
rect 250479 995256 250545 995259
rect 243567 995254 250545 995256
rect 243567 995198 243572 995254
rect 243628 995198 250484 995254
rect 250540 995198 250545 995254
rect 243567 995196 250545 995198
rect 211023 995193 211089 995196
rect 243567 995193 243633 995196
rect 250479 995193 250545 995196
rect 250671 995256 250737 995259
rect 258498 995256 258558 995818
rect 260463 995790 260468 995846
rect 260524 995790 261024 995846
rect 268623 995846 268896 995848
rect 260463 995788 261024 995790
rect 260463 995785 260529 995788
rect 264066 995407 264126 995818
rect 268002 995700 268062 995818
rect 268623 995790 268628 995846
rect 268684 995790 268896 995846
rect 268623 995788 268896 995790
rect 269664 995846 273681 995848
rect 269664 995790 273620 995846
rect 273676 995790 273681 995846
rect 269664 995788 273681 995790
rect 268623 995785 268689 995788
rect 273615 995785 273681 995788
rect 292431 995848 292497 995851
rect 293442 995848 293502 995936
rect 299727 995933 299793 995936
rect 292431 995846 293502 995848
rect 292431 995790 292436 995846
rect 292492 995790 293502 995846
rect 292431 995788 293502 995790
rect 293583 995848 293649 995851
rect 298287 995848 298353 995851
rect 293583 995846 298353 995848
rect 293583 995790 293588 995846
rect 293644 995790 298292 995846
rect 298348 995790 298353 995846
rect 293583 995788 298353 995790
rect 292431 995785 292497 995788
rect 293583 995785 293649 995788
rect 298287 995785 298353 995788
rect 273711 995700 273777 995703
rect 268002 995698 273777 995700
rect 268002 995642 273716 995698
rect 273772 995642 273777 995698
rect 268002 995640 273777 995642
rect 273711 995637 273777 995640
rect 291087 995700 291153 995703
rect 299535 995700 299601 995703
rect 291087 995698 299601 995700
rect 291087 995642 291092 995698
rect 291148 995642 299540 995698
rect 299596 995642 299601 995698
rect 291087 995640 299601 995642
rect 303042 995700 303102 1002300
rect 304719 1002302 304724 1002358
rect 304780 1002302 305376 1002358
rect 304719 1002300 305376 1002302
rect 306543 1002358 307008 1002360
rect 306543 1002302 306548 1002358
rect 306604 1002302 307008 1002358
rect 306543 1002300 307008 1002302
rect 504960 1002358 505137 1002360
rect 504960 1002302 505076 1002358
rect 505132 1002302 505137 1002358
rect 504960 1002300 505137 1002302
rect 304719 1002297 304785 1002300
rect 306543 1002297 306609 1002300
rect 505071 1002297 505137 1002300
rect 544239 1002360 544305 1002363
rect 560463 1002360 560529 1002363
rect 561519 1002360 561585 1002363
rect 544239 1002358 549216 1002360
rect 544239 1002302 544244 1002358
rect 544300 1002330 549216 1002358
rect 560256 1002358 560529 1002360
rect 544300 1002302 549246 1002330
rect 544239 1002300 549246 1002302
rect 560256 1002302 560468 1002358
rect 560524 1002302 560529 1002358
rect 560256 1002300 560529 1002302
rect 561120 1002358 561585 1002360
rect 561120 1002302 561524 1002358
rect 561580 1002302 561585 1002358
rect 561120 1002300 561585 1002302
rect 544239 1002297 544305 1002300
rect 511023 1001324 511089 1001327
rect 510528 1001322 511089 1001324
rect 510528 1001266 511028 1001322
rect 511084 1001266 511089 1001322
rect 510528 1001264 511089 1001266
rect 511023 1001261 511089 1001264
rect 516687 1001324 516753 1001327
rect 523599 1001324 523665 1001327
rect 516687 1001322 523665 1001324
rect 516687 1001266 516692 1001322
rect 516748 1001266 523604 1001322
rect 523660 1001266 523665 1001322
rect 516687 1001264 523665 1001266
rect 516687 1001261 516753 1001264
rect 523599 1001261 523665 1001264
rect 434127 1001176 434193 1001179
rect 433536 1001174 434193 1001176
rect 433536 1001118 434132 1001174
rect 434188 1001118 434193 1001174
rect 433536 1001116 434193 1001118
rect 434127 1001113 434193 1001116
rect 432495 1001028 432561 1001031
rect 509391 1001028 509457 1001031
rect 431904 1001026 432561 1001028
rect 431904 1000970 432500 1001026
rect 432556 1000970 432561 1001026
rect 431904 1000968 432561 1000970
rect 508896 1001026 509457 1001028
rect 508896 1000970 509396 1001026
rect 509452 1000970 509457 1001026
rect 508896 1000968 509457 1000970
rect 432495 1000965 432561 1000968
rect 509391 1000965 509457 1000968
rect 516687 1001028 516753 1001031
rect 523695 1001028 523761 1001031
rect 516687 1001026 523761 1001028
rect 516687 1000970 516692 1001026
rect 516748 1000970 523700 1001026
rect 523756 1000970 523761 1001026
rect 516687 1000968 523761 1000970
rect 516687 1000965 516753 1000968
rect 523695 1000965 523761 1000968
rect 361551 1000880 361617 1000883
rect 427311 1000880 427377 1000883
rect 428943 1000880 429009 1000883
rect 361344 1000878 361617 1000880
rect 361344 1000822 361556 1000878
rect 361612 1000822 361617 1000878
rect 361344 1000820 361617 1000822
rect 427104 1000878 427377 1000880
rect 427104 1000822 427316 1000878
rect 427372 1000822 427377 1000878
rect 427104 1000820 427377 1000822
rect 428736 1000878 429009 1000880
rect 428736 1000822 428948 1000878
rect 429004 1000822 429009 1000878
rect 428736 1000820 429009 1000822
rect 361551 1000817 361617 1000820
rect 427311 1000817 427377 1000820
rect 428943 1000817 429009 1000820
rect 507759 1000732 507825 1000735
rect 507360 1000730 507825 1000732
rect 507360 1000674 507764 1000730
rect 507820 1000674 507825 1000730
rect 507360 1000672 507825 1000674
rect 507759 1000669 507825 1000672
rect 516687 1000732 516753 1000735
rect 523503 1000732 523569 1000735
rect 516687 1000730 523569 1000732
rect 516687 1000674 516692 1000730
rect 516748 1000674 523508 1000730
rect 523564 1000674 523569 1000730
rect 516687 1000672 523569 1000674
rect 516687 1000669 516753 1000672
rect 523503 1000669 523569 1000672
rect 521583 999992 521649 999995
rect 523887 999992 523953 999995
rect 521583 999990 523953 999992
rect 521583 999934 521588 999990
rect 521644 999934 523892 999990
rect 523948 999934 523953 999990
rect 521583 999932 523953 999934
rect 521583 999929 521649 999932
rect 523887 999929 523953 999932
rect 516687 999844 516753 999847
rect 523311 999844 523377 999847
rect 516687 999842 523377 999844
rect 516687 999786 516692 999842
rect 516748 999786 523316 999842
rect 523372 999786 523377 999842
rect 516687 999784 523377 999786
rect 516687 999781 516753 999784
rect 523311 999781 523377 999784
rect 521391 999696 521457 999699
rect 523983 999696 524049 999699
rect 521391 999694 524049 999696
rect 521391 999638 521396 999694
rect 521452 999638 523988 999694
rect 524044 999638 524049 999694
rect 521391 999636 524049 999638
rect 521391 999633 521457 999636
rect 523983 999633 524049 999636
rect 311151 999548 311217 999551
rect 488847 999548 488913 999551
rect 497583 999548 497649 999551
rect 506319 999548 506385 999551
rect 311151 999546 311712 999548
rect 311151 999490 311156 999546
rect 311212 999490 311712 999546
rect 311151 999488 311712 999490
rect 488847 999546 497649 999548
rect 488847 999490 488852 999546
rect 488908 999490 497588 999546
rect 497644 999490 497649 999546
rect 488847 999488 497649 999490
rect 505728 999546 506385 999548
rect 505728 999490 506324 999546
rect 506380 999490 506385 999546
rect 505728 999488 506385 999490
rect 311151 999485 311217 999488
rect 488847 999485 488913 999488
rect 497583 999485 497649 999488
rect 506319 999485 506385 999488
rect 516783 999548 516849 999551
rect 521487 999548 521553 999551
rect 524079 999548 524145 999551
rect 516783 999546 521406 999548
rect 516783 999490 516788 999546
rect 516844 999490 521406 999546
rect 516783 999488 521406 999490
rect 516783 999485 516849 999488
rect 310287 999400 310353 999403
rect 502383 999400 502449 999403
rect 310287 999398 310944 999400
rect 310287 999342 310292 999398
rect 310348 999342 310944 999398
rect 310287 999340 310944 999342
rect 501792 999398 502449 999400
rect 501792 999342 502388 999398
rect 502444 999342 502449 999398
rect 501792 999340 502449 999342
rect 310287 999337 310353 999340
rect 502383 999337 502449 999340
rect 516687 999400 516753 999403
rect 521103 999400 521169 999403
rect 516687 999398 521169 999400
rect 516687 999342 516692 999398
rect 516748 999342 521108 999398
rect 521164 999342 521169 999398
rect 516687 999340 521169 999342
rect 521346 999400 521406 999488
rect 521487 999546 524145 999548
rect 521487 999490 521492 999546
rect 521548 999490 524084 999546
rect 524140 999490 524145 999546
rect 521487 999488 524145 999490
rect 521487 999485 521553 999488
rect 524079 999485 524145 999488
rect 523791 999400 523857 999403
rect 521346 999398 523857 999400
rect 521346 999342 523796 999398
rect 523852 999342 523857 999398
rect 521346 999340 523857 999342
rect 516687 999337 516753 999340
rect 521103 999337 521169 999340
rect 523791 999337 523857 999340
rect 356271 998068 356337 998071
rect 357039 998068 357105 998071
rect 355776 998066 356337 998068
rect 355776 998010 356276 998066
rect 356332 998010 356337 998066
rect 355776 998008 356337 998010
rect 356640 998066 357105 998068
rect 356640 998010 357044 998066
rect 357100 998010 357105 998066
rect 356640 998008 357105 998010
rect 356271 998005 356337 998008
rect 357039 998005 357105 998008
rect 367887 997920 367953 997923
rect 367776 997918 367953 997920
rect 367776 997862 367892 997918
rect 367948 997862 367953 997918
rect 367776 997860 367953 997862
rect 367887 997857 367953 997860
rect 369039 997920 369105 997923
rect 369039 997918 369216 997920
rect 369039 997862 369044 997918
rect 369100 997862 369216 997918
rect 369039 997860 369216 997862
rect 369039 997857 369105 997860
rect 508623 996588 508689 996591
rect 510255 996588 510321 996591
rect 508032 996586 508689 996588
rect 508032 996530 508628 996586
rect 508684 996530 508689 996586
rect 508032 996528 508689 996530
rect 509664 996586 510321 996588
rect 509664 996530 510260 996586
rect 510316 996530 510321 996586
rect 509664 996528 510321 996530
rect 508623 996525 508689 996528
rect 510255 996525 510321 996528
rect 436335 996292 436401 996295
rect 436335 996290 436608 996292
rect 436335 996234 436340 996290
rect 436396 996234 436608 996290
rect 436335 996232 436608 996234
rect 436335 996229 436401 996232
rect 317103 996144 317169 996147
rect 318639 996144 318705 996147
rect 436431 996144 436497 996147
rect 317103 996142 317280 996144
rect 317103 996086 317108 996142
rect 317164 996086 317280 996142
rect 317103 996084 317280 996086
rect 318639 996142 318816 996144
rect 318639 996086 318644 996142
rect 318700 996086 318816 996142
rect 318639 996084 318816 996086
rect 435840 996142 436497 996144
rect 435840 996086 436436 996142
rect 436492 996086 436497 996142
rect 435840 996084 436497 996086
rect 317103 996081 317169 996084
rect 318639 996081 318705 996084
rect 436431 996081 436497 996084
rect 513423 996144 513489 996147
rect 513423 996142 513696 996144
rect 513423 996086 513428 996142
rect 513484 996086 513696 996142
rect 513423 996084 513696 996086
rect 513423 996081 513489 996084
rect 313839 995996 313905 995999
rect 316335 995996 316401 995999
rect 326799 995996 326865 995999
rect 362319 995996 362385 995999
rect 367119 995996 367185 995999
rect 370575 995996 370641 995999
rect 377295 995996 377361 995999
rect 429711 995996 429777 995999
rect 313839 995994 314016 995996
rect 313839 995938 313844 995994
rect 313900 995938 314016 995994
rect 313839 995936 314016 995938
rect 316335 995994 316512 995996
rect 316335 995938 316340 995994
rect 316396 995938 316512 995994
rect 316335 995936 316512 995938
rect 321312 995994 326865 995996
rect 321312 995938 326804 995994
rect 326860 995938 326865 995994
rect 321312 995936 326865 995938
rect 362208 995994 362385 995996
rect 362208 995938 362324 995994
rect 362380 995938 362385 995994
rect 362208 995936 362385 995938
rect 366912 995994 367185 995996
rect 366912 995938 367124 995994
rect 367180 995938 367185 995994
rect 366912 995936 367185 995938
rect 370080 995994 370641 995996
rect 370080 995938 370580 995994
rect 370636 995938 370641 995994
rect 370080 995936 370641 995938
rect 371712 995994 377361 995996
rect 371712 995938 377300 995994
rect 377356 995938 377361 995994
rect 371712 995936 377361 995938
rect 429600 995994 429777 995996
rect 429600 995938 429716 995994
rect 429772 995938 429777 995994
rect 429600 995936 429777 995938
rect 313839 995933 313905 995936
rect 316335 995933 316401 995936
rect 326799 995933 326865 995936
rect 362319 995933 362385 995936
rect 367119 995933 367185 995936
rect 370575 995933 370641 995936
rect 377295 995933 377361 995936
rect 429711 995933 429777 995936
rect 434127 995996 434193 995999
rect 445071 995996 445137 995999
rect 434127 995994 434304 995996
rect 434127 995938 434132 995994
rect 434188 995938 434304 995994
rect 434127 995936 434304 995938
rect 439104 995994 445137 995996
rect 439104 995938 445076 995994
rect 445132 995938 445137 995994
rect 439104 995936 445137 995938
rect 434127 995933 434193 995936
rect 445071 995933 445137 995936
rect 471951 995996 472017 995999
rect 511119 995996 511185 995999
rect 513423 995996 513489 995999
rect 521295 995996 521361 995999
rect 471951 995994 481278 995996
rect 471951 995938 471956 995994
rect 472012 995938 481278 995994
rect 471951 995936 481278 995938
rect 471951 995933 472017 995936
rect 371343 995848 371409 995851
rect 304002 995788 304608 995848
rect 304002 995700 304062 995788
rect 303042 995640 304062 995700
rect 310287 995700 310353 995703
rect 312546 995700 312606 995818
rect 310287 995698 312606 995700
rect 310287 995642 310292 995698
rect 310348 995642 312606 995698
rect 310287 995640 312606 995642
rect 291087 995637 291153 995640
rect 299535 995637 299601 995640
rect 310287 995637 310353 995640
rect 291759 995552 291825 995555
rect 299631 995552 299697 995555
rect 291759 995550 299697 995552
rect 291759 995494 291764 995550
rect 291820 995494 299636 995550
rect 299692 995494 299697 995550
rect 291759 995492 299697 995494
rect 291759 995489 291825 995492
rect 299631 995489 299697 995492
rect 264015 995402 264126 995407
rect 264015 995346 264020 995402
rect 264076 995346 264126 995402
rect 264015 995344 264126 995346
rect 264015 995341 264081 995344
rect 250671 995254 258558 995256
rect 250671 995198 250676 995254
rect 250732 995198 258558 995254
rect 250671 995196 258558 995198
rect 311055 995256 311121 995259
rect 313218 995256 313278 995818
rect 311055 995254 313278 995256
rect 311055 995198 311060 995254
rect 311116 995198 313278 995254
rect 311055 995196 313278 995198
rect 250671 995193 250737 995196
rect 311055 995193 311121 995196
rect 207279 995106 210270 995108
rect 207279 995050 207284 995106
rect 207340 995050 210270 995106
rect 207279 995048 210270 995050
rect 237423 995108 237489 995111
rect 288783 995108 288849 995111
rect 237423 995106 288849 995108
rect 237423 995050 237428 995106
rect 237484 995050 288788 995106
rect 288844 995050 288849 995106
rect 237423 995048 288849 995050
rect 207279 995045 207345 995048
rect 237423 995045 237489 995048
rect 288783 995045 288849 995048
rect 198639 994960 198705 994963
rect 188610 994958 198705 994960
rect 188610 994902 198644 994958
rect 198700 994902 198705 994958
rect 188610 994900 198705 994902
rect 198639 994897 198705 994900
rect 134607 994812 134673 994815
rect 134607 994810 141054 994812
rect 134607 994754 134612 994810
rect 134668 994754 141054 994810
rect 134607 994752 141054 994754
rect 134607 994749 134673 994752
rect 84495 994664 84561 994667
rect 106575 994664 106641 994667
rect 84495 994662 106641 994664
rect 84495 994606 84500 994662
rect 84556 994606 106580 994662
rect 106636 994606 106641 994662
rect 84495 994604 106641 994606
rect 84495 994601 84561 994604
rect 106575 994601 106641 994604
rect 140994 994516 141054 994752
rect 146991 994664 147057 994667
rect 158415 994664 158481 994667
rect 146991 994662 158481 994664
rect 146991 994606 146996 994662
rect 147052 994606 158420 994662
rect 158476 994606 158481 994662
rect 146991 994604 158481 994606
rect 146991 994601 147057 994604
rect 158415 994601 158481 994604
rect 178479 994664 178545 994667
rect 185775 994664 185841 994667
rect 178479 994662 185841 994664
rect 178479 994606 178484 994662
rect 178540 994606 185780 994662
rect 185836 994606 185841 994662
rect 178479 994604 185841 994606
rect 178479 994601 178545 994604
rect 185775 994601 185841 994604
rect 238671 994664 238737 994667
rect 260463 994664 260529 994667
rect 238671 994662 260529 994664
rect 238671 994606 238676 994662
rect 238732 994606 260468 994662
rect 260524 994606 260529 994662
rect 238671 994604 260529 994606
rect 238671 994601 238737 994604
rect 260463 994601 260529 994604
rect 141231 994516 141297 994519
rect 140994 994514 141297 994516
rect 140994 994458 141236 994514
rect 141292 994458 141297 994514
rect 140994 994456 141297 994458
rect 141231 994453 141297 994456
rect 290319 994516 290385 994519
rect 310287 994516 310353 994519
rect 290319 994514 310353 994516
rect 290319 994458 290324 994514
rect 290380 994458 310292 994514
rect 310348 994458 310353 994514
rect 290319 994456 310353 994458
rect 290319 994453 290385 994456
rect 310287 994453 310353 994456
rect 295407 994368 295473 994371
rect 314850 994368 314910 995818
rect 319650 995700 319710 995818
rect 323919 995700 323985 995703
rect 319650 995698 323985 995700
rect 319650 995642 323924 995698
rect 323980 995642 323985 995698
rect 319650 995640 323985 995642
rect 323919 995637 323985 995640
rect 343887 995700 343953 995703
rect 353442 995700 353502 995818
rect 354912 995788 355134 995848
rect 370848 995846 371409 995848
rect 355074 995700 355134 995788
rect 343887 995698 355134 995700
rect 343887 995642 343892 995698
rect 343948 995642 355134 995698
rect 343887 995640 355134 995642
rect 368418 995700 368478 995818
rect 370848 995790 371348 995846
rect 371404 995790 371409 995846
rect 370848 995788 371409 995790
rect 371343 995785 371409 995788
rect 380175 995848 380241 995851
rect 388815 995848 388881 995851
rect 422511 995848 422577 995851
rect 438735 995848 438801 995851
rect 380175 995846 388881 995848
rect 380175 995790 380180 995846
rect 380236 995790 388820 995846
rect 388876 995790 388881 995846
rect 422304 995846 422656 995848
rect 380175 995788 388881 995790
rect 380175 995785 380241 995788
rect 388815 995785 388881 995788
rect 371535 995700 371601 995703
rect 368418 995698 371601 995700
rect 368418 995642 371540 995698
rect 371596 995642 371601 995698
rect 368418 995640 371601 995642
rect 343887 995637 343953 995640
rect 371535 995637 371601 995640
rect 380271 995700 380337 995703
rect 396687 995700 396753 995703
rect 380271 995698 396753 995700
rect 380271 995642 380276 995698
rect 380332 995642 396692 995698
rect 396748 995642 396753 995698
rect 380271 995640 396753 995642
rect 420834 995700 420894 995818
rect 422304 995790 422516 995846
rect 422572 995790 422656 995846
rect 438240 995846 438801 995848
rect 422304 995788 422656 995790
rect 422466 995785 422577 995788
rect 422466 995700 422526 995785
rect 420834 995640 422526 995700
rect 437442 995700 437502 995818
rect 438240 995790 438740 995846
rect 438796 995790 438801 995846
rect 438240 995788 438801 995790
rect 438735 995785 438801 995788
rect 472239 995848 472305 995851
rect 480975 995848 481041 995851
rect 472239 995846 481041 995848
rect 472239 995790 472244 995846
rect 472300 995790 480980 995846
rect 481036 995790 481041 995846
rect 472239 995788 481041 995790
rect 481218 995848 481278 995936
rect 511119 995994 511296 995996
rect 511119 995938 511124 995994
rect 511180 995938 511296 995994
rect 511119 995936 511296 995938
rect 512832 995994 513489 995996
rect 512832 995938 513428 995994
rect 513484 995938 513489 995994
rect 512832 995936 513489 995938
rect 516096 995994 521361 995996
rect 516096 995938 521300 995994
rect 521356 995938 521361 995994
rect 516096 995936 521361 995938
rect 511119 995933 511185 995936
rect 513423 995933 513489 995936
rect 521295 995933 521361 995936
rect 523503 995996 523569 995999
rect 523503 995994 528126 995996
rect 523503 995938 523508 995994
rect 523564 995938 528126 995994
rect 523503 995936 528126 995938
rect 523503 995933 523569 995936
rect 485679 995848 485745 995851
rect 499983 995848 500049 995851
rect 481218 995846 485745 995848
rect 481218 995790 485684 995846
rect 485740 995790 485745 995846
rect 499296 995846 500049 995848
rect 481218 995788 485745 995790
rect 472239 995785 472305 995788
rect 480975 995785 481041 995788
rect 485679 995785 485745 995788
rect 440655 995700 440721 995703
rect 437442 995698 440721 995700
rect 437442 995642 440660 995698
rect 440716 995642 440721 995698
rect 437442 995640 440721 995642
rect 380271 995637 380337 995640
rect 396687 995637 396753 995640
rect 440655 995637 440721 995640
rect 472047 995700 472113 995703
rect 477039 995700 477105 995703
rect 472047 995698 477105 995700
rect 472047 995642 472052 995698
rect 472108 995642 477044 995698
rect 477100 995642 477105 995698
rect 472047 995640 477105 995642
rect 472047 995637 472113 995640
rect 477039 995637 477105 995640
rect 479919 995700 479985 995703
rect 488847 995700 488913 995703
rect 479919 995698 488913 995700
rect 479919 995642 479924 995698
rect 479980 995642 488852 995698
rect 488908 995642 488913 995698
rect 479919 995640 488913 995642
rect 497826 995700 497886 995818
rect 499296 995790 499988 995846
rect 500044 995790 500049 995846
rect 511887 995848 511953 995851
rect 521199 995848 521265 995851
rect 527919 995848 527985 995851
rect 511887 995846 512160 995848
rect 499296 995788 500049 995790
rect 499458 995700 499518 995788
rect 499983 995785 500049 995788
rect 497826 995640 499518 995700
rect 479919 995637 479985 995640
rect 488847 995637 488913 995640
rect 471471 995552 471537 995555
rect 482031 995552 482097 995555
rect 471471 995550 482097 995552
rect 471471 995494 471476 995550
rect 471532 995494 482036 995550
rect 482092 995494 482097 995550
rect 471471 995492 482097 995494
rect 471471 995489 471537 995492
rect 482031 995489 482097 995492
rect 466479 995404 466545 995407
rect 476463 995404 476529 995407
rect 466479 995402 476529 995404
rect 466479 995346 466484 995402
rect 466540 995346 476468 995402
rect 476524 995346 476529 995402
rect 466479 995344 476529 995346
rect 466479 995341 466545 995344
rect 476463 995341 476529 995344
rect 506562 995259 506622 995818
rect 511887 995790 511892 995846
rect 511948 995790 512160 995846
rect 511887 995788 512160 995790
rect 511887 995785 511953 995788
rect 514434 995552 514494 995818
rect 515232 995788 515454 995848
rect 515394 995700 515454 995788
rect 521199 995846 527985 995848
rect 521199 995790 521204 995846
rect 521260 995790 527924 995846
rect 527980 995790 527985 995846
rect 521199 995788 527985 995790
rect 528066 995848 528126 995936
rect 532239 995848 532305 995851
rect 528066 995846 532305 995848
rect 528066 995790 532244 995846
rect 532300 995790 532305 995846
rect 549186 995848 549246 1002300
rect 560463 1002297 560529 1002300
rect 561519 1002297 561585 1002300
rect 555279 998068 555345 998071
rect 554688 998066 555345 998068
rect 554688 998010 555284 998066
rect 555340 998010 555345 998066
rect 554688 998008 555345 998010
rect 555279 998005 555345 998008
rect 557295 997920 557361 997923
rect 557088 997918 557361 997920
rect 557088 997862 557300 997918
rect 557356 997862 557361 997918
rect 557088 997860 557361 997862
rect 557295 997857 557361 997860
rect 564783 995996 564849 995999
rect 564783 995994 565056 995996
rect 564783 995938 564788 995994
rect 564844 995938 565056 995994
rect 564783 995936 565056 995938
rect 564783 995933 564849 995936
rect 573135 995848 573201 995851
rect 549186 995818 549630 995848
rect 567456 995846 573201 995848
rect 528066 995788 532305 995790
rect 549216 995788 549630 995818
rect 521199 995785 521265 995788
rect 527919 995785 527985 995788
rect 532239 995785 532305 995788
rect 518415 995700 518481 995703
rect 515394 995698 518481 995700
rect 515394 995642 518420 995698
rect 518476 995642 518481 995698
rect 515394 995640 518481 995642
rect 518415 995637 518481 995640
rect 523599 995700 523665 995703
rect 526095 995700 526161 995703
rect 523599 995698 526161 995700
rect 523599 995642 523604 995698
rect 523660 995642 526100 995698
rect 526156 995642 526161 995698
rect 523599 995640 526161 995642
rect 549570 995700 549630 995788
rect 550722 995700 550782 995818
rect 549570 995640 550782 995700
rect 523599 995637 523665 995640
rect 526095 995637 526161 995640
rect 518607 995552 518673 995555
rect 514434 995550 518673 995552
rect 514434 995494 518612 995550
rect 518668 995494 518673 995550
rect 514434 995492 518673 995494
rect 518607 995489 518673 995492
rect 520911 995552 520977 995555
rect 535311 995552 535377 995555
rect 520911 995550 535377 995552
rect 520911 995494 520916 995550
rect 520972 995494 535316 995550
rect 535372 995494 535377 995550
rect 520911 995492 535377 995494
rect 520911 995489 520977 995492
rect 535311 995489 535377 995492
rect 557922 995407 557982 995818
rect 562722 995703 562782 995818
rect 563490 995703 563550 995818
rect 562722 995698 562833 995703
rect 562722 995642 562772 995698
rect 562828 995642 562833 995698
rect 562722 995640 562833 995642
rect 563490 995698 563601 995703
rect 563490 995642 563540 995698
rect 563596 995642 563601 995698
rect 563490 995640 563601 995642
rect 562767 995637 562833 995640
rect 563535 995637 563601 995640
rect 565794 995552 565854 995818
rect 566658 995700 566718 995818
rect 567456 995790 573140 995846
rect 573196 995790 573201 995846
rect 567456 995788 573201 995790
rect 573135 995785 573201 995788
rect 570351 995700 570417 995703
rect 566658 995698 570417 995700
rect 566658 995642 570356 995698
rect 570412 995642 570417 995698
rect 566658 995640 570417 995642
rect 570351 995637 570417 995640
rect 570543 995552 570609 995555
rect 565794 995550 570609 995552
rect 565794 995494 570548 995550
rect 570604 995494 570609 995550
rect 565794 995492 570609 995494
rect 570543 995489 570609 995492
rect 523311 995404 523377 995407
rect 530895 995404 530961 995407
rect 523311 995402 530961 995404
rect 523311 995346 523316 995402
rect 523372 995346 530900 995402
rect 530956 995346 530961 995402
rect 523311 995344 530961 995346
rect 557922 995402 558033 995407
rect 557922 995346 557972 995402
rect 558028 995346 558033 995402
rect 557922 995344 558033 995346
rect 523311 995341 523377 995344
rect 530895 995341 530961 995344
rect 557967 995341 558033 995344
rect 506562 995254 506673 995259
rect 506562 995198 506612 995254
rect 506668 995198 506673 995254
rect 506562 995196 506673 995198
rect 506607 995193 506673 995196
rect 573231 994664 573297 994667
rect 631791 994664 631857 994667
rect 573231 994662 631857 994664
rect 573231 994606 573236 994662
rect 573292 994606 631796 994662
rect 631852 994606 631857 994662
rect 573231 994604 631857 994606
rect 573231 994601 573297 994604
rect 631791 994601 631857 994604
rect 567567 994516 567633 994519
rect 628143 994516 628209 994519
rect 567567 994514 628209 994516
rect 567567 994458 567572 994514
rect 567628 994458 628148 994514
rect 628204 994458 628209 994514
rect 567567 994456 628209 994458
rect 567567 994453 567633 994456
rect 628143 994453 628209 994456
rect 295407 994366 314910 994368
rect 295407 994310 295412 994366
rect 295468 994310 314910 994366
rect 295407 994308 314910 994310
rect 570447 994368 570513 994371
rect 634287 994368 634353 994371
rect 570447 994366 634353 994368
rect 570447 994310 570452 994366
rect 570508 994310 634292 994366
rect 634348 994310 634353 994366
rect 570447 994308 634353 994310
rect 295407 994305 295473 994308
rect 570447 994305 570513 994308
rect 634287 994305 634353 994308
rect 187311 994220 187377 994223
rect 207375 994220 207441 994223
rect 187311 994218 207441 994220
rect 187311 994162 187316 994218
rect 187372 994162 207380 994218
rect 207436 994162 207441 994218
rect 187311 994160 207441 994162
rect 187311 994157 187377 994160
rect 207375 994157 207441 994160
rect 231471 994220 231537 994223
rect 261807 994220 261873 994223
rect 231471 994218 261873 994220
rect 231471 994162 231476 994218
rect 231532 994162 261812 994218
rect 261868 994162 261873 994218
rect 231471 994160 261873 994162
rect 231471 994157 231537 994160
rect 261807 994157 261873 994160
rect 285999 994220 286065 994223
rect 311055 994220 311121 994223
rect 285999 994218 311121 994220
rect 285999 994162 286004 994218
rect 286060 994162 311060 994218
rect 311116 994162 311121 994218
rect 285999 994160 311121 994162
rect 285999 994157 286065 994160
rect 311055 994157 311121 994160
rect 531183 994220 531249 994223
rect 631023 994220 631089 994223
rect 632751 994220 632817 994223
rect 531183 994218 632817 994220
rect 531183 994162 531188 994218
rect 531244 994162 631028 994218
rect 631084 994162 632756 994218
rect 632812 994162 632817 994218
rect 531183 994160 632817 994162
rect 531183 994157 531249 994160
rect 631023 994157 631089 994160
rect 632751 994157 632817 994160
rect 136143 994072 136209 994075
rect 156687 994072 156753 994075
rect 136143 994070 156753 994072
rect 136143 994014 136148 994070
rect 136204 994014 156692 994070
rect 156748 994014 156753 994070
rect 136143 994012 156753 994014
rect 136143 994009 136209 994012
rect 156687 994009 156753 994012
rect 185775 994072 185841 994075
rect 237423 994072 237489 994075
rect 185775 994070 237489 994072
rect 185775 994014 185780 994070
rect 185836 994014 237428 994070
rect 237484 994014 237489 994070
rect 185775 994012 237489 994014
rect 185775 994009 185841 994012
rect 237423 994009 237489 994012
rect 288783 994072 288849 994075
rect 390831 994072 390897 994075
rect 479823 994072 479889 994075
rect 288783 994070 479889 994072
rect 288783 994014 288788 994070
rect 288844 994014 390836 994070
rect 390892 994014 479828 994070
rect 479884 994014 479889 994070
rect 288783 994012 479889 994014
rect 288783 994009 288849 994012
rect 390831 994009 390897 994012
rect 479823 994009 479889 994012
rect 485583 994072 485649 994075
rect 604719 994072 604785 994075
rect 485583 994070 604785 994072
rect 485583 994014 485588 994070
rect 485644 994014 604724 994070
rect 604780 994014 604785 994070
rect 485583 994012 604785 994014
rect 485583 994009 485649 994012
rect 604719 994009 604785 994012
rect 61839 993924 61905 993927
rect 82575 993924 82641 993927
rect 61839 993922 82641 993924
rect 61839 993866 61844 993922
rect 61900 993866 82580 993922
rect 82636 993866 82641 993922
rect 61839 993864 82641 993866
rect 61839 993861 61905 993864
rect 82575 993861 82641 993864
rect 191535 993924 191601 993927
rect 649551 993924 649617 993927
rect 191535 993922 649617 993924
rect 191535 993866 191540 993922
rect 191596 993866 649556 993922
rect 649612 993866 649617 993922
rect 191535 993864 649617 993866
rect 191535 993861 191601 993864
rect 649551 993861 649617 993864
rect 78351 993776 78417 993779
rect 108399 993776 108465 993779
rect 78351 993774 108465 993776
rect 78351 993718 78356 993774
rect 78412 993718 108404 993774
rect 108460 993718 108465 993774
rect 78351 993716 108465 993718
rect 78351 993713 78417 993716
rect 108399 993713 108465 993716
rect 140367 993776 140433 993779
rect 621999 993776 622065 993779
rect 140367 993774 622065 993776
rect 140367 993718 140372 993774
rect 140428 993718 622004 993774
rect 622060 993718 622065 993774
rect 140367 993716 622065 993718
rect 140367 993713 140433 993716
rect 621999 993713 622065 993716
rect 83439 993628 83505 993631
rect 93039 993628 93105 993631
rect 83439 993626 93105 993628
rect 83439 993570 83444 993626
rect 83500 993570 93044 993626
rect 93100 993570 93105 993626
rect 83439 993568 93105 993570
rect 83439 993565 83505 993568
rect 93039 993565 93105 993568
rect 279279 993628 279345 993631
rect 288399 993628 288465 993631
rect 279279 993626 288465 993628
rect 279279 993570 279284 993626
rect 279340 993570 288404 993626
rect 288460 993570 288465 993626
rect 279279 993568 288465 993570
rect 279279 993565 279345 993568
rect 288399 993565 288465 993568
rect 390159 993628 390225 993631
rect 469455 993628 469521 993631
rect 390159 993626 469521 993628
rect 390159 993570 390164 993626
rect 390220 993570 469460 993626
rect 469516 993570 469521 993626
rect 390159 993568 469521 993570
rect 390159 993565 390225 993568
rect 469455 993565 469521 993568
rect 62031 992148 62097 992151
rect 83439 992148 83505 992151
rect 62031 992146 83505 992148
rect 62031 992090 62036 992146
rect 62092 992090 83444 992146
rect 83500 992090 83505 992146
rect 62031 992088 83505 992090
rect 62031 992085 62097 992088
rect 83439 992085 83505 992088
rect 288399 992148 288465 992151
rect 390159 992148 390225 992151
rect 288399 992146 390225 992148
rect 288399 992090 288404 992146
rect 288460 992090 390164 992146
rect 390220 992090 390225 992146
rect 288399 992088 390225 992090
rect 288399 992085 288465 992088
rect 390159 992085 390225 992088
rect 100815 985488 100881 985491
rect 120879 985488 120945 985491
rect 100815 985486 120945 985488
rect 100815 985430 100820 985486
rect 100876 985430 120884 985486
rect 120940 985430 120945 985486
rect 100815 985428 120945 985430
rect 100815 985425 100881 985428
rect 120879 985425 120945 985428
rect 239055 985340 239121 985343
rect 239535 985340 239601 985343
rect 239055 985338 239601 985340
rect 239055 985282 239060 985338
rect 239116 985282 239540 985338
rect 239596 985282 239601 985338
rect 239055 985280 239601 985282
rect 239055 985277 239121 985280
rect 239535 985277 239601 985280
rect 239151 985192 239217 985195
rect 239727 985192 239793 985195
rect 239151 985190 239793 985192
rect 239151 985134 239156 985190
rect 239212 985134 239732 985190
rect 239788 985134 239793 985190
rect 239151 985132 239793 985134
rect 239151 985129 239217 985132
rect 239727 985129 239793 985132
rect 161295 981048 161361 981051
rect 171279 981048 171345 981051
rect 161295 981046 171345 981048
rect 161295 980990 161300 981046
rect 161356 980990 171284 981046
rect 171340 980990 171345 981046
rect 161295 980988 171345 980990
rect 161295 980985 161361 980988
rect 171279 980985 171345 980988
rect 218895 980752 218961 980755
rect 238959 980752 239025 980755
rect 218895 980750 239025 980752
rect 218895 980694 218900 980750
rect 218956 980694 238964 980750
rect 239020 980694 239025 980750
rect 218895 980692 239025 980694
rect 218895 980689 218961 980692
rect 238959 980689 239025 980692
rect 655119 974684 655185 974687
rect 650208 974682 655185 974684
rect 650208 974626 655124 974682
rect 655180 974626 655185 974682
rect 650208 974624 655185 974626
rect 655119 974621 655185 974624
rect 59535 973204 59601 973207
rect 59535 973202 64416 973204
rect 59535 973146 59540 973202
rect 59596 973146 64416 973202
rect 59535 973144 64416 973146
rect 59535 973141 59601 973144
rect 42063 968766 42129 968767
rect 42063 968762 42112 968766
rect 42176 968764 42182 968766
rect 42063 968706 42068 968762
rect 42063 968702 42112 968706
rect 42176 968704 42220 968764
rect 42176 968702 42182 968704
rect 42063 968701 42129 968702
rect 40378 967074 40384 967138
rect 40448 967136 40454 967138
rect 41775 967136 41841 967139
rect 40448 967134 41841 967136
rect 40448 967078 41780 967134
rect 41836 967078 41841 967134
rect 40448 967076 41841 967078
rect 40448 967074 40454 967076
rect 41775 967073 41841 967076
rect 674362 966334 674368 966398
rect 674432 966396 674438 966398
rect 675375 966396 675441 966399
rect 674432 966394 675441 966396
rect 674432 966338 675380 966394
rect 675436 966338 675441 966394
rect 674432 966336 675441 966338
rect 674432 966334 674438 966336
rect 675375 966333 675441 966336
rect 675759 965804 675825 965807
rect 676474 965804 676480 965806
rect 675759 965802 676480 965804
rect 675759 965746 675764 965802
rect 675820 965746 676480 965802
rect 675759 965744 676480 965746
rect 675759 965741 675825 965744
rect 676474 965742 676480 965744
rect 676544 965742 676550 965806
rect 40954 965002 40960 965066
rect 41024 965064 41030 965066
rect 41775 965064 41841 965067
rect 41024 965062 41841 965064
rect 41024 965006 41780 965062
rect 41836 965006 41841 965062
rect 41024 965004 41841 965006
rect 41024 965002 41030 965004
rect 41775 965001 41841 965004
rect 675759 965064 675825 965067
rect 675898 965064 675904 965066
rect 675759 965062 675904 965064
rect 675759 965006 675764 965062
rect 675820 965006 675904 965062
rect 675759 965004 675904 965006
rect 675759 965001 675825 965004
rect 675898 965002 675904 965004
rect 675968 965002 675974 965066
rect 42159 964028 42225 964031
rect 42490 964028 42496 964030
rect 42159 964026 42496 964028
rect 42159 963970 42164 964026
rect 42220 963970 42496 964026
rect 42159 963968 42496 963970
rect 42159 963965 42225 963968
rect 42490 963966 42496 963968
rect 42560 963966 42566 964030
rect 41338 963374 41344 963438
rect 41408 963436 41414 963438
rect 41775 963436 41841 963439
rect 41408 963434 41841 963436
rect 41408 963378 41780 963434
rect 41836 963378 41841 963434
rect 41408 963376 41841 963378
rect 41408 963374 41414 963376
rect 41775 963373 41841 963376
rect 675375 963290 675441 963291
rect 675322 963288 675328 963290
rect 675284 963228 675328 963288
rect 675392 963286 675441 963290
rect 675436 963230 675441 963286
rect 675322 963226 675328 963228
rect 675392 963226 675441 963230
rect 675375 963225 675441 963226
rect 42159 962844 42225 962847
rect 42298 962844 42304 962846
rect 42159 962842 42304 962844
rect 42159 962786 42164 962842
rect 42220 962786 42304 962842
rect 42159 962784 42304 962786
rect 42159 962781 42225 962784
rect 42298 962782 42304 962784
rect 42368 962782 42374 962846
rect 655215 962844 655281 962847
rect 650208 962842 655281 962844
rect 650208 962786 655220 962842
rect 655276 962786 655281 962842
rect 650208 962784 655281 962786
rect 655215 962781 655281 962784
rect 674746 962634 674752 962698
rect 674816 962696 674822 962698
rect 675471 962696 675537 962699
rect 674816 962694 675537 962696
rect 674816 962638 675476 962694
rect 675532 962638 675537 962694
rect 674816 962636 675537 962638
rect 674816 962634 674822 962636
rect 675471 962633 675537 962636
rect 42543 962548 42609 962551
rect 62031 962548 62097 962551
rect 42543 962546 62097 962548
rect 42543 962490 42548 962546
rect 42604 962490 62036 962546
rect 62092 962490 62097 962546
rect 42543 962488 62097 962490
rect 42543 962485 42609 962488
rect 62031 962485 62097 962488
rect 674554 962190 674560 962254
rect 674624 962252 674630 962254
rect 675375 962252 675441 962255
rect 674624 962250 675441 962252
rect 674624 962194 675380 962250
rect 675436 962194 675441 962250
rect 674624 962192 675441 962194
rect 674624 962190 674630 962192
rect 675375 962189 675441 962192
rect 41722 962042 41728 962106
rect 41792 962104 41798 962106
rect 41871 962104 41937 962107
rect 41792 962102 41937 962104
rect 41792 962046 41876 962102
rect 41932 962046 41937 962102
rect 41792 962044 41937 962046
rect 41792 962042 41798 962044
rect 41871 962041 41937 962044
rect 42351 962104 42417 962107
rect 61839 962104 61905 962107
rect 42351 962102 61905 962104
rect 42351 962046 42356 962102
rect 42412 962046 61844 962102
rect 61900 962046 61905 962102
rect 42351 962044 61905 962046
rect 42351 962041 42417 962044
rect 61839 962041 61905 962044
rect 675759 961364 675825 961367
rect 676090 961364 676096 961366
rect 675759 961362 676096 961364
rect 675759 961306 675764 961362
rect 675820 961306 676096 961362
rect 675759 961304 676096 961306
rect 675759 961301 675825 961304
rect 676090 961302 676096 961304
rect 676160 961302 676166 961366
rect 675663 960774 675729 960775
rect 675663 960772 675712 960774
rect 675620 960770 675712 960772
rect 675620 960714 675668 960770
rect 675620 960712 675712 960714
rect 675663 960710 675712 960712
rect 675776 960710 675782 960774
rect 675663 960709 675729 960710
rect 675471 960182 675537 960183
rect 675471 960180 675520 960182
rect 675428 960178 675520 960180
rect 675428 960122 675476 960178
rect 675428 960120 675520 960122
rect 675471 960118 675520 960120
rect 675584 960118 675590 960182
rect 675471 960117 675537 960118
rect 41146 959674 41152 959738
rect 41216 959736 41222 959738
rect 41775 959736 41841 959739
rect 41216 959734 41841 959736
rect 41216 959678 41780 959734
rect 41836 959678 41841 959734
rect 41216 959676 41841 959678
rect 41216 959674 41222 959676
rect 41775 959673 41841 959676
rect 41530 959082 41536 959146
rect 41600 959144 41606 959146
rect 41775 959144 41841 959147
rect 41600 959142 41841 959144
rect 41600 959086 41780 959142
rect 41836 959086 41841 959142
rect 41600 959084 41841 959086
rect 41600 959082 41606 959084
rect 41775 959081 41841 959084
rect 59535 958848 59601 958851
rect 59535 958846 64416 958848
rect 59535 958790 59540 958846
rect 59596 958790 64416 958846
rect 59535 958788 64416 958790
rect 59535 958785 59601 958788
rect 41967 958406 42033 958407
rect 41914 958404 41920 958406
rect 41876 958344 41920 958404
rect 41984 958402 42033 958406
rect 42028 958346 42033 958402
rect 41914 958342 41920 958344
rect 41984 958342 42033 958346
rect 41967 958341 42033 958342
rect 40762 957750 40768 957814
rect 40832 957812 40838 957814
rect 41775 957812 41841 957815
rect 40832 957810 41841 957812
rect 40832 957754 41780 957810
rect 41836 957754 41841 957810
rect 40832 957752 41841 957754
rect 40832 957750 40838 957752
rect 41775 957749 41841 957752
rect 674938 957602 674944 957666
rect 675008 957664 675014 957666
rect 675375 957664 675441 957667
rect 675008 957662 675441 957664
rect 675008 957606 675380 957662
rect 675436 957606 675441 957662
rect 675008 957604 675441 957606
rect 675008 957602 675014 957604
rect 675375 957601 675441 957604
rect 40570 956122 40576 956186
rect 40640 956184 40646 956186
rect 41775 956184 41841 956187
rect 40640 956182 41841 956184
rect 40640 956126 41780 956182
rect 41836 956126 41841 956182
rect 40640 956124 41841 956126
rect 40640 956122 40646 956124
rect 41775 956121 41841 956124
rect 675130 955974 675136 956038
rect 675200 956036 675206 956038
rect 675471 956036 675537 956039
rect 675200 956034 675537 956036
rect 675200 955978 675476 956034
rect 675532 955978 675537 956034
rect 675200 955976 675537 955978
rect 675200 955974 675206 955976
rect 675471 955973 675537 955976
rect 675087 953520 675153 953523
rect 677050 953520 677056 953522
rect 675087 953518 677056 953520
rect 675087 953462 675092 953518
rect 675148 953462 677056 953518
rect 675087 953460 677056 953462
rect 675087 953457 675153 953460
rect 677050 953458 677056 953460
rect 677120 953458 677126 953522
rect 675183 953372 675249 953375
rect 676858 953372 676864 953374
rect 675183 953370 676864 953372
rect 675183 953314 675188 953370
rect 675244 953314 676864 953370
rect 675183 953312 676864 953314
rect 675183 953309 675249 953312
rect 676858 953310 676864 953312
rect 676928 953310 676934 953374
rect 42543 953224 42609 953227
rect 42874 953224 42880 953226
rect 42543 953222 42880 953224
rect 42543 953166 42548 953222
rect 42604 953166 42880 953222
rect 42543 953164 42880 953166
rect 42543 953161 42609 953164
rect 42874 953162 42880 953164
rect 42944 953162 42950 953226
rect 654351 951152 654417 951155
rect 650208 951150 654417 951152
rect 650208 951094 654356 951150
rect 654412 951094 654417 951150
rect 650208 951092 654417 951094
rect 654351 951089 654417 951092
rect 42114 949379 42174 949494
rect 42114 949374 42225 949379
rect 42114 949318 42164 949374
rect 42220 949318 42225 949374
rect 42114 949316 42225 949318
rect 42159 949313 42225 949316
rect 42306 948491 42366 948680
rect 42306 948486 42417 948491
rect 42306 948430 42356 948486
rect 42412 948430 42417 948486
rect 42306 948428 42417 948430
rect 42351 948425 42417 948428
rect 43119 947896 43185 947899
rect 42336 947894 43185 947896
rect 42336 947838 43124 947894
rect 43180 947838 43185 947894
rect 42336 947836 43185 947838
rect 43119 947833 43185 947836
rect 42639 947602 42705 947603
rect 42639 947598 42688 947602
rect 42752 947600 42758 947602
rect 42639 947542 42644 947598
rect 42639 947538 42688 947542
rect 42752 947540 42796 947600
rect 42752 947538 42758 947540
rect 42639 947537 42705 947538
rect 42682 947390 42688 947454
rect 42752 947390 42758 947454
rect 42874 947390 42880 947454
rect 42944 947452 42950 947454
rect 42944 947392 43134 947452
rect 42944 947390 42950 947392
rect 40386 946567 40446 947052
rect 42690 947008 42750 947390
rect 43074 947306 43134 947392
rect 43066 947242 43072 947306
rect 43136 947242 43142 947306
rect 43023 947008 43089 947011
rect 42690 947006 43089 947008
rect 42690 946950 43028 947006
rect 43084 946950 43089 947006
rect 42690 946948 43089 946950
rect 43023 946945 43089 946948
rect 40335 946562 40446 946567
rect 40335 946506 40340 946562
rect 40396 946506 40446 946562
rect 40335 946504 40446 946506
rect 40335 946501 40401 946504
rect 47439 946268 47505 946271
rect 42336 946266 47505 946268
rect 42336 946210 47444 946266
rect 47500 946210 47505 946266
rect 42336 946208 47505 946210
rect 47439 946205 47505 946208
rect 44751 945676 44817 945679
rect 42306 945674 44817 945676
rect 42306 945618 44756 945674
rect 44812 945618 44817 945674
rect 42306 945616 44817 945618
rect 42306 945602 42366 945616
rect 44751 945613 44817 945616
rect 40224 945572 42366 945602
rect 40194 945542 42336 945572
rect 40047 945084 40113 945087
rect 40194 945084 40254 945542
rect 674754 945383 674814 945942
rect 674703 945378 674814 945383
rect 674703 945322 674708 945378
rect 674764 945322 674814 945378
rect 674703 945320 674814 945322
rect 674703 945317 674769 945320
rect 40047 945082 40254 945084
rect 40047 945026 40052 945082
rect 40108 945026 40254 945082
rect 40047 945024 40254 945026
rect 40047 945021 40113 945024
rect 674754 944791 674814 945054
rect 42682 944788 42688 944790
rect 42336 944728 42688 944788
rect 42682 944726 42688 944728
rect 42752 944788 42758 944790
rect 44559 944788 44625 944791
rect 42752 944786 44625 944788
rect 42752 944730 44564 944786
rect 44620 944730 44625 944786
rect 42752 944728 44625 944730
rect 42752 944726 42758 944728
rect 44559 944725 44625 944728
rect 674703 944786 674814 944791
rect 674703 944730 674708 944786
rect 674764 944730 674814 944786
rect 674703 944728 674814 944730
rect 674703 944725 674769 944728
rect 59535 944640 59601 944643
rect 59535 944638 64416 944640
rect 59535 944582 59540 944638
rect 59596 944582 64416 944638
rect 59535 944580 64416 944582
rect 59535 944577 59601 944580
rect 40570 944430 40576 944494
rect 40640 944430 40646 944494
rect 40578 943944 40638 944430
rect 674607 944048 674673 944051
rect 674754 944048 674814 944240
rect 674607 944046 674814 944048
rect 674607 943990 674612 944046
rect 674668 943990 674814 944046
rect 674607 943988 674814 943990
rect 674607 943985 674673 943988
rect 40378 943690 40384 943754
rect 40448 943690 40454 943754
rect 40386 943130 40446 943690
rect 674754 943311 674814 943426
rect 674754 943306 674865 943311
rect 674754 943250 674804 943306
rect 674860 943250 674865 943306
rect 674754 943248 674865 943250
rect 674799 943245 674865 943248
rect 674754 942423 674814 942612
rect 674703 942418 674814 942423
rect 674703 942362 674708 942418
rect 674764 942362 674814 942418
rect 674703 942360 674814 942362
rect 674703 942357 674769 942360
rect 42831 942272 42897 942275
rect 42336 942270 42897 942272
rect 42336 942214 42836 942270
rect 42892 942214 42897 942270
rect 42336 942212 42897 942214
rect 42831 942209 42897 942212
rect 674703 942124 674769 942127
rect 674703 942122 674814 942124
rect 674703 942066 674708 942122
rect 674764 942066 674814 942122
rect 674703 942061 674814 942066
rect 674754 941946 674814 942061
rect 40762 941618 40768 941682
rect 40832 941618 40838 941682
rect 40770 941502 40830 941618
rect 41722 941174 41728 941238
rect 41792 941174 41798 941238
rect 41730 940762 41790 941174
rect 674754 940795 674814 941132
rect 675898 940878 675904 940942
rect 675968 940878 675974 940942
rect 674703 940790 674814 940795
rect 674703 940734 674708 940790
rect 674764 940734 674814 940790
rect 674703 940732 674814 940734
rect 674703 940729 674769 940732
rect 42106 940582 42112 940646
rect 42176 940582 42182 940646
rect 42114 940022 42174 940582
rect 675906 940318 675966 940878
rect 674127 939608 674193 939611
rect 674127 939606 674814 939608
rect 674127 939550 674132 939606
rect 674188 939550 674814 939606
rect 674127 939548 674814 939550
rect 674127 939545 674193 939548
rect 674754 939504 674814 939548
rect 653775 939460 653841 939463
rect 650208 939458 653841 939460
rect 650208 939402 653780 939458
rect 653836 939402 653841 939458
rect 650208 939400 653841 939402
rect 653775 939397 653841 939400
rect 42927 939164 42993 939167
rect 42336 939162 42993 939164
rect 42336 939106 42932 939162
rect 42988 939106 42993 939162
rect 42336 939104 42993 939106
rect 42927 939101 42993 939104
rect 41914 938806 41920 938870
rect 41984 938806 41990 938870
rect 41922 938394 41982 938806
rect 674362 938658 674368 938722
rect 674432 938720 674438 938722
rect 674432 938660 674784 938720
rect 674432 938658 674438 938660
rect 675322 938362 675328 938426
rect 675392 938362 675398 938426
rect 41530 938066 41536 938130
rect 41600 938066 41606 938130
rect 41538 937506 41598 938066
rect 675330 937802 675390 938362
rect 40954 937326 40960 937390
rect 41024 937326 41030 937390
rect 40962 936766 41022 937326
rect 673935 937240 674001 937243
rect 673935 937238 674784 937240
rect 673935 937182 673940 937238
rect 673996 937182 674784 937238
rect 673935 937180 674784 937182
rect 673935 937177 674001 937180
rect 41338 936438 41344 936502
rect 41408 936438 41414 936502
rect 41346 936026 41406 936438
rect 674031 936352 674097 936355
rect 674031 936350 674784 936352
rect 674031 936294 674036 936350
rect 674092 936294 674784 936350
rect 674031 936292 674784 936294
rect 674031 936289 674097 936292
rect 41146 935846 41152 935910
rect 41216 935846 41222 935910
rect 676474 935846 676480 935910
rect 676544 935846 676550 935910
rect 41154 935286 41214 935846
rect 676482 935582 676542 935846
rect 674746 935254 674752 935318
rect 674816 935254 674822 935318
rect 42298 934958 42304 935022
rect 42368 934958 42374 935022
rect 42306 934398 42366 934958
rect 674754 934694 674814 935254
rect 674554 934514 674560 934578
rect 674624 934576 674630 934578
rect 674624 934516 674814 934576
rect 674624 934514 674630 934516
rect 42490 934132 42496 934134
rect 42306 934072 42496 934132
rect 42306 933584 42366 934072
rect 42490 934070 42496 934072
rect 42560 934070 42566 934134
rect 674754 933954 674814 934516
rect 675130 933330 675136 933394
rect 675200 933330 675206 933394
rect 43023 933098 43089 933099
rect 43023 933096 43072 933098
rect 42980 933094 43072 933096
rect 42980 933038 43028 933094
rect 42980 933036 43072 933038
rect 43023 933034 43072 933036
rect 43136 933034 43142 933098
rect 675138 933066 675198 933330
rect 43023 933033 43089 933034
rect 674938 932886 674944 932950
rect 675008 932886 675014 932950
rect 42306 932655 42366 932770
rect 42306 932650 42417 932655
rect 42306 932594 42356 932650
rect 42412 932594 42417 932650
rect 42306 932592 42417 932594
rect 42351 932589 42417 932592
rect 674946 932474 675006 932886
rect 676090 932146 676096 932210
rect 676160 932146 676166 932210
rect 676098 931586 676158 932146
rect 677050 931406 677056 931470
rect 677120 931406 677126 931470
rect 42306 931027 42366 931290
rect 42306 931022 42417 931027
rect 42306 930966 42356 931022
rect 42412 930966 42417 931022
rect 42306 930964 42417 930966
rect 42351 930961 42417 930964
rect 677058 930846 677118 931406
rect 676858 930222 676864 930286
rect 676928 930222 676934 930286
rect 59535 930136 59601 930139
rect 59535 930134 64416 930136
rect 59535 930078 59540 930134
rect 59596 930078 64416 930134
rect 59535 930076 64416 930078
rect 59535 930073 59601 930076
rect 676866 929958 676926 930222
rect 679746 928659 679806 929144
rect 679746 928654 679857 928659
rect 679746 928598 679796 928654
rect 679852 928598 679857 928654
rect 679746 928596 679857 928598
rect 679791 928593 679857 928596
rect 679791 928064 679857 928067
rect 679746 928062 679857 928064
rect 679746 928006 679796 928062
rect 679852 928006 679857 928062
rect 679746 928001 679857 928006
rect 679746 927664 679806 928001
rect 654447 927620 654513 927623
rect 650208 927618 654513 927620
rect 650208 927562 654452 927618
rect 654508 927562 654513 927618
rect 650208 927560 654513 927562
rect 654447 927557 654513 927560
rect 654447 915928 654513 915931
rect 650208 915926 654513 915928
rect 650208 915870 654452 915926
rect 654508 915870 654513 915926
rect 650208 915868 654513 915870
rect 654447 915865 654513 915868
rect 59535 915780 59601 915783
rect 59535 915778 64416 915780
rect 59535 915722 59540 915778
rect 59596 915722 64416 915778
rect 59535 915720 64416 915722
rect 59535 915717 59601 915720
rect 42490 912906 42496 912970
rect 42560 912968 42566 912970
rect 43066 912968 43072 912970
rect 42560 912908 43072 912968
rect 42560 912906 42566 912908
rect 43066 912906 43072 912908
rect 43136 912906 43142 912970
rect 42490 907134 42496 907198
rect 42560 907196 42566 907198
rect 43119 907196 43185 907199
rect 42560 907194 43185 907196
rect 42560 907138 43124 907194
rect 43180 907138 43185 907194
rect 42560 907136 43185 907138
rect 42560 907134 42566 907136
rect 43119 907133 43185 907136
rect 654447 904236 654513 904239
rect 650208 904234 654513 904236
rect 650208 904178 654452 904234
rect 654508 904178 654513 904234
rect 650208 904176 654513 904178
rect 654447 904173 654513 904176
rect 58191 901572 58257 901575
rect 58191 901570 64416 901572
rect 58191 901514 58196 901570
rect 58252 901514 64416 901570
rect 58191 901512 64416 901514
rect 58191 901509 58257 901512
rect 650031 892840 650097 892843
rect 649986 892838 650097 892840
rect 649986 892782 650036 892838
rect 650092 892782 650097 892838
rect 649986 892777 650097 892782
rect 649986 892514 650046 892777
rect 43119 887218 43185 887219
rect 43066 887154 43072 887218
rect 43136 887216 43185 887218
rect 43136 887214 43228 887216
rect 43180 887158 43228 887214
rect 43136 887156 43228 887158
rect 43136 887154 43185 887156
rect 43119 887153 43185 887154
rect 59535 887068 59601 887071
rect 59535 887066 64416 887068
rect 59535 887010 59540 887066
rect 59596 887010 64416 887066
rect 59535 887008 64416 887010
rect 59535 887005 59601 887008
rect 654447 880704 654513 880707
rect 650208 880702 654513 880704
rect 650208 880646 654452 880702
rect 654508 880646 654513 880702
rect 650208 880644 654513 880646
rect 654447 880641 654513 880644
rect 674554 876350 674560 876414
rect 674624 876412 674630 876414
rect 675087 876412 675153 876415
rect 674624 876410 675153 876412
rect 674624 876354 675092 876410
rect 675148 876354 675153 876410
rect 674624 876352 675153 876354
rect 674624 876350 674630 876352
rect 675087 876349 675153 876352
rect 675759 876412 675825 876415
rect 676090 876412 676096 876414
rect 675759 876410 676096 876412
rect 675759 876354 675764 876410
rect 675820 876354 676096 876410
rect 675759 876352 676096 876354
rect 675759 876349 675825 876352
rect 676090 876350 676096 876352
rect 676160 876350 676166 876414
rect 674938 876202 674944 876266
rect 675008 876264 675014 876266
rect 675087 876264 675153 876267
rect 675008 876262 675153 876264
rect 675008 876206 675092 876262
rect 675148 876206 675153 876262
rect 675008 876204 675153 876206
rect 675008 876202 675014 876204
rect 675087 876201 675153 876204
rect 675279 875820 675345 875823
rect 675514 875820 675520 875822
rect 675279 875818 675520 875820
rect 675279 875762 675284 875818
rect 675340 875762 675520 875818
rect 675279 875760 675520 875762
rect 675279 875757 675345 875760
rect 675514 875758 675520 875760
rect 675584 875758 675590 875822
rect 675183 875672 675249 875675
rect 675706 875672 675712 875674
rect 675183 875670 675712 875672
rect 675183 875614 675188 875670
rect 675244 875614 675712 875670
rect 675183 875612 675712 875614
rect 675183 875609 675249 875612
rect 675706 875610 675712 875612
rect 675776 875610 675782 875674
rect 674746 873982 674752 874046
rect 674816 874044 674822 874046
rect 675471 874044 675537 874047
rect 674816 874042 675537 874044
rect 674816 873986 675476 874042
rect 675532 873986 675537 874042
rect 674816 873984 675537 873986
rect 674816 873982 674822 873984
rect 675471 873981 675537 873984
rect 674362 873390 674368 873454
rect 674432 873452 674438 873454
rect 675375 873452 675441 873455
rect 674432 873450 675441 873452
rect 674432 873394 675380 873450
rect 675436 873394 675441 873450
rect 674432 873392 675441 873394
rect 674432 873390 674438 873392
rect 675375 873389 675441 873392
rect 674170 872798 674176 872862
rect 674240 872860 674246 872862
rect 675375 872860 675441 872863
rect 674240 872858 675441 872860
rect 674240 872802 675380 872858
rect 675436 872802 675441 872858
rect 674240 872800 675441 872802
rect 674240 872798 674246 872800
rect 675375 872797 675441 872800
rect 42490 872502 42496 872566
rect 42560 872564 42566 872566
rect 43066 872564 43072 872566
rect 42560 872504 43072 872564
rect 42560 872502 42566 872504
rect 43066 872502 43072 872504
rect 43136 872502 43142 872566
rect 58959 872564 59025 872567
rect 58959 872562 64416 872564
rect 58959 872506 58964 872562
rect 59020 872506 64416 872562
rect 58959 872504 64416 872506
rect 58959 872501 59025 872504
rect 675375 869902 675441 869903
rect 675322 869900 675328 869902
rect 675284 869840 675328 869900
rect 675392 869898 675441 869902
rect 675436 869842 675441 869898
rect 675322 869838 675328 869840
rect 675392 869838 675441 869842
rect 675375 869837 675441 869838
rect 654447 869012 654513 869015
rect 650208 869010 654513 869012
rect 650208 868954 654452 869010
rect 654508 868954 654513 869010
rect 650208 868952 654513 868954
rect 654447 868949 654513 868952
rect 675130 866878 675136 866942
rect 675200 866940 675206 866942
rect 675375 866940 675441 866943
rect 675200 866938 675441 866940
rect 675200 866882 675380 866938
rect 675436 866882 675441 866938
rect 675200 866880 675441 866882
rect 675200 866878 675206 866880
rect 675375 866877 675441 866880
rect 675663 864722 675729 864723
rect 675663 864718 675712 864722
rect 675776 864720 675782 864722
rect 675663 864662 675668 864718
rect 675663 864658 675712 864662
rect 675776 864660 675820 864720
rect 675776 864658 675782 864660
rect 675663 864657 675729 864658
rect 675471 862946 675537 862947
rect 675471 862942 675520 862946
rect 675584 862944 675590 862946
rect 675471 862886 675476 862942
rect 675471 862882 675520 862886
rect 675584 862884 675628 862944
rect 675584 862882 675590 862884
rect 675471 862881 675537 862882
rect 59535 858356 59601 858359
rect 59535 858354 64416 858356
rect 59535 858298 59540 858354
rect 59596 858298 64416 858354
rect 59535 858296 64416 858298
rect 59535 858293 59601 858296
rect 654447 857320 654513 857323
rect 650208 857318 654513 857320
rect 650208 857262 654452 857318
rect 654508 857262 654513 857318
rect 650208 857260 654513 857262
rect 654447 857257 654513 857260
rect 42490 846750 42496 846814
rect 42560 846812 42566 846814
rect 43066 846812 43072 846814
rect 42560 846752 43072 846812
rect 42560 846750 42566 846752
rect 43066 846750 43072 846752
rect 43136 846750 43142 846814
rect 649935 846220 650001 846223
rect 649935 846218 650046 846220
rect 649935 846162 649940 846218
rect 649996 846162 650046 846218
rect 649935 846157 650046 846162
rect 649986 845598 650046 846157
rect 59535 844000 59601 844003
rect 59535 843998 64416 844000
rect 59535 843942 59540 843998
rect 59596 843942 64416 843998
rect 59535 843940 64416 843942
rect 59535 843937 59601 843940
rect 654447 833788 654513 833791
rect 650208 833786 654513 833788
rect 650208 833730 654452 833786
rect 654508 833730 654513 833786
rect 650208 833728 654513 833730
rect 654447 833725 654513 833728
rect 41914 832246 41920 832310
rect 41984 832308 41990 832310
rect 43066 832308 43072 832310
rect 41984 832248 43072 832308
rect 41984 832246 41990 832248
rect 43066 832246 43072 832248
rect 43136 832246 43142 832310
rect 59535 829644 59601 829647
rect 59535 829642 64416 829644
rect 59535 829586 59540 829642
rect 59596 829586 64416 829642
rect 59535 829584 64416 829586
rect 59535 829581 59601 829584
rect 674799 826684 674865 826687
rect 674799 826682 675006 826684
rect 674799 826626 674804 826682
rect 674860 826626 675006 826682
rect 674799 826624 675006 826626
rect 674799 826621 674865 826624
rect 674946 826539 675006 826624
rect 674895 826534 675006 826539
rect 674895 826478 674900 826534
rect 674956 826478 675006 826534
rect 674895 826476 675006 826478
rect 674895 826473 674961 826476
rect 42351 823872 42417 823875
rect 42306 823870 42417 823872
rect 42306 823814 42356 823870
rect 42412 823814 42417 823870
rect 42306 823809 42417 823814
rect 42306 823694 42366 823809
rect 42306 822688 42366 822880
rect 42447 822688 42513 822691
rect 42306 822686 42513 822688
rect 42306 822630 42452 822686
rect 42508 822630 42513 822686
rect 42306 822628 42513 822630
rect 42447 822625 42513 822628
rect 42351 822244 42417 822247
rect 42306 822242 42417 822244
rect 42306 822186 42356 822242
rect 42412 822186 42417 822242
rect 42306 822181 42417 822186
rect 42306 822066 42366 822181
rect 654447 822096 654513 822099
rect 650208 822094 654513 822096
rect 650208 822038 654452 822094
rect 654508 822038 654513 822094
rect 650208 822036 654513 822038
rect 654447 822033 654513 822036
rect 43215 821208 43281 821211
rect 42336 821206 43281 821208
rect 42336 821150 43220 821206
rect 43276 821150 43281 821206
rect 42336 821148 43281 821150
rect 43215 821145 43281 821148
rect 40335 820764 40401 820767
rect 40335 820762 40446 820764
rect 40335 820706 40340 820762
rect 40396 820706 40446 820762
rect 40335 820701 40446 820706
rect 40386 820438 40446 820701
rect 40047 820172 40113 820175
rect 40002 820170 40113 820172
rect 40002 820114 40052 820170
rect 40108 820114 40113 820170
rect 40002 820109 40113 820114
rect 37455 819136 37521 819139
rect 40002 819136 40062 820109
rect 42106 819518 42112 819582
rect 42176 819518 42182 819582
rect 37455 819134 40062 819136
rect 37455 819078 37460 819134
rect 37516 819078 40062 819134
rect 37455 819076 40062 819078
rect 37455 819073 37521 819076
rect 42114 818988 42174 819518
rect 40800 818958 42174 818988
rect 40770 818928 42144 818958
rect 40770 818694 40830 818928
rect 40762 818630 40768 818694
rect 40832 818630 40838 818694
rect 41730 817955 41790 818070
rect 41679 817950 41790 817955
rect 41679 817894 41684 817950
rect 41740 817894 41790 817950
rect 41679 817892 41790 817894
rect 41679 817889 41745 817892
rect 40194 816771 40254 817330
rect 40143 816766 40254 816771
rect 40143 816710 40148 816766
rect 40204 816710 40254 816766
rect 40143 816708 40254 816710
rect 40143 816705 40209 816708
rect 40194 815883 40254 816442
rect 41914 816262 41920 816326
rect 41984 816324 41990 816326
rect 42682 816324 42688 816326
rect 41984 816264 42688 816324
rect 41984 816262 41990 816264
rect 42682 816262 42688 816264
rect 42752 816262 42758 816326
rect 40194 815878 40305 815883
rect 40194 815822 40244 815878
rect 40300 815822 40305 815878
rect 40194 815820 40305 815822
rect 40239 815817 40305 815820
rect 41538 815291 41598 815702
rect 41538 815286 41649 815291
rect 41538 815230 41588 815286
rect 41644 815230 41649 815286
rect 41538 815228 41649 815230
rect 41583 815225 41649 815228
rect 59535 815288 59601 815291
rect 59535 815286 64416 815288
rect 59535 815230 59540 815286
rect 59596 815230 64416 815286
rect 59535 815228 64416 815230
rect 59535 815225 59601 815228
rect 41922 814403 41982 814962
rect 41922 814398 42033 814403
rect 41922 814342 41972 814398
rect 42028 814342 42033 814398
rect 41922 814340 42033 814342
rect 41967 814337 42033 814340
rect 41922 813663 41982 814222
rect 41871 813658 41982 813663
rect 41871 813602 41876 813658
rect 41932 813602 41982 813658
rect 41871 813600 41982 813602
rect 41871 813597 41937 813600
rect 37314 812775 37374 813334
rect 37314 812770 37425 812775
rect 37314 812714 37364 812770
rect 37420 812714 37425 812770
rect 37314 812712 37425 812714
rect 37359 812709 37425 812712
rect 42306 812331 42366 812520
rect 42306 812326 42417 812331
rect 42306 812270 42356 812326
rect 42412 812270 42417 812326
rect 42306 812268 42417 812270
rect 42351 812265 42417 812268
rect 42490 811970 42496 812034
rect 42560 812032 42566 812034
rect 42874 812032 42880 812034
rect 42560 811972 42880 812032
rect 42560 811970 42566 811972
rect 42874 811970 42880 811972
rect 42944 811970 42950 812034
rect 42114 811147 42174 811706
rect 42063 811142 42174 811147
rect 42063 811086 42068 811142
rect 42124 811086 42174 811142
rect 42063 811084 42174 811086
rect 42063 811081 42129 811084
rect 42306 810404 42366 810892
rect 43119 810404 43185 810407
rect 654447 810404 654513 810407
rect 42306 810402 43185 810404
rect 42306 810346 43124 810402
rect 43180 810346 43185 810402
rect 42306 810344 43185 810346
rect 650208 810402 654513 810404
rect 650208 810346 654452 810402
rect 654508 810346 654513 810402
rect 650208 810344 654513 810346
rect 43119 810341 43185 810344
rect 654447 810341 654513 810344
rect 41730 809667 41790 810226
rect 41730 809662 41841 809667
rect 41730 809606 41780 809662
rect 41836 809606 41841 809662
rect 41730 809604 41841 809606
rect 41775 809601 41841 809604
rect 42306 809368 42366 809412
rect 43023 809368 43089 809371
rect 42306 809366 43089 809368
rect 42306 809310 43028 809366
rect 43084 809310 43089 809366
rect 42306 809308 43089 809310
rect 43023 809305 43089 809308
rect 42114 808335 42174 808598
rect 42114 808330 42225 808335
rect 42114 808274 42164 808330
rect 42220 808274 42225 808330
rect 42114 808272 42225 808274
rect 42159 808269 42225 808272
rect 42306 807592 42366 807784
rect 42447 807592 42513 807595
rect 42306 807590 42513 807592
rect 42306 807534 42452 807590
rect 42508 807534 42513 807590
rect 42306 807532 42513 807534
rect 42447 807529 42513 807532
rect 42306 806408 42366 806970
rect 42306 806348 42750 806408
rect 42690 805964 42750 806348
rect 42306 805904 42750 805964
rect 42306 805227 42366 805904
rect 42255 805222 42366 805227
rect 42255 805166 42260 805222
rect 42316 805166 42366 805222
rect 42255 805164 42366 805166
rect 42255 805161 42321 805164
rect 42447 803598 42513 803599
rect 42447 803596 42496 803598
rect 42404 803594 42496 803596
rect 42404 803538 42452 803594
rect 42404 803536 42496 803538
rect 42447 803534 42496 803536
rect 42560 803534 42566 803598
rect 42447 803533 42513 803534
rect 37359 802264 37425 802267
rect 41338 802264 41344 802266
rect 37359 802262 41344 802264
rect 37359 802206 37364 802262
rect 37420 802206 41344 802262
rect 37359 802204 41344 802206
rect 37359 802201 37425 802204
rect 41338 802202 41344 802204
rect 41408 802202 41414 802266
rect 37263 802116 37329 802119
rect 40378 802116 40384 802118
rect 37263 802114 40384 802116
rect 37263 802058 37268 802114
rect 37324 802058 40384 802114
rect 37263 802056 40384 802058
rect 37263 802053 37329 802056
rect 40378 802054 40384 802056
rect 40448 802054 40454 802118
rect 40239 801968 40305 801971
rect 41530 801968 41536 801970
rect 40239 801966 41536 801968
rect 40239 801910 40244 801966
rect 40300 801910 41536 801966
rect 40239 801908 41536 801910
rect 40239 801905 40305 801908
rect 41530 801906 41536 801908
rect 41600 801906 41606 801970
rect 59535 800784 59601 800787
rect 59535 800782 64416 800784
rect 59535 800726 59540 800782
rect 59596 800726 64416 800782
rect 59535 800724 64416 800726
rect 59535 800721 59601 800724
rect 41775 800342 41841 800343
rect 41722 800340 41728 800342
rect 41684 800280 41728 800340
rect 41792 800338 41841 800342
rect 41836 800282 41841 800338
rect 41722 800278 41728 800280
rect 41792 800278 41841 800282
rect 41775 800277 41841 800278
rect 42063 800340 42129 800343
rect 42490 800340 42496 800342
rect 42063 800338 42496 800340
rect 42063 800282 42068 800338
rect 42124 800282 42496 800338
rect 42063 800280 42496 800282
rect 42063 800277 42129 800280
rect 42490 800278 42496 800280
rect 42560 800278 42566 800342
rect 42255 800046 42321 800047
rect 42255 800042 42304 800046
rect 42368 800044 42374 800046
rect 42255 799986 42260 800042
rect 42255 799982 42304 799986
rect 42368 799984 42412 800044
rect 42368 799982 42374 799984
rect 42255 799981 42321 799982
rect 653775 798712 653841 798715
rect 650208 798710 653841 798712
rect 650208 798654 653780 798710
rect 653836 798654 653841 798710
rect 650208 798652 653841 798654
rect 653775 798649 653841 798652
rect 42298 797910 42304 797974
rect 42368 797972 42374 797974
rect 42447 797972 42513 797975
rect 42368 797970 42513 797972
rect 42368 797914 42452 797970
rect 42508 797914 42513 797970
rect 42368 797912 42513 797914
rect 42368 797910 42374 797912
rect 42447 797909 42513 797912
rect 42490 794802 42496 794866
rect 42560 794864 42566 794866
rect 42735 794864 42801 794867
rect 42560 794862 42801 794864
rect 42560 794806 42740 794862
rect 42796 794806 42801 794862
rect 42560 794804 42801 794806
rect 42560 794802 42566 794804
rect 42735 794801 42801 794804
rect 41775 794274 41841 794275
rect 41722 794210 41728 794274
rect 41792 794272 41841 794274
rect 41792 794270 41884 794272
rect 41836 794214 41884 794270
rect 41792 794212 41884 794214
rect 41792 794210 41841 794212
rect 41775 794209 41841 794210
rect 41530 791842 41536 791906
rect 41600 791904 41606 791906
rect 42447 791904 42513 791907
rect 41600 791902 42513 791904
rect 41600 791846 42452 791902
rect 42508 791846 42513 791902
rect 41600 791844 42513 791846
rect 41600 791842 41606 791844
rect 42447 791841 42513 791844
rect 41338 791694 41344 791758
rect 41408 791756 41414 791758
rect 42735 791756 42801 791759
rect 41408 791754 42801 791756
rect 41408 791698 42740 791754
rect 42796 791698 42801 791754
rect 41408 791696 42801 791698
rect 41408 791694 41414 791696
rect 42735 791693 42801 791696
rect 41775 791314 41841 791315
rect 41722 791312 41728 791314
rect 41684 791252 41728 791312
rect 41792 791310 41841 791314
rect 41836 791254 41841 791310
rect 41722 791250 41728 791252
rect 41792 791250 41841 791254
rect 41775 791249 41841 791250
rect 41914 790954 41920 791018
rect 41984 791016 41990 791018
rect 42159 791016 42225 791019
rect 42490 791016 42496 791018
rect 41984 791014 42496 791016
rect 41984 790958 42164 791014
rect 42220 790958 42496 791014
rect 41984 790956 42496 790958
rect 41984 790954 41990 790956
rect 42159 790953 42225 790956
rect 42490 790954 42496 790956
rect 42560 790954 42566 791018
rect 675759 787908 675825 787911
rect 676282 787908 676288 787910
rect 675759 787906 676288 787908
rect 675759 787850 675764 787906
rect 675820 787850 676288 787906
rect 675759 787848 676288 787850
rect 675759 787845 675825 787848
rect 676282 787846 676288 787848
rect 676352 787846 676358 787910
rect 673978 787402 673984 787466
rect 674048 787464 674054 787466
rect 675471 787464 675537 787467
rect 674048 787462 675537 787464
rect 674048 787406 675476 787462
rect 675532 787406 675537 787462
rect 674048 787404 675537 787406
rect 674048 787402 674054 787404
rect 675471 787401 675537 787404
rect 654447 786872 654513 786875
rect 650208 786870 654513 786872
rect 650208 786814 654452 786870
rect 654508 786814 654513 786870
rect 650208 786812 654513 786814
rect 654447 786809 654513 786812
rect 675759 786724 675825 786727
rect 676474 786724 676480 786726
rect 675759 786722 676480 786724
rect 675759 786666 675764 786722
rect 675820 786666 676480 786722
rect 675759 786664 676480 786666
rect 675759 786661 675825 786664
rect 676474 786662 676480 786664
rect 676544 786662 676550 786726
rect 58959 786576 59025 786579
rect 58959 786574 64416 786576
rect 58959 786518 58964 786574
rect 59020 786518 64416 786574
rect 58959 786516 64416 786518
rect 58959 786513 59025 786516
rect 675759 784208 675825 784211
rect 675898 784208 675904 784210
rect 675759 784206 675904 784208
rect 675759 784150 675764 784206
rect 675820 784150 675904 784206
rect 675759 784148 675904 784150
rect 675759 784145 675825 784148
rect 675898 784146 675904 784148
rect 675968 784146 675974 784210
rect 675759 781988 675825 781991
rect 676666 781988 676672 781990
rect 675759 781986 676672 781988
rect 675759 781930 675764 781986
rect 675820 781930 676672 781986
rect 675759 781928 676672 781930
rect 675759 781925 675825 781928
rect 676666 781926 676672 781928
rect 676736 781926 676742 781990
rect 42735 780508 42801 780511
rect 42336 780506 42801 780508
rect 42336 780450 42740 780506
rect 42796 780450 42801 780506
rect 42336 780448 42801 780450
rect 42735 780445 42801 780448
rect 674223 780508 674289 780511
rect 677050 780508 677056 780510
rect 674223 780506 677056 780508
rect 674223 780450 674228 780506
rect 674284 780450 677056 780506
rect 674223 780448 677056 780450
rect 674223 780445 674289 780448
rect 677050 780446 677056 780448
rect 677120 780446 677126 780510
rect 42447 779916 42513 779919
rect 42306 779914 42513 779916
rect 42306 779858 42452 779914
rect 42508 779858 42513 779914
rect 42306 779856 42513 779858
rect 42306 779664 42366 779856
rect 42447 779853 42513 779856
rect 42735 778880 42801 778883
rect 42336 778878 42801 778880
rect 42336 778822 42740 778878
rect 42796 778822 42801 778878
rect 42336 778820 42801 778822
rect 42735 778817 42801 778820
rect 42306 777992 42366 778036
rect 43311 777992 43377 777995
rect 42306 777990 43377 777992
rect 42306 777934 43316 777990
rect 43372 777934 43377 777990
rect 42306 777932 43377 777934
rect 43311 777929 43377 777932
rect 674991 777548 675057 777551
rect 677050 777548 677056 777550
rect 674991 777546 677056 777548
rect 674991 777490 674996 777546
rect 675052 777490 677056 777546
rect 674991 777488 677056 777490
rect 674991 777485 675057 777488
rect 677050 777486 677056 777488
rect 677120 777486 677126 777550
rect 674703 777400 674769 777403
rect 676858 777400 676864 777402
rect 674703 777398 676864 777400
rect 674703 777342 674708 777398
rect 674764 777342 676864 777398
rect 674703 777340 676864 777342
rect 674703 777337 674769 777340
rect 676858 777338 676864 777340
rect 676928 777338 676934 777402
rect 43215 777252 43281 777255
rect 42336 777250 43281 777252
rect 42336 777194 43220 777250
rect 43276 777194 43281 777250
rect 42336 777192 43281 777194
rect 43215 777189 43281 777192
rect 40378 776746 40384 776810
rect 40448 776746 40454 776810
rect 40386 776512 40446 776746
rect 40386 776482 41376 776512
rect 40416 776452 41406 776482
rect 41346 775922 41406 776452
rect 41338 775858 41344 775922
rect 41408 775858 41414 775922
rect 40770 775182 40830 775742
rect 40762 775118 40768 775182
rect 40832 775118 40838 775182
rect 654447 775180 654513 775183
rect 650208 775178 654513 775180
rect 650208 775122 654452 775178
rect 654508 775122 654513 775178
rect 650208 775120 654513 775122
rect 654447 775117 654513 775120
rect 42831 774884 42897 774887
rect 42336 774882 42897 774884
rect 42336 774826 42836 774882
rect 42892 774826 42897 774882
rect 42336 774824 42897 774826
rect 42831 774821 42897 774824
rect 39042 773555 39102 774114
rect 38991 773550 39102 773555
rect 38991 773494 38996 773550
rect 39052 773494 39102 773550
rect 38991 773492 39102 773494
rect 38991 773489 39057 773492
rect 38850 772667 38910 773226
rect 676858 773046 676864 773110
rect 676928 773108 676934 773110
rect 677818 773108 677824 773110
rect 676928 773048 677824 773108
rect 676928 773046 676934 773048
rect 677818 773046 677824 773048
rect 677888 773046 677894 773110
rect 676858 772898 676864 772962
rect 676928 772960 676934 772962
rect 677242 772960 677248 772962
rect 676928 772900 677248 772960
rect 676928 772898 676934 772900
rect 677242 772898 677248 772900
rect 677312 772898 677318 772962
rect 38799 772662 38910 772667
rect 38799 772606 38804 772662
rect 38860 772606 38910 772662
rect 38799 772604 38910 772606
rect 674415 772664 674481 772667
rect 677242 772664 677248 772666
rect 674415 772662 677248 772664
rect 674415 772606 674420 772662
rect 674476 772606 677248 772662
rect 674415 772604 677248 772606
rect 38799 772601 38865 772604
rect 674415 772601 674481 772604
rect 677242 772602 677248 772604
rect 677312 772602 677318 772666
rect 42927 772516 42993 772519
rect 42336 772514 42993 772516
rect 42336 772458 42932 772514
rect 42988 772458 42993 772514
rect 42336 772456 42993 772458
rect 42927 772453 42993 772456
rect 59535 772072 59601 772075
rect 59535 772070 64416 772072
rect 59535 772014 59540 772070
rect 59596 772014 64416 772070
rect 59535 772012 64416 772014
rect 59535 772009 59601 772012
rect 42306 771184 42366 771746
rect 42447 771184 42513 771187
rect 42306 771182 42513 771184
rect 42306 771126 42452 771182
rect 42508 771126 42513 771182
rect 42306 771124 42513 771126
rect 42447 771121 42513 771124
rect 41730 770447 41790 771006
rect 41730 770442 41841 770447
rect 41730 770386 41780 770442
rect 41836 770386 41841 770442
rect 41730 770384 41841 770386
rect 41775 770381 41841 770384
rect 37314 769559 37374 770118
rect 37314 769554 37425 769559
rect 37314 769498 37364 769554
rect 37420 769498 37425 769554
rect 37314 769496 37425 769498
rect 37359 769493 37425 769496
rect 41922 769115 41982 769378
rect 41871 769110 41982 769115
rect 41871 769054 41876 769110
rect 41932 769054 41982 769110
rect 41871 769052 41982 769054
rect 41871 769049 41937 769052
rect 41922 767931 41982 768490
rect 41922 767926 42033 767931
rect 41922 767870 41972 767926
rect 42028 767870 42033 767926
rect 41922 767868 42033 767870
rect 41967 767865 42033 767868
rect 43119 767780 43185 767783
rect 42336 767778 43185 767780
rect 42336 767722 43124 767778
rect 43180 767722 43185 767778
rect 42336 767720 43185 767722
rect 43119 767717 43185 767720
rect 674415 767484 674481 767487
rect 674415 767482 674784 767484
rect 674415 767426 674420 767482
rect 674476 767426 674784 767482
rect 674415 767424 674784 767426
rect 674415 767421 674481 767424
rect 43023 767040 43089 767043
rect 42336 767038 43089 767040
rect 42336 766982 43028 767038
rect 43084 766982 43089 767038
rect 42336 766980 43089 766982
rect 43023 766977 43089 766980
rect 674703 766892 674769 766895
rect 674703 766890 674814 766892
rect 674703 766834 674708 766890
rect 674764 766834 674814 766890
rect 674703 766829 674814 766834
rect 674754 766714 674814 766829
rect 42114 766006 42174 766196
rect 42106 765942 42112 766006
rect 42176 765942 42182 766006
rect 674415 765856 674481 765859
rect 674415 765854 674784 765856
rect 674415 765798 674420 765854
rect 674476 765798 674784 765854
rect 674415 765796 674784 765798
rect 674415 765793 674481 765796
rect 42114 765267 42174 765382
rect 42063 765262 42174 765267
rect 42063 765206 42068 765262
rect 42124 765206 42174 765262
rect 42063 765204 42174 765206
rect 674703 765264 674769 765267
rect 674703 765262 674814 765264
rect 674703 765206 674708 765262
rect 674764 765206 674814 765262
rect 42063 765201 42129 765204
rect 674703 765201 674814 765206
rect 674754 765086 674814 765201
rect 41538 764082 41598 764568
rect 673743 764228 673809 764231
rect 673743 764226 674784 764228
rect 673743 764170 673748 764226
rect 673804 764170 674784 764226
rect 673743 764168 674784 764170
rect 673743 764165 673809 764168
rect 41530 764018 41536 764082
rect 41600 764018 41606 764082
rect 42735 763784 42801 763787
rect 42336 763782 42801 763784
rect 42336 763726 42740 763782
rect 42796 763726 42801 763782
rect 42336 763724 42801 763726
rect 42735 763721 42801 763724
rect 674754 763343 674814 763532
rect 654447 763340 654513 763343
rect 650208 763338 654513 763340
rect 650208 763282 654452 763338
rect 654508 763282 654513 763338
rect 650208 763280 654513 763282
rect 654447 763277 654513 763280
rect 674703 763338 674814 763343
rect 674703 763282 674708 763338
rect 674764 763282 674814 763338
rect 674703 763280 674814 763282
rect 674703 763277 674769 763280
rect 674754 762603 674814 762718
rect 674703 762598 674814 762603
rect 674703 762542 674708 762598
rect 674764 762542 674814 762598
rect 674703 762540 674814 762542
rect 674703 762537 674769 762540
rect 674938 762390 674944 762454
rect 675008 762390 675014 762454
rect 42735 762304 42801 762307
rect 42336 762302 42801 762304
rect 42336 762246 42740 762302
rect 42796 762246 42801 762302
rect 42336 762244 42801 762246
rect 42735 762241 42801 762244
rect 674946 761904 675006 762390
rect 675706 761650 675712 761714
rect 675776 761650 675782 761714
rect 675714 761090 675774 761650
rect 674554 760466 674560 760530
rect 674624 760528 674630 760530
rect 674624 760468 674814 760528
rect 674624 760466 674630 760468
rect 674754 760276 674814 760468
rect 38799 760232 38865 760235
rect 40954 760232 40960 760234
rect 38799 760230 40960 760232
rect 38799 760174 38804 760230
rect 38860 760174 40960 760230
rect 38799 760172 40960 760174
rect 38799 760169 38865 760172
rect 40954 760170 40960 760172
rect 41024 760170 41030 760234
rect 674746 760022 674752 760086
rect 674816 760022 674822 760086
rect 674754 759462 674814 760022
rect 675322 759134 675328 759198
rect 675392 759134 675398 759198
rect 675330 758722 675390 759134
rect 37359 758604 37425 758607
rect 40378 758604 40384 758606
rect 37359 758602 40384 758604
rect 37359 758546 37364 758602
rect 37420 758546 40384 758602
rect 37359 758544 40384 758546
rect 37359 758541 37425 758544
rect 40378 758542 40384 758544
rect 40448 758542 40454 758606
rect 675514 758542 675520 758606
rect 675584 758542 675590 758606
rect 675522 757982 675582 758542
rect 59535 757716 59601 757719
rect 59535 757714 64416 757716
rect 59535 757658 59540 757714
rect 59596 757658 64416 757714
rect 59535 757656 64416 757658
rect 59535 757653 59601 757656
rect 676090 757358 676096 757422
rect 676160 757358 676166 757422
rect 676098 757094 676158 757358
rect 674362 756322 674368 756386
rect 674432 756384 674438 756386
rect 674432 756324 674784 756384
rect 674432 756322 674438 756324
rect 674170 755434 674176 755498
rect 674240 755496 674246 755498
rect 674240 755436 674784 755496
rect 674240 755434 674246 755436
rect 675130 755286 675136 755350
rect 675200 755286 675206 755350
rect 675138 754726 675198 755286
rect 676858 754398 676864 754462
rect 676928 754398 676934 754462
rect 676866 753986 676926 754398
rect 677818 753806 677824 753870
rect 677888 753806 677894 753870
rect 677826 753246 677886 753806
rect 677242 752918 677248 752982
rect 677312 752918 677318 752982
rect 649647 752388 649713 752391
rect 649602 752386 649713 752388
rect 649602 752330 649652 752386
rect 649708 752330 649713 752386
rect 677250 752358 677310 752918
rect 649602 752325 649713 752330
rect 42831 751946 42897 751947
rect 42831 751944 42880 751946
rect 42788 751942 42880 751944
rect 42788 751886 42836 751942
rect 42788 751884 42880 751886
rect 42831 751882 42880 751884
rect 42944 751882 42950 751946
rect 42831 751881 42897 751882
rect 41530 751734 41536 751798
rect 41600 751796 41606 751798
rect 41775 751796 41841 751799
rect 41600 751794 41841 751796
rect 41600 751738 41780 751794
rect 41836 751738 41841 751794
rect 649602 751766 649662 752325
rect 41600 751736 41841 751738
rect 41600 751734 41606 751736
rect 41775 751733 41841 751736
rect 42831 751650 42897 751651
rect 42831 751648 42880 751650
rect 42788 751646 42880 751648
rect 42788 751590 42836 751646
rect 42788 751588 42880 751590
rect 42831 751586 42880 751588
rect 42944 751586 42950 751650
rect 673647 751648 673713 751651
rect 673647 751646 674784 751648
rect 673647 751590 673652 751646
rect 673708 751590 674784 751646
rect 673647 751588 674784 751590
rect 42831 751585 42897 751586
rect 673647 751585 673713 751588
rect 679746 750171 679806 750730
rect 679695 750166 679806 750171
rect 679695 750110 679700 750166
rect 679756 750110 679806 750166
rect 679695 750108 679806 750110
rect 679695 750105 679761 750108
rect 679695 749576 679761 749579
rect 679695 749574 679806 749576
rect 679695 749518 679700 749574
rect 679756 749518 679806 749574
rect 679695 749513 679806 749518
rect 679746 749250 679806 749513
rect 41775 748690 41841 748691
rect 41722 748626 41728 748690
rect 41792 748688 41841 748690
rect 41792 748686 41884 748688
rect 41836 748630 41884 748686
rect 41792 748628 41884 748630
rect 41792 748626 41841 748628
rect 41775 748625 41841 748626
rect 42159 747506 42225 747507
rect 42106 747504 42112 747506
rect 42068 747444 42112 747504
rect 42176 747502 42225 747506
rect 42220 747446 42225 747502
rect 42106 747442 42112 747444
rect 42176 747442 42225 747446
rect 42159 747441 42225 747442
rect 41967 747358 42033 747359
rect 41914 747294 41920 747358
rect 41984 747356 42033 747358
rect 41984 747354 42076 747356
rect 42028 747298 42076 747354
rect 41984 747296 42076 747298
rect 41984 747294 42033 747296
rect 41967 747293 42033 747294
rect 40378 747146 40384 747210
rect 40448 747208 40454 747210
rect 42927 747208 42993 747211
rect 40448 747206 42993 747208
rect 40448 747150 42932 747206
rect 42988 747150 42993 747206
rect 40448 747148 42993 747150
rect 40448 747146 40454 747148
rect 42927 747145 42993 747148
rect 40954 746850 40960 746914
rect 41024 746912 41030 746914
rect 42735 746912 42801 746915
rect 41024 746910 42801 746912
rect 41024 746854 42740 746910
rect 42796 746854 42801 746910
rect 41024 746852 42801 746854
rect 41024 746850 41030 746852
rect 42735 746849 42801 746852
rect 41914 745814 41920 745878
rect 41984 745814 41990 745878
rect 41922 745432 41982 745814
rect 42106 745432 42112 745434
rect 41922 745372 42112 745432
rect 42106 745370 42112 745372
rect 42176 745370 42182 745434
rect 59535 743360 59601 743363
rect 59535 743358 64416 743360
rect 59535 743302 59540 743358
rect 59596 743302 64416 743358
rect 59535 743300 64416 743302
rect 59535 743297 59601 743300
rect 674554 743298 674560 743362
rect 674624 743360 674630 743362
rect 675087 743360 675153 743363
rect 674624 743358 675153 743360
rect 674624 743302 675092 743358
rect 675148 743302 675153 743358
rect 674624 743300 675153 743302
rect 674624 743298 674630 743300
rect 675087 743297 675153 743300
rect 674170 742114 674176 742178
rect 674240 742176 674246 742178
rect 675087 742176 675153 742179
rect 674240 742174 675153 742176
rect 674240 742118 675092 742174
rect 675148 742118 675153 742174
rect 674240 742116 675153 742118
rect 674240 742114 674246 742116
rect 675087 742113 675153 742116
rect 674746 740190 674752 740254
rect 674816 740252 674822 740254
rect 675087 740252 675153 740255
rect 674816 740250 675153 740252
rect 674816 740194 675092 740250
rect 675148 740194 675153 740250
rect 674816 740192 675153 740194
rect 674816 740190 674822 740192
rect 675087 740189 675153 740192
rect 674362 740042 674368 740106
rect 674432 740104 674438 740106
rect 675375 740104 675441 740107
rect 674432 740102 675441 740104
rect 674432 740046 675380 740102
rect 675436 740046 675441 740102
rect 674432 740044 675441 740046
rect 674432 740042 674438 740044
rect 675375 740041 675441 740044
rect 654447 739956 654513 739959
rect 650208 739954 654513 739956
rect 650208 739898 654452 739954
rect 654508 739898 654513 739954
rect 650208 739896 654513 739898
rect 654447 739893 654513 739896
rect 675471 739218 675537 739219
rect 675471 739214 675520 739218
rect 675584 739216 675590 739218
rect 675471 739158 675476 739214
rect 675471 739154 675520 739158
rect 675584 739156 675628 739216
rect 675584 739154 675590 739156
rect 675471 739153 675537 739154
rect 675759 738772 675825 738775
rect 676090 738772 676096 738774
rect 675759 738770 676096 738772
rect 675759 738714 675764 738770
rect 675820 738714 676096 738770
rect 675759 738712 676096 738714
rect 675759 738709 675825 738712
rect 676090 738710 676096 738712
rect 676160 738710 676166 738774
rect 674938 737674 674944 737738
rect 675008 737736 675014 737738
rect 675759 737736 675825 737739
rect 676666 737736 676672 737738
rect 675008 737734 676672 737736
rect 675008 737678 675764 737734
rect 675820 737678 676672 737734
rect 675008 737676 676672 737678
rect 675008 737674 675014 737676
rect 675759 737673 675825 737676
rect 676666 737674 676672 737676
rect 676736 737674 676742 737738
rect 42639 737292 42705 737295
rect 42336 737290 42705 737292
rect 42336 737234 42644 737290
rect 42700 737234 42705 737290
rect 42336 737232 42705 737234
rect 42639 737229 42705 737232
rect 42351 736700 42417 736703
rect 42306 736698 42417 736700
rect 42306 736642 42356 736698
rect 42412 736642 42417 736698
rect 42306 736637 42417 736642
rect 42306 736522 42366 736637
rect 42063 735962 42129 735963
rect 42063 735958 42112 735962
rect 42176 735960 42182 735962
rect 42063 735902 42068 735958
rect 42063 735898 42112 735902
rect 42176 735900 42220 735960
rect 42176 735898 42182 735900
rect 42063 735897 42129 735898
rect 42306 735519 42366 735634
rect 42306 735514 42417 735519
rect 42306 735458 42356 735514
rect 42412 735458 42417 735514
rect 42306 735456 42417 735458
rect 42351 735453 42417 735456
rect 43215 734924 43281 734927
rect 42336 734922 43281 734924
rect 42336 734866 43220 734922
rect 43276 734866 43281 734922
rect 42336 734864 43281 734866
rect 43215 734861 43281 734864
rect 675759 734924 675825 734927
rect 676858 734924 676864 734926
rect 675759 734922 676864 734924
rect 675759 734866 675764 734922
rect 675820 734866 676864 734922
rect 675759 734864 676864 734866
rect 675759 734861 675825 734864
rect 676858 734862 676864 734864
rect 676928 734862 676934 734926
rect 675130 734122 675136 734186
rect 675200 734184 675206 734186
rect 675375 734184 675441 734187
rect 675200 734182 675441 734184
rect 675200 734126 675380 734182
rect 675436 734126 675441 734182
rect 675200 734124 675441 734126
rect 675200 734122 675206 734124
rect 675375 734121 675441 734124
rect 43311 734036 43377 734039
rect 42336 734034 43377 734036
rect 42336 733978 43316 734034
rect 43372 733978 43377 734034
rect 42336 733976 43377 733978
rect 43311 733973 43377 733976
rect 41338 733826 41344 733890
rect 41408 733826 41414 733890
rect 41346 733370 41406 733826
rect 40608 733340 41406 733370
rect 40578 733310 41376 733340
rect 40578 733150 40638 733310
rect 40570 733086 40576 733150
rect 40640 733086 40646 733150
rect 40762 733086 40768 733150
rect 40832 733086 40838 733150
rect 40770 732556 40830 733086
rect 40770 732526 40992 732556
rect 40800 732496 41022 732526
rect 40962 732262 41022 732496
rect 40954 732198 40960 732262
rect 41024 732198 41030 732262
rect 42306 731668 42366 731712
rect 42927 731668 42993 731671
rect 42306 731666 42993 731668
rect 42306 731610 42932 731666
rect 42988 731610 42993 731666
rect 42306 731608 42993 731610
rect 42927 731605 42993 731608
rect 40194 730339 40254 730898
rect 40143 730334 40254 730339
rect 40143 730278 40148 730334
rect 40204 730278 40254 730334
rect 40143 730276 40254 730278
rect 40143 730273 40209 730276
rect 40194 729599 40254 730084
rect 40194 729594 40305 729599
rect 40194 729538 40244 729594
rect 40300 729538 40305 729594
rect 40194 729536 40305 729538
rect 40239 729533 40305 729536
rect 41730 728859 41790 729270
rect 58383 729004 58449 729007
rect 58383 729002 64416 729004
rect 58383 728946 58388 729002
rect 58444 728946 64416 729002
rect 58383 728944 64416 728946
rect 58383 728941 58449 728944
rect 41679 728854 41790 728859
rect 41679 728798 41684 728854
rect 41740 728798 41790 728854
rect 41679 728796 41790 728798
rect 41679 728793 41745 728796
rect 41922 727971 41982 728530
rect 655215 728264 655281 728267
rect 650208 728262 655281 728264
rect 650208 728206 655220 728262
rect 655276 728206 655281 728262
rect 650208 728204 655281 728206
rect 655215 728201 655281 728204
rect 41922 727966 42033 727971
rect 41922 727910 41972 727966
rect 42028 727910 42033 727966
rect 41922 727908 42033 727910
rect 41967 727905 42033 727908
rect 41538 727231 41598 727790
rect 41538 727226 41649 727231
rect 41538 727170 41588 727226
rect 41644 727170 41649 727226
rect 41538 727168 41649 727170
rect 41583 727165 41649 727168
rect 37314 726343 37374 726902
rect 37314 726338 37425 726343
rect 37314 726282 37364 726338
rect 37420 726282 37425 726338
rect 37314 726280 37425 726282
rect 37359 726277 37425 726280
rect 41730 725899 41790 726162
rect 41730 725894 41841 725899
rect 42063 725898 42129 725899
rect 42063 725896 42112 725898
rect 41730 725838 41780 725894
rect 41836 725838 41841 725894
rect 41730 725836 41841 725838
rect 42020 725894 42112 725896
rect 42020 725838 42068 725894
rect 42020 725836 42112 725838
rect 41775 725833 41841 725836
rect 42063 725834 42112 725836
rect 42176 725834 42182 725898
rect 42063 725833 42129 725834
rect 42114 724715 42174 725274
rect 42063 724710 42174 724715
rect 42063 724654 42068 724710
rect 42124 724654 42174 724710
rect 42063 724652 42174 724654
rect 42063 724649 42129 724652
rect 42114 724123 42174 724534
rect 42114 724118 42225 724123
rect 42114 724062 42164 724118
rect 42220 724062 42225 724118
rect 42114 724060 42225 724062
rect 42159 724057 42225 724060
rect 42682 723824 42688 723826
rect 42336 723764 42688 723824
rect 42682 723762 42688 723764
rect 42752 723762 42758 723826
rect 42306 722642 42366 723054
rect 42298 722578 42304 722642
rect 42368 722578 42374 722642
rect 674415 722492 674481 722495
rect 674415 722490 674784 722492
rect 674415 722434 674420 722490
rect 674476 722434 674784 722490
rect 674415 722432 674784 722434
rect 674415 722429 674481 722432
rect 43023 722196 43089 722199
rect 42336 722194 43089 722196
rect 42336 722138 43028 722194
rect 43084 722138 43089 722194
rect 42336 722136 43089 722138
rect 43023 722133 43089 722136
rect 674415 721752 674481 721755
rect 674415 721750 674784 721752
rect 674415 721694 674420 721750
rect 674476 721694 674784 721750
rect 674415 721692 674784 721694
rect 674415 721689 674481 721692
rect 41346 720866 41406 721426
rect 41338 720802 41344 720866
rect 41408 720802 41414 720866
rect 674415 720864 674481 720867
rect 674415 720862 674784 720864
rect 674415 720806 674420 720862
rect 674476 720806 674784 720862
rect 674415 720804 674784 720806
rect 674415 720801 674481 720804
rect 43311 720568 43377 720571
rect 42336 720566 43377 720568
rect 42336 720510 43316 720566
rect 43372 720510 43377 720566
rect 42336 720508 43377 720510
rect 43311 720505 43377 720508
rect 673743 720568 673809 720571
rect 673743 720566 674814 720568
rect 673743 720510 673748 720566
rect 673804 720510 674814 720566
rect 673743 720508 674814 720510
rect 673743 720505 673809 720508
rect 674754 720094 674814 720508
rect 674415 719236 674481 719239
rect 674415 719234 674784 719236
rect 674415 719178 674420 719234
rect 674476 719178 674784 719234
rect 674415 719176 674784 719178
rect 674415 719173 674481 719176
rect 43311 719088 43377 719091
rect 42336 719086 43377 719088
rect 42336 719030 43316 719086
rect 43372 719030 43377 719086
rect 42336 719028 43377 719030
rect 43311 719025 43377 719028
rect 672687 718496 672753 718499
rect 673647 718496 673713 718499
rect 674754 718496 674814 718540
rect 672687 718494 674814 718496
rect 672687 718438 672692 718494
rect 672748 718438 673652 718494
rect 673708 718438 674814 718494
rect 672687 718436 674814 718438
rect 672687 718433 672753 718436
rect 673647 718433 673713 718436
rect 674415 717756 674481 717759
rect 674415 717754 674784 717756
rect 674415 717698 674420 717754
rect 674476 717698 674784 717754
rect 674415 717696 674784 717698
rect 674415 717693 674481 717696
rect 676474 717102 676480 717166
rect 676544 717102 676550 717166
rect 37359 717016 37425 717019
rect 40378 717016 40384 717018
rect 37359 717014 40384 717016
rect 37359 716958 37364 717014
rect 37420 716958 40384 717014
rect 37359 716956 40384 716958
rect 37359 716953 37425 716956
rect 40378 716954 40384 716956
rect 40448 716954 40454 717018
rect 676482 716912 676542 717102
rect 40239 716720 40305 716723
rect 41146 716720 41152 716722
rect 40239 716718 41152 716720
rect 40239 716662 40244 716718
rect 40300 716662 41152 716718
rect 40239 716660 41152 716662
rect 40239 716657 40305 716660
rect 41146 716658 41152 716660
rect 41216 716658 41222 716722
rect 654447 716424 654513 716427
rect 650208 716422 654513 716424
rect 650208 716366 654452 716422
rect 654508 716366 654513 716422
rect 650208 716364 654513 716366
rect 654447 716361 654513 716364
rect 41530 716066 41536 716130
rect 41600 716128 41606 716130
rect 41967 716128 42033 716131
rect 41600 716126 42033 716128
rect 41600 716070 41972 716126
rect 42028 716070 42033 716126
rect 41600 716068 42033 716070
rect 41600 716066 41606 716068
rect 41967 716065 42033 716068
rect 674223 716128 674289 716131
rect 674223 716126 674784 716128
rect 674223 716070 674228 716126
rect 674284 716070 674784 716126
rect 674223 716068 674784 716070
rect 674223 716065 674289 716068
rect 676282 715770 676288 715834
rect 676352 715770 676358 715834
rect 676290 715284 676350 715770
rect 58383 714648 58449 714651
rect 58383 714646 64416 714648
rect 58383 714590 58388 714646
rect 58444 714590 64416 714646
rect 58383 714588 64416 714590
rect 58383 714585 58449 714588
rect 674031 714500 674097 714503
rect 674031 714498 674784 714500
rect 674031 714442 674036 714498
rect 674092 714442 674784 714498
rect 674031 714440 674784 714442
rect 674031 714437 674097 714440
rect 674991 714056 675057 714059
rect 674946 714054 675057 714056
rect 674946 713998 674996 714054
rect 675052 713998 675057 714054
rect 674946 713993 675057 713998
rect 41871 713910 41937 713911
rect 41871 713908 41920 713910
rect 41828 713906 41920 713908
rect 41828 713850 41876 713906
rect 41828 713848 41920 713850
rect 41871 713846 41920 713848
rect 41984 713846 41990 713910
rect 42063 713908 42129 713911
rect 42490 713908 42496 713910
rect 42063 713906 42496 713908
rect 42063 713850 42068 713906
rect 42124 713850 42496 713906
rect 42063 713848 42496 713850
rect 41871 713845 41937 713846
rect 42063 713845 42129 713848
rect 42490 713846 42496 713848
rect 42560 713846 42566 713910
rect 674946 713730 675006 713993
rect 674319 713020 674385 713023
rect 674319 713018 674784 713020
rect 674319 712962 674324 713018
rect 674380 712962 674784 713018
rect 674319 712960 674784 712962
rect 674319 712957 674385 712960
rect 673978 712070 673984 712134
rect 674048 712132 674054 712134
rect 674048 712072 674784 712132
rect 674048 712070 674054 712072
rect 675898 711922 675904 711986
rect 675968 711922 675974 711986
rect 41871 711690 41937 711691
rect 41871 711688 41920 711690
rect 41828 711686 41920 711688
rect 41828 711630 41876 711686
rect 41828 711628 41920 711630
rect 41871 711626 41920 711628
rect 41984 711626 41990 711690
rect 41871 711625 41937 711626
rect 675906 711362 675966 711922
rect 42490 710738 42496 710802
rect 42560 710800 42566 710802
rect 42831 710800 42897 710803
rect 42560 710798 42897 710800
rect 42560 710742 42836 710798
rect 42892 710742 42897 710798
rect 42560 710740 42897 710742
rect 42560 710738 42566 710740
rect 42831 710737 42897 710740
rect 674415 710504 674481 710507
rect 674415 710502 674784 710504
rect 674415 710446 674420 710502
rect 674476 710446 674784 710502
rect 674415 710444 674784 710446
rect 674415 710441 674481 710444
rect 674799 709912 674865 709915
rect 674754 709910 674865 709912
rect 674754 709854 674804 709910
rect 674860 709854 674865 709910
rect 674754 709849 674865 709854
rect 674754 709734 674814 709849
rect 674415 709024 674481 709027
rect 674415 709022 674784 709024
rect 674415 708966 674420 709022
rect 674476 708966 674784 709022
rect 674415 708964 674784 708966
rect 674415 708961 674481 708964
rect 41338 708518 41344 708582
rect 41408 708580 41414 708582
rect 41775 708580 41841 708583
rect 41408 708578 41841 708580
rect 41408 708522 41780 708578
rect 41836 708522 41841 708578
rect 41408 708520 41841 708522
rect 41408 708518 41414 708520
rect 41775 708517 41841 708520
rect 677050 708370 677056 708434
rect 677120 708370 677126 708434
rect 677058 708254 677118 708370
rect 42159 707840 42225 707843
rect 42682 707840 42688 707842
rect 42159 707838 42688 707840
rect 42159 707782 42164 707838
rect 42220 707782 42688 707838
rect 42159 707780 42688 707782
rect 42159 707777 42225 707780
rect 42682 707778 42688 707780
rect 42752 707778 42758 707842
rect 674415 707396 674481 707399
rect 674415 707394 674784 707396
rect 674415 707338 674420 707394
rect 674476 707338 674784 707394
rect 674415 707336 674784 707338
rect 674415 707333 674481 707336
rect 41530 706742 41536 706806
rect 41600 706804 41606 706806
rect 41775 706804 41841 706807
rect 674799 706804 674865 706807
rect 41600 706802 41841 706804
rect 41600 706746 41780 706802
rect 41836 706746 41841 706802
rect 41600 706744 41841 706746
rect 41600 706742 41606 706744
rect 41775 706741 41841 706744
rect 674754 706802 674865 706804
rect 674754 706746 674804 706802
rect 674860 706746 674865 706802
rect 674754 706741 674865 706746
rect 674754 706626 674814 706741
rect 42159 706212 42225 706215
rect 42298 706212 42304 706214
rect 42159 706210 42304 706212
rect 42159 706154 42164 706210
rect 42220 706154 42304 706210
rect 42159 706152 42304 706154
rect 42159 706149 42225 706152
rect 42298 706150 42304 706152
rect 42368 706150 42374 706214
rect 650223 705472 650289 705475
rect 650178 705470 650289 705472
rect 650178 705414 650228 705470
rect 650284 705414 650289 705470
rect 650178 705409 650289 705414
rect 650178 704850 650238 705409
rect 679746 705179 679806 705738
rect 679695 705174 679806 705179
rect 679695 705118 679700 705174
rect 679756 705118 679806 705174
rect 679695 705116 679806 705118
rect 679695 705113 679761 705116
rect 41775 704734 41841 704735
rect 41338 704670 41344 704734
rect 41408 704732 41414 704734
rect 41722 704732 41728 704734
rect 41408 704672 41728 704732
rect 41792 704730 41841 704734
rect 41836 704674 41841 704730
rect 41408 704670 41414 704672
rect 41722 704670 41728 704672
rect 41792 704670 41841 704674
rect 41775 704669 41841 704670
rect 679695 704584 679761 704587
rect 679695 704582 679806 704584
rect 679695 704526 679700 704582
rect 679756 704526 679806 704582
rect 679695 704521 679806 704526
rect 679746 704258 679806 704521
rect 41530 704078 41536 704142
rect 41600 704140 41606 704142
rect 41775 704140 41841 704143
rect 42106 704140 42112 704142
rect 41600 704138 42112 704140
rect 41600 704082 41780 704138
rect 41836 704082 42112 704138
rect 41600 704080 42112 704082
rect 41600 704078 41606 704080
rect 41775 704077 41841 704080
rect 42106 704078 42112 704080
rect 42176 704078 42182 704142
rect 41146 703634 41152 703698
rect 41216 703696 41222 703698
rect 42255 703696 42321 703699
rect 41216 703694 42321 703696
rect 41216 703638 42260 703694
rect 42316 703638 42321 703694
rect 41216 703636 42321 703638
rect 41216 703634 41222 703636
rect 42255 703633 42321 703636
rect 40378 703486 40384 703550
rect 40448 703548 40454 703550
rect 42831 703548 42897 703551
rect 40448 703546 42897 703548
rect 40448 703490 42836 703546
rect 42892 703490 42897 703546
rect 40448 703488 42897 703490
rect 40448 703486 40454 703488
rect 42831 703485 42897 703488
rect 675898 703042 675904 703106
rect 675968 703104 675974 703106
rect 676282 703104 676288 703106
rect 675968 703044 676288 703104
rect 675968 703042 675974 703044
rect 676282 703042 676288 703044
rect 676352 703042 676358 703106
rect 674991 702512 675057 702515
rect 676090 702512 676096 702514
rect 674991 702510 676096 702512
rect 674991 702454 674996 702510
rect 675052 702454 676096 702510
rect 674991 702452 676096 702454
rect 674991 702449 675057 702452
rect 676090 702450 676096 702452
rect 676160 702450 676166 702514
rect 42255 700884 42321 700887
rect 42255 700882 42366 700884
rect 42255 700826 42260 700882
rect 42316 700826 42366 700882
rect 42255 700821 42366 700826
rect 42306 700591 42366 700821
rect 42255 700586 42366 700591
rect 42255 700530 42260 700586
rect 42316 700530 42366 700586
rect 42255 700528 42366 700530
rect 42255 700525 42321 700528
rect 57807 700292 57873 700295
rect 57807 700290 64416 700292
rect 57807 700234 57812 700290
rect 57868 700234 64416 700290
rect 57807 700232 64416 700234
rect 57807 700229 57873 700232
rect 675375 697926 675441 697927
rect 675322 697924 675328 697926
rect 675284 697864 675328 697924
rect 675392 697922 675441 697926
rect 675436 697866 675441 697922
rect 675322 697862 675328 697864
rect 675392 697862 675441 697866
rect 675375 697861 675441 697862
rect 673978 697270 673984 697334
rect 674048 697332 674054 697334
rect 675471 697332 675537 697335
rect 674048 697330 675537 697332
rect 674048 697274 675476 697330
rect 675532 697274 675537 697330
rect 674048 697272 675537 697274
rect 674048 697270 674054 697272
rect 675471 697269 675537 697272
rect 675759 697184 675825 697187
rect 675898 697184 675904 697186
rect 675759 697182 675904 697184
rect 675759 697126 675764 697182
rect 675820 697126 675904 697182
rect 675759 697124 675904 697126
rect 675759 697121 675825 697124
rect 675898 697122 675904 697124
rect 675968 697122 675974 697186
rect 675471 694818 675537 694819
rect 675471 694814 675520 694818
rect 675584 694816 675590 694818
rect 675471 694758 675476 694814
rect 675471 694754 675520 694758
rect 675584 694756 675628 694816
rect 675584 694754 675590 694756
rect 675471 694753 675537 694754
rect 674938 694310 674944 694374
rect 675008 694372 675014 694374
rect 675279 694372 675345 694375
rect 675008 694370 675345 694372
rect 675008 694314 675284 694370
rect 675340 694314 675345 694370
rect 675008 694312 675345 694314
rect 675008 694310 675014 694312
rect 675279 694309 675345 694312
rect 675759 694372 675825 694375
rect 676666 694372 676672 694374
rect 675759 694370 676672 694372
rect 675759 694314 675764 694370
rect 675820 694314 676672 694370
rect 675759 694312 676672 694314
rect 675759 694309 675825 694312
rect 676666 694310 676672 694312
rect 676736 694310 676742 694374
rect 42639 694076 42705 694079
rect 42336 694074 42705 694076
rect 42336 694018 42644 694074
rect 42700 694018 42705 694074
rect 42336 694016 42705 694018
rect 42639 694013 42705 694016
rect 42351 693484 42417 693487
rect 42306 693482 42417 693484
rect 42306 693426 42356 693482
rect 42412 693426 42417 693482
rect 42306 693421 42417 693426
rect 674938 693422 674944 693486
rect 675008 693484 675014 693486
rect 675471 693484 675537 693487
rect 675008 693482 675537 693484
rect 675008 693426 675476 693482
rect 675532 693426 675537 693482
rect 675008 693424 675537 693426
rect 675008 693422 675014 693424
rect 675471 693421 675537 693424
rect 42306 693306 42366 693421
rect 654447 693040 654513 693043
rect 650208 693038 654513 693040
rect 650208 692982 654452 693038
rect 654508 692982 654513 693038
rect 650208 692980 654513 692982
rect 654447 692977 654513 692980
rect 41391 692746 41457 692747
rect 41338 692744 41344 692746
rect 41300 692684 41344 692744
rect 41408 692742 41457 692746
rect 41452 692686 41457 692742
rect 41338 692682 41344 692684
rect 41408 692682 41457 692686
rect 41391 692681 41457 692682
rect 42639 692448 42705 692451
rect 42336 692446 42705 692448
rect 42336 692390 42644 692446
rect 42700 692390 42705 692446
rect 42336 692388 42705 692390
rect 42639 692385 42705 692388
rect 675375 692004 675441 692007
rect 676282 692004 676288 692006
rect 675375 692002 676288 692004
rect 675375 691946 675380 692002
rect 675436 691946 676288 692002
rect 675375 691944 676288 691946
rect 675375 691941 675441 691944
rect 676282 691942 676288 691944
rect 676352 691942 676358 692006
rect 43503 691708 43569 691711
rect 42336 691706 43569 691708
rect 42336 691650 43508 691706
rect 43564 691650 43569 691706
rect 42336 691648 43569 691650
rect 43503 691645 43569 691648
rect 43215 690820 43281 690823
rect 42336 690818 43281 690820
rect 42336 690762 43220 690818
rect 43276 690762 43281 690818
rect 42336 690760 43281 690762
rect 43215 690757 43281 690760
rect 40570 690314 40576 690378
rect 40640 690314 40646 690378
rect 40578 690228 40638 690314
rect 40578 690198 42336 690228
rect 40608 690168 42366 690198
rect 42306 689638 42366 690168
rect 40954 689574 40960 689638
rect 41024 689574 41030 689638
rect 42298 689574 42304 689638
rect 42368 689574 42374 689638
rect 40962 689340 41022 689574
rect 674170 689426 674176 689490
rect 674240 689488 674246 689490
rect 675706 689488 675712 689490
rect 674240 689428 675712 689488
rect 674240 689426 674246 689428
rect 675706 689426 675712 689428
rect 675776 689426 675782 689490
rect 40962 689310 42144 689340
rect 40992 689280 42174 689310
rect 42114 688750 42174 689280
rect 42106 688686 42112 688750
rect 42176 688686 42182 688750
rect 41922 688307 41982 688496
rect 41871 688302 41982 688307
rect 41871 688246 41876 688302
rect 41932 688246 41982 688302
rect 41871 688244 41982 688246
rect 674895 688304 674961 688307
rect 677050 688304 677056 688306
rect 674895 688302 677056 688304
rect 674895 688246 674900 688302
rect 674956 688246 677056 688302
rect 674895 688244 677056 688246
rect 41871 688241 41937 688244
rect 674895 688241 674961 688244
rect 677050 688242 677056 688244
rect 677120 688242 677126 688306
rect 40194 687123 40254 687682
rect 40194 687118 40305 687123
rect 40194 687062 40244 687118
rect 40300 687062 40305 687118
rect 40194 687060 40305 687062
rect 40239 687057 40305 687060
rect 40578 686382 40638 686868
rect 40570 686318 40576 686382
rect 40640 686318 40646 686382
rect 42735 686084 42801 686087
rect 42336 686082 42801 686084
rect 42336 686026 42740 686082
rect 42796 686026 42801 686082
rect 42336 686024 42801 686026
rect 42735 686021 42801 686024
rect 59535 685936 59601 685939
rect 59535 685934 64416 685936
rect 59535 685878 59540 685934
rect 59596 685878 64416 685934
rect 59535 685876 64416 685878
rect 59535 685873 59601 685876
rect 675087 685640 675153 685643
rect 677050 685640 677056 685642
rect 675087 685638 677056 685640
rect 675087 685582 675092 685638
rect 675148 685582 677056 685638
rect 675087 685580 677056 685582
rect 675087 685577 675153 685580
rect 677050 685578 677056 685580
rect 677120 685578 677126 685642
rect 42114 684903 42174 685388
rect 42063 684898 42174 684903
rect 42063 684842 42068 684898
rect 42124 684842 42174 684898
rect 42063 684840 42174 684842
rect 42063 684837 42129 684840
rect 41730 684015 41790 684574
rect 41730 684010 41841 684015
rect 41730 683954 41780 684010
rect 41836 683954 41841 684010
rect 41730 683952 41841 683954
rect 41775 683949 41841 683952
rect 40962 683274 41022 683760
rect 40954 683210 40960 683274
rect 41024 683210 41030 683274
rect 42114 682683 42174 682946
rect 42114 682678 42225 682683
rect 42114 682622 42164 682678
rect 42220 682622 42225 682678
rect 42114 682620 42225 682622
rect 42159 682617 42225 682620
rect 42306 681499 42366 682058
rect 42255 681494 42366 681499
rect 42255 681438 42260 681494
rect 42316 681438 42366 681494
rect 42255 681436 42366 681438
rect 42255 681433 42321 681436
rect 655407 681348 655473 681351
rect 650208 681346 655473 681348
rect 41730 680906 41790 681318
rect 650208 681290 655412 681346
rect 655468 681290 655473 681346
rect 650208 681288 655473 681290
rect 655407 681285 655473 681288
rect 41722 680842 41728 680906
rect 41792 680842 41798 680906
rect 41346 680019 41406 680578
rect 41295 680014 41406 680019
rect 41295 679958 41300 680014
rect 41356 679958 41406 680014
rect 41295 679956 41406 679958
rect 41295 679953 41361 679956
rect 41922 679575 41982 679838
rect 674170 679658 674176 679722
rect 674240 679720 674246 679722
rect 674415 679720 674481 679723
rect 674240 679718 674481 679720
rect 674240 679662 674420 679718
rect 674476 679662 674481 679718
rect 674240 679660 674481 679662
rect 674240 679658 674246 679660
rect 674415 679657 674481 679660
rect 674991 679720 675057 679723
rect 676474 679720 676480 679722
rect 674991 679718 676480 679720
rect 674991 679662 674996 679718
rect 675052 679662 676480 679718
rect 674991 679660 676480 679662
rect 674991 679657 675057 679660
rect 676474 679658 676480 679660
rect 676544 679658 676550 679722
rect 41922 679570 42033 679575
rect 41922 679514 41972 679570
rect 42028 679514 42033 679570
rect 41922 679512 42033 679514
rect 41967 679509 42033 679512
rect 674031 679572 674097 679575
rect 674991 679574 675057 679575
rect 674170 679572 674176 679574
rect 674031 679570 674176 679572
rect 674031 679514 674036 679570
rect 674092 679514 674176 679570
rect 674031 679512 674176 679514
rect 674031 679509 674097 679512
rect 674170 679510 674176 679512
rect 674240 679510 674246 679574
rect 674938 679572 674944 679574
rect 674900 679512 674944 679572
rect 675008 679570 675057 679574
rect 675855 679574 675921 679575
rect 675855 679572 675904 679574
rect 675052 679514 675057 679570
rect 674938 679510 674944 679512
rect 675008 679510 675057 679514
rect 675812 679570 675904 679572
rect 675812 679514 675860 679570
rect 675812 679512 675904 679514
rect 674991 679509 675057 679510
rect 675855 679510 675904 679512
rect 675968 679510 675974 679574
rect 675855 679509 675921 679510
rect 42306 678388 42366 678950
rect 42490 678388 42496 678390
rect 42306 678328 42496 678388
rect 42490 678326 42496 678328
rect 42560 678326 42566 678390
rect 43119 678240 43185 678243
rect 42336 678238 43185 678240
rect 42336 678182 43124 678238
rect 43180 678182 43185 678238
rect 42336 678180 43185 678182
rect 43119 678177 43185 678180
rect 674415 677352 674481 677355
rect 674415 677350 674784 677352
rect 42306 677207 42366 677322
rect 674415 677294 674420 677350
rect 674476 677294 674784 677350
rect 674415 677292 674784 677294
rect 674415 677289 674481 677292
rect 42306 677202 42417 677207
rect 42306 677146 42356 677202
rect 42412 677146 42417 677202
rect 42306 677144 42417 677146
rect 42351 677141 42417 677144
rect 674415 676464 674481 676467
rect 674415 676462 674784 676464
rect 674415 676406 674420 676462
rect 674476 676406 674784 676462
rect 674415 676404 674784 676406
rect 674415 676401 674481 676404
rect 42306 675727 42366 675842
rect 42306 675722 42417 675727
rect 42306 675666 42356 675722
rect 42412 675666 42417 675722
rect 42306 675664 42417 675666
rect 42351 675661 42417 675664
rect 674415 675724 674481 675727
rect 674415 675722 674784 675724
rect 674415 675666 674420 675722
rect 674476 675666 674784 675722
rect 674415 675664 674784 675666
rect 674415 675661 674481 675664
rect 674938 675366 674944 675430
rect 675008 675428 675014 675430
rect 675322 675428 675328 675430
rect 675008 675368 675328 675428
rect 675008 675366 675014 675368
rect 675322 675366 675328 675368
rect 675392 675366 675398 675430
rect 674415 674836 674481 674839
rect 674415 674834 674784 674836
rect 674415 674778 674420 674834
rect 674476 674778 674784 674834
rect 674415 674776 674784 674778
rect 674415 674773 674481 674776
rect 674415 674096 674481 674099
rect 674415 674094 674784 674096
rect 674415 674038 674420 674094
rect 674476 674038 674784 674094
rect 674415 674036 674784 674038
rect 674415 674033 674481 674036
rect 672687 673356 672753 673359
rect 672687 673354 674784 673356
rect 672687 673298 672692 673354
rect 672748 673298 674784 673354
rect 672687 673296 674784 673298
rect 672687 673293 672753 673296
rect 675138 672323 675198 672512
rect 674746 672258 674752 672322
rect 674816 672258 674822 672322
rect 675138 672318 675249 672323
rect 675138 672262 675188 672318
rect 675244 672262 675249 672318
rect 675138 672260 675249 672262
rect 674754 671698 674814 672258
rect 675183 672257 675249 672260
rect 59439 671580 59505 671583
rect 59439 671578 64416 671580
rect 59439 671522 59444 671578
rect 59500 671522 64416 671578
rect 59439 671520 64416 671522
rect 59439 671517 59505 671520
rect 674746 671518 674752 671582
rect 674816 671580 674822 671582
rect 674991 671580 675057 671583
rect 674816 671578 675057 671580
rect 674816 671522 674996 671578
rect 675052 671522 675057 671578
rect 674816 671520 675057 671522
rect 674816 671518 674822 671520
rect 674991 671517 675057 671520
rect 675087 671286 675153 671287
rect 675087 671284 675136 671286
rect 675044 671282 675136 671284
rect 675044 671226 675092 671282
rect 675044 671224 675136 671226
rect 675087 671222 675136 671224
rect 675200 671222 675206 671286
rect 675087 671221 675153 671222
rect 674703 671136 674769 671139
rect 674703 671134 674814 671136
rect 674703 671078 674708 671134
rect 674764 671078 674814 671134
rect 674703 671073 674814 671078
rect 41391 670990 41457 670991
rect 41338 670926 41344 670990
rect 41408 670988 41457 670990
rect 42639 670988 42705 670991
rect 42874 670988 42880 670990
rect 41408 670986 41500 670988
rect 41452 670930 41500 670986
rect 41408 670928 41500 670930
rect 42639 670986 42880 670988
rect 42639 670930 42644 670986
rect 42700 670930 42880 670986
rect 42639 670928 42880 670930
rect 41408 670926 41457 670928
rect 41391 670925 41457 670926
rect 42639 670925 42705 670928
rect 42874 670926 42880 670928
rect 42944 670926 42950 670990
rect 674754 670884 674814 671073
rect 41914 670778 41920 670842
rect 41984 670840 41990 670842
rect 42682 670840 42688 670842
rect 41984 670780 42688 670840
rect 41984 670778 41990 670780
rect 42682 670778 42688 670780
rect 42752 670778 42758 670842
rect 42159 670692 42225 670695
rect 675087 670694 675153 670695
rect 42682 670692 42688 670694
rect 42159 670690 42688 670692
rect 42159 670634 42164 670690
rect 42220 670634 42688 670690
rect 42159 670632 42688 670634
rect 42159 670629 42225 670632
rect 42682 670630 42688 670632
rect 42752 670630 42758 670694
rect 675087 670690 675136 670694
rect 675200 670692 675206 670694
rect 675087 670634 675092 670690
rect 675087 670630 675136 670634
rect 675200 670632 675244 670692
rect 675200 670630 675206 670632
rect 675322 670630 675328 670694
rect 675392 670692 675398 670694
rect 675855 670692 675921 670695
rect 675392 670690 675921 670692
rect 675392 670634 675860 670690
rect 675916 670634 675921 670690
rect 675392 670632 675921 670634
rect 675392 670630 675398 670632
rect 675087 670629 675153 670630
rect 675855 670629 675921 670632
rect 674554 670482 674560 670546
rect 674624 670544 674630 670546
rect 674624 670484 674814 670544
rect 674624 670482 674630 670484
rect 674031 670396 674097 670399
rect 674554 670396 674560 670398
rect 674031 670394 674560 670396
rect 674031 670338 674036 670394
rect 674092 670338 674560 670394
rect 674031 670336 674560 670338
rect 674031 670333 674097 670336
rect 674554 670334 674560 670336
rect 674624 670334 674630 670398
rect 674754 670070 674814 670484
rect 654447 669508 654513 669511
rect 650208 669506 654513 669508
rect 650208 669450 654452 669506
rect 654508 669450 654513 669506
rect 650208 669448 654513 669450
rect 654447 669445 654513 669448
rect 42447 669360 42513 669363
rect 42447 669358 42558 669360
rect 42447 669302 42452 669358
rect 42508 669302 42558 669358
rect 42447 669297 42558 669302
rect 42498 668919 42558 669297
rect 674362 669224 674368 669288
rect 674432 669286 674438 669288
rect 674432 669226 674784 669286
rect 674432 669224 674438 669226
rect 42498 668914 42609 668919
rect 42498 668858 42548 668914
rect 42604 668858 42609 668914
rect 42498 668856 42609 668858
rect 42543 668853 42609 668856
rect 42543 668770 42609 668771
rect 42490 668706 42496 668770
rect 42560 668768 42609 668770
rect 674511 668768 674577 668771
rect 42560 668766 42652 668768
rect 42604 668710 42652 668766
rect 42560 668708 42652 668710
rect 674511 668766 674814 668768
rect 674511 668710 674516 668766
rect 674572 668710 674814 668766
rect 674511 668708 674814 668710
rect 42560 668706 42609 668708
rect 42543 668705 42609 668706
rect 674511 668705 674577 668708
rect 674754 668590 674814 668708
rect 674607 668028 674673 668031
rect 674607 668026 674814 668028
rect 674607 667970 674612 668026
rect 674668 667970 674814 668026
rect 674607 667968 674814 667970
rect 674607 667965 674673 667968
rect 674754 667776 674814 667968
rect 675706 667522 675712 667586
rect 675776 667522 675782 667586
rect 675714 666962 675774 667522
rect 41775 666698 41841 666699
rect 41722 666634 41728 666698
rect 41792 666696 41841 666698
rect 41792 666694 41884 666696
rect 41836 666638 41884 666694
rect 41792 666636 41884 666638
rect 41792 666634 41841 666636
rect 676090 666634 676096 666698
rect 676160 666634 676166 666698
rect 41775 666633 41841 666634
rect 42682 666486 42688 666550
rect 42752 666548 42758 666550
rect 42831 666548 42897 666551
rect 42752 666546 42897 666548
rect 42752 666490 42836 666546
rect 42892 666490 42897 666546
rect 42752 666488 42897 666490
rect 42752 666486 42758 666488
rect 42831 666485 42897 666488
rect 676098 666074 676158 666634
rect 676474 665894 676480 665958
rect 676544 665894 676550 665958
rect 41338 665450 41344 665514
rect 41408 665512 41414 665514
rect 41408 665452 41598 665512
rect 41408 665450 41414 665452
rect 41538 665366 41598 665452
rect 41530 665302 41536 665366
rect 41600 665302 41606 665366
rect 676482 665334 676542 665894
rect 41530 665006 41536 665070
rect 41600 665068 41606 665070
rect 42682 665068 42688 665070
rect 41600 665008 42688 665068
rect 41600 665006 41606 665008
rect 42682 665006 42688 665008
rect 42752 665006 42758 665070
rect 42874 664710 42880 664774
rect 42944 664772 42950 664774
rect 43023 664772 43089 664775
rect 42944 664770 43089 664772
rect 42944 664714 43028 664770
rect 43084 664714 43089 664770
rect 42944 664712 43089 664714
rect 42944 664710 42950 664712
rect 43023 664709 43089 664712
rect 674127 664476 674193 664479
rect 674127 664474 674784 664476
rect 674127 664418 674132 664474
rect 674188 664418 674784 664474
rect 674127 664416 674784 664418
rect 674127 664413 674193 664416
rect 675130 664266 675136 664330
rect 675200 664266 675206 664330
rect 675138 663854 675198 664266
rect 677242 663526 677248 663590
rect 677312 663526 677318 663590
rect 677250 662966 677310 663526
rect 676858 662342 676864 662406
rect 676928 662342 676934 662406
rect 676866 662226 676926 662342
rect 42159 661516 42225 661519
rect 42682 661516 42688 661518
rect 42159 661514 42688 661516
rect 42159 661458 42164 661514
rect 42220 661458 42688 661514
rect 42159 661456 42688 661458
rect 42159 661453 42225 661456
rect 42682 661454 42688 661456
rect 42752 661454 42758 661518
rect 674415 661368 674481 661371
rect 674415 661366 674784 661368
rect 674415 661310 674420 661366
rect 674476 661310 674784 661366
rect 674415 661308 674784 661310
rect 674415 661305 674481 661308
rect 41871 660778 41937 660779
rect 41871 660776 41920 660778
rect 41828 660774 41920 660776
rect 41828 660718 41876 660774
rect 41828 660716 41920 660718
rect 41871 660714 41920 660716
rect 41984 660714 41990 660778
rect 41871 660713 41937 660714
rect 679746 660039 679806 660598
rect 679695 660034 679806 660039
rect 679695 659978 679700 660034
rect 679756 659978 679806 660034
rect 679695 659976 679806 659978
rect 679695 659973 679761 659976
rect 679695 659296 679761 659299
rect 679695 659294 679806 659296
rect 679695 659238 679700 659294
rect 679756 659238 679806 659294
rect 679695 659233 679806 659238
rect 679746 659118 679806 659233
rect 652239 658556 652305 658559
rect 650178 658554 652305 658556
rect 650178 658498 652244 658554
rect 652300 658498 652305 658554
rect 650178 658496 652305 658498
rect 650178 657934 650238 658496
rect 652239 658493 652305 658496
rect 674746 658346 674752 658410
rect 674816 658408 674822 658410
rect 676474 658408 676480 658410
rect 674816 658348 676480 658408
rect 674816 658346 674822 658348
rect 676474 658346 676480 658348
rect 676544 658346 676550 658410
rect 59535 657224 59601 657227
rect 59535 657222 64416 657224
rect 59535 657166 59540 657222
rect 59596 657166 64416 657222
rect 59535 657164 64416 657166
rect 59535 657161 59601 657164
rect 40954 656718 40960 656782
rect 41024 656780 41030 656782
rect 41775 656780 41841 656783
rect 41024 656778 41841 656780
rect 41024 656722 41780 656778
rect 41836 656722 41841 656778
rect 41024 656720 41841 656722
rect 41024 656718 41030 656720
rect 41775 656717 41841 656720
rect 40570 656126 40576 656190
rect 40640 656188 40646 656190
rect 41775 656188 41841 656191
rect 40640 656186 41841 656188
rect 40640 656130 41780 656186
rect 41836 656130 41841 656186
rect 40640 656128 41841 656130
rect 40640 656126 40646 656128
rect 41775 656125 41841 656128
rect 675759 652636 675825 652639
rect 675898 652636 675904 652638
rect 675759 652634 675904 652636
rect 675759 652578 675764 652634
rect 675820 652578 675904 652634
rect 675759 652576 675904 652578
rect 675759 652573 675825 652576
rect 675898 652574 675904 652576
rect 675968 652574 675974 652638
rect 674170 652130 674176 652194
rect 674240 652192 674246 652194
rect 675471 652192 675537 652195
rect 674240 652190 675537 652192
rect 674240 652134 675476 652190
rect 675532 652134 675537 652190
rect 674240 652132 675537 652134
rect 674240 652130 674246 652132
rect 675471 652129 675537 652132
rect 675130 651390 675136 651454
rect 675200 651452 675206 651454
rect 675471 651452 675537 651455
rect 675200 651450 675537 651452
rect 675200 651394 675476 651450
rect 675532 651394 675537 651450
rect 675200 651392 675537 651394
rect 675200 651390 675206 651392
rect 675471 651389 675537 651392
rect 675183 651008 675249 651011
rect 676282 651008 676288 651010
rect 675183 651006 676288 651008
rect 675183 650950 675188 651006
rect 675244 650950 676288 651006
rect 675183 650948 676288 650950
rect 675183 650945 675249 650948
rect 676282 650946 676288 650948
rect 676352 650946 676358 651010
rect 42831 650860 42897 650863
rect 42336 650858 42897 650860
rect 42336 650802 42836 650858
rect 42892 650802 42897 650858
rect 42336 650800 42897 650802
rect 42831 650797 42897 650800
rect 42306 649824 42366 650090
rect 42447 649824 42513 649827
rect 42306 649822 42513 649824
rect 42306 649766 42452 649822
rect 42508 649766 42513 649822
rect 42306 649764 42513 649766
rect 42447 649761 42513 649764
rect 675759 649676 675825 649679
rect 676090 649676 676096 649678
rect 675759 649674 676096 649676
rect 675759 649618 675764 649674
rect 675820 649618 676096 649674
rect 675759 649616 676096 649618
rect 675759 649613 675825 649616
rect 676090 649614 676096 649616
rect 676160 649614 676166 649678
rect 42447 649528 42513 649531
rect 42306 649526 42513 649528
rect 42306 649470 42452 649526
rect 42508 649470 42513 649526
rect 42306 649468 42513 649470
rect 42306 649202 42366 649468
rect 42447 649465 42513 649468
rect 43215 648492 43281 648495
rect 42336 648490 43281 648492
rect 42336 648434 43220 648490
rect 43276 648434 43281 648490
rect 42336 648432 43281 648434
rect 43215 648429 43281 648432
rect 674938 647986 674944 648050
rect 675008 648048 675014 648050
rect 675183 648048 675249 648051
rect 675008 648046 675249 648048
rect 675008 647990 675188 648046
rect 675244 647990 675249 648046
rect 675008 647988 675249 647990
rect 675008 647986 675014 647988
rect 675183 647985 675249 647988
rect 43503 647604 43569 647607
rect 42336 647602 43569 647604
rect 42336 647546 43508 647602
rect 43564 647546 43569 647602
rect 42336 647544 43569 647546
rect 43503 647541 43569 647544
rect 42298 647394 42304 647458
rect 42368 647394 42374 647458
rect 42306 647012 42366 647394
rect 43791 647012 43857 647015
rect 42306 647010 43857 647012
rect 42306 646982 43796 647010
rect 42336 646954 43796 646982
rect 43852 646954 43857 647010
rect 42336 646952 43857 646954
rect 43791 646949 43857 646952
rect 42106 646654 42112 646718
rect 42176 646654 42182 646718
rect 42114 646124 42174 646654
rect 43599 646124 43665 646127
rect 654447 646124 654513 646127
rect 42114 646122 43665 646124
rect 42114 646094 43604 646122
rect 42144 646066 43604 646094
rect 43660 646066 43665 646122
rect 42144 646064 43665 646066
rect 650208 646122 654513 646124
rect 650208 646066 654452 646122
rect 654508 646066 654513 646122
rect 650208 646064 654513 646066
rect 43599 646061 43665 646064
rect 654447 646061 654513 646064
rect 43119 645384 43185 645387
rect 42336 645382 43185 645384
rect 42336 645326 43124 645382
rect 43180 645326 43185 645382
rect 42336 645324 43185 645326
rect 43119 645321 43185 645324
rect 674362 645322 674368 645386
rect 674432 645384 674438 645386
rect 675471 645384 675537 645387
rect 674432 645382 675537 645384
rect 674432 645326 675476 645382
rect 675532 645326 675537 645382
rect 674432 645324 675537 645326
rect 674432 645322 674438 645324
rect 675471 645321 675537 645324
rect 40002 643907 40062 644466
rect 40002 643902 40113 643907
rect 40002 643846 40052 643902
rect 40108 643846 40113 643902
rect 40002 643844 40113 643846
rect 40047 643841 40113 643844
rect 40578 643166 40638 643726
rect 40570 643102 40576 643166
rect 40640 643102 40646 643166
rect 59247 642868 59313 642871
rect 59247 642866 64416 642868
rect 41922 642427 41982 642838
rect 59247 642810 59252 642866
rect 59308 642810 64416 642866
rect 59247 642808 64416 642810
rect 59247 642805 59313 642808
rect 675514 642510 675520 642574
rect 675584 642572 675590 642574
rect 676282 642572 676288 642574
rect 675584 642512 676288 642572
rect 675584 642510 675590 642512
rect 676282 642510 676288 642512
rect 676352 642510 676358 642574
rect 41871 642422 41982 642427
rect 41871 642366 41876 642422
rect 41932 642366 41982 642422
rect 41871 642364 41982 642366
rect 41871 642361 41937 642364
rect 42114 641687 42174 642172
rect 42114 641682 42225 641687
rect 42114 641626 42164 641682
rect 42220 641626 42225 641682
rect 42114 641624 42225 641626
rect 42159 641621 42225 641624
rect 41730 640799 41790 641358
rect 674746 641178 674752 641242
rect 674816 641178 674822 641242
rect 41730 640794 41841 640799
rect 41730 640738 41780 640794
rect 41836 640738 41841 640794
rect 41730 640736 41841 640738
rect 674754 640796 674814 641178
rect 675322 640882 675328 640946
rect 675392 640944 675398 640946
rect 675898 640944 675904 640946
rect 675392 640884 675904 640944
rect 675392 640882 675398 640884
rect 675898 640882 675904 640884
rect 675968 640882 675974 640946
rect 675514 640796 675520 640798
rect 674754 640736 675520 640796
rect 41775 640733 41841 640736
rect 675514 640734 675520 640736
rect 675584 640734 675590 640798
rect 674554 640586 674560 640650
rect 674624 640648 674630 640650
rect 674938 640648 674944 640650
rect 674624 640588 674944 640648
rect 674624 640586 674630 640588
rect 674938 640586 674944 640588
rect 675008 640586 675014 640650
rect 40770 640058 40830 640544
rect 676474 640500 676480 640502
rect 674946 640440 676480 640500
rect 674946 640206 675006 640440
rect 676474 640438 676480 640440
rect 676544 640438 676550 640502
rect 675759 640352 675825 640355
rect 676474 640352 676480 640354
rect 675759 640350 676480 640352
rect 675759 640294 675764 640350
rect 675820 640294 676480 640350
rect 675759 640292 676480 640294
rect 675759 640289 675825 640292
rect 676474 640290 676480 640292
rect 676544 640290 676550 640354
rect 674938 640142 674944 640206
rect 675008 640142 675014 640206
rect 40762 639994 40768 640058
rect 40832 639994 40838 640058
rect 41922 639467 41982 639730
rect 41922 639462 42033 639467
rect 41922 639406 41972 639462
rect 42028 639406 42033 639462
rect 41922 639404 42033 639406
rect 41967 639401 42033 639404
rect 41538 638431 41598 638916
rect 675375 638578 675441 638579
rect 675322 638576 675328 638578
rect 675284 638516 675328 638576
rect 675392 638574 675441 638578
rect 675436 638518 675441 638574
rect 675322 638514 675328 638516
rect 675392 638514 675441 638518
rect 675375 638513 675441 638514
rect 41487 638426 41598 638431
rect 41487 638370 41492 638426
rect 41548 638370 41598 638426
rect 41487 638368 41598 638370
rect 41487 638365 41553 638368
rect 42306 637690 42366 638102
rect 42298 637626 42304 637690
rect 42368 637626 42374 637690
rect 42114 636803 42174 637362
rect 42063 636798 42174 636803
rect 42063 636742 42068 636798
rect 42124 636742 42174 636798
rect 42063 636740 42174 636742
rect 42063 636737 42129 636740
rect 43023 636652 43089 636655
rect 42336 636650 43089 636652
rect 42336 636594 43028 636650
rect 43084 636594 43089 636650
rect 42336 636592 43089 636594
rect 43023 636589 43089 636592
rect 42639 635764 42705 635767
rect 42336 635762 42705 635764
rect 42336 635706 42644 635762
rect 42700 635706 42705 635762
rect 42336 635704 42705 635706
rect 42639 635701 42705 635704
rect 42927 635024 42993 635027
rect 42336 635022 42993 635024
rect 42336 634966 42932 635022
rect 42988 634966 42993 635022
rect 42336 634964 42993 634966
rect 42927 634961 42993 634964
rect 655311 634432 655377 634435
rect 650208 634430 655377 634432
rect 650208 634374 655316 634430
rect 655372 634374 655377 634430
rect 650208 634372 655377 634374
rect 655311 634369 655377 634372
rect 42306 633544 42366 634106
rect 42306 633484 42750 633544
rect 42690 633100 42750 633484
rect 42306 633040 42750 633100
rect 42306 632508 42366 633040
rect 42447 632508 42513 632511
rect 42306 632506 42513 632508
rect 42306 632450 42452 632506
rect 42508 632450 42513 632506
rect 42306 632448 42513 632450
rect 42447 632445 42513 632448
rect 674703 632508 674769 632511
rect 674703 632506 674814 632508
rect 674703 632450 674708 632506
rect 674764 632450 674814 632506
rect 674703 632445 674814 632450
rect 674754 632330 674814 632445
rect 674703 631768 674769 631771
rect 674703 631766 674814 631768
rect 674703 631710 674708 631766
rect 674764 631710 674814 631766
rect 674703 631705 674814 631710
rect 674754 631442 674814 631705
rect 674127 630732 674193 630735
rect 674127 630730 674784 630732
rect 674127 630674 674132 630730
rect 674188 630674 674784 630730
rect 674127 630672 674784 630674
rect 674127 630669 674193 630672
rect 673839 629844 673905 629847
rect 673839 629842 674784 629844
rect 673839 629786 673844 629842
rect 673900 629786 674784 629842
rect 673839 629784 674784 629786
rect 673839 629781 673905 629784
rect 673839 629104 673905 629107
rect 673839 629102 674784 629104
rect 673839 629046 673844 629102
rect 673900 629046 674784 629102
rect 673839 629044 674784 629046
rect 673839 629041 673905 629044
rect 57999 628512 58065 628515
rect 57999 628510 64416 628512
rect 57999 628454 58004 628510
rect 58060 628454 64416 628510
rect 57999 628452 64416 628454
rect 57999 628449 58065 628452
rect 673839 628364 673905 628367
rect 673839 628362 674784 628364
rect 673839 628306 673844 628362
rect 673900 628306 674784 628362
rect 673839 628304 674784 628306
rect 673839 628301 673905 628304
rect 675183 628068 675249 628071
rect 675138 628066 675249 628068
rect 675138 628010 675188 628066
rect 675244 628010 675249 628066
rect 675138 628005 675249 628010
rect 43119 627922 43185 627923
rect 43066 627920 43072 627922
rect 43028 627860 43072 627920
rect 43136 627918 43185 627922
rect 43180 627862 43185 627918
rect 43066 627858 43072 627860
rect 43136 627858 43185 627862
rect 43119 627857 43185 627858
rect 675138 627520 675198 628005
rect 41871 627478 41937 627479
rect 42159 627478 42225 627479
rect 41871 627476 41920 627478
rect 41828 627474 41920 627476
rect 41828 627418 41876 627474
rect 41828 627416 41920 627418
rect 41871 627414 41920 627416
rect 41984 627414 41990 627478
rect 42106 627476 42112 627478
rect 42068 627416 42112 627476
rect 42176 627474 42225 627478
rect 42220 627418 42225 627474
rect 42106 627414 42112 627416
rect 42176 627414 42225 627418
rect 41871 627413 41937 627414
rect 42159 627413 42225 627414
rect 675898 627266 675904 627330
rect 675968 627266 675974 627330
rect 675906 626706 675966 627266
rect 674799 626144 674865 626147
rect 674754 626142 674865 626144
rect 674754 626086 674804 626142
rect 674860 626086 674865 626142
rect 674754 626081 674865 626086
rect 674754 625892 674814 626081
rect 675514 625638 675520 625702
rect 675584 625638 675590 625702
rect 675522 625078 675582 625638
rect 676282 624750 676288 624814
rect 676352 624750 676358 624814
rect 676290 624264 676350 624750
rect 42447 623924 42513 623927
rect 42682 623924 42688 623926
rect 42447 623922 42688 623924
rect 42447 623866 42452 623922
rect 42508 623866 42688 623922
rect 42447 623864 42688 623866
rect 42447 623861 42513 623864
rect 42682 623862 42688 623864
rect 42752 623862 42758 623926
rect 674319 623628 674385 623631
rect 674319 623626 674784 623628
rect 674319 623570 674324 623626
rect 674380 623570 674784 623626
rect 674319 623568 674784 623570
rect 674319 623565 674385 623568
rect 42159 623480 42225 623483
rect 42298 623480 42304 623482
rect 42159 623478 42304 623480
rect 42159 623422 42164 623478
rect 42220 623422 42304 623478
rect 42159 623420 42304 623422
rect 42159 623417 42225 623420
rect 42298 623418 42304 623420
rect 42368 623418 42374 623482
rect 41914 623270 41920 623334
rect 41984 623332 41990 623334
rect 42447 623332 42513 623335
rect 41984 623330 42513 623332
rect 41984 623274 42452 623330
rect 42508 623274 42513 623330
rect 41984 623272 42513 623274
rect 41984 623270 41990 623272
rect 42447 623269 42513 623272
rect 674415 622740 674481 622743
rect 674415 622738 674784 622740
rect 674415 622682 674420 622738
rect 674476 622682 674784 622738
rect 674415 622680 674784 622682
rect 674415 622677 674481 622680
rect 656367 622592 656433 622595
rect 650208 622590 656433 622592
rect 650208 622534 656372 622590
rect 656428 622534 656433 622590
rect 650208 622532 656433 622534
rect 656367 622529 656433 622532
rect 673978 621938 673984 622002
rect 674048 622000 674054 622002
rect 674048 621940 674784 622000
rect 674048 621938 674054 621940
rect 676666 621642 676672 621706
rect 676736 621642 676742 621706
rect 676674 621082 676734 621642
rect 674938 620902 674944 620966
rect 675008 620902 675014 620966
rect 42927 620816 42993 620819
rect 43066 620816 43072 620818
rect 42927 620814 43072 620816
rect 42927 620758 42932 620814
rect 42988 620758 43072 620814
rect 42927 620756 43072 620758
rect 42927 620753 42993 620756
rect 43066 620754 43072 620756
rect 43136 620754 43142 620818
rect 674946 620342 675006 620902
rect 42063 620226 42129 620227
rect 42063 620224 42112 620226
rect 42020 620222 42112 620224
rect 42020 620166 42068 620222
rect 42020 620164 42112 620166
rect 42063 620162 42112 620164
rect 42176 620162 42182 620226
rect 42063 620161 42129 620162
rect 674223 619484 674289 619487
rect 674223 619482 674784 619484
rect 674223 619426 674228 619482
rect 674284 619426 674784 619482
rect 674223 619424 674784 619426
rect 674223 619421 674289 619424
rect 674746 619126 674752 619190
rect 674816 619126 674822 619190
rect 674754 618862 674814 619126
rect 41967 618450 42033 618451
rect 41914 618448 41920 618450
rect 41876 618388 41920 618448
rect 41984 618446 42033 618450
rect 42028 618390 42033 618446
rect 41914 618386 41920 618388
rect 41984 618386 42033 618390
rect 41967 618385 42033 618386
rect 40762 618238 40768 618302
rect 40832 618300 40838 618302
rect 42735 618300 42801 618303
rect 40832 618298 42801 618300
rect 40832 618242 42740 618298
rect 42796 618242 42801 618298
rect 40832 618240 42801 618242
rect 40832 618238 40838 618240
rect 42735 618237 42801 618240
rect 40570 618090 40576 618154
rect 40640 618152 40646 618154
rect 42831 618152 42897 618155
rect 40640 618150 42897 618152
rect 40640 618094 42836 618150
rect 42892 618094 42897 618150
rect 40640 618092 42897 618094
rect 40640 618090 40646 618092
rect 42831 618089 42897 618092
rect 673839 618004 673905 618007
rect 673839 618002 674784 618004
rect 673839 617946 673844 618002
rect 673900 617946 674784 618002
rect 673839 617944 674784 617946
rect 673839 617941 673905 617944
rect 41775 617858 41841 617859
rect 41722 617794 41728 617858
rect 41792 617856 41841 617858
rect 41792 617854 41884 617856
rect 41836 617798 41884 617854
rect 41792 617796 41884 617798
rect 41792 617794 41841 617796
rect 677050 617794 677056 617858
rect 677120 617794 677126 617858
rect 41775 617793 41841 617794
rect 677058 617234 677118 617794
rect 673839 616376 673905 616379
rect 673839 616374 674784 616376
rect 673839 616318 673844 616374
rect 673900 616318 674784 616374
rect 673839 616316 674784 616318
rect 673839 616313 673905 616316
rect 679746 615047 679806 615606
rect 679695 615042 679806 615047
rect 679695 614986 679700 615042
rect 679756 614986 679806 615042
rect 679695 614984 679806 614986
rect 679695 614981 679761 614984
rect 679695 614452 679761 614455
rect 679695 614450 679806 614452
rect 679695 614394 679700 614450
rect 679756 614394 679806 614450
rect 679695 614389 679806 614394
rect 679746 614052 679806 614389
rect 59439 614008 59505 614011
rect 59439 614006 64416 614008
rect 59439 613950 59444 614006
rect 59500 613950 64416 614006
rect 59439 613948 64416 613950
rect 59439 613945 59505 613948
rect 654447 611048 654513 611051
rect 650208 611046 654513 611048
rect 650208 610990 654452 611046
rect 654508 610990 654513 611046
rect 650208 610988 654513 610990
rect 654447 610985 654513 610988
rect 674746 607730 674752 607794
rect 674816 607792 674822 607794
rect 675087 607792 675153 607795
rect 674816 607790 675153 607792
rect 674816 607734 675092 607790
rect 675148 607734 675153 607790
rect 674816 607732 675153 607734
rect 674816 607730 674822 607732
rect 675087 607729 675153 607732
rect 42735 607718 42801 607721
rect 42336 607716 42801 607718
rect 42336 607660 42740 607716
rect 42796 607660 42801 607716
rect 42336 607658 42801 607660
rect 42735 607655 42801 607658
rect 673978 607434 673984 607498
rect 674048 607496 674054 607498
rect 675087 607496 675153 607499
rect 674048 607494 675153 607496
rect 674048 607438 675092 607494
rect 675148 607438 675153 607494
rect 674048 607436 675153 607438
rect 674048 607434 674054 607436
rect 675087 607433 675153 607436
rect 42735 606904 42801 606907
rect 42336 606902 42801 606904
rect 42336 606846 42740 606902
rect 42796 606846 42801 606902
rect 42336 606844 42801 606846
rect 42735 606841 42801 606844
rect 675471 606462 675537 606463
rect 675471 606458 675520 606462
rect 675584 606460 675590 606462
rect 675471 606402 675476 606458
rect 675471 606398 675520 606402
rect 675584 606400 675628 606460
rect 675584 606398 675590 606400
rect 675471 606397 675537 606398
rect 42447 606312 42513 606315
rect 42306 606310 42513 606312
rect 42306 606254 42452 606310
rect 42508 606254 42513 606310
rect 42306 606252 42513 606254
rect 42306 606060 42366 606252
rect 42447 606249 42513 606252
rect 43503 605276 43569 605279
rect 42336 605274 43569 605276
rect 42336 605218 43508 605274
rect 43564 605218 43569 605274
rect 42336 605216 43569 605218
rect 43503 605213 43569 605216
rect 674895 604980 674961 604983
rect 674754 604978 674961 604980
rect 674754 604922 674900 604978
rect 674956 604922 674961 604978
rect 674754 604920 674961 604922
rect 674754 604835 674814 604920
rect 674895 604917 674961 604920
rect 674703 604830 674814 604835
rect 674703 604774 674708 604830
rect 674764 604774 674814 604830
rect 674703 604772 674814 604774
rect 674703 604769 674769 604772
rect 674938 604770 674944 604834
rect 675008 604832 675014 604834
rect 675087 604832 675153 604835
rect 675008 604830 675153 604832
rect 675008 604774 675092 604830
rect 675148 604774 675153 604830
rect 675008 604772 675153 604774
rect 675008 604770 675014 604772
rect 675087 604769 675153 604772
rect 43215 604684 43281 604687
rect 42306 604682 43281 604684
rect 42306 604626 43220 604682
rect 43276 604626 43281 604682
rect 42306 604624 43281 604626
rect 42306 604432 42366 604624
rect 43215 604621 43281 604624
rect 43407 603796 43473 603799
rect 43791 603796 43857 603799
rect 42336 603794 43857 603796
rect 42336 603738 43412 603794
rect 43468 603738 43796 603794
rect 43852 603738 43857 603794
rect 42336 603736 43857 603738
rect 43407 603733 43473 603736
rect 43791 603733 43857 603736
rect 43599 602908 43665 602911
rect 42336 602906 43665 602908
rect 42336 602850 43604 602906
rect 43660 602850 43665 602906
rect 42336 602848 43665 602850
rect 43599 602845 43665 602848
rect 43119 602168 43185 602171
rect 42336 602166 43185 602168
rect 42336 602110 43124 602166
rect 43180 602110 43185 602166
rect 42336 602108 43185 602110
rect 43119 602105 43185 602108
rect 40002 600691 40062 601250
rect 40002 600686 40113 600691
rect 40002 600630 40052 600686
rect 40108 600630 40113 600686
rect 40002 600628 40113 600630
rect 40047 600625 40113 600628
rect 40578 599950 40638 600510
rect 675759 600244 675825 600247
rect 675898 600244 675904 600246
rect 675759 600242 675904 600244
rect 675759 600186 675764 600242
rect 675820 600186 675904 600242
rect 675759 600184 675904 600186
rect 675759 600181 675825 600184
rect 675898 600182 675904 600184
rect 675968 600182 675974 600246
rect 40570 599886 40576 599950
rect 40640 599886 40646 599950
rect 59535 599800 59601 599803
rect 59535 599798 64416 599800
rect 59535 599742 59540 599798
rect 59596 599742 64416 599798
rect 59535 599740 64416 599742
rect 59535 599737 59601 599740
rect 43023 599652 43089 599655
rect 42336 599650 43089 599652
rect 42336 599594 43028 599650
rect 43084 599594 43089 599650
rect 42336 599592 43089 599594
rect 43023 599589 43089 599592
rect 654447 599208 654513 599211
rect 650208 599206 654513 599208
rect 650208 599150 654452 599206
rect 654508 599150 654513 599206
rect 650208 599148 654513 599150
rect 654447 599145 654513 599148
rect 41922 598471 41982 599030
rect 41871 598466 41982 598471
rect 41871 598410 41876 598466
rect 41932 598410 41982 598466
rect 41871 598408 41982 598410
rect 41871 598405 41937 598408
rect 41730 597583 41790 598142
rect 41730 597578 41841 597583
rect 41730 597522 41780 597578
rect 41836 597522 41841 597578
rect 41730 597520 41841 597522
rect 41775 597517 41841 597520
rect 40962 596842 41022 597402
rect 40954 596778 40960 596842
rect 41024 596778 41030 596842
rect 42114 596251 42174 596514
rect 42063 596246 42174 596251
rect 42063 596190 42068 596246
rect 42124 596190 42174 596246
rect 42063 596188 42174 596190
rect 42063 596185 42129 596188
rect 41922 595215 41982 595774
rect 675759 595360 675825 595363
rect 676666 595360 676672 595362
rect 675759 595358 676672 595360
rect 675759 595302 675764 595358
rect 675820 595302 676672 595358
rect 675759 595300 676672 595302
rect 675759 595297 675825 595300
rect 676666 595298 676672 595300
rect 676736 595298 676742 595362
rect 41922 595210 42033 595215
rect 41922 595154 41972 595210
rect 42028 595154 42033 595210
rect 41922 595152 42033 595154
rect 41967 595149 42033 595152
rect 42831 594916 42897 594919
rect 42336 594914 42897 594916
rect 42336 594858 42836 594914
rect 42892 594858 42897 594914
rect 42336 594856 42897 594858
rect 42831 594853 42897 594856
rect 42114 593735 42174 594220
rect 42114 593730 42225 593735
rect 42114 593674 42164 593730
rect 42220 593674 42225 593730
rect 42114 593672 42225 593674
rect 42159 593669 42225 593672
rect 42543 593584 42609 593587
rect 42306 593582 42609 593584
rect 42306 593526 42548 593582
rect 42604 593526 42609 593582
rect 42306 593524 42609 593526
rect 42306 593406 42366 593524
rect 42543 593521 42609 593524
rect 675759 593436 675825 593439
rect 676282 593436 676288 593438
rect 675759 593434 676288 593436
rect 675759 593378 675764 593434
rect 675820 593378 676288 593434
rect 675759 593376 676288 593378
rect 675759 593373 675825 593376
rect 676282 593374 676288 593376
rect 676352 593374 676358 593438
rect 42306 592400 42366 592592
rect 42543 592400 42609 592403
rect 42306 592398 42609 592400
rect 42306 592342 42548 592398
rect 42604 592342 42609 592398
rect 42306 592340 42609 592342
rect 42543 592337 42609 592340
rect 42927 591808 42993 591811
rect 42336 591806 42993 591808
rect 42336 591750 42932 591806
rect 42988 591750 42993 591806
rect 42336 591748 42993 591750
rect 42927 591745 42993 591748
rect 42306 590624 42366 590964
rect 42447 590624 42513 590627
rect 42306 590622 42513 590624
rect 42306 590566 42452 590622
rect 42508 590566 42513 590622
rect 42306 590564 42513 590566
rect 42447 590561 42513 590564
rect 42306 589292 42366 589410
rect 42447 589292 42513 589295
rect 42306 589290 42513 589292
rect 42306 589234 42452 589290
rect 42508 589234 42513 589290
rect 42306 589232 42513 589234
rect 42447 589229 42513 589232
rect 655119 587368 655185 587371
rect 650208 587366 655185 587368
rect 650208 587310 655124 587366
rect 655180 587310 655185 587366
rect 650208 587308 655185 587310
rect 655119 587305 655185 587308
rect 674754 586483 674814 587042
rect 674703 586478 674814 586483
rect 674703 586422 674708 586478
rect 674764 586422 674814 586478
rect 674703 586420 674814 586422
rect 674703 586417 674769 586420
rect 674415 586332 674481 586335
rect 674415 586330 674784 586332
rect 674415 586274 674420 586330
rect 674476 586274 674784 586330
rect 674415 586272 674784 586274
rect 674415 586269 674481 586272
rect 42874 585382 42880 585446
rect 42944 585444 42950 585446
rect 43023 585444 43089 585447
rect 42944 585442 43089 585444
rect 42944 585386 43028 585442
rect 43084 585386 43089 585442
rect 42944 585384 43089 585386
rect 42944 585382 42950 585384
rect 43023 585381 43089 585384
rect 59535 585444 59601 585447
rect 674415 585444 674481 585447
rect 59535 585442 64416 585444
rect 59535 585386 59540 585442
rect 59596 585386 64416 585442
rect 59535 585384 64416 585386
rect 674415 585442 674784 585444
rect 674415 585386 674420 585442
rect 674476 585386 674784 585442
rect 674415 585384 674784 585386
rect 59535 585381 59601 585384
rect 674415 585381 674481 585384
rect 674607 584852 674673 584855
rect 674607 584850 674814 584852
rect 674607 584794 674612 584850
rect 674668 584794 674814 584850
rect 674607 584792 674814 584794
rect 674607 584789 674673 584792
rect 42543 584706 42609 584707
rect 42490 584704 42496 584706
rect 42452 584644 42496 584704
rect 42560 584702 42609 584706
rect 42604 584646 42609 584702
rect 674754 584674 674814 584792
rect 42490 584642 42496 584644
rect 42560 584642 42609 584646
rect 42543 584641 42609 584642
rect 42447 584554 42513 584559
rect 42447 584498 42452 584554
rect 42508 584498 42513 584554
rect 42447 584493 42513 584498
rect 42450 584263 42510 584493
rect 41530 584198 41536 584262
rect 41600 584260 41606 584262
rect 41871 584260 41937 584263
rect 41600 584258 41937 584260
rect 41600 584202 41876 584258
rect 41932 584202 41937 584258
rect 41600 584200 41937 584202
rect 41600 584198 41606 584200
rect 41871 584197 41937 584200
rect 42063 584260 42129 584263
rect 42298 584260 42304 584262
rect 42063 584258 42304 584260
rect 42063 584202 42068 584258
rect 42124 584202 42304 584258
rect 42063 584200 42304 584202
rect 42063 584197 42129 584200
rect 42298 584198 42304 584200
rect 42368 584198 42374 584262
rect 42447 584258 42513 584263
rect 42447 584202 42452 584258
rect 42508 584202 42513 584258
rect 42447 584197 42513 584202
rect 674754 583671 674814 583786
rect 674703 583666 674814 583671
rect 674703 583610 674708 583666
rect 674764 583610 674814 583666
rect 674703 583608 674814 583610
rect 674703 583605 674769 583608
rect 670959 583224 671025 583227
rect 674415 583224 674481 583227
rect 670959 583222 674784 583224
rect 670959 583166 670964 583222
rect 671020 583166 674420 583222
rect 674476 583166 674784 583222
rect 670959 583164 674784 583166
rect 670959 583161 671025 583164
rect 674415 583161 674481 583164
rect 676815 582632 676881 582635
rect 676815 582630 676926 582632
rect 676815 582574 676820 582630
rect 676876 582574 676926 582630
rect 676815 582569 676926 582574
rect 676866 582306 676926 582569
rect 675130 581682 675136 581746
rect 675200 581682 675206 581746
rect 675138 581566 675198 581682
rect 676474 581238 676480 581302
rect 676544 581238 676550 581302
rect 676482 580678 676542 581238
rect 675706 580350 675712 580414
rect 675776 580350 675782 580414
rect 42298 580054 42304 580118
rect 42368 580116 42374 580118
rect 43023 580116 43089 580119
rect 42368 580114 43089 580116
rect 42368 580058 43028 580114
rect 43084 580058 43089 580114
rect 42368 580056 43089 580058
rect 42368 580054 42374 580056
rect 43023 580053 43089 580056
rect 675714 579864 675774 580350
rect 676090 579610 676096 579674
rect 676160 579610 676166 579674
rect 676098 579050 676158 579610
rect 674415 578932 674481 578935
rect 676090 578932 676096 578934
rect 674415 578930 676096 578932
rect 674415 578874 674420 578930
rect 674476 578874 676096 578930
rect 674415 578872 676096 578874
rect 674415 578869 674481 578872
rect 676090 578870 676096 578872
rect 676160 578870 676166 578934
rect 674362 578352 674368 578416
rect 674432 578414 674438 578416
rect 674432 578354 674784 578414
rect 674432 578352 674438 578354
rect 42927 578342 42993 578343
rect 42874 578278 42880 578342
rect 42944 578340 42993 578342
rect 42944 578338 43036 578340
rect 42988 578282 43036 578338
rect 42944 578280 43036 578282
rect 42944 578278 42993 578280
rect 42927 578277 42993 578278
rect 675322 578130 675328 578194
rect 675392 578130 675398 578194
rect 675330 577570 675390 578130
rect 41530 577094 41536 577158
rect 41600 577156 41606 577158
rect 41775 577156 41841 577159
rect 41600 577154 41841 577156
rect 41600 577098 41780 577154
rect 41836 577098 41841 577154
rect 41600 577096 41841 577098
rect 41600 577094 41606 577096
rect 41775 577093 41841 577096
rect 674170 576724 674176 576788
rect 674240 576786 674246 576788
rect 674240 576726 674784 576786
rect 674240 576724 674246 576726
rect 674554 576058 674560 576122
rect 674624 576120 674630 576122
rect 674624 576060 674814 576120
rect 674624 576058 674630 576060
rect 42255 575972 42321 575975
rect 42490 575972 42496 575974
rect 42255 575970 42496 575972
rect 42255 575914 42260 575970
rect 42316 575914 42496 575970
rect 42255 575912 42496 575914
rect 42255 575909 42321 575912
rect 42490 575910 42496 575912
rect 42560 575910 42566 575974
rect 674754 575942 674814 576060
rect 654447 575676 654513 575679
rect 650208 575674 654513 575676
rect 650208 575618 654452 575674
rect 654508 575618 654513 575674
rect 650208 575616 654513 575618
rect 654447 575613 654513 575616
rect 674703 575380 674769 575383
rect 674703 575378 674814 575380
rect 674703 575322 674708 575378
rect 674764 575322 674814 575378
rect 674703 575317 674814 575322
rect 41967 575234 42033 575235
rect 41914 575170 41920 575234
rect 41984 575232 42033 575234
rect 41984 575230 42076 575232
rect 42028 575174 42076 575230
rect 41984 575172 42076 575174
rect 41984 575170 42033 575172
rect 41967 575169 42033 575170
rect 674754 575128 674814 575317
rect 41775 574642 41841 574643
rect 41722 574578 41728 574642
rect 41792 574640 41841 574642
rect 41792 574638 41884 574640
rect 41836 574582 41884 574638
rect 41792 574580 41884 574582
rect 41792 574578 41841 574580
rect 41775 574577 41841 574578
rect 674703 574492 674769 574495
rect 674703 574490 674814 574492
rect 674703 574434 674708 574490
rect 674764 574434 674814 574490
rect 674703 574429 674814 574434
rect 674754 574314 674814 574429
rect 40954 573986 40960 574050
rect 41024 574048 41030 574050
rect 42447 574048 42513 574051
rect 41024 574046 42513 574048
rect 41024 573990 42452 574046
rect 42508 573990 42513 574046
rect 41024 573988 42513 573990
rect 41024 573986 41030 573988
rect 42447 573985 42513 573988
rect 40570 573838 40576 573902
rect 40640 573900 40646 573902
rect 42831 573900 42897 573903
rect 40640 573898 42897 573900
rect 40640 573842 42836 573898
rect 42892 573842 42897 573898
rect 40640 573840 42897 573842
rect 40640 573838 40646 573840
rect 42831 573837 42897 573840
rect 674415 573604 674481 573607
rect 674415 573602 674784 573604
rect 674415 573546 674420 573602
rect 674476 573546 674784 573602
rect 674415 573544 674784 573546
rect 674415 573541 674481 573544
rect 674703 573012 674769 573015
rect 674703 573010 674814 573012
rect 674703 572954 674708 573010
rect 674764 572954 674814 573010
rect 674703 572949 674814 572954
rect 674754 572834 674814 572949
rect 674415 571976 674481 571979
rect 674415 571974 674784 571976
rect 674415 571918 674420 571974
rect 674476 571918 674784 571974
rect 674415 571916 674784 571918
rect 674415 571913 674481 571916
rect 674703 571384 674769 571387
rect 674703 571382 674814 571384
rect 674703 571326 674708 571382
rect 674764 571326 674814 571382
rect 674703 571321 674814 571326
rect 674754 571206 674814 571321
rect 59535 570940 59601 570943
rect 59535 570938 64416 570940
rect 59535 570882 59540 570938
rect 59596 570882 64416 570938
rect 59535 570880 64416 570882
rect 59535 570877 59601 570880
rect 679746 569759 679806 570318
rect 679746 569754 679857 569759
rect 679746 569698 679796 569754
rect 679852 569698 679857 569754
rect 679746 569696 679857 569698
rect 679791 569693 679857 569696
rect 679791 569164 679857 569167
rect 679746 569162 679857 569164
rect 679746 569106 679796 569162
rect 679852 569106 679857 569162
rect 679746 569101 679857 569106
rect 679746 568838 679806 569101
rect 34479 564724 34545 564727
rect 34434 564722 34545 564724
rect 34434 564666 34484 564722
rect 34540 564666 34545 564722
rect 34434 564661 34545 564666
rect 34434 564472 34494 564661
rect 654447 564132 654513 564135
rect 650208 564130 654513 564132
rect 650208 564074 654452 564130
rect 654508 564074 654513 564130
rect 650208 564072 654513 564074
rect 654447 564069 654513 564072
rect 42306 563540 42366 563658
rect 42447 563540 42513 563543
rect 42306 563538 42513 563540
rect 42306 563482 42452 563538
rect 42508 563482 42513 563538
rect 42306 563480 42513 563482
rect 42447 563477 42513 563480
rect 42351 563096 42417 563099
rect 42306 563094 42417 563096
rect 42306 563038 42356 563094
rect 42412 563038 42417 563094
rect 42306 563033 42417 563038
rect 42306 562844 42366 563033
rect 675279 562950 675345 562951
rect 675279 562946 675328 562950
rect 675392 562948 675398 562950
rect 675279 562890 675284 562946
rect 675279 562886 675328 562890
rect 675392 562888 675436 562948
rect 675392 562886 675398 562888
rect 675279 562885 675345 562886
rect 43215 562060 43281 562063
rect 42336 562058 43281 562060
rect 42336 562002 43220 562058
rect 43276 562002 43281 562058
rect 42336 562000 43281 562002
rect 43215 561997 43281 562000
rect 674170 561702 674176 561766
rect 674240 561764 674246 561766
rect 675087 561764 675153 561767
rect 674240 561762 675153 561764
rect 674240 561706 675092 561762
rect 675148 561706 675153 561762
rect 674240 561704 675153 561706
rect 674240 561702 674246 561704
rect 675087 561701 675153 561704
rect 43503 561616 43569 561619
rect 42306 561614 43569 561616
rect 42306 561558 43508 561614
rect 43564 561558 43569 561614
rect 42306 561556 43569 561558
rect 42306 561216 42366 561556
rect 43503 561553 43569 561556
rect 674554 561554 674560 561618
rect 674624 561616 674630 561618
rect 675279 561616 675345 561619
rect 674624 561614 675345 561616
rect 674624 561558 675284 561614
rect 675340 561558 675345 561614
rect 674624 561556 675345 561558
rect 674624 561554 674630 561556
rect 675279 561553 675345 561556
rect 43407 560580 43473 560583
rect 42336 560578 43473 560580
rect 42336 560522 43412 560578
rect 43468 560522 43473 560578
rect 42336 560520 43473 560522
rect 43407 560517 43473 560520
rect 43599 559840 43665 559843
rect 42306 559838 43665 559840
rect 42306 559782 43604 559838
rect 43660 559782 43665 559838
rect 42306 559780 43665 559782
rect 42306 559736 42366 559780
rect 43599 559777 43665 559780
rect 41730 558656 41790 558922
rect 675130 558890 675136 558954
rect 675200 558952 675206 558954
rect 675471 558952 675537 558955
rect 675200 558950 675537 558952
rect 675200 558894 675476 558950
rect 675532 558894 675537 558950
rect 675200 558892 675537 558894
rect 675200 558890 675206 558892
rect 675471 558889 675537 558892
rect 41967 558656 42033 558659
rect 41730 558654 42033 558656
rect 41730 558598 41972 558654
rect 42028 558598 42033 558654
rect 41730 558596 42033 558598
rect 41967 558593 42033 558596
rect 40002 557475 40062 558034
rect 674362 557706 674368 557770
rect 674432 557768 674438 557770
rect 675375 557768 675441 557771
rect 674432 557766 675441 557768
rect 674432 557710 675380 557766
rect 675436 557710 675441 557766
rect 674432 557708 675441 557710
rect 674432 557706 674438 557708
rect 675375 557705 675441 557708
rect 40002 557470 40113 557475
rect 40002 557414 40052 557470
rect 40108 557414 40113 557470
rect 40002 557412 40113 557414
rect 40047 557409 40113 557412
rect 40194 556735 40254 557294
rect 40143 556730 40254 556735
rect 40143 556674 40148 556730
rect 40204 556674 40254 556730
rect 40143 556672 40254 556674
rect 59535 556732 59601 556735
rect 59535 556730 64416 556732
rect 59535 556674 59540 556730
rect 59596 556674 64416 556730
rect 59535 556672 64416 556674
rect 40143 556669 40209 556672
rect 59535 556669 59601 556672
rect 41922 555995 41982 556406
rect 41871 555990 41982 555995
rect 41871 555934 41876 555990
rect 41932 555934 41982 555990
rect 41871 555932 41982 555934
rect 41871 555929 41937 555932
rect 41730 555255 41790 555814
rect 41679 555250 41790 555255
rect 41679 555194 41684 555250
rect 41740 555194 41790 555250
rect 41679 555192 41790 555194
rect 41679 555189 41745 555192
rect 41730 554367 41790 554926
rect 41730 554362 41841 554367
rect 41730 554306 41780 554362
rect 41836 554306 41841 554362
rect 41730 554304 41841 554306
rect 41775 554301 41841 554304
rect 37314 553627 37374 554186
rect 37314 553622 37425 553627
rect 37314 553566 37364 553622
rect 37420 553566 37425 553622
rect 37314 553564 37425 553566
rect 37359 553561 37425 553564
rect 42114 553035 42174 553298
rect 42063 553030 42174 553035
rect 42063 552974 42068 553030
rect 42124 552974 42174 553030
rect 42063 552972 42174 552974
rect 42063 552969 42129 552972
rect 42306 551999 42366 552558
rect 654447 552292 654513 552295
rect 650208 552290 654513 552292
rect 650208 552234 654452 552290
rect 654508 552234 654513 552290
rect 650208 552232 654513 552234
rect 654447 552229 654513 552232
rect 42306 551994 42417 551999
rect 42306 551938 42356 551994
rect 42412 551938 42417 551994
rect 42306 551936 42417 551938
rect 42351 551933 42417 551936
rect 43023 551700 43089 551703
rect 42336 551698 43089 551700
rect 42336 551642 43028 551698
rect 43084 551642 43089 551698
rect 42336 551640 43089 551642
rect 43023 551637 43089 551640
rect 42927 551108 42993 551111
rect 42336 551106 42993 551108
rect 42336 551050 42932 551106
rect 42988 551050 42993 551106
rect 42336 551048 42993 551050
rect 42927 551045 42993 551048
rect 674991 550220 675057 550223
rect 675706 550220 675712 550222
rect 674991 550218 675712 550220
rect 42114 550075 42174 550190
rect 674991 550162 674996 550218
rect 675052 550162 675712 550218
rect 674991 550160 675712 550162
rect 674991 550157 675057 550160
rect 675706 550158 675712 550160
rect 675776 550158 675782 550222
rect 42114 550070 42225 550075
rect 42114 550014 42164 550070
rect 42220 550014 42225 550070
rect 42114 550012 42225 550014
rect 42159 550009 42225 550012
rect 42306 549332 42366 549376
rect 43119 549332 43185 549335
rect 42306 549330 43185 549332
rect 42306 549274 43124 549330
rect 43180 549274 43185 549330
rect 42306 549272 43185 549274
rect 43119 549269 43185 549272
rect 42831 548592 42897 548595
rect 42336 548590 42897 548592
rect 42336 548534 42836 548590
rect 42892 548534 42897 548590
rect 42336 548532 42897 548534
rect 42831 548529 42897 548532
rect 42306 547260 42366 547748
rect 42306 547200 42750 547260
rect 42690 546816 42750 547200
rect 676090 547050 676096 547114
rect 676160 547112 676166 547114
rect 676527 547112 676593 547115
rect 676160 547110 676593 547112
rect 676160 547054 676532 547110
rect 676588 547054 676593 547110
rect 676160 547052 676593 547054
rect 676160 547050 676166 547052
rect 676527 547049 676593 547052
rect 675706 546902 675712 546966
rect 675776 546964 675782 546966
rect 676623 546964 676689 546967
rect 675776 546962 676689 546964
rect 675776 546906 676628 546962
rect 676684 546906 676689 546962
rect 675776 546904 676689 546906
rect 675776 546902 675782 546904
rect 676623 546901 676689 546904
rect 42306 546756 42750 546816
rect 42306 546298 42366 546756
rect 42639 546298 42705 546301
rect 42306 546296 42705 546298
rect 42306 546268 42644 546296
rect 42336 546240 42644 546268
rect 42700 546240 42705 546296
rect 42336 546238 42705 546240
rect 42639 546235 42705 546238
rect 40143 544300 40209 544303
rect 41146 544300 41152 544302
rect 40143 544298 41152 544300
rect 40143 544242 40148 544298
rect 40204 544242 41152 544298
rect 40143 544240 41152 544242
rect 40143 544237 40209 544240
rect 41146 544238 41152 544240
rect 41216 544238 41222 544302
rect 37359 542968 37425 542971
rect 40954 542968 40960 542970
rect 37359 542966 40960 542968
rect 37359 542910 37364 542966
rect 37420 542910 40960 542966
rect 37359 542908 40960 542910
rect 37359 542905 37425 542908
rect 40954 542906 40960 542908
rect 41024 542906 41030 542970
rect 59535 542376 59601 542379
rect 59535 542374 64416 542376
rect 59535 542318 59540 542374
rect 59596 542318 64416 542374
rect 59535 542316 64416 542318
rect 59535 542313 59601 542316
rect 674754 541639 674814 542050
rect 674703 541634 674814 541639
rect 674703 541578 674708 541634
rect 674764 541578 674814 541634
rect 674703 541576 674814 541578
rect 674703 541573 674769 541576
rect 41679 541340 41745 541343
rect 42106 541340 42112 541342
rect 41679 541338 42112 541340
rect 41679 541282 41684 541338
rect 41740 541282 42112 541338
rect 41679 541280 42112 541282
rect 41679 541277 41745 541280
rect 42106 541278 42112 541280
rect 42176 541278 42182 541342
rect 674223 541340 674289 541343
rect 674223 541338 674784 541340
rect 674223 541282 674228 541338
rect 674284 541282 674784 541338
rect 674223 541280 674784 541282
rect 674223 541277 674289 541280
rect 41871 541192 41937 541195
rect 42874 541192 42880 541194
rect 41871 541190 42880 541192
rect 41871 541134 41876 541190
rect 41932 541134 42880 541190
rect 41871 541132 42880 541134
rect 41871 541129 41937 541132
rect 42874 541130 42880 541132
rect 42944 541130 42950 541194
rect 42063 541044 42129 541047
rect 43066 541044 43072 541046
rect 42063 541042 43072 541044
rect 42063 540986 42068 541042
rect 42124 540986 43072 541042
rect 42063 540984 43072 540986
rect 42063 540981 42129 540984
rect 43066 540982 43072 540984
rect 43136 540982 43142 541046
rect 654447 540452 654513 540455
rect 650208 540450 654513 540452
rect 650208 540394 654452 540450
rect 654508 540394 654513 540450
rect 650208 540392 654513 540394
rect 654447 540389 654513 540392
rect 674223 540452 674289 540455
rect 674223 540450 674784 540452
rect 674223 540394 674228 540450
rect 674284 540394 674784 540450
rect 674223 540392 674784 540394
rect 674223 540389 674289 540392
rect 673839 539712 673905 539715
rect 673839 539710 674784 539712
rect 673839 539654 673844 539710
rect 673900 539654 674784 539710
rect 673839 539652 674784 539654
rect 673839 539649 673905 539652
rect 42106 538762 42112 538826
rect 42176 538824 42182 538826
rect 43023 538824 43089 538827
rect 42176 538822 43089 538824
rect 42176 538766 43028 538822
rect 43084 538766 43089 538822
rect 42176 538764 43089 538766
rect 42176 538762 42182 538764
rect 43023 538761 43089 538764
rect 676674 538679 676734 538794
rect 676674 538674 676785 538679
rect 676674 538618 676724 538674
rect 676780 538618 676785 538674
rect 676674 538616 676785 538618
rect 676719 538613 676785 538616
rect 676482 537939 676542 538128
rect 676482 537934 676593 537939
rect 676482 537878 676532 537934
rect 676588 537878 676593 537934
rect 676482 537876 676593 537878
rect 676527 537873 676593 537876
rect 676674 537199 676734 537314
rect 676623 537194 676734 537199
rect 676623 537138 676628 537194
rect 676684 537138 676734 537194
rect 676623 537136 676734 537138
rect 676623 537133 676689 537136
rect 675514 536986 675520 537050
rect 675584 536986 675590 537050
rect 42927 536902 42993 536903
rect 42874 536838 42880 536902
rect 42944 536900 42993 536902
rect 42944 536898 43036 536900
rect 42988 536842 43036 536898
rect 42944 536840 43036 536842
rect 42944 536838 42993 536840
rect 42927 536837 42993 536838
rect 675522 536500 675582 536986
rect 676666 536246 676672 536310
rect 676736 536246 676742 536310
rect 42831 535716 42897 535719
rect 43066 535716 43072 535718
rect 42831 535714 43072 535716
rect 42831 535658 42836 535714
rect 42892 535658 43072 535714
rect 42831 535656 43072 535658
rect 42831 535653 42897 535656
rect 43066 535654 43072 535656
rect 43136 535654 43142 535718
rect 676674 535686 676734 536246
rect 674746 535358 674752 535422
rect 674816 535358 674822 535422
rect 674754 534872 674814 535358
rect 674938 534618 674944 534682
rect 675008 534618 675014 534682
rect 674946 534058 675006 534618
rect 675898 533730 675904 533794
rect 675968 533730 675974 533794
rect 675906 533392 675966 533730
rect 676282 532694 676288 532758
rect 676352 532694 676358 532758
rect 40954 532546 40960 532610
rect 41024 532608 41030 532610
rect 42735 532608 42801 532611
rect 41024 532606 42801 532608
rect 41024 532550 42740 532606
rect 42796 532550 42801 532606
rect 676290 532578 676350 532694
rect 41024 532548 42801 532550
rect 41024 532546 41030 532548
rect 42735 532545 42801 532548
rect 41146 532250 41152 532314
rect 41216 532312 41222 532314
rect 42639 532312 42705 532315
rect 41216 532310 42705 532312
rect 41216 532254 42644 532310
rect 42700 532254 42705 532310
rect 41216 532252 42705 532254
rect 41216 532250 41222 532252
rect 42639 532249 42705 532252
rect 41871 532018 41937 532019
rect 41871 532016 41920 532018
rect 41828 532014 41920 532016
rect 41828 531958 41876 532014
rect 41828 531956 41920 531958
rect 41871 531954 41920 531956
rect 41984 531954 41990 532018
rect 41871 531953 41937 531954
rect 673978 531658 673984 531722
rect 674048 531720 674054 531722
rect 674048 531660 674784 531720
rect 674048 531658 674054 531660
rect 41775 531278 41841 531279
rect 41722 531214 41728 531278
rect 41792 531276 41841 531278
rect 41792 531274 41884 531276
rect 41836 531218 41884 531274
rect 41792 531216 41884 531218
rect 41792 531214 41841 531216
rect 41775 531213 41841 531214
rect 673743 530980 673809 530983
rect 673743 530978 674784 530980
rect 673743 530922 673748 530978
rect 673804 530922 674784 530978
rect 673743 530920 674784 530922
rect 673743 530917 673809 530920
rect 673839 530092 673905 530095
rect 673839 530090 674784 530092
rect 673839 530034 673844 530090
rect 673900 530034 674784 530090
rect 673839 530032 674784 530034
rect 673839 530029 673905 530032
rect 673839 529352 673905 529355
rect 673839 529350 674784 529352
rect 673839 529294 673844 529350
rect 673900 529294 674784 529350
rect 673839 529292 674784 529294
rect 673839 529289 673905 529292
rect 654447 528760 654513 528763
rect 650208 528758 654513 528760
rect 650208 528702 654452 528758
rect 654508 528702 654513 528758
rect 650208 528700 654513 528702
rect 654447 528697 654513 528700
rect 673839 528612 673905 528615
rect 673839 528610 674784 528612
rect 673839 528554 673844 528610
rect 673900 528554 674784 528610
rect 673839 528552 674784 528554
rect 673839 528549 673905 528552
rect 59535 527872 59601 527875
rect 673167 527872 673233 527875
rect 59535 527870 64416 527872
rect 59535 527814 59540 527870
rect 59596 527814 64416 527870
rect 59535 527812 64416 527814
rect 673167 527870 674784 527872
rect 673167 527814 673172 527870
rect 673228 527814 674784 527870
rect 673167 527812 674784 527814
rect 59535 527809 59601 527812
rect 673167 527809 673233 527812
rect 673839 526984 673905 526987
rect 673839 526982 674784 526984
rect 673839 526926 673844 526982
rect 673900 526926 674784 526982
rect 673839 526924 674784 526926
rect 673839 526921 673905 526924
rect 673839 526244 673905 526247
rect 673839 526242 674784 526244
rect 673839 526186 673844 526242
rect 673900 526186 674784 526242
rect 673839 526184 674784 526186
rect 673839 526181 673905 526184
rect 679746 524767 679806 525326
rect 679746 524762 679857 524767
rect 679746 524706 679796 524762
rect 679852 524706 679857 524762
rect 679746 524704 679857 524706
rect 679791 524701 679857 524704
rect 679791 524172 679857 524175
rect 679746 524170 679857 524172
rect 679746 524114 679796 524170
rect 679852 524114 679857 524170
rect 679746 524109 679857 524114
rect 679746 523846 679806 524109
rect 654063 517216 654129 517219
rect 650208 517214 654129 517216
rect 650208 517158 654068 517214
rect 654124 517158 654129 517214
rect 650208 517156 654129 517158
rect 654063 517153 654129 517156
rect 59343 513516 59409 513519
rect 59343 513514 64416 513516
rect 59343 513458 59348 513514
rect 59404 513458 64416 513514
rect 59343 513456 64416 513458
rect 59343 513453 59409 513456
rect 654927 505376 654993 505379
rect 650208 505374 654993 505376
rect 650208 505318 654932 505374
rect 654988 505318 654993 505374
rect 650208 505316 654993 505318
rect 654927 505313 654993 505316
rect 57807 499160 57873 499163
rect 57807 499158 64416 499160
rect 57807 499102 57812 499158
rect 57868 499102 64416 499158
rect 57807 499100 64416 499102
rect 57807 499097 57873 499100
rect 674754 497831 674814 498094
rect 674703 497826 674814 497831
rect 674703 497770 674708 497826
rect 674764 497770 674814 497826
rect 674703 497768 674814 497770
rect 674703 497765 674769 497768
rect 674511 497532 674577 497535
rect 674511 497530 674814 497532
rect 674511 497474 674516 497530
rect 674572 497474 674814 497530
rect 674511 497472 674814 497474
rect 674511 497469 674577 497472
rect 674754 497280 674814 497472
rect 674511 496644 674577 496647
rect 674511 496642 674814 496644
rect 674511 496586 674516 496642
rect 674572 496586 674814 496642
rect 674511 496584 674814 496586
rect 674511 496581 674577 496584
rect 674754 496466 674814 496584
rect 676719 495904 676785 495907
rect 676674 495902 676785 495904
rect 676674 495846 676724 495902
rect 676780 495846 676785 495902
rect 676674 495841 676785 495846
rect 676674 495578 676734 495841
rect 676674 494575 676734 494838
rect 676674 494570 676785 494575
rect 676674 494514 676724 494570
rect 676780 494514 676785 494570
rect 676674 494512 676785 494514
rect 676719 494509 676785 494512
rect 676482 493983 676542 494098
rect 676482 493978 676593 493983
rect 676482 493922 676532 493978
rect 676588 493922 676593 493978
rect 676482 493920 676593 493922
rect 676527 493917 676593 493920
rect 655215 493536 655281 493539
rect 650208 493534 655281 493536
rect 650208 493478 655220 493534
rect 655276 493478 655281 493534
rect 650208 493476 655281 493478
rect 655215 493473 655281 493476
rect 676674 493095 676734 493358
rect 676623 493090 676734 493095
rect 676623 493034 676628 493090
rect 676684 493034 676734 493090
rect 676623 493032 676734 493034
rect 676623 493029 676689 493032
rect 674554 492290 674560 492354
rect 674624 492352 674630 492354
rect 674754 492352 674814 492470
rect 674624 492292 674814 492352
rect 674624 492290 674630 492292
rect 674799 491908 674865 491911
rect 674754 491906 674865 491908
rect 674754 491850 674804 491906
rect 674860 491850 674865 491906
rect 674754 491845 674865 491850
rect 674754 491730 674814 491845
rect 675322 491402 675328 491466
rect 675392 491402 675398 491466
rect 675330 490842 675390 491402
rect 674319 490132 674385 490135
rect 674319 490130 674784 490132
rect 674319 490074 674324 490130
rect 674380 490074 674784 490130
rect 674319 490072 674784 490074
rect 674319 490069 674385 490072
rect 674415 489392 674481 489395
rect 674415 489390 674784 489392
rect 674415 489334 674420 489390
rect 674476 489334 674784 489390
rect 674415 489332 674784 489334
rect 674415 489329 674481 489332
rect 674607 488800 674673 488803
rect 674607 488798 674814 488800
rect 674607 488742 674612 488798
rect 674668 488742 674814 488798
rect 674607 488740 674814 488742
rect 674607 488737 674673 488740
rect 674754 488622 674814 488740
rect 674170 487702 674176 487766
rect 674240 487764 674246 487766
rect 674240 487704 674784 487764
rect 674240 487702 674246 487704
rect 675130 487406 675136 487470
rect 675200 487406 675206 487470
rect 675138 486920 675198 487406
rect 673935 486136 674001 486139
rect 673935 486134 674784 486136
rect 673935 486078 673940 486134
rect 673996 486078 674784 486134
rect 673935 486076 674784 486078
rect 673935 486073 674001 486076
rect 674223 485322 674289 485325
rect 674223 485320 674784 485322
rect 674223 485264 674228 485320
rect 674284 485264 674784 485320
rect 674223 485262 674784 485264
rect 674223 485259 674289 485262
rect 59535 484804 59601 484807
rect 59535 484802 64416 484804
rect 59535 484746 59540 484802
rect 59596 484746 64416 484802
rect 59535 484744 64416 484746
rect 59535 484741 59601 484744
rect 674127 484656 674193 484659
rect 674127 484654 674784 484656
rect 674127 484598 674132 484654
rect 674188 484598 674784 484654
rect 674127 484596 674784 484598
rect 674127 484593 674193 484596
rect 674362 483780 674368 483844
rect 674432 483842 674438 483844
rect 674432 483782 674784 483842
rect 674432 483780 674438 483782
rect 674031 483028 674097 483031
rect 674031 483026 674784 483028
rect 674031 482970 674036 483026
rect 674092 482970 674784 483026
rect 674031 482968 674784 482970
rect 674031 482965 674097 482968
rect 674895 482436 674961 482439
rect 674895 482434 675006 482436
rect 674895 482378 674900 482434
rect 674956 482378 675006 482434
rect 674895 482373 675006 482378
rect 674946 482184 675006 482373
rect 654447 481844 654513 481847
rect 650208 481842 654513 481844
rect 650208 481786 654452 481842
rect 654508 481786 654513 481842
rect 650208 481784 654513 481786
rect 654447 481781 654513 481784
rect 679746 480811 679806 481370
rect 679746 480806 679857 480811
rect 679746 480750 679796 480806
rect 679852 480750 679857 480806
rect 679746 480748 679857 480750
rect 679791 480745 679857 480748
rect 679791 480068 679857 480071
rect 679746 480066 679857 480068
rect 679746 480010 679796 480066
rect 679852 480010 679857 480066
rect 679746 480005 679857 480010
rect 679746 479890 679806 480005
rect 59535 470448 59601 470451
rect 59535 470446 64416 470448
rect 59535 470390 59540 470446
rect 59596 470390 64416 470446
rect 59535 470388 64416 470390
rect 59535 470385 59601 470388
rect 654447 470300 654513 470303
rect 650208 470298 654513 470300
rect 650208 470242 654452 470298
rect 654508 470242 654513 470298
rect 650208 470240 654513 470242
rect 654447 470237 654513 470240
rect 656367 458460 656433 458463
rect 650208 458458 656433 458460
rect 650208 458402 656372 458458
rect 656428 458402 656433 458458
rect 650208 458400 656433 458402
rect 656367 458397 656433 458400
rect 59535 456092 59601 456095
rect 59535 456090 64416 456092
rect 59535 456034 59540 456090
rect 59596 456034 64416 456090
rect 59535 456032 64416 456034
rect 59535 456029 59601 456032
rect 654447 446620 654513 446623
rect 650208 446618 654513 446620
rect 650208 446562 654452 446618
rect 654508 446562 654513 446618
rect 650208 446560 654513 446562
rect 654447 446557 654513 446560
rect 57807 441588 57873 441591
rect 57807 441586 64416 441588
rect 57807 441530 57812 441586
rect 57868 441530 64416 441586
rect 57807 441528 64416 441530
rect 57807 441525 57873 441528
rect 42639 436926 42705 436929
rect 42336 436924 42705 436926
rect 42336 436868 42644 436924
rect 42700 436868 42705 436924
rect 42336 436866 42705 436868
rect 42639 436863 42705 436866
rect 42639 436112 42705 436115
rect 42336 436110 42705 436112
rect 42336 436054 42644 436110
rect 42700 436054 42705 436110
rect 42336 436052 42705 436054
rect 42639 436049 42705 436052
rect 42351 435520 42417 435523
rect 42306 435518 42417 435520
rect 42306 435462 42356 435518
rect 42412 435462 42417 435518
rect 42306 435457 42417 435462
rect 42306 435194 42366 435457
rect 654447 434928 654513 434931
rect 650208 434926 654513 434928
rect 650208 434870 654452 434926
rect 654508 434870 654513 434926
rect 650208 434868 654513 434870
rect 654447 434865 654513 434868
rect 43503 434484 43569 434487
rect 42336 434482 43569 434484
rect 42336 434426 43508 434482
rect 43564 434426 43569 434482
rect 42336 434424 43569 434426
rect 43503 434421 43569 434424
rect 43215 433596 43281 433599
rect 42336 433594 43281 433596
rect 42336 433538 43220 433594
rect 43276 433538 43281 433594
rect 42336 433536 43281 433538
rect 43215 433533 43281 433536
rect 43407 433004 43473 433007
rect 40608 433002 43473 433004
rect 40608 432974 43412 433002
rect 40578 432946 43412 432974
rect 43468 432946 43473 433002
rect 40578 432944 43473 432946
rect 40578 432710 40638 432944
rect 43407 432941 43473 432944
rect 40570 432646 40576 432710
rect 40640 432646 40646 432710
rect 43599 432116 43665 432119
rect 40416 432114 43665 432116
rect 40416 432086 43604 432114
rect 40386 432058 43604 432086
rect 43660 432058 43665 432114
rect 40386 432056 43665 432058
rect 40386 431970 40446 432056
rect 43599 432053 43665 432056
rect 40378 431906 40384 431970
rect 40448 431906 40454 431970
rect 40770 430786 40830 431346
rect 40762 430722 40768 430786
rect 40832 430722 40838 430786
rect 42114 429899 42174 430458
rect 42114 429894 42225 429899
rect 42114 429838 42164 429894
rect 42220 429838 42225 429894
rect 42114 429836 42225 429838
rect 42159 429833 42225 429836
rect 40962 429454 41022 429718
rect 40954 429390 40960 429454
rect 41024 429390 41030 429454
rect 41346 428418 41406 428830
rect 41338 428354 41344 428418
rect 41408 428354 41414 428418
rect 41538 427678 41598 428238
rect 41530 427614 41536 427678
rect 41600 427614 41606 427678
rect 59535 427380 59601 427383
rect 59535 427378 64416 427380
rect 41730 426791 41790 427350
rect 59535 427322 59540 427378
rect 59596 427322 64416 427378
rect 59535 427320 64416 427322
rect 59535 427317 59601 427320
rect 41730 426786 41841 426791
rect 41730 426730 41780 426786
rect 41836 426730 41841 426786
rect 41730 426728 41841 426730
rect 41775 426725 41841 426728
rect 41154 426346 41214 426536
rect 41146 426282 41152 426346
rect 41216 426282 41222 426346
rect 42114 425162 42174 425722
rect 42106 425098 42112 425162
rect 42176 425098 42182 425162
rect 37314 424423 37374 424908
rect 37314 424418 37425 424423
rect 37314 424362 37364 424418
rect 37420 424362 37425 424418
rect 37314 424360 37425 424362
rect 37359 424357 37425 424360
rect 42735 424124 42801 424127
rect 42336 424122 42801 424124
rect 42336 424066 42740 424122
rect 42796 424066 42801 424122
rect 42336 424064 42801 424066
rect 42735 424061 42801 424064
rect 40194 423239 40254 423428
rect 654447 423384 654513 423387
rect 650208 423382 654513 423384
rect 650208 423326 654452 423382
rect 654508 423326 654513 423382
rect 650208 423324 654513 423326
rect 654447 423321 654513 423324
rect 40143 423234 40254 423239
rect 40143 423178 40148 423234
rect 40204 423178 40254 423234
rect 40143 423176 40254 423178
rect 40143 423173 40209 423176
rect 37314 422055 37374 422614
rect 37263 422050 37374 422055
rect 37263 421994 37268 422050
rect 37324 421994 37374 422050
rect 37263 421992 37374 421994
rect 37263 421989 37329 421992
rect 42306 421312 42366 421800
rect 43023 421312 43089 421315
rect 42306 421310 43089 421312
rect 42306 421254 43028 421310
rect 43084 421254 43089 421310
rect 42306 421252 43089 421254
rect 43023 421249 43089 421252
rect 40194 420575 40254 420986
rect 40194 420570 40305 420575
rect 40194 420514 40244 420570
rect 40300 420514 40305 420570
rect 40194 420512 40305 420514
rect 40239 420509 40305 420512
rect 42639 420128 42705 420131
rect 42336 420126 42705 420128
rect 42336 420070 42644 420126
rect 42700 420070 42705 420126
rect 42336 420068 42705 420070
rect 42639 420065 42705 420068
rect 42639 418648 42705 418651
rect 42336 418646 42705 418648
rect 42336 418590 42644 418646
rect 42700 418590 42705 418646
rect 42336 418588 42705 418590
rect 42639 418585 42705 418588
rect 59535 412876 59601 412879
rect 59535 412874 64416 412876
rect 59535 412818 59540 412874
rect 59596 412818 64416 412874
rect 59535 412816 64416 412818
rect 59535 412813 59601 412816
rect 676527 412138 676593 412139
rect 676474 412136 676480 412138
rect 676436 412076 676480 412136
rect 676544 412134 676593 412138
rect 676588 412078 676593 412134
rect 676474 412074 676480 412076
rect 676544 412074 676593 412078
rect 676527 412073 676593 412074
rect 676623 411990 676689 411991
rect 676623 411986 676672 411990
rect 676736 411988 676742 411990
rect 676623 411930 676628 411986
rect 676623 411926 676672 411930
rect 676736 411928 676780 411988
rect 676736 411926 676742 411928
rect 676623 411925 676689 411926
rect 654447 411396 654513 411399
rect 650208 411394 654513 411396
rect 650208 411338 654452 411394
rect 654508 411338 654513 411394
rect 650208 411336 654513 411338
rect 654447 411333 654513 411336
rect 674754 409327 674814 409886
rect 674703 409322 674814 409327
rect 674703 409266 674708 409322
rect 674764 409266 674814 409322
rect 674703 409264 674814 409266
rect 674703 409261 674769 409264
rect 674415 409102 674481 409105
rect 674415 409100 674784 409102
rect 674415 409044 674420 409100
rect 674476 409044 674784 409100
rect 674415 409042 674784 409044
rect 674415 409039 674481 409042
rect 674703 408436 674769 408439
rect 674703 408434 674814 408436
rect 674703 408378 674708 408434
rect 674764 408378 674814 408434
rect 674703 408373 674814 408378
rect 674754 408258 674814 408373
rect 676719 407696 676785 407699
rect 676674 407694 676785 407696
rect 676674 407638 676724 407694
rect 676780 407638 676785 407694
rect 676674 407633 676785 407638
rect 676674 407444 676734 407633
rect 673839 406660 673905 406663
rect 673839 406658 674784 406660
rect 673839 406602 673844 406658
rect 673900 406602 674784 406658
rect 673839 406600 674784 406602
rect 673839 406597 673905 406600
rect 676474 406154 676480 406218
rect 676544 406154 676550 406218
rect 41530 406006 41536 406070
rect 41600 406068 41606 406070
rect 41775 406068 41841 406071
rect 41600 406066 41841 406068
rect 41600 406010 41780 406066
rect 41836 406010 41841 406066
rect 41600 406008 41841 406010
rect 41600 406006 41606 406008
rect 41775 406005 41841 406008
rect 674170 405858 674176 405922
rect 674240 405920 674246 405922
rect 676482 405920 676542 406154
rect 674240 405890 676542 405920
rect 674240 405860 676512 405890
rect 674240 405858 674246 405860
rect 675514 405266 675520 405330
rect 675584 405328 675590 405330
rect 676666 405328 676672 405330
rect 675584 405268 676672 405328
rect 675584 405266 675590 405268
rect 676666 405266 676672 405268
rect 676736 405266 676742 405330
rect 676674 405150 676734 405266
rect 41967 404886 42033 404887
rect 41914 404884 41920 404886
rect 41876 404824 41920 404884
rect 41984 404882 42033 404886
rect 42028 404826 42033 404882
rect 41914 404822 41920 404824
rect 41984 404822 42033 404826
rect 41967 404821 42033 404822
rect 674946 404147 675006 404262
rect 674895 404142 675006 404147
rect 674895 404086 674900 404142
rect 674956 404086 675006 404142
rect 674895 404084 675006 404086
rect 674895 404081 674961 404084
rect 41775 403850 41841 403851
rect 41722 403786 41728 403850
rect 41792 403848 41841 403850
rect 41792 403846 41884 403848
rect 41836 403790 41884 403846
rect 41792 403788 41884 403790
rect 41792 403786 41841 403788
rect 41775 403785 41841 403786
rect 674946 403258 675006 403522
rect 674938 403194 674944 403258
rect 675008 403194 675014 403258
rect 42159 402666 42225 402667
rect 42106 402664 42112 402666
rect 42068 402604 42112 402664
rect 42176 402662 42225 402666
rect 42220 402606 42225 402662
rect 42106 402602 42112 402604
rect 42176 402602 42225 402606
rect 42159 402601 42225 402602
rect 675330 402519 675390 402634
rect 675279 402514 675390 402519
rect 675279 402458 675284 402514
rect 675340 402458 675390 402514
rect 675279 402456 675390 402458
rect 675279 402453 675345 402456
rect 41338 401862 41344 401926
rect 41408 401924 41414 401926
rect 41775 401924 41841 401927
rect 41408 401922 41841 401924
rect 41408 401866 41780 401922
rect 41836 401866 41841 401922
rect 41408 401864 41841 401866
rect 41408 401862 41414 401864
rect 41775 401861 41841 401864
rect 674031 401924 674097 401927
rect 674031 401922 674784 401924
rect 674031 401866 674036 401922
rect 674092 401866 674784 401922
rect 674031 401864 674784 401866
rect 674031 401861 674097 401864
rect 674554 400530 674560 400594
rect 674624 400592 674630 400594
rect 674754 400592 674814 401154
rect 674624 400532 674814 400592
rect 674624 400530 674630 400532
rect 674362 400382 674368 400446
rect 674432 400444 674438 400446
rect 674432 400384 674784 400444
rect 674432 400382 674438 400384
rect 40762 400086 40768 400150
rect 40832 400148 40838 400150
rect 41775 400148 41841 400151
rect 40832 400146 41841 400148
rect 40832 400090 41780 400146
rect 41836 400090 41841 400146
rect 40832 400088 41841 400090
rect 40832 400086 40838 400088
rect 41775 400085 41841 400088
rect 41914 399938 41920 400002
rect 41984 400000 41990 400002
rect 42255 400000 42321 400003
rect 41984 399998 42321 400000
rect 41984 399942 42260 399998
rect 42316 399942 42321 399998
rect 41984 399940 42321 399942
rect 41984 399938 41990 399940
rect 42255 399937 42321 399940
rect 654639 399704 654705 399707
rect 650208 399702 654705 399704
rect 650208 399646 654644 399702
rect 654700 399646 654705 399702
rect 650208 399644 654705 399646
rect 654639 399641 654705 399644
rect 41146 399494 41152 399558
rect 41216 399556 41222 399558
rect 41775 399556 41841 399559
rect 41216 399554 41841 399556
rect 41216 399498 41780 399554
rect 41836 399498 41841 399554
rect 41216 399496 41841 399498
rect 41216 399494 41222 399496
rect 41775 399493 41841 399496
rect 675138 399411 675198 399526
rect 675138 399406 675249 399411
rect 675138 399350 675188 399406
rect 675244 399350 675249 399406
rect 675138 399348 675249 399350
rect 675183 399345 675249 399348
rect 40954 398754 40960 398818
rect 41024 398816 41030 398818
rect 41775 398816 41841 398819
rect 41024 398814 41841 398816
rect 41024 398758 41780 398814
rect 41836 398758 41841 398814
rect 41024 398756 41841 398758
rect 41024 398754 41030 398756
rect 41775 398753 41841 398756
rect 58959 398668 59025 398671
rect 58959 398666 64416 398668
rect 58959 398610 58964 398666
rect 59020 398610 64416 398666
rect 58959 398608 64416 398610
rect 58959 398605 59025 398608
rect 674946 398523 675006 398786
rect 674946 398518 675057 398523
rect 674946 398462 674996 398518
rect 675052 398462 675057 398518
rect 674946 398460 675057 398462
rect 674991 398457 675057 398460
rect 674511 397780 674577 397783
rect 674754 397780 674814 397898
rect 674511 397778 674814 397780
rect 674511 397722 674516 397778
rect 674572 397722 674814 397778
rect 674511 397720 674814 397722
rect 674511 397717 674577 397720
rect 673935 397188 674001 397191
rect 673935 397186 674784 397188
rect 673935 397130 673940 397186
rect 673996 397130 674784 397186
rect 673935 397128 674784 397130
rect 673935 397125 674001 397128
rect 674415 396448 674481 396451
rect 674415 396446 674784 396448
rect 674415 396390 674420 396446
rect 674476 396390 674784 396446
rect 674415 396388 674784 396390
rect 674415 396385 674481 396388
rect 674754 395415 674814 395604
rect 674754 395410 674865 395415
rect 674754 395354 674804 395410
rect 674860 395354 674865 395410
rect 674754 395352 674865 395354
rect 674799 395349 674865 395352
rect 674754 394527 674814 394790
rect 674703 394522 674814 394527
rect 674703 394466 674708 394522
rect 674764 394466 674814 394522
rect 674703 394464 674814 394466
rect 674703 394461 674769 394464
rect 674319 394006 674385 394009
rect 674319 394004 674784 394006
rect 674319 393948 674324 394004
rect 674380 393948 674784 394004
rect 674319 393946 674784 393948
rect 674319 393943 674385 393946
rect 42351 393932 42417 393935
rect 42306 393930 42417 393932
rect 42306 393874 42356 393930
rect 42412 393874 42417 393930
rect 42306 393869 42417 393874
rect 42306 393680 42366 393869
rect 42351 393192 42417 393195
rect 42306 393190 42417 393192
rect 42306 393134 42356 393190
rect 42412 393134 42417 393190
rect 42306 393129 42417 393134
rect 42306 392866 42366 393129
rect 679746 392603 679806 393162
rect 679695 392598 679806 392603
rect 679695 392542 679700 392598
rect 679756 392542 679806 392598
rect 679695 392540 679806 392542
rect 679695 392537 679761 392540
rect 42351 392304 42417 392307
rect 42306 392302 42417 392304
rect 42306 392246 42356 392302
rect 42412 392246 42417 392302
rect 42306 392241 42417 392246
rect 42306 392052 42366 392241
rect 679695 392156 679761 392159
rect 679695 392154 679806 392156
rect 679695 392098 679700 392154
rect 679756 392098 679806 392154
rect 679695 392093 679806 392098
rect 679746 391682 679806 392093
rect 43215 391268 43281 391271
rect 42336 391266 43281 391268
rect 42336 391210 43220 391266
rect 43276 391210 43281 391266
rect 42336 391208 43281 391210
rect 43215 391205 43281 391208
rect 43119 390972 43185 390975
rect 42306 390970 43185 390972
rect 42306 390914 43124 390970
rect 43180 390914 43185 390970
rect 42306 390912 43185 390914
rect 42306 390424 42366 390912
rect 43119 390909 43185 390912
rect 40570 390170 40576 390234
rect 40640 390170 40646 390234
rect 40578 389758 40638 390170
rect 40378 389134 40384 389198
rect 40448 389134 40454 389198
rect 40386 388870 40446 389134
rect 40770 387570 40830 388130
rect 654447 388012 654513 388015
rect 650208 388010 654513 388012
rect 650208 387954 654452 388010
rect 654508 387954 654513 388010
rect 650208 387952 654513 387954
rect 654447 387949 654513 387952
rect 40762 387506 40768 387570
rect 40832 387506 40838 387570
rect 43023 387272 43089 387275
rect 42336 387270 43089 387272
rect 42336 387214 43028 387270
rect 43084 387214 43089 387270
rect 42336 387212 43089 387214
rect 43023 387209 43089 387212
rect 40962 386090 41022 386502
rect 40954 386026 40960 386090
rect 41024 386026 41030 386090
rect 41346 385202 41406 385614
rect 41338 385138 41344 385202
rect 41408 385138 41414 385202
rect 35970 384463 36030 385022
rect 35919 384458 36030 384463
rect 35919 384402 35924 384458
rect 35980 384402 36030 384458
rect 35919 384400 36030 384402
rect 35919 384397 35985 384400
rect 59535 384164 59601 384167
rect 59535 384162 64416 384164
rect 41730 383575 41790 384134
rect 59535 384106 59540 384162
rect 59596 384106 64416 384162
rect 59535 384104 64416 384106
rect 59535 384101 59601 384104
rect 41730 383570 41841 383575
rect 41730 383514 41780 383570
rect 41836 383514 41841 383570
rect 41730 383512 41841 383514
rect 41775 383509 41841 383512
rect 41154 383130 41214 383394
rect 41146 383066 41152 383130
rect 41216 383066 41222 383130
rect 41538 381946 41598 382506
rect 41530 381882 41536 381946
rect 41600 381882 41606 381946
rect 37122 381207 37182 381766
rect 37122 381202 37233 381207
rect 37122 381146 37172 381202
rect 37228 381146 37233 381202
rect 37122 381144 37233 381146
rect 37167 381141 37233 381144
rect 40002 380467 40062 380878
rect 40002 380462 40113 380467
rect 40002 380406 40052 380462
rect 40108 380406 40113 380462
rect 40002 380404 40113 380406
rect 40047 380401 40113 380404
rect 42927 380316 42993 380319
rect 42306 380314 42993 380316
rect 42306 380258 42932 380314
rect 42988 380258 42993 380314
rect 42306 380256 42993 380258
rect 42306 380212 42366 380256
rect 42927 380253 42993 380256
rect 37314 378839 37374 379398
rect 37263 378834 37374 378839
rect 37263 378778 37268 378834
rect 37324 378778 37374 378834
rect 37263 378776 37374 378778
rect 37263 378773 37329 378776
rect 674554 378774 674560 378838
rect 674624 378836 674630 378838
rect 675471 378836 675537 378839
rect 674624 378834 675537 378836
rect 674624 378778 675476 378834
rect 675532 378778 675537 378834
rect 674624 378776 675537 378778
rect 674624 378774 674630 378776
rect 675471 378773 675537 378776
rect 37314 378099 37374 378584
rect 37314 378094 37425 378099
rect 37314 378038 37364 378094
rect 37420 378038 37425 378094
rect 37314 378036 37425 378038
rect 37359 378033 37425 378036
rect 40194 377507 40254 377770
rect 40143 377502 40254 377507
rect 40143 377446 40148 377502
rect 40204 377446 40254 377502
rect 40143 377444 40254 377446
rect 40143 377441 40209 377444
rect 42306 376767 42366 376956
rect 42306 376762 42417 376767
rect 42306 376706 42356 376762
rect 42412 376706 42417 376762
rect 42306 376704 42417 376706
rect 42351 376701 42417 376704
rect 654447 376468 654513 376471
rect 650208 376466 654513 376468
rect 650208 376410 654452 376466
rect 654508 376410 654513 376466
rect 650208 376408 654513 376410
rect 654447 376405 654513 376408
rect 42306 375287 42366 375402
rect 42306 375282 42417 375287
rect 42306 375226 42356 375282
rect 42412 375226 42417 375282
rect 42306 375224 42417 375226
rect 42351 375221 42417 375224
rect 675087 374544 675153 374547
rect 675322 374544 675328 374546
rect 675087 374542 675328 374544
rect 675087 374486 675092 374542
rect 675148 374486 675328 374542
rect 675087 374484 675328 374486
rect 675087 374481 675153 374484
rect 675322 374482 675328 374484
rect 675392 374482 675398 374546
rect 674938 373890 674944 373954
rect 675008 373952 675014 373954
rect 675471 373952 675537 373955
rect 675008 373950 675537 373952
rect 675008 373894 675476 373950
rect 675532 373894 675537 373950
rect 675008 373892 675537 373894
rect 675008 373890 675014 373892
rect 675471 373889 675537 373892
rect 674362 371966 674368 372030
rect 674432 372028 674438 372030
rect 675375 372028 675441 372031
rect 674432 372026 675441 372028
rect 674432 371970 675380 372026
rect 675436 371970 675441 372026
rect 674432 371968 675441 371970
rect 674432 371966 674438 371968
rect 675375 371965 675441 371968
rect 675183 371732 675249 371735
rect 675706 371732 675712 371734
rect 675183 371730 675712 371732
rect 675183 371674 675188 371730
rect 675244 371674 675712 371730
rect 675183 371672 675712 371674
rect 675183 371669 675249 371672
rect 675706 371670 675712 371672
rect 675776 371670 675782 371734
rect 35919 371584 35985 371587
rect 42106 371584 42112 371586
rect 35919 371582 42112 371584
rect 35919 371526 35924 371582
rect 35980 371526 42112 371582
rect 35919 371524 42112 371526
rect 35919 371521 35985 371524
rect 42106 371522 42112 371524
rect 42176 371522 42182 371586
rect 59535 369808 59601 369811
rect 59535 369806 64416 369808
rect 59535 369750 59540 369806
rect 59596 369750 64416 369806
rect 59535 369748 64416 369750
rect 59535 369745 59601 369748
rect 674703 364924 674769 364927
rect 674703 364922 674814 364924
rect 674703 364866 674708 364922
rect 674764 364866 674814 364922
rect 674703 364861 674814 364866
rect 674754 364672 674814 364861
rect 654447 364480 654513 364483
rect 650208 364478 654513 364480
rect 650208 364422 654452 364478
rect 654508 364422 654513 364478
rect 650208 364420 654513 364422
rect 654447 364417 654513 364420
rect 674415 363888 674481 363891
rect 674415 363886 674784 363888
rect 674415 363830 674420 363886
rect 674476 363830 674784 363886
rect 674415 363828 674784 363830
rect 674415 363825 674481 363828
rect 674703 363296 674769 363299
rect 674703 363294 674814 363296
rect 674703 363238 674708 363294
rect 674764 363238 674814 363294
rect 674703 363233 674814 363238
rect 674754 363044 674814 363233
rect 42063 362854 42129 362855
rect 42063 362850 42112 362854
rect 42176 362852 42182 362854
rect 42063 362794 42068 362850
rect 42063 362790 42112 362794
rect 42176 362792 42220 362852
rect 42176 362790 42182 362792
rect 42063 362789 42129 362790
rect 673839 362260 673905 362263
rect 673839 362258 674784 362260
rect 673839 362202 673844 362258
rect 673900 362202 674784 362258
rect 673839 362200 674784 362202
rect 673839 362197 673905 362200
rect 41871 361966 41937 361967
rect 41871 361964 41920 361966
rect 41828 361962 41920 361964
rect 41828 361906 41876 361962
rect 41828 361904 41920 361906
rect 41871 361902 41920 361904
rect 41984 361902 41990 361966
rect 41871 361901 41937 361902
rect 674362 361384 674368 361448
rect 674432 361446 674438 361448
rect 674432 361386 674784 361446
rect 674432 361384 674438 361386
rect 41775 361374 41841 361375
rect 41722 361310 41728 361374
rect 41792 361372 41841 361374
rect 41792 361370 41884 361372
rect 41836 361314 41884 361370
rect 41792 361312 41884 361314
rect 41792 361310 41841 361312
rect 41775 361309 41841 361310
rect 674170 360718 674176 360782
rect 674240 360780 674246 360782
rect 674240 360720 674784 360780
rect 674240 360718 674246 360720
rect 675514 360126 675520 360190
rect 675584 360126 675590 360190
rect 673978 359978 673984 360042
rect 674048 360040 674054 360042
rect 675522 360040 675582 360126
rect 674048 359980 675582 360040
rect 674048 359978 674054 359980
rect 675522 359936 675582 359980
rect 41530 359386 41536 359450
rect 41600 359448 41606 359450
rect 41775 359448 41841 359451
rect 41600 359446 41841 359448
rect 41600 359390 41780 359446
rect 41836 359390 41841 359446
rect 41600 359388 41841 359390
rect 41600 359386 41606 359388
rect 41775 359385 41841 359388
rect 674031 359152 674097 359155
rect 674031 359150 674784 359152
rect 674031 359094 674036 359150
rect 674092 359094 674784 359150
rect 674031 359092 674784 359094
rect 674031 359089 674097 359092
rect 41338 358646 41344 358710
rect 41408 358708 41414 358710
rect 41775 358708 41841 358711
rect 41408 358706 41841 358708
rect 41408 358650 41780 358706
rect 41836 358650 41841 358706
rect 41408 358648 41841 358650
rect 41408 358646 41414 358648
rect 41775 358645 41841 358648
rect 677058 358119 677118 358234
rect 677058 358114 677169 358119
rect 677058 358058 677108 358114
rect 677164 358058 677169 358114
rect 677058 358056 677169 358058
rect 677103 358053 677169 358056
rect 674607 357228 674673 357231
rect 674754 357228 674814 357494
rect 674607 357226 674814 357228
rect 674607 357170 674612 357226
rect 674668 357170 674814 357226
rect 674607 357168 674814 357170
rect 674607 357165 674673 357168
rect 40762 356870 40768 356934
rect 40832 356932 40838 356934
rect 41871 356932 41937 356935
rect 40832 356930 41937 356932
rect 40832 356874 41876 356930
rect 41932 356874 41937 356930
rect 40832 356872 41937 356874
rect 40832 356870 40838 356872
rect 41871 356869 41937 356872
rect 675138 356491 675198 356606
rect 41146 356426 41152 356490
rect 41216 356488 41222 356490
rect 41775 356488 41841 356491
rect 41216 356486 41841 356488
rect 41216 356430 41780 356486
rect 41836 356430 41841 356486
rect 41216 356428 41841 356430
rect 675138 356486 675249 356491
rect 675138 356430 675188 356486
rect 675244 356430 675249 356486
rect 675138 356428 675249 356430
rect 41216 356426 41222 356428
rect 41775 356425 41841 356428
rect 675183 356425 675249 356428
rect 676866 355751 676926 356014
rect 676866 355746 676977 355751
rect 676866 355690 676916 355746
rect 676972 355690 676977 355746
rect 676866 355688 676977 355690
rect 676911 355685 676977 355688
rect 40954 355538 40960 355602
rect 41024 355600 41030 355602
rect 41775 355600 41841 355603
rect 41024 355598 41841 355600
rect 41024 355542 41780 355598
rect 41836 355542 41841 355598
rect 41024 355540 41841 355542
rect 41024 355538 41030 355540
rect 41775 355537 41841 355540
rect 59535 355600 59601 355603
rect 59535 355598 64416 355600
rect 59535 355542 59540 355598
rect 59596 355542 64416 355598
rect 59535 355540 64416 355542
rect 59535 355537 59601 355540
rect 677058 355011 677118 355126
rect 677007 355006 677118 355011
rect 677007 354950 677012 355006
rect 677068 354950 677118 355006
rect 677007 354948 677118 354950
rect 677007 354945 677073 354948
rect 675330 354123 675390 354386
rect 675279 354118 675390 354123
rect 675279 354062 675284 354118
rect 675340 354062 675390 354118
rect 675279 354060 675390 354062
rect 675279 354057 675345 354060
rect 675138 353383 675198 353498
rect 675087 353378 675198 353383
rect 675087 353322 675092 353378
rect 675148 353322 675198 353378
rect 675087 353320 675198 353322
rect 675087 353317 675153 353320
rect 655311 352788 655377 352791
rect 650208 352786 655377 352788
rect 650208 352730 655316 352786
rect 655372 352730 655377 352786
rect 650208 352728 655377 352730
rect 655311 352725 655377 352728
rect 674511 352492 674577 352495
rect 674754 352492 674814 352758
rect 674511 352490 674814 352492
rect 674511 352434 674516 352490
rect 674572 352434 674814 352490
rect 674511 352432 674814 352434
rect 674511 352429 674577 352432
rect 676866 351755 676926 351870
rect 676815 351750 676926 351755
rect 676815 351694 676820 351750
rect 676876 351694 676926 351750
rect 676815 351692 676926 351694
rect 676815 351689 676881 351692
rect 674223 351308 674289 351311
rect 674223 351306 674784 351308
rect 674223 351250 674228 351306
rect 674284 351250 674784 351306
rect 674223 351248 674784 351250
rect 674223 351245 674289 351248
rect 42351 350716 42417 350719
rect 42306 350714 42417 350716
rect 42306 350658 42356 350714
rect 42412 350658 42417 350714
rect 42306 350653 42417 350658
rect 42306 350538 42366 350653
rect 674754 350275 674814 350390
rect 674754 350270 674865 350275
rect 674754 350214 674804 350270
rect 674860 350214 674865 350270
rect 674754 350212 674865 350214
rect 674799 350209 674865 350212
rect 42639 349680 42705 349683
rect 42336 349678 42705 349680
rect 42336 349622 42644 349678
rect 42700 349622 42705 349678
rect 42336 349620 42705 349622
rect 42639 349617 42705 349620
rect 674319 349606 674385 349609
rect 674319 349604 674784 349606
rect 674319 349548 674324 349604
rect 674380 349548 674784 349604
rect 674319 349546 674784 349548
rect 674319 349543 674385 349546
rect 42351 349088 42417 349091
rect 42306 349086 42417 349088
rect 42306 349030 42356 349086
rect 42412 349030 42417 349086
rect 42306 349025 42417 349030
rect 42306 348910 42366 349025
rect 674127 348792 674193 348795
rect 674127 348790 674784 348792
rect 674127 348734 674132 348790
rect 674188 348734 674784 348790
rect 674127 348732 674784 348734
rect 674127 348729 674193 348732
rect 42306 347904 42366 348022
rect 42306 347844 43518 347904
rect 43215 347756 43281 347759
rect 42306 347754 43281 347756
rect 42306 347698 43220 347754
rect 43276 347698 43281 347754
rect 42306 347696 43281 347698
rect 42306 347208 42366 347696
rect 43215 347693 43281 347696
rect 43215 347608 43281 347611
rect 43458 347608 43518 347844
rect 43215 347606 43518 347608
rect 43215 347550 43220 347606
rect 43276 347550 43518 347606
rect 43215 347548 43518 347550
rect 43215 347545 43281 347548
rect 679746 347463 679806 347948
rect 679746 347458 679857 347463
rect 679746 347402 679796 347458
rect 679852 347402 679857 347458
rect 679746 347400 679857 347402
rect 679791 347397 679857 347400
rect 40570 346806 40576 346870
rect 40640 346806 40646 346870
rect 40578 346572 40638 346806
rect 679791 346720 679857 346723
rect 679746 346718 679857 346720
rect 679746 346662 679796 346718
rect 679852 346662 679857 346718
rect 679746 346657 679857 346662
rect 40578 346542 42144 346572
rect 40608 346512 42174 346542
rect 42114 346278 42174 346512
rect 679746 346468 679806 346657
rect 42106 346214 42112 346278
rect 42176 346214 42182 346278
rect 40378 345918 40384 345982
rect 40448 345980 40454 345982
rect 42298 345980 42304 345982
rect 40448 345920 42304 345980
rect 40448 345918 40454 345920
rect 42298 345918 42304 345920
rect 42368 345918 42374 345982
rect 42306 345728 42366 345918
rect 676666 345474 676672 345538
rect 676736 345536 676742 345538
rect 677103 345536 677169 345539
rect 676736 345534 677169 345536
rect 676736 345478 677108 345534
rect 677164 345478 677169 345534
rect 676736 345476 677169 345478
rect 676736 345474 676742 345476
rect 677103 345473 677169 345476
rect 676090 345326 676096 345390
rect 676160 345388 676166 345390
rect 676911 345388 676977 345391
rect 676160 345386 676977 345388
rect 676160 345330 676916 345386
rect 676972 345330 676977 345386
rect 676160 345328 676977 345330
rect 676160 345326 676166 345328
rect 676911 345325 676977 345328
rect 676474 345178 676480 345242
rect 676544 345240 676550 345242
rect 677007 345240 677073 345243
rect 676544 345238 677073 345240
rect 676544 345182 677012 345238
rect 677068 345182 677073 345238
rect 676544 345180 677073 345182
rect 676544 345178 676550 345180
rect 677007 345177 677073 345180
rect 40962 344354 41022 344914
rect 676282 344438 676288 344502
rect 676352 344500 676358 344502
rect 676815 344500 676881 344503
rect 676352 344498 676881 344500
rect 676352 344442 676820 344498
rect 676876 344442 676881 344498
rect 676352 344440 676881 344442
rect 676352 344438 676358 344440
rect 676815 344437 676881 344440
rect 40954 344290 40960 344354
rect 41024 344290 41030 344354
rect 42735 344130 42801 344133
rect 42336 344128 42801 344130
rect 42336 344072 42740 344128
rect 42796 344072 42801 344128
rect 42336 344070 42801 344072
rect 42735 344067 42801 344070
rect 40770 342874 40830 343286
rect 40762 342810 40768 342874
rect 40832 342810 40838 342874
rect 41346 341986 41406 342472
rect 41338 341922 41344 341986
rect 41408 341922 41414 341986
rect 40386 341246 40446 341806
rect 40378 341182 40384 341246
rect 40448 341182 40454 341246
rect 59535 341096 59601 341099
rect 654447 341096 654513 341099
rect 59535 341094 64416 341096
rect 59535 341038 59540 341094
rect 59596 341038 64416 341094
rect 59535 341036 64416 341038
rect 650208 341094 654513 341096
rect 650208 341038 654452 341094
rect 654508 341038 654513 341094
rect 650208 341036 654513 341038
rect 59535 341033 59601 341036
rect 654447 341033 654513 341036
rect 40002 340359 40062 340918
rect 39951 340354 40062 340359
rect 39951 340298 39956 340354
rect 40012 340298 40062 340354
rect 39951 340296 40062 340298
rect 39951 340293 40017 340296
rect 41154 339914 41214 340178
rect 41146 339850 41152 339914
rect 41216 339850 41222 339914
rect 41538 338730 41598 339290
rect 41530 338666 41536 338730
rect 41600 338666 41606 338730
rect 42306 337991 42366 338550
rect 42306 337986 42417 337991
rect 42306 337930 42356 337986
rect 42412 337930 42417 337986
rect 42306 337928 42417 337930
rect 42351 337925 42417 337928
rect 37122 337399 37182 337662
rect 37122 337394 37233 337399
rect 37122 337338 37172 337394
rect 37228 337338 37233 337394
rect 37122 337336 37233 337338
rect 37167 337333 37233 337336
rect 40047 337248 40113 337251
rect 40002 337246 40113 337248
rect 40002 337190 40052 337246
rect 40108 337190 40113 337246
rect 40002 337185 40113 337190
rect 40002 337070 40062 337185
rect 42682 336212 42688 336214
rect 42336 336152 42688 336212
rect 42682 336150 42688 336152
rect 42752 336150 42758 336214
rect 43119 335472 43185 335475
rect 42336 335470 43185 335472
rect 42336 335414 43124 335470
rect 43180 335414 43185 335470
rect 42336 335412 43185 335414
rect 43119 335409 43185 335412
rect 675279 335030 675345 335031
rect 675279 335026 675328 335030
rect 675392 335028 675398 335030
rect 675279 334970 675284 335026
rect 675279 334966 675328 334970
rect 675392 334968 675436 335028
rect 675392 334966 675398 334968
rect 675279 334965 675345 334966
rect 40194 334143 40254 334554
rect 40194 334138 40305 334143
rect 40194 334082 40244 334138
rect 40300 334082 40305 334138
rect 40194 334080 40305 334082
rect 40239 334077 40305 334080
rect 675567 333846 675633 333847
rect 42114 333551 42174 333814
rect 675514 333782 675520 333846
rect 675584 333844 675633 333846
rect 675584 333842 675676 333844
rect 675628 333786 675676 333842
rect 675584 333784 675676 333786
rect 675584 333782 675633 333784
rect 675567 333781 675633 333782
rect 42114 333546 42225 333551
rect 42114 333490 42164 333546
rect 42220 333490 42225 333546
rect 42114 333488 42225 333490
rect 42159 333485 42225 333488
rect 675759 333548 675825 333551
rect 676090 333548 676096 333550
rect 675759 333546 676096 333548
rect 675759 333490 675764 333546
rect 675820 333490 676096 333546
rect 675759 333488 676096 333490
rect 675759 333485 675825 333488
rect 676090 333486 676096 333488
rect 676160 333486 676166 333550
rect 42114 332071 42174 332260
rect 42114 332066 42225 332071
rect 42114 332010 42164 332066
rect 42220 332010 42225 332066
rect 42114 332008 42225 332010
rect 42159 332005 42225 332008
rect 675759 330588 675825 330591
rect 676282 330588 676288 330590
rect 675759 330586 676288 330588
rect 675759 330530 675764 330586
rect 675820 330530 676288 330586
rect 675759 330528 676288 330530
rect 675759 330525 675825 330528
rect 676282 330526 676288 330528
rect 676352 330526 676358 330590
rect 654063 329552 654129 329555
rect 650208 329550 654129 329552
rect 650208 329494 654068 329550
rect 654124 329494 654129 329550
rect 650208 329492 654129 329494
rect 654063 329489 654129 329492
rect 675183 329552 675249 329555
rect 675322 329552 675328 329554
rect 675183 329550 675328 329552
rect 675183 329494 675188 329550
rect 675244 329494 675328 329550
rect 675183 329492 675328 329494
rect 675183 329489 675249 329492
rect 675322 329490 675328 329492
rect 675392 329490 675398 329554
rect 675759 328072 675825 328075
rect 676666 328072 676672 328074
rect 675759 328070 676672 328072
rect 675759 328014 675764 328070
rect 675820 328014 676672 328070
rect 675759 328012 676672 328014
rect 675759 328009 675825 328012
rect 676666 328010 676672 328012
rect 676736 328010 676742 328074
rect 42351 327480 42417 327483
rect 42490 327480 42496 327482
rect 42351 327478 42496 327480
rect 42351 327422 42356 327478
rect 42412 327422 42496 327478
rect 42351 327420 42496 327422
rect 42351 327417 42417 327420
rect 42490 327418 42496 327420
rect 42560 327418 42566 327482
rect 675759 326888 675825 326891
rect 676474 326888 676480 326890
rect 675759 326886 676480 326888
rect 675759 326830 675764 326886
rect 675820 326830 676480 326886
rect 675759 326828 676480 326830
rect 675759 326825 675825 326828
rect 676474 326826 676480 326828
rect 676544 326826 676550 326890
rect 59535 326740 59601 326743
rect 59535 326738 64416 326740
rect 59535 326682 59540 326738
rect 59596 326682 64416 326738
rect 59535 326680 64416 326682
rect 59535 326677 59601 326680
rect 42351 323040 42417 323043
rect 42490 323040 42496 323042
rect 42351 323038 42496 323040
rect 42351 322982 42356 323038
rect 42412 322982 42496 323038
rect 42351 322980 42496 322982
rect 42351 322977 42417 322980
rect 42490 322978 42496 322980
rect 42560 322978 42566 323042
rect 40378 319722 40384 319786
rect 40448 319784 40454 319786
rect 41775 319784 41841 319787
rect 40448 319782 41841 319784
rect 40448 319726 41780 319782
rect 41836 319726 41841 319782
rect 40448 319724 41841 319726
rect 40448 319722 40454 319724
rect 41775 319721 41841 319724
rect 674415 319710 674481 319713
rect 674415 319708 674784 319710
rect 674415 319652 674420 319708
rect 674476 319652 674784 319708
rect 674415 319650 674784 319652
rect 674415 319647 674481 319650
rect 674415 318896 674481 318899
rect 674415 318894 674784 318896
rect 674415 318838 674420 318894
rect 674476 318838 674784 318894
rect 674415 318836 674784 318838
rect 674415 318833 674481 318836
rect 41871 318750 41937 318751
rect 41871 318748 41920 318750
rect 41828 318746 41920 318748
rect 41828 318690 41876 318746
rect 41828 318688 41920 318690
rect 41871 318686 41920 318688
rect 41984 318686 41990 318750
rect 41871 318685 41937 318686
rect 674703 318304 674769 318307
rect 674703 318302 674814 318304
rect 674703 318246 674708 318302
rect 674764 318246 674814 318302
rect 674703 318241 674814 318246
rect 674754 318052 674814 318241
rect 41775 318010 41841 318011
rect 41722 317946 41728 318010
rect 41792 318008 41841 318010
rect 41792 318006 41884 318008
rect 41836 317950 41884 318006
rect 41792 317948 41884 317950
rect 41792 317946 41841 317948
rect 41775 317945 41841 317946
rect 655119 317564 655185 317567
rect 650208 317562 655185 317564
rect 650208 317506 655124 317562
rect 655180 317506 655185 317562
rect 650208 317504 655185 317506
rect 655119 317501 655185 317504
rect 42159 317416 42225 317419
rect 42682 317416 42688 317418
rect 42159 317414 42688 317416
rect 42159 317358 42164 317414
rect 42220 317358 42688 317414
rect 42159 317356 42688 317358
rect 42159 317353 42225 317356
rect 42682 317354 42688 317356
rect 42752 317354 42758 317418
rect 674362 317206 674368 317270
rect 674432 317268 674438 317270
rect 674432 317208 674784 317268
rect 674432 317206 674438 317208
rect 674362 316392 674368 316456
rect 674432 316454 674438 316456
rect 674432 316394 674784 316454
rect 674432 316392 674438 316394
rect 41530 316170 41536 316234
rect 41600 316232 41606 316234
rect 41775 316232 41841 316235
rect 41600 316230 41841 316232
rect 41600 316174 41780 316230
rect 41836 316174 41841 316230
rect 41600 316172 41841 316174
rect 41600 316170 41606 316172
rect 41775 316169 41841 316172
rect 674170 315726 674176 315790
rect 674240 315788 674246 315790
rect 674240 315728 674784 315788
rect 674240 315726 674246 315728
rect 41338 315430 41344 315494
rect 41408 315492 41414 315494
rect 41775 315492 41841 315495
rect 41408 315490 41841 315492
rect 41408 315434 41780 315490
rect 41836 315434 41841 315490
rect 41408 315432 41841 315434
rect 41408 315430 41414 315432
rect 41775 315429 41841 315432
rect 673978 314838 673984 314902
rect 674048 314900 674054 314902
rect 674048 314840 674784 314900
rect 674048 314838 674054 314840
rect 673935 314160 674001 314163
rect 673935 314158 674784 314160
rect 673935 314102 673940 314158
rect 673996 314102 674784 314158
rect 673935 314100 674784 314102
rect 673935 314097 674001 314100
rect 40954 313654 40960 313718
rect 41024 313716 41030 313718
rect 41775 313716 41841 313719
rect 41024 313714 41841 313716
rect 41024 313658 41780 313714
rect 41836 313658 41841 313714
rect 41024 313656 41841 313658
rect 41024 313654 41030 313656
rect 41775 313653 41841 313656
rect 41146 313210 41152 313274
rect 41216 313272 41222 313274
rect 41775 313272 41841 313275
rect 41216 313270 41841 313272
rect 41216 313214 41780 313270
rect 41836 313214 41841 313270
rect 41216 313212 41841 313214
rect 41216 313210 41222 313212
rect 41775 313209 41841 313212
rect 674554 312618 674560 312682
rect 674624 312680 674630 312682
rect 674754 312680 674814 313242
rect 674624 312620 674814 312680
rect 674624 312618 674630 312620
rect 674319 312532 674385 312535
rect 674319 312530 674784 312532
rect 674319 312474 674324 312530
rect 674380 312474 674784 312530
rect 674319 312472 674784 312474
rect 674319 312469 674385 312472
rect 40762 312322 40768 312386
rect 40832 312384 40838 312386
rect 41775 312384 41841 312387
rect 40832 312382 41841 312384
rect 40832 312326 41780 312382
rect 41836 312326 41841 312382
rect 40832 312324 41841 312326
rect 40832 312322 40838 312324
rect 41775 312321 41841 312324
rect 59535 312384 59601 312387
rect 59535 312382 64416 312384
rect 59535 312326 59540 312382
rect 59596 312326 64416 312382
rect 59535 312324 64416 312326
rect 59535 312321 59601 312324
rect 677058 311499 677118 311614
rect 677058 311494 677169 311499
rect 677058 311438 677108 311494
rect 677164 311438 677169 311494
rect 677058 311436 677169 311438
rect 677103 311433 677169 311436
rect 676866 310759 676926 311022
rect 676866 310754 676977 310759
rect 676866 310698 676916 310754
rect 676972 310698 676977 310754
rect 676866 310696 676977 310698
rect 676911 310693 676977 310696
rect 677250 310019 677310 310134
rect 677199 310014 677310 310019
rect 677199 309958 677204 310014
rect 677260 309958 677310 310014
rect 677199 309956 677310 309958
rect 677199 309953 677265 309956
rect 674511 309128 674577 309131
rect 674754 309128 674814 309394
rect 674511 309126 674814 309128
rect 674511 309070 674516 309126
rect 674572 309070 674814 309126
rect 674511 309068 674814 309070
rect 674511 309065 674577 309068
rect 675138 308391 675198 308506
rect 675087 308386 675198 308391
rect 675087 308330 675092 308386
rect 675148 308330 675198 308386
rect 675087 308328 675198 308330
rect 675087 308325 675153 308328
rect 674946 307503 675006 307766
rect 42255 307500 42321 307503
rect 42255 307498 42366 307500
rect 42255 307442 42260 307498
rect 42316 307442 42366 307498
rect 42255 307437 42366 307442
rect 674946 307498 675057 307503
rect 674946 307442 674996 307498
rect 675052 307442 675057 307498
rect 674946 307440 675057 307442
rect 674991 307437 675057 307440
rect 42306 307322 42366 307437
rect 677058 306763 677118 306878
rect 42255 306760 42321 306763
rect 42255 306758 42366 306760
rect 42255 306702 42260 306758
rect 42316 306702 42366 306758
rect 42255 306697 42366 306702
rect 677007 306758 677118 306763
rect 677007 306702 677012 306758
rect 677068 306702 677118 306758
rect 677007 306700 677118 306702
rect 677007 306697 677073 306700
rect 42306 306434 42366 306697
rect 676866 306023 676926 306212
rect 676815 306018 676926 306023
rect 676815 305962 676820 306018
rect 676876 305962 676926 306018
rect 676815 305960 676926 305962
rect 676815 305957 676881 305960
rect 655215 305872 655281 305875
rect 650208 305870 655281 305872
rect 650208 305814 655220 305870
rect 655276 305814 655281 305870
rect 650208 305812 655281 305814
rect 655215 305809 655281 305812
rect 42831 305724 42897 305727
rect 42336 305722 42897 305724
rect 42336 305666 42836 305722
rect 42892 305666 42897 305722
rect 42336 305664 42897 305666
rect 42831 305661 42897 305664
rect 674415 305428 674481 305431
rect 674415 305426 674784 305428
rect 674415 305370 674420 305426
rect 674476 305370 674784 305426
rect 674415 305368 674784 305370
rect 674415 305365 674481 305368
rect 42306 304244 42366 304806
rect 674223 304614 674289 304617
rect 674223 304612 674784 304614
rect 674223 304556 674228 304612
rect 674284 304556 674784 304612
rect 674223 304554 674784 304556
rect 674223 304551 674289 304554
rect 42306 304184 43518 304244
rect 43215 304096 43281 304099
rect 42336 304094 43281 304096
rect 42336 304038 43220 304094
rect 43276 304038 43281 304094
rect 42336 304036 43281 304038
rect 43215 304033 43281 304036
rect 43215 303948 43281 303951
rect 43458 303948 43518 304184
rect 43215 303946 43518 303948
rect 43215 303890 43220 303946
rect 43276 303890 43518 303946
rect 43215 303888 43518 303890
rect 43215 303885 43281 303888
rect 42106 303738 42112 303802
rect 42176 303738 42182 303802
rect 674127 303800 674193 303803
rect 674127 303798 674784 303800
rect 674127 303742 674132 303798
rect 674188 303742 674784 303798
rect 674127 303740 674784 303742
rect 42114 303326 42174 303738
rect 674127 303737 674193 303740
rect 42298 302998 42304 303062
rect 42368 302998 42374 303062
rect 42306 302542 42366 302998
rect 40800 302512 42366 302542
rect 40770 302482 42336 302512
rect 40770 302322 40830 302482
rect 679746 302471 679806 302956
rect 679746 302466 679857 302471
rect 679746 302410 679796 302466
rect 679852 302410 679857 302466
rect 679746 302408 679857 302410
rect 679791 302405 679857 302408
rect 40762 302258 40768 302322
rect 40832 302258 40838 302322
rect 679791 301728 679857 301731
rect 679746 301726 679857 301728
rect 40962 301138 41022 301698
rect 679746 301670 679796 301726
rect 679852 301670 679857 301726
rect 679746 301665 679857 301670
rect 679746 301402 679806 301665
rect 40954 301074 40960 301138
rect 41024 301074 41030 301138
rect 41922 300399 41982 300884
rect 41922 300394 42033 300399
rect 41922 300338 41972 300394
rect 42028 300338 42033 300394
rect 41922 300336 42033 300338
rect 41967 300333 42033 300336
rect 41154 299658 41214 300070
rect 41146 299594 41152 299658
rect 41216 299594 41222 299658
rect 675706 299446 675712 299510
rect 675776 299508 675782 299510
rect 677007 299508 677073 299511
rect 675776 299506 677073 299508
rect 675776 299450 677012 299506
rect 677068 299450 677073 299506
rect 675776 299448 677073 299450
rect 675776 299446 675782 299448
rect 677007 299445 677073 299448
rect 676666 299298 676672 299362
rect 676736 299360 676742 299362
rect 677199 299360 677265 299363
rect 676736 299358 677265 299360
rect 676736 299302 677204 299358
rect 677260 299302 677265 299358
rect 676736 299300 677265 299302
rect 676736 299298 676742 299300
rect 677199 299297 677265 299300
rect 40578 298770 40638 299256
rect 40570 298706 40576 298770
rect 40640 298706 40646 298770
rect 40386 298030 40446 298590
rect 40378 297966 40384 298030
rect 40448 297966 40454 298030
rect 59535 298028 59601 298031
rect 59535 298026 64416 298028
rect 59535 297970 59540 298026
rect 59596 297970 64416 298026
rect 59535 297968 64416 297970
rect 59535 297965 59601 297968
rect 40002 297291 40062 297776
rect 39951 297286 40062 297291
rect 39951 297230 39956 297286
rect 40012 297230 40062 297286
rect 39951 297228 40062 297230
rect 39951 297225 40017 297228
rect 41346 296698 41406 296962
rect 40570 296634 40576 296698
rect 40640 296696 40646 296698
rect 40640 296636 41214 296696
rect 40640 296634 40646 296636
rect 41154 296548 41214 296636
rect 41338 296634 41344 296698
rect 41408 296634 41414 296698
rect 41530 296634 41536 296698
rect 41600 296634 41606 296698
rect 41538 296548 41598 296634
rect 41154 296488 41598 296548
rect 40578 295514 40638 296074
rect 40570 295450 40576 295514
rect 40640 295450 40646 295514
rect 42114 294775 42174 295334
rect 42114 294770 42225 294775
rect 42114 294714 42164 294770
rect 42220 294714 42225 294770
rect 42114 294712 42225 294714
rect 42159 294709 42225 294712
rect 37314 294035 37374 294446
rect 655407 294180 655473 294183
rect 650208 294178 655473 294180
rect 650208 294122 655412 294178
rect 655468 294122 655473 294178
rect 650208 294120 655473 294122
rect 655407 294117 655473 294120
rect 37314 294030 37425 294035
rect 37314 293974 37364 294030
rect 37420 293974 37425 294030
rect 37314 293972 37425 293974
rect 37359 293969 37425 293972
rect 40143 294032 40209 294035
rect 40143 294030 40254 294032
rect 40143 293974 40148 294030
rect 40204 293974 40254 294030
rect 40143 293969 40254 293974
rect 40194 293854 40254 293969
rect 42306 292703 42366 292966
rect 42255 292698 42366 292703
rect 42255 292642 42260 292698
rect 42316 292642 42366 292698
rect 42255 292640 42366 292642
rect 42255 292637 42321 292640
rect 42831 292256 42897 292259
rect 42336 292254 42897 292256
rect 42336 292198 42836 292254
rect 42892 292198 42897 292254
rect 42336 292196 42897 292198
rect 42831 292193 42897 292196
rect 40194 290927 40254 291338
rect 40194 290922 40305 290927
rect 40194 290866 40244 290922
rect 40300 290866 40305 290922
rect 40194 290864 40305 290866
rect 40239 290861 40305 290864
rect 42306 290332 42366 290598
rect 42543 290332 42609 290335
rect 42306 290330 42609 290332
rect 42306 290274 42548 290330
rect 42604 290274 42609 290330
rect 42306 290272 42609 290274
rect 42543 290269 42609 290272
rect 675279 290038 675345 290039
rect 675279 290034 675328 290038
rect 675392 290036 675398 290038
rect 675279 289978 675284 290034
rect 675279 289974 675328 289978
rect 675392 289976 675436 290036
rect 675392 289974 675398 289976
rect 675279 289973 675345 289974
rect 675471 289594 675537 289595
rect 675471 289590 675520 289594
rect 675584 289592 675590 289594
rect 675471 289534 675476 289590
rect 675471 289530 675520 289534
rect 675584 289532 675628 289592
rect 675584 289530 675590 289532
rect 675471 289529 675537 289530
rect 42639 289148 42705 289151
rect 42336 289146 42705 289148
rect 42336 289090 42644 289146
rect 42700 289090 42705 289146
rect 42336 289088 42705 289090
rect 42639 289085 42705 289088
rect 675663 285302 675729 285303
rect 675663 285298 675712 285302
rect 675776 285300 675782 285302
rect 675663 285242 675668 285298
rect 675663 285238 675712 285242
rect 675776 285240 675820 285300
rect 675776 285238 675782 285240
rect 675663 285237 675729 285238
rect 674991 285004 675057 285007
rect 675130 285004 675136 285006
rect 674991 285002 675136 285004
rect 674991 284946 674996 285002
rect 675052 284946 675136 285002
rect 674991 284944 675136 284946
rect 674991 284941 675057 284944
rect 675130 284942 675136 284944
rect 675200 284942 675206 285006
rect 674127 284856 674193 284859
rect 675087 284856 675153 284859
rect 674127 284854 675153 284856
rect 674127 284798 674132 284854
rect 674188 284798 675092 284854
rect 675148 284798 675153 284854
rect 674127 284796 675153 284798
rect 674127 284793 674193 284796
rect 675087 284793 675153 284796
rect 42255 283674 42321 283675
rect 42255 283670 42304 283674
rect 42368 283672 42374 283674
rect 59535 283672 59601 283675
rect 42255 283614 42260 283670
rect 42255 283610 42304 283614
rect 42368 283612 42412 283672
rect 59535 283670 64416 283672
rect 59535 283614 59540 283670
rect 59596 283614 64416 283670
rect 59535 283612 64416 283614
rect 42368 283610 42374 283612
rect 42255 283609 42321 283610
rect 59535 283609 59601 283612
rect 674554 283610 674560 283674
rect 674624 283672 674630 283674
rect 675375 283672 675441 283675
rect 674624 283670 675441 283672
rect 674624 283614 675380 283670
rect 675436 283614 675441 283670
rect 674624 283612 675441 283614
rect 674624 283610 674630 283612
rect 675375 283609 675441 283612
rect 654447 282636 654513 282639
rect 650208 282634 654513 282636
rect 650208 282578 654452 282634
rect 654508 282578 654513 282634
rect 650208 282576 654513 282578
rect 654447 282573 654513 282576
rect 675759 281896 675825 281899
rect 676666 281896 676672 281898
rect 675759 281894 676672 281896
rect 675759 281838 675764 281894
rect 675820 281838 676672 281894
rect 675759 281836 676672 281838
rect 675759 281833 675825 281836
rect 676666 281834 676672 281836
rect 676736 281834 676742 281898
rect 42298 281538 42304 281602
rect 42368 281600 42374 281602
rect 42543 281600 42609 281603
rect 42368 281598 42609 281600
rect 42368 281542 42548 281598
rect 42604 281542 42609 281598
rect 42368 281540 42609 281542
rect 42368 281538 42374 281540
rect 42543 281537 42609 281540
rect 40378 276506 40384 276570
rect 40448 276568 40454 276570
rect 41775 276568 41841 276571
rect 40448 276566 41841 276568
rect 40448 276510 41780 276566
rect 41836 276510 41841 276566
rect 40448 276508 41841 276510
rect 40448 276506 40454 276508
rect 41775 276505 41841 276508
rect 674127 275384 674193 275387
rect 674938 275384 674944 275386
rect 674127 275382 674944 275384
rect 674127 275326 674132 275382
rect 674188 275326 674944 275382
rect 674127 275324 674944 275326
rect 674127 275321 674193 275324
rect 674938 275322 674944 275324
rect 675008 275322 675014 275386
rect 41967 275238 42033 275239
rect 41914 275236 41920 275238
rect 41876 275176 41920 275236
rect 41984 275234 42033 275238
rect 42028 275178 42033 275234
rect 41914 275174 41920 275176
rect 41984 275174 42033 275178
rect 41967 275173 42033 275174
rect 674703 274940 674769 274943
rect 674703 274938 674814 274940
rect 674703 274882 674708 274938
rect 674764 274882 674814 274938
rect 674703 274877 674814 274882
rect 674754 274688 674814 274877
rect 41775 274646 41841 274647
rect 41722 274644 41728 274646
rect 41684 274584 41728 274644
rect 41792 274642 41841 274646
rect 41836 274586 41841 274642
rect 41722 274582 41728 274584
rect 41792 274582 41841 274586
rect 41775 274581 41841 274582
rect 41914 273990 41920 274054
rect 41984 274052 41990 274054
rect 674127 274052 674193 274055
rect 41984 274050 674193 274052
rect 41984 273994 674132 274050
rect 674188 273994 674193 274050
rect 41984 273992 674193 273994
rect 41984 273990 41990 273992
rect 674127 273989 674193 273992
rect 674703 274052 674769 274055
rect 674703 274050 674814 274052
rect 674703 273994 674708 274050
rect 674764 273994 674814 274050
rect 674703 273989 674814 273994
rect 674754 273874 674814 273989
rect 268239 273608 268305 273611
rect 605487 273608 605553 273611
rect 268239 273606 605553 273608
rect 268239 273550 268244 273606
rect 268300 273550 605492 273606
rect 605548 273550 605553 273606
rect 268239 273548 605553 273550
rect 268239 273545 268305 273548
rect 605487 273545 605553 273548
rect 267759 273460 267825 273463
rect 602223 273460 602289 273463
rect 267759 273458 602289 273460
rect 267759 273402 267764 273458
rect 267820 273402 602228 273458
rect 602284 273402 602289 273458
rect 267759 273400 602289 273402
rect 267759 273397 267825 273400
rect 602223 273397 602289 273400
rect 268719 273312 268785 273315
rect 609423 273312 609489 273315
rect 268719 273310 609489 273312
rect 268719 273254 268724 273310
rect 268780 273254 609428 273310
rect 609484 273254 609489 273310
rect 268719 273252 609489 273254
rect 268719 273249 268785 273252
rect 609423 273249 609489 273252
rect 674703 273312 674769 273315
rect 674703 273310 674814 273312
rect 674703 273254 674708 273310
rect 674764 273254 674814 273310
rect 674703 273249 674814 273254
rect 269103 273164 269169 273167
rect 612975 273164 613041 273167
rect 269103 273162 613041 273164
rect 269103 273106 269108 273162
rect 269164 273106 612980 273162
rect 613036 273106 613041 273162
rect 269103 273104 613041 273106
rect 269103 273101 269169 273104
rect 612975 273101 613041 273104
rect 674754 273060 674814 273249
rect 269775 273016 269841 273019
rect 616527 273016 616593 273019
rect 269775 273014 616593 273016
rect 269775 272958 269780 273014
rect 269836 272958 616532 273014
rect 616588 272958 616593 273014
rect 269775 272956 616593 272958
rect 269775 272953 269841 272956
rect 616527 272953 616593 272956
rect 40570 272806 40576 272870
rect 40640 272868 40646 272870
rect 41775 272868 41841 272871
rect 40640 272866 41841 272868
rect 40640 272810 41780 272866
rect 41836 272810 41841 272866
rect 40640 272808 41841 272810
rect 40640 272806 40646 272808
rect 41775 272805 41841 272808
rect 270255 272868 270321 272871
rect 620079 272868 620145 272871
rect 270255 272866 620145 272868
rect 270255 272810 270260 272866
rect 270316 272810 620084 272866
rect 620140 272810 620145 272866
rect 270255 272808 620145 272810
rect 270255 272805 270321 272808
rect 620079 272805 620145 272808
rect 270447 272720 270513 272723
rect 623631 272720 623697 272723
rect 270447 272718 623697 272720
rect 270447 272662 270452 272718
rect 270508 272662 623636 272718
rect 623692 272662 623697 272718
rect 270447 272660 623697 272662
rect 270447 272657 270513 272660
rect 623631 272657 623697 272660
rect 270831 272572 270897 272575
rect 627279 272572 627345 272575
rect 270831 272570 627345 272572
rect 270831 272514 270836 272570
rect 270892 272514 627284 272570
rect 627340 272514 627345 272570
rect 270831 272512 627345 272514
rect 270831 272509 270897 272512
rect 627279 272509 627345 272512
rect 41530 272362 41536 272426
rect 41600 272424 41606 272426
rect 41775 272424 41841 272427
rect 41600 272422 41841 272424
rect 41600 272366 41780 272422
rect 41836 272366 41841 272422
rect 41600 272364 41841 272366
rect 41600 272362 41606 272364
rect 41775 272361 41841 272364
rect 271311 272424 271377 272427
rect 630831 272424 630897 272427
rect 271311 272422 630897 272424
rect 271311 272366 271316 272422
rect 271372 272366 630836 272422
rect 630892 272366 630897 272422
rect 271311 272364 630897 272366
rect 271311 272361 271377 272364
rect 630831 272361 630897 272364
rect 272559 272276 272625 272279
rect 641487 272276 641553 272279
rect 272559 272274 641553 272276
rect 272559 272218 272564 272274
rect 272620 272218 641492 272274
rect 641548 272218 641553 272274
rect 272559 272216 641553 272218
rect 272559 272213 272625 272216
rect 641487 272213 641553 272216
rect 674362 272214 674368 272278
rect 674432 272276 674438 272278
rect 674432 272216 674784 272276
rect 674432 272214 674438 272216
rect 273039 272128 273105 272131
rect 645135 272128 645201 272131
rect 273039 272126 645201 272128
rect 273039 272070 273044 272126
rect 273100 272070 645140 272126
rect 645196 272070 645201 272126
rect 273039 272068 645201 272070
rect 273039 272065 273105 272068
rect 645135 272065 645201 272068
rect 267567 271980 267633 271983
rect 598767 271980 598833 271983
rect 267567 271978 598833 271980
rect 267567 271922 267572 271978
rect 267628 271922 598772 271978
rect 598828 271922 598833 271978
rect 267567 271920 598833 271922
rect 267567 271917 267633 271920
rect 598767 271917 598833 271920
rect 675714 270946 675774 271432
rect 675706 270882 675712 270946
rect 675776 270882 675782 270946
rect 40954 270586 40960 270650
rect 41024 270648 41030 270650
rect 41775 270648 41841 270651
rect 41024 270646 41841 270648
rect 41024 270590 41780 270646
rect 41836 270590 41841 270646
rect 41024 270588 41841 270590
rect 41024 270586 41030 270588
rect 41775 270585 41841 270588
rect 129231 270648 129297 270651
rect 392175 270648 392241 270651
rect 129231 270646 392241 270648
rect 129231 270590 129236 270646
rect 129292 270590 392180 270646
rect 392236 270590 392241 270646
rect 129231 270588 392241 270590
rect 129231 270585 129297 270588
rect 392175 270585 392241 270588
rect 41914 270438 41920 270502
rect 41984 270500 41990 270502
rect 42255 270500 42321 270503
rect 41984 270498 42321 270500
rect 41984 270442 42260 270498
rect 42316 270442 42321 270498
rect 41984 270440 42321 270442
rect 41984 270438 41990 270440
rect 42255 270437 42321 270440
rect 121743 270500 121809 270503
rect 398991 270500 399057 270503
rect 121743 270498 399057 270500
rect 121743 270442 121748 270498
rect 121804 270442 398996 270498
rect 399052 270442 399057 270498
rect 121743 270440 399057 270442
rect 121743 270437 121809 270440
rect 398991 270437 399057 270440
rect 111087 270352 111153 270355
rect 390639 270352 390705 270355
rect 111087 270350 390705 270352
rect 111087 270294 111092 270350
rect 111148 270294 390644 270350
rect 390700 270294 390705 270350
rect 111087 270292 390705 270294
rect 111087 270289 111153 270292
rect 390639 270289 390705 270292
rect 109839 270204 109905 270207
rect 395919 270204 395985 270207
rect 109839 270202 395985 270204
rect 109839 270146 109844 270202
rect 109900 270146 395924 270202
rect 395980 270146 395985 270202
rect 109839 270144 395985 270146
rect 109839 270141 109905 270144
rect 395919 270141 395985 270144
rect 674170 270142 674176 270206
rect 674240 270204 674246 270206
rect 674554 270204 674560 270206
rect 674240 270144 674560 270204
rect 674240 270142 674246 270144
rect 674554 270142 674560 270144
rect 674624 270204 674630 270206
rect 674946 270204 675006 270766
rect 674624 270144 675006 270204
rect 674624 270142 674630 270144
rect 41338 269994 41344 270058
rect 41408 270056 41414 270058
rect 41775 270056 41841 270059
rect 41408 270054 41841 270056
rect 41408 269998 41780 270054
rect 41836 269998 41841 270054
rect 41408 269996 41841 269998
rect 41408 269994 41414 269996
rect 41775 269993 41841 269996
rect 102639 270056 102705 270059
rect 389007 270056 389073 270059
rect 102639 270054 389073 270056
rect 102639 269998 102644 270054
rect 102700 269998 389012 270054
rect 389068 269998 389073 270054
rect 102639 269996 389073 269998
rect 102639 269993 102705 269996
rect 389007 269993 389073 269996
rect 103887 269908 103953 269911
rect 395055 269908 395121 269911
rect 103887 269906 395121 269908
rect 103887 269850 103892 269906
rect 103948 269850 395060 269906
rect 395116 269850 395121 269906
rect 103887 269848 395121 269850
rect 103887 269845 103953 269848
rect 395055 269845 395121 269848
rect 673978 269846 673984 269910
rect 674048 269908 674054 269910
rect 674048 269878 675360 269908
rect 674048 269848 675390 269878
rect 674048 269846 674054 269848
rect 95631 269760 95697 269763
rect 391599 269760 391665 269763
rect 675330 269762 675390 269848
rect 95631 269758 391665 269760
rect 95631 269702 95636 269758
rect 95692 269702 391604 269758
rect 391660 269702 391665 269758
rect 95631 269700 391665 269702
rect 95631 269697 95697 269700
rect 391599 269697 391665 269700
rect 675322 269698 675328 269762
rect 675392 269698 675398 269762
rect 96783 269612 96849 269615
rect 392559 269612 392625 269615
rect 96783 269610 392625 269612
rect 96783 269554 96788 269610
rect 96844 269554 392564 269610
rect 392620 269554 392625 269610
rect 96783 269552 392625 269554
rect 96783 269549 96849 269552
rect 392559 269549 392625 269552
rect 88431 269464 88497 269467
rect 386127 269464 386193 269467
rect 88431 269462 386193 269464
rect 88431 269406 88436 269462
rect 88492 269406 386132 269462
rect 386188 269406 386193 269462
rect 88431 269404 386193 269406
rect 88431 269401 88497 269404
rect 386127 269401 386193 269404
rect 77775 269316 77841 269319
rect 387663 269316 387729 269319
rect 77775 269314 387729 269316
rect 77775 269258 77780 269314
rect 77836 269258 387668 269314
rect 387724 269258 387729 269314
rect 77775 269256 387729 269258
rect 77775 269253 77841 269256
rect 387663 269253 387729 269256
rect 388527 269316 388593 269319
rect 391791 269316 391857 269319
rect 388527 269314 391857 269316
rect 388527 269258 388532 269314
rect 388588 269258 391796 269314
rect 391852 269258 391857 269314
rect 388527 269256 391857 269258
rect 388527 269253 388593 269256
rect 391791 269253 391857 269256
rect 41146 269106 41152 269170
rect 41216 269168 41222 269170
rect 41775 269168 41841 269171
rect 41216 269166 41841 269168
rect 41216 269110 41780 269166
rect 41836 269110 41841 269166
rect 41216 269108 41841 269110
rect 41216 269106 41222 269108
rect 41775 269105 41841 269108
rect 135951 269168 136017 269171
rect 402255 269168 402321 269171
rect 135951 269166 402321 269168
rect 135951 269110 135956 269166
rect 136012 269110 402260 269166
rect 402316 269110 402321 269166
rect 135951 269108 402321 269110
rect 135951 269105 136017 269108
rect 402255 269105 402321 269108
rect 384783 269020 384849 269023
rect 647535 269020 647601 269023
rect 384783 269018 647601 269020
rect 384783 268962 384788 269018
rect 384844 268962 647540 269018
rect 647596 268962 647601 269018
rect 384783 268960 647601 268962
rect 384783 268957 384849 268960
rect 647535 268957 647601 268960
rect 143151 268872 143217 268875
rect 398607 268872 398673 268875
rect 143151 268870 398673 268872
rect 143151 268814 143156 268870
rect 143212 268814 398612 268870
rect 398668 268814 398673 268870
rect 143151 268812 398673 268814
rect 143151 268809 143217 268812
rect 398607 268809 398673 268812
rect 326799 268724 326865 268727
rect 548751 268724 548817 268727
rect 326799 268722 548817 268724
rect 326799 268666 326804 268722
rect 326860 268666 548756 268722
rect 548812 268666 548817 268722
rect 326799 268664 548817 268666
rect 326799 268661 326865 268664
rect 548751 268661 548817 268664
rect 383631 268576 383697 268579
rect 395343 268576 395409 268579
rect 674754 268578 674814 269138
rect 383631 268574 395409 268576
rect 383631 268518 383636 268574
rect 383692 268518 395348 268574
rect 395404 268518 395409 268574
rect 383631 268516 395409 268518
rect 383631 268513 383697 268516
rect 395343 268513 395409 268516
rect 674746 268514 674752 268578
rect 674816 268514 674822 268578
rect 674362 268218 674368 268282
rect 674432 268280 674438 268282
rect 674432 268220 674784 268280
rect 674432 268218 674438 268220
rect 256143 267836 256209 267839
rect 505935 267836 506001 267839
rect 256143 267834 506001 267836
rect 256143 267778 256148 267834
rect 256204 267778 505940 267834
rect 505996 267778 506001 267834
rect 256143 267776 506001 267778
rect 256143 267773 256209 267776
rect 505935 267773 506001 267776
rect 319215 267688 319281 267691
rect 567759 267688 567825 267691
rect 319215 267686 567825 267688
rect 319215 267630 319220 267686
rect 319276 267630 567764 267686
rect 567820 267630 567825 267686
rect 319215 267628 567825 267630
rect 319215 267625 319281 267628
rect 567759 267625 567825 267628
rect 320271 267540 320337 267543
rect 574575 267540 574641 267543
rect 320271 267538 574641 267540
rect 320271 267482 320276 267538
rect 320332 267482 574580 267538
rect 574636 267482 574641 267538
rect 320271 267480 574641 267482
rect 320271 267477 320337 267480
rect 574575 267477 574641 267480
rect 673935 267540 674001 267543
rect 673935 267538 674784 267540
rect 673935 267482 673940 267538
rect 673996 267482 674784 267538
rect 673935 267480 674784 267482
rect 673935 267477 674001 267480
rect 256911 267392 256977 267395
rect 512751 267392 512817 267395
rect 256911 267390 512817 267392
rect 256911 267334 256916 267390
rect 256972 267334 512756 267390
rect 512812 267334 512817 267390
rect 256911 267332 512817 267334
rect 256911 267329 256977 267332
rect 512751 267329 512817 267332
rect 257295 267244 257361 267247
rect 516591 267244 516657 267247
rect 257295 267242 516657 267244
rect 257295 267186 257300 267242
rect 257356 267186 516596 267242
rect 516652 267186 516657 267242
rect 257295 267184 516657 267186
rect 257295 267181 257361 267184
rect 516591 267181 516657 267184
rect 257775 267096 257841 267099
rect 520143 267096 520209 267099
rect 257775 267094 520209 267096
rect 257775 267038 257780 267094
rect 257836 267038 520148 267094
rect 520204 267038 520209 267094
rect 257775 267036 520209 267038
rect 257775 267033 257841 267036
rect 520143 267033 520209 267036
rect 252015 266948 252081 266951
rect 256527 266948 256593 266951
rect 252015 266946 256593 266948
rect 252015 266890 252020 266946
rect 252076 266890 256532 266946
rect 256588 266890 256593 266946
rect 252015 266888 256593 266890
rect 252015 266885 252081 266888
rect 256527 266885 256593 266888
rect 258447 266948 258513 266951
rect 523791 266948 523857 266951
rect 258447 266946 523857 266948
rect 258447 266890 258452 266946
rect 258508 266890 523796 266946
rect 523852 266890 523857 266946
rect 258447 266888 523857 266890
rect 258447 266885 258513 266888
rect 523791 266885 523857 266888
rect 258927 266800 258993 266803
rect 527343 266800 527409 266803
rect 258927 266798 527409 266800
rect 258927 266742 258932 266798
rect 258988 266742 527348 266798
rect 527404 266742 527409 266798
rect 258927 266740 527409 266742
rect 258927 266737 258993 266740
rect 527343 266737 527409 266740
rect 259023 266652 259089 266655
rect 530895 266652 530961 266655
rect 259023 266650 530961 266652
rect 259023 266594 259028 266650
rect 259084 266594 530900 266650
rect 530956 266594 530961 266650
rect 259023 266592 530961 266594
rect 259023 266589 259089 266592
rect 530895 266589 530961 266592
rect 678210 266507 678270 266622
rect 259503 266504 259569 266507
rect 534447 266504 534513 266507
rect 259503 266502 534513 266504
rect 259503 266446 259508 266502
rect 259564 266446 534452 266502
rect 534508 266446 534513 266502
rect 259503 266444 534513 266446
rect 678210 266502 678321 266507
rect 678210 266446 678260 266502
rect 678316 266446 678321 266502
rect 678210 266444 678321 266446
rect 259503 266441 259569 266444
rect 534447 266441 534513 266444
rect 678255 266441 678321 266444
rect 259983 266356 260049 266359
rect 537999 266356 538065 266359
rect 259983 266354 538065 266356
rect 259983 266298 259988 266354
rect 260044 266298 538004 266354
rect 538060 266298 538065 266354
rect 259983 266296 538065 266298
rect 259983 266293 260049 266296
rect 537999 266293 538065 266296
rect 256719 266208 256785 266211
rect 509487 266208 509553 266211
rect 256719 266206 509553 266208
rect 256719 266150 256724 266206
rect 256780 266150 509492 266206
rect 509548 266150 509553 266206
rect 256719 266148 509553 266150
rect 256719 266145 256785 266148
rect 509487 266145 509553 266148
rect 255663 266060 255729 266063
rect 502287 266060 502353 266063
rect 255663 266058 502353 266060
rect 255663 266002 255668 266058
rect 255724 266002 502292 266058
rect 502348 266002 502353 266058
rect 255663 266000 502353 266002
rect 255663 265997 255729 266000
rect 502287 265997 502353 266000
rect 319599 265912 319665 265915
rect 321903 265912 321969 265915
rect 319599 265910 321969 265912
rect 319599 265854 319604 265910
rect 319660 265854 321908 265910
rect 321964 265854 321969 265910
rect 319599 265852 321969 265854
rect 319599 265849 319665 265852
rect 321903 265849 321969 265852
rect 678210 265767 678270 266030
rect 678159 265762 678270 265767
rect 678159 265706 678164 265762
rect 678220 265706 678270 265762
rect 678159 265704 678270 265706
rect 678159 265701 678225 265704
rect 380079 265320 380145 265323
rect 382383 265320 382449 265323
rect 380079 265318 382449 265320
rect 380079 265262 380084 265318
rect 380140 265262 382388 265318
rect 382444 265262 382449 265318
rect 380079 265260 382449 265262
rect 380079 265257 380145 265260
rect 382383 265257 382449 265260
rect 678402 265027 678462 265142
rect 678351 265022 678462 265027
rect 678351 264966 678356 265022
rect 678412 264966 678462 265022
rect 678351 264964 678462 264966
rect 678351 264961 678417 264964
rect 118095 264876 118161 264879
rect 397839 264876 397905 264879
rect 118095 264874 397905 264876
rect 118095 264818 118100 264874
rect 118156 264818 397844 264874
rect 397900 264818 397905 264874
rect 118095 264816 397905 264818
rect 118095 264813 118161 264816
rect 397839 264813 397905 264816
rect 106287 264728 106353 264731
rect 394767 264728 394833 264731
rect 106287 264726 394833 264728
rect 106287 264670 106292 264726
rect 106348 264670 394772 264726
rect 394828 264670 394833 264726
rect 106287 264668 394833 264670
rect 106287 264665 106353 264668
rect 394767 264665 394833 264668
rect 99183 264580 99249 264583
rect 393039 264580 393105 264583
rect 99183 264578 393105 264580
rect 99183 264522 99188 264578
rect 99244 264522 393044 264578
rect 393100 264522 393105 264578
rect 99183 264520 393105 264522
rect 99183 264517 99249 264520
rect 393039 264517 393105 264520
rect 100239 264432 100305 264435
rect 393711 264432 393777 264435
rect 100239 264430 393777 264432
rect 100239 264374 100244 264430
rect 100300 264374 393716 264430
rect 393772 264374 393777 264430
rect 100239 264372 393777 264374
rect 100239 264369 100305 264372
rect 393711 264369 393777 264372
rect 42255 264284 42321 264287
rect 93231 264284 93297 264287
rect 391983 264284 392049 264287
rect 42255 264282 42366 264284
rect 42255 264226 42260 264282
rect 42316 264226 42366 264282
rect 42255 264221 42366 264226
rect 93231 264282 392049 264284
rect 93231 264226 93236 264282
rect 93292 264226 391988 264282
rect 392044 264226 392049 264282
rect 93231 264224 392049 264226
rect 93231 264221 93297 264224
rect 391983 264221 392049 264224
rect 42306 264106 42366 264221
rect 83631 264136 83697 264139
rect 389391 264136 389457 264139
rect 83631 264134 389457 264136
rect 83631 264078 83636 264134
rect 83692 264078 389396 264134
rect 389452 264078 389457 264134
rect 83631 264076 389457 264078
rect 83631 264073 83697 264076
rect 389391 264073 389457 264076
rect 392175 264136 392241 264139
rect 400719 264136 400785 264139
rect 392175 264134 400785 264136
rect 392175 264078 392180 264134
rect 392236 264078 400724 264134
rect 400780 264078 400785 264134
rect 392175 264076 400785 264078
rect 392175 264073 392241 264076
rect 400719 264073 400785 264076
rect 674607 264136 674673 264139
rect 674754 264136 674814 264402
rect 674607 264134 674814 264136
rect 674607 264078 674612 264134
rect 674668 264078 674814 264134
rect 674607 264076 674814 264078
rect 674607 264073 674673 264076
rect 86031 263988 86097 263991
rect 389775 263988 389841 263991
rect 86031 263986 389841 263988
rect 86031 263930 86036 263986
rect 86092 263930 389780 263986
rect 389836 263930 389841 263986
rect 86031 263928 389841 263930
rect 86031 263925 86097 263928
rect 389775 263925 389841 263928
rect 82863 263840 82929 263843
rect 388815 263840 388881 263843
rect 82863 263838 388881 263840
rect 82863 263782 82868 263838
rect 82924 263782 388820 263838
rect 388876 263782 388881 263838
rect 82863 263780 388881 263782
rect 82863 263777 82929 263780
rect 388815 263777 388881 263780
rect 42255 263544 42321 263547
rect 216591 263544 216657 263547
rect 648687 263544 648753 263547
rect 42255 263542 42366 263544
rect 42255 263486 42260 263542
rect 42316 263486 42366 263542
rect 42255 263481 42366 263486
rect 216591 263542 648753 263544
rect 216591 263486 216596 263542
rect 216652 263486 648692 263542
rect 648748 263486 648753 263542
rect 216591 263484 648753 263486
rect 216591 263481 216657 263484
rect 648687 263481 648753 263484
rect 674319 263544 674385 263547
rect 674319 263542 674784 263544
rect 674319 263486 674324 263542
rect 674380 263486 674784 263542
rect 674319 263484 674784 263486
rect 674319 263481 674385 263484
rect 42306 263218 42366 263481
rect 125295 263396 125361 263399
rect 399567 263396 399633 263399
rect 125295 263394 399633 263396
rect 125295 263338 125300 263394
rect 125356 263338 399572 263394
rect 399628 263338 399633 263394
rect 125295 263336 399633 263338
rect 125295 263333 125361 263336
rect 399567 263333 399633 263336
rect 139215 263248 139281 263251
rect 403311 263248 403377 263251
rect 139215 263246 403377 263248
rect 139215 263190 139220 263246
rect 139276 263190 403316 263246
rect 403372 263190 403377 263246
rect 139215 263188 403377 263190
rect 139215 263185 139281 263188
rect 403311 263185 403377 263188
rect 279279 263100 279345 263103
rect 401103 263100 401169 263103
rect 279279 263098 401169 263100
rect 279279 263042 279284 263098
rect 279340 263042 401108 263098
rect 401164 263042 401169 263098
rect 279279 263040 401169 263042
rect 279279 263037 279345 263040
rect 401103 263037 401169 263040
rect 367983 262952 368049 262955
rect 386511 262952 386577 262955
rect 367983 262950 386577 262952
rect 367983 262894 367988 262950
rect 368044 262894 386516 262950
rect 386572 262894 386577 262950
rect 367983 262892 386577 262894
rect 367983 262889 368049 262892
rect 386511 262889 386577 262892
rect 70575 262804 70641 262807
rect 385455 262804 385521 262807
rect 70575 262802 385521 262804
rect 70575 262746 70580 262802
rect 70636 262746 385460 262802
rect 385516 262746 385521 262802
rect 70575 262744 385521 262746
rect 70575 262741 70641 262744
rect 385455 262741 385521 262744
rect 674415 262804 674481 262807
rect 674415 262802 674784 262804
rect 674415 262746 674420 262802
rect 674476 262746 674784 262802
rect 674415 262744 674784 262746
rect 674415 262741 674481 262744
rect 42255 262656 42321 262659
rect 42255 262654 42366 262656
rect 42255 262598 42260 262654
rect 42316 262598 42366 262654
rect 42255 262593 42366 262598
rect 42306 262478 42366 262593
rect 394479 262360 394545 262363
rect 397071 262360 397137 262363
rect 394479 262358 397137 262360
rect 394479 262302 394484 262358
rect 394540 262302 397076 262358
rect 397132 262302 397137 262358
rect 394479 262300 397137 262302
rect 394479 262297 394545 262300
rect 397071 262297 397137 262300
rect 382575 262212 382641 262215
rect 386703 262212 386769 262215
rect 382575 262210 386769 262212
rect 382575 262154 382580 262210
rect 382636 262154 386708 262210
rect 386764 262154 386769 262210
rect 382575 262152 386769 262154
rect 382575 262149 382641 262152
rect 386703 262149 386769 262152
rect 263439 262064 263505 262067
rect 566511 262064 566577 262067
rect 263439 262062 566577 262064
rect 263439 262006 263444 262062
rect 263500 262006 566516 262062
rect 566572 262006 566577 262062
rect 263439 262004 566577 262006
rect 263439 262001 263505 262004
rect 566511 262001 566577 262004
rect 326895 261916 326961 261919
rect 628431 261916 628497 261919
rect 326895 261914 628497 261916
rect 326895 261858 326900 261914
rect 326956 261858 628436 261914
rect 628492 261858 628497 261914
rect 326895 261856 628497 261858
rect 326895 261853 326961 261856
rect 628431 261853 628497 261856
rect 676866 261771 676926 261886
rect 263919 261768 263985 261771
rect 570159 261768 570225 261771
rect 263919 261766 570225 261768
rect 263919 261710 263924 261766
rect 263980 261710 570164 261766
rect 570220 261710 570225 261766
rect 263919 261708 570225 261710
rect 676866 261766 676977 261771
rect 676866 261710 676916 261766
rect 676972 261710 676977 261766
rect 676866 261708 676977 261710
rect 263919 261705 263985 261708
rect 570159 261705 570225 261708
rect 676911 261705 676977 261708
rect 43407 261620 43473 261623
rect 42336 261618 43473 261620
rect 42336 261562 43412 261618
rect 43468 261562 43473 261618
rect 42336 261560 43473 261562
rect 43407 261557 43473 261560
rect 327471 261620 327537 261623
rect 635535 261620 635601 261623
rect 327471 261618 635601 261620
rect 327471 261562 327476 261618
rect 327532 261562 635540 261618
rect 635596 261562 635601 261618
rect 327471 261560 635601 261562
rect 327471 261557 327537 261560
rect 635535 261557 635601 261560
rect 264303 261472 264369 261475
rect 573711 261472 573777 261475
rect 264303 261470 573777 261472
rect 264303 261414 264308 261470
rect 264364 261414 573716 261470
rect 573772 261414 573777 261470
rect 264303 261412 573777 261414
rect 264303 261409 264369 261412
rect 573711 261409 573777 261412
rect 264879 261324 264945 261327
rect 577263 261324 577329 261327
rect 264879 261322 577329 261324
rect 264879 261266 264884 261322
rect 264940 261266 577268 261322
rect 577324 261266 577329 261322
rect 264879 261264 577329 261266
rect 264879 261261 264945 261264
rect 577263 261261 577329 261264
rect 265455 261176 265521 261179
rect 580911 261176 580977 261179
rect 265455 261174 580977 261176
rect 265455 261118 265460 261174
rect 265516 261118 580916 261174
rect 580972 261118 580977 261174
rect 265455 261116 580977 261118
rect 265455 261113 265521 261116
rect 580911 261113 580977 261116
rect 676866 261031 676926 261220
rect 265839 261028 265905 261031
rect 584367 261028 584433 261031
rect 265839 261026 584433 261028
rect 265839 260970 265844 261026
rect 265900 260970 584372 261026
rect 584428 260970 584433 261026
rect 265839 260968 584433 260970
rect 265839 260965 265905 260968
rect 584367 260965 584433 260968
rect 676815 261026 676926 261031
rect 676815 260970 676820 261026
rect 676876 260970 676926 261026
rect 676815 260968 676926 260970
rect 676815 260965 676881 260968
rect 43215 260880 43281 260883
rect 42336 260878 43281 260880
rect 42336 260822 43220 260878
rect 43276 260822 43281 260878
rect 42336 260820 43281 260822
rect 43215 260817 43281 260820
rect 266031 260880 266097 260883
rect 588015 260880 588081 260883
rect 266031 260878 588081 260880
rect 266031 260822 266036 260878
rect 266092 260822 588020 260878
rect 588076 260822 588081 260878
rect 266031 260820 588081 260822
rect 266031 260817 266097 260820
rect 588015 260817 588081 260820
rect 271983 260732 272049 260735
rect 634383 260732 634449 260735
rect 271983 260730 634449 260732
rect 271983 260674 271988 260730
rect 272044 260674 634388 260730
rect 634444 260674 634449 260730
rect 271983 260672 634449 260674
rect 271983 260669 272049 260672
rect 634383 260669 634449 260672
rect 272367 260584 272433 260587
rect 637935 260584 638001 260587
rect 272367 260582 638001 260584
rect 272367 260526 272372 260582
rect 272428 260526 637940 260582
rect 637996 260526 638001 260582
rect 272367 260524 638001 260526
rect 272367 260521 272433 260524
rect 637935 260521 638001 260524
rect 42106 260374 42112 260438
rect 42176 260374 42182 260438
rect 263247 260436 263313 260439
rect 563055 260436 563121 260439
rect 263247 260434 563121 260436
rect 263247 260378 263252 260434
rect 263308 260378 563060 260434
rect 563116 260378 563121 260434
rect 263247 260376 563121 260378
rect 42114 260140 42174 260374
rect 263247 260373 263313 260376
rect 563055 260373 563121 260376
rect 262767 260288 262833 260291
rect 559119 260288 559185 260291
rect 262767 260286 559185 260288
rect 262767 260230 262772 260286
rect 262828 260230 559124 260286
rect 559180 260230 559185 260286
rect 262767 260228 559185 260230
rect 262767 260225 262833 260228
rect 559119 260225 559185 260228
rect 41760 260110 42174 260140
rect 41730 260080 42144 260110
rect 41730 259551 41790 260080
rect 674754 259847 674814 260406
rect 674703 259842 674814 259847
rect 674703 259786 674708 259842
rect 674764 259786 674814 259842
rect 674703 259784 674814 259786
rect 674703 259781 674769 259784
rect 40762 259486 40768 259550
rect 40832 259486 40838 259550
rect 41730 259546 41841 259551
rect 41730 259490 41780 259546
rect 41836 259490 41841 259546
rect 41730 259488 41841 259490
rect 40770 259400 40830 259486
rect 41775 259485 41841 259488
rect 675138 259403 675198 259592
rect 43023 259400 43089 259403
rect 40770 259398 43089 259400
rect 40770 259370 43028 259398
rect 40800 259342 43028 259370
rect 43084 259342 43089 259398
rect 40800 259340 43089 259342
rect 43023 259337 43089 259340
rect 675087 259398 675198 259403
rect 675087 259342 675092 259398
rect 675148 259342 675198 259398
rect 675087 259340 675198 259342
rect 675087 259337 675153 259340
rect 674127 258808 674193 258811
rect 674127 258806 674784 258808
rect 674127 258750 674132 258806
rect 674188 258750 674784 258806
rect 674127 258748 674784 258750
rect 674127 258745 674193 258748
rect 40386 257922 40446 258482
rect 40378 257858 40384 257922
rect 40448 257858 40454 257922
rect 41922 257183 41982 257742
rect 679746 257479 679806 257964
rect 679746 257474 679857 257479
rect 679746 257418 679796 257474
rect 679852 257418 679857 257474
rect 679746 257416 679857 257418
rect 679791 257413 679857 257416
rect 41922 257178 42033 257183
rect 41922 257122 41972 257178
rect 42028 257122 42033 257178
rect 41922 257120 42033 257122
rect 41967 257117 42033 257120
rect 679791 256884 679857 256887
rect 679746 256882 679857 256884
rect 40578 256442 40638 256854
rect 679746 256826 679796 256882
rect 679852 256826 679857 256882
rect 679746 256821 679857 256826
rect 40570 256378 40576 256442
rect 40640 256378 40646 256442
rect 210159 256440 210225 256443
rect 215490 256440 215550 256484
rect 210159 256438 215550 256440
rect 210159 256382 210164 256438
rect 210220 256382 215550 256438
rect 679746 256410 679806 256821
rect 210159 256380 215550 256382
rect 210159 256377 210225 256380
rect 675130 256230 675136 256294
rect 675200 256292 675206 256294
rect 676282 256292 676288 256294
rect 675200 256232 676288 256292
rect 675200 256230 675206 256232
rect 676282 256230 676288 256232
rect 676352 256230 676358 256294
rect 40962 255702 41022 256114
rect 40954 255638 40960 255702
rect 41024 255638 41030 255702
rect 41346 254814 41406 255374
rect 41338 254750 41344 254814
rect 41408 254750 41414 254814
rect 40194 254075 40254 254560
rect 40194 254070 40305 254075
rect 40194 254014 40244 254070
rect 40300 254014 40305 254070
rect 40194 254012 40305 254014
rect 40239 254009 40305 254012
rect 40770 253482 40830 253746
rect 676090 253566 676096 253630
rect 676160 253628 676166 253630
rect 678351 253628 678417 253631
rect 676160 253626 678417 253628
rect 676160 253570 678356 253626
rect 678412 253570 678417 253626
rect 676160 253568 678417 253570
rect 676160 253566 676166 253568
rect 678351 253565 678417 253568
rect 40762 253418 40768 253482
rect 40832 253418 40838 253482
rect 675898 253418 675904 253482
rect 675968 253480 675974 253482
rect 678159 253480 678225 253483
rect 675968 253478 678225 253480
rect 675968 253422 678164 253478
rect 678220 253422 678225 253478
rect 675968 253420 678225 253422
rect 675968 253418 675974 253420
rect 678159 253417 678225 253420
rect 41154 252446 41214 252932
rect 41146 252382 41152 252446
rect 41216 252382 41222 252446
rect 215490 252151 215550 252784
rect 215490 252146 215601 252151
rect 42114 251559 42174 252118
rect 215490 252090 215540 252146
rect 215596 252090 215601 252146
rect 215490 252088 215601 252090
rect 215535 252085 215601 252088
rect 42063 251554 42174 251559
rect 42063 251498 42068 251554
rect 42124 251498 42174 251554
rect 42063 251496 42174 251498
rect 42063 251493 42129 251496
rect 37314 250819 37374 251304
rect 37314 250814 37425 250819
rect 40047 250816 40113 250819
rect 37314 250758 37364 250814
rect 37420 250758 37425 250814
rect 37314 250756 37425 250758
rect 37359 250753 37425 250756
rect 40002 250814 40113 250816
rect 40002 250758 40052 250814
rect 40108 250758 40113 250814
rect 40002 250753 40113 250758
rect 40002 250638 40062 250753
rect 674746 250458 674752 250522
rect 674816 250520 674822 250522
rect 675279 250520 675345 250523
rect 674816 250518 675345 250520
rect 674816 250462 675284 250518
rect 675340 250462 675345 250518
rect 674816 250460 675345 250462
rect 674816 250458 674822 250460
rect 675279 250457 675345 250460
rect 37314 249191 37374 249750
rect 37263 249186 37374 249191
rect 37263 249130 37268 249186
rect 37324 249130 37374 249186
rect 37263 249128 37374 249130
rect 37263 249125 37329 249128
rect 42306 248451 42366 249010
rect 215490 248596 215550 249158
rect 215631 248596 215697 248599
rect 215490 248594 215697 248596
rect 215490 248538 215636 248594
rect 215692 248538 215697 248594
rect 215490 248536 215697 248538
rect 215631 248533 215697 248536
rect 42255 248446 42366 248451
rect 42255 248390 42260 248446
rect 42316 248390 42366 248446
rect 42255 248388 42366 248390
rect 42255 248385 42321 248388
rect 40194 248007 40254 248122
rect 40143 248002 40254 248007
rect 40143 247946 40148 248002
rect 40204 247946 40254 248002
rect 40143 247944 40254 247946
rect 40143 247941 40209 247944
rect 40570 247794 40576 247858
rect 40640 247794 40646 247858
rect 40578 247708 40638 247794
rect 41530 247708 41536 247710
rect 40578 247648 41536 247708
rect 41530 247646 41536 247648
rect 41600 247646 41606 247710
rect 42306 246820 42366 247382
rect 42306 246760 42750 246820
rect 42690 246376 42750 246760
rect 42306 246316 42750 246376
rect 65199 246376 65265 246379
rect 210682 246376 210688 246378
rect 65199 246374 210688 246376
rect 65199 246318 65204 246374
rect 65260 246318 210688 246374
rect 65199 246316 210688 246318
rect 42306 245491 42366 246316
rect 65199 246313 65265 246316
rect 210682 246314 210688 246316
rect 210752 246314 210758 246378
rect 65007 246228 65073 246231
rect 210298 246228 210304 246230
rect 65007 246226 210304 246228
rect 65007 246170 65012 246226
rect 65068 246170 210304 246226
rect 65007 246168 210304 246170
rect 65007 246165 65073 246168
rect 210298 246166 210304 246168
rect 210368 246166 210374 246230
rect 463599 245636 463665 245639
rect 443586 245634 463665 245636
rect 443586 245578 463604 245634
rect 463660 245578 463665 245634
rect 443586 245576 463665 245578
rect 42306 245486 42417 245491
rect 42306 245430 42356 245486
rect 42412 245430 42417 245486
rect 42306 245428 42417 245430
rect 42351 245425 42417 245428
rect 43119 245340 43185 245343
rect 80655 245340 80721 245343
rect 43119 245338 80721 245340
rect 43119 245282 43124 245338
rect 43180 245282 80660 245338
rect 80716 245282 80721 245338
rect 43119 245280 80721 245282
rect 43119 245277 43185 245280
rect 80655 245277 80721 245280
rect 224463 245340 224529 245343
rect 440559 245340 440625 245343
rect 443586 245340 443646 245576
rect 463599 245573 463665 245576
rect 224463 245338 241854 245340
rect 224463 245282 224468 245338
rect 224524 245282 241854 245338
rect 224463 245280 241854 245282
rect 224463 245277 224529 245280
rect 100719 245192 100785 245195
rect 126543 245192 126609 245195
rect 100719 245190 106494 245192
rect 100719 245134 100724 245190
rect 100780 245134 106494 245190
rect 100719 245132 106494 245134
rect 100719 245129 100785 245132
rect 106434 244896 106494 245132
rect 106626 245190 126609 245192
rect 106626 245134 126548 245190
rect 126604 245134 126609 245190
rect 106626 245132 126609 245134
rect 106626 244896 106686 245132
rect 126543 245129 126609 245132
rect 126735 245192 126801 245195
rect 126735 245190 141054 245192
rect 126735 245134 126740 245190
rect 126796 245134 141054 245190
rect 126735 245132 141054 245134
rect 126735 245129 126801 245132
rect 140994 245044 141054 245132
rect 158415 245044 158481 245047
rect 140994 245042 158481 245044
rect 140994 244986 158420 245042
rect 158476 244986 158481 245042
rect 140994 244984 158481 244986
rect 241794 245044 241854 245280
rect 440559 245338 443646 245340
rect 440559 245282 440564 245338
rect 440620 245282 443646 245338
rect 440559 245280 443646 245282
rect 440559 245277 440625 245280
rect 259215 245192 259281 245195
rect 279279 245192 279345 245195
rect 337018 245192 337024 245194
rect 259215 245190 279345 245192
rect 259215 245134 259220 245190
rect 259276 245134 279284 245190
rect 279340 245134 279345 245190
rect 259215 245132 279345 245134
rect 259215 245129 259281 245132
rect 279279 245129 279345 245132
rect 316674 245132 337024 245192
rect 259215 245044 259281 245047
rect 241794 245042 259281 245044
rect 241794 244986 259220 245042
rect 259276 244986 259281 245042
rect 241794 244984 259281 244986
rect 158415 244981 158481 244984
rect 259215 244981 259281 244984
rect 296655 245044 296721 245047
rect 316674 245044 316734 245132
rect 337018 245130 337024 245132
rect 337088 245130 337094 245194
rect 339855 245192 339921 245195
rect 463599 245192 463665 245195
rect 675759 245192 675825 245195
rect 676282 245192 676288 245194
rect 339855 245190 348606 245192
rect 339855 245134 339860 245190
rect 339916 245134 348606 245190
rect 339855 245132 348606 245134
rect 339855 245129 339921 245132
rect 296655 245042 316734 245044
rect 296655 244986 296660 245042
rect 296716 244986 316734 245042
rect 296655 244984 316734 244986
rect 296655 244981 296721 244984
rect 337018 244982 337024 245046
rect 337088 245044 337094 245046
rect 339759 245044 339825 245047
rect 337088 245042 339825 245044
rect 337088 244986 339764 245042
rect 339820 244986 339825 245042
rect 337088 244984 339825 244986
rect 348546 245044 348606 245132
rect 463599 245190 469374 245192
rect 463599 245134 463604 245190
rect 463660 245134 469374 245190
rect 463599 245132 469374 245134
rect 463599 245129 463665 245132
rect 403023 245044 403089 245047
rect 348546 244984 390078 245044
rect 337088 244982 337094 244984
rect 339759 244981 339825 244984
rect 106434 244836 106686 244896
rect 168495 244896 168561 244899
rect 279279 244896 279345 244899
rect 296655 244896 296721 244899
rect 168495 244894 221886 244896
rect 168495 244838 168500 244894
rect 168556 244838 221886 244894
rect 168495 244836 221886 244838
rect 168495 244833 168561 244836
rect 221826 244748 221886 244836
rect 279279 244894 296721 244896
rect 279279 244838 279284 244894
rect 279340 244838 296660 244894
rect 296716 244838 296721 244894
rect 279279 244836 296721 244838
rect 390018 244896 390078 244984
rect 390402 245042 403089 245044
rect 390402 244986 403028 245042
rect 403084 244986 403089 245042
rect 390402 244984 403089 244986
rect 390402 244896 390462 244984
rect 403023 244981 403089 244984
rect 403215 245044 403281 245047
rect 403215 245042 410430 245044
rect 403215 244986 403220 245042
rect 403276 244986 410430 245042
rect 403215 244984 410430 244986
rect 403215 244981 403281 244984
rect 390018 244836 390462 244896
rect 410370 244896 410430 244984
rect 420495 244896 420561 244899
rect 410370 244894 420561 244896
rect 410370 244838 420500 244894
rect 420556 244838 420561 244894
rect 410370 244836 420561 244838
rect 469314 244896 469374 245132
rect 478146 245132 498174 245192
rect 478146 244896 478206 245132
rect 469314 244836 478206 244896
rect 498114 244896 498174 245132
rect 518466 245132 538494 245192
rect 518466 244896 518526 245132
rect 498114 244836 518526 244896
rect 538434 244896 538494 245132
rect 558786 245132 578814 245192
rect 558786 244896 558846 245132
rect 538434 244836 558846 244896
rect 578754 244896 578814 245132
rect 599106 245132 619134 245192
rect 599106 244896 599166 245132
rect 578754 244836 599166 244896
rect 619074 244896 619134 245132
rect 675759 245190 676288 245192
rect 675759 245134 675764 245190
rect 675820 245134 676288 245190
rect 675759 245132 676288 245134
rect 675759 245129 675825 245132
rect 676282 245130 676288 245132
rect 676352 245130 676358 245194
rect 675087 245044 675153 245047
rect 619266 245042 675153 245044
rect 619266 244986 675092 245042
rect 675148 244986 675153 245042
rect 619266 244984 675153 244986
rect 619266 244896 619326 244984
rect 675087 244981 675153 244984
rect 619074 244836 619326 244896
rect 279279 244833 279345 244836
rect 296655 244833 296721 244836
rect 420495 244833 420561 244836
rect 224463 244748 224529 244751
rect 221826 244746 224529 244748
rect 221826 244690 224468 244746
rect 224524 244690 224529 244746
rect 221826 244688 224529 244690
rect 224463 244685 224529 244688
rect 224655 244748 224721 244751
rect 342543 244748 342609 244751
rect 224655 244746 342609 244748
rect 224655 244690 224660 244746
rect 224716 244690 342548 244746
rect 342604 244690 342609 244746
rect 224655 244688 342609 244690
rect 224655 244685 224721 244688
rect 342543 244685 342609 244688
rect 228111 244600 228177 244603
rect 343983 244600 344049 244603
rect 228111 244598 344049 244600
rect 228111 244542 228116 244598
rect 228172 244542 343988 244598
rect 344044 244542 344049 244598
rect 228111 244540 344049 244542
rect 228111 244537 228177 244540
rect 343983 244537 344049 244540
rect 229647 244452 229713 244455
rect 344751 244452 344817 244455
rect 229647 244450 344817 244452
rect 229647 244394 229652 244450
rect 229708 244394 344756 244450
rect 344812 244394 344817 244450
rect 229647 244392 344817 244394
rect 229647 244389 229713 244392
rect 344751 244389 344817 244392
rect 232911 244304 232977 244307
rect 346191 244304 346257 244307
rect 675183 244306 675249 244307
rect 675130 244304 675136 244306
rect 232911 244302 346257 244304
rect 232911 244246 232916 244302
rect 232972 244246 346196 244302
rect 346252 244246 346257 244302
rect 232911 244244 346257 244246
rect 675092 244244 675136 244304
rect 675200 244302 675249 244306
rect 675244 244246 675249 244302
rect 232911 244241 232977 244244
rect 346191 244241 346257 244244
rect 675130 244242 675136 244244
rect 675200 244242 675249 244246
rect 675183 244241 675249 244242
rect 216015 244156 216081 244159
rect 335151 244156 335217 244159
rect 216015 244154 335217 244156
rect 216015 244098 216020 244154
rect 216076 244098 335156 244154
rect 335212 244098 335217 244154
rect 216015 244096 335217 244098
rect 216015 244093 216081 244096
rect 335151 244093 335217 244096
rect 223599 244008 223665 244011
rect 341775 244008 341841 244011
rect 223599 244006 341841 244008
rect 223599 243950 223604 244006
rect 223660 243950 341780 244006
rect 341836 243950 341841 244006
rect 223599 243948 341841 243950
rect 223599 243945 223665 243948
rect 341775 243945 341841 243948
rect 226383 243860 226449 243863
rect 343023 243860 343089 243863
rect 226383 243858 343089 243860
rect 226383 243802 226388 243858
rect 226444 243802 343028 243858
rect 343084 243802 343089 243858
rect 226383 243800 343089 243802
rect 226383 243797 226449 243800
rect 343023 243797 343089 243800
rect 221583 243712 221649 243715
rect 340815 243712 340881 243715
rect 221583 243710 340881 243712
rect 221583 243654 221588 243710
rect 221644 243654 340820 243710
rect 340876 243654 340881 243710
rect 221583 243652 340881 243654
rect 221583 243649 221649 243652
rect 340815 243649 340881 243652
rect 217647 243564 217713 243567
rect 348399 243564 348465 243567
rect 217647 243562 348465 243564
rect 217647 243506 217652 243562
rect 217708 243506 348404 243562
rect 348460 243506 348465 243562
rect 217647 243504 348465 243506
rect 217647 243501 217713 243504
rect 348399 243501 348465 243504
rect 675759 243564 675825 243567
rect 675898 243564 675904 243566
rect 675759 243562 675904 243564
rect 675759 243506 675764 243562
rect 675820 243506 675904 243562
rect 675759 243504 675904 243506
rect 675759 243501 675825 243504
rect 675898 243502 675904 243504
rect 675968 243502 675974 243566
rect 41722 243354 41728 243418
rect 41792 243416 41798 243418
rect 43119 243416 43185 243419
rect 41792 243414 43185 243416
rect 41792 243358 43124 243414
rect 43180 243358 43185 243414
rect 41792 243356 43185 243358
rect 41792 243354 41798 243356
rect 43119 243353 43185 243356
rect 215535 243416 215601 243419
rect 385071 243416 385137 243419
rect 215535 243414 385137 243416
rect 215535 243358 215540 243414
rect 215596 243358 385076 243414
rect 385132 243358 385137 243414
rect 215535 243356 385137 243358
rect 215535 243353 215601 243356
rect 385071 243353 385137 243356
rect 494511 243416 494577 243419
rect 521295 243416 521361 243419
rect 494511 243414 521361 243416
rect 494511 243358 494516 243414
rect 494572 243358 521300 243414
rect 521356 243358 521361 243414
rect 494511 243356 521361 243358
rect 494511 243353 494577 243356
rect 521295 243353 521361 243356
rect 235983 243268 236049 243271
rect 347439 243268 347505 243271
rect 235983 243266 347505 243268
rect 235983 243210 235988 243266
rect 236044 243210 347444 243266
rect 347500 243210 347505 243266
rect 235983 243208 347505 243210
rect 235983 243205 236049 243208
rect 347439 243205 347505 243208
rect 231183 243120 231249 243123
rect 345231 243120 345297 243123
rect 231183 243118 345297 243120
rect 231183 243062 231188 243118
rect 231244 243062 345236 243118
rect 345292 243062 345297 243118
rect 231183 243060 345297 243062
rect 231183 243057 231249 243060
rect 345231 243057 345297 243060
rect 234351 242972 234417 242975
rect 346959 242972 347025 242975
rect 234351 242970 347025 242972
rect 234351 242914 234356 242970
rect 234412 242914 346964 242970
rect 347020 242914 347025 242970
rect 234351 242912 347025 242914
rect 234351 242909 234417 242912
rect 346959 242909 347025 242912
rect 140802 242084 140862 242276
rect 209967 242232 210033 242235
rect 421839 242232 421905 242235
rect 209967 242230 421905 242232
rect 209967 242174 209972 242230
rect 210028 242174 421844 242230
rect 421900 242174 421905 242230
rect 209967 242172 421905 242174
rect 209967 242169 210033 242172
rect 421839 242169 421905 242172
rect 145402 242084 145408 242086
rect 140802 242024 145408 242084
rect 145402 242022 145408 242024
rect 145472 242022 145478 242086
rect 208335 242084 208401 242087
rect 494511 242084 494577 242087
rect 208335 242082 494577 242084
rect 208335 242026 208340 242082
rect 208396 242026 494516 242082
rect 494572 242026 494577 242082
rect 208335 242024 494577 242026
rect 208335 242021 208401 242024
rect 494511 242021 494577 242024
rect 207279 241936 207345 241939
rect 208719 241936 208785 241939
rect 207279 241934 208785 241936
rect 207279 241878 207284 241934
rect 207340 241878 208724 241934
rect 208780 241878 208785 241934
rect 207279 241876 208785 241878
rect 207279 241873 207345 241876
rect 208719 241873 208785 241876
rect 240591 241936 240657 241939
rect 331215 241936 331281 241939
rect 240591 241934 331281 241936
rect 240591 241878 240596 241934
rect 240652 241878 331220 241934
rect 331276 241878 331281 241934
rect 240591 241876 331281 241878
rect 240591 241873 240657 241876
rect 331215 241873 331281 241876
rect 365679 241936 365745 241939
rect 409839 241936 409905 241939
rect 365679 241934 409905 241936
rect 365679 241878 365684 241934
rect 365740 241878 409844 241934
rect 409900 241878 409905 241934
rect 365679 241876 409905 241878
rect 365679 241873 365745 241876
rect 409839 241873 409905 241876
rect 215055 241788 215121 241791
rect 325455 241788 325521 241791
rect 215055 241786 325521 241788
rect 215055 241730 215060 241786
rect 215116 241730 325460 241786
rect 325516 241730 325521 241786
rect 215055 241728 325521 241730
rect 215055 241725 215121 241728
rect 325455 241725 325521 241728
rect 365583 241788 365649 241791
rect 408975 241788 409041 241791
rect 365583 241786 409041 241788
rect 365583 241730 365588 241786
rect 365644 241730 408980 241786
rect 409036 241730 409041 241786
rect 365583 241728 409041 241730
rect 365583 241725 365649 241728
rect 408975 241725 409041 241728
rect 243375 241640 243441 241643
rect 365391 241640 365457 241643
rect 243375 241638 365457 241640
rect 243375 241582 243380 241638
rect 243436 241582 365396 241638
rect 365452 241582 365457 241638
rect 243375 241580 365457 241582
rect 243375 241577 243441 241580
rect 365391 241577 365457 241580
rect 365775 241640 365841 241643
rect 367599 241640 367665 241643
rect 365775 241638 367665 241640
rect 365775 241582 365780 241638
rect 365836 241582 367604 241638
rect 367660 241582 367665 241638
rect 365775 241580 367665 241582
rect 365775 241577 365841 241580
rect 367599 241577 367665 241580
rect 367791 241640 367857 241643
rect 413103 241640 413169 241643
rect 367791 241638 413169 241640
rect 367791 241582 367796 241638
rect 367852 241582 413108 241638
rect 413164 241582 413169 241638
rect 367791 241580 413169 241582
rect 367791 241577 367857 241580
rect 413103 241577 413169 241580
rect 242799 241492 242865 241495
rect 366063 241492 366129 241495
rect 366447 241492 366513 241495
rect 242799 241490 366129 241492
rect 242799 241434 242804 241490
rect 242860 241434 366068 241490
rect 366124 241434 366129 241490
rect 242799 241432 366129 241434
rect 242799 241429 242865 241432
rect 366063 241429 366129 241432
rect 366210 241490 366513 241492
rect 366210 241434 366452 241490
rect 366508 241434 366513 241490
rect 366210 241432 366513 241434
rect 242415 241344 242481 241347
rect 366210 241344 366270 241432
rect 366447 241429 366513 241432
rect 379215 241492 379281 241495
rect 412623 241492 412689 241495
rect 379215 241490 412689 241492
rect 379215 241434 379220 241490
rect 379276 241434 412628 241490
rect 412684 241434 412689 241490
rect 379215 241432 412689 241434
rect 379215 241429 379281 241432
rect 412623 241429 412689 241432
rect 242415 241342 366270 241344
rect 242415 241286 242420 241342
rect 242476 241286 366270 241342
rect 242415 241284 366270 241286
rect 366447 241344 366513 241347
rect 411567 241344 411633 241347
rect 366447 241342 411633 241344
rect 366447 241286 366452 241342
rect 366508 241286 411572 241342
rect 411628 241286 411633 241342
rect 366447 241284 411633 241286
rect 242415 241281 242481 241284
rect 366447 241281 366513 241284
rect 411567 241281 411633 241284
rect 675087 241344 675153 241347
rect 675514 241344 675520 241346
rect 675087 241342 675520 241344
rect 675087 241286 675092 241342
rect 675148 241286 675520 241342
rect 675087 241284 675520 241286
rect 675087 241281 675153 241284
rect 675514 241282 675520 241284
rect 675584 241282 675590 241346
rect 242319 241196 242385 241199
rect 365775 241196 365841 241199
rect 242319 241194 365841 241196
rect 242319 241138 242324 241194
rect 242380 241138 365780 241194
rect 365836 241138 365841 241194
rect 242319 241136 365841 241138
rect 242319 241133 242385 241136
rect 365775 241133 365841 241136
rect 366063 241196 366129 241199
rect 410511 241196 410577 241199
rect 366063 241194 410577 241196
rect 366063 241138 366068 241194
rect 366124 241138 410516 241194
rect 410572 241138 410577 241194
rect 366063 241136 410577 241138
rect 366063 241133 366129 241136
rect 410511 241133 410577 241136
rect 42063 240754 42129 240755
rect 42063 240752 42112 240754
rect 42020 240750 42112 240752
rect 42020 240694 42068 240750
rect 42020 240692 42112 240694
rect 42063 240690 42112 240692
rect 42176 240690 42182 240754
rect 42351 240752 42417 240755
rect 42490 240752 42496 240754
rect 42351 240750 42496 240752
rect 42351 240694 42356 240750
rect 42412 240694 42496 240750
rect 42351 240692 42496 240694
rect 42063 240689 42129 240690
rect 42351 240689 42417 240692
rect 42490 240690 42496 240692
rect 42560 240690 42566 240754
rect 140802 240604 140862 241092
rect 285423 241048 285489 241051
rect 286671 241048 286737 241051
rect 285423 241046 286737 241048
rect 285423 240990 285428 241046
rect 285484 240990 286676 241046
rect 286732 240990 286737 241046
rect 285423 240988 286737 240990
rect 285423 240985 285489 240988
rect 286671 240985 286737 240988
rect 289839 241048 289905 241051
rect 294447 241048 294513 241051
rect 289839 241046 294513 241048
rect 289839 240990 289844 241046
rect 289900 240990 294452 241046
rect 294508 240990 294513 241046
rect 289839 240988 294513 240990
rect 289839 240985 289905 240988
rect 294447 240985 294513 240988
rect 367407 241048 367473 241051
rect 412527 241048 412593 241051
rect 367407 241046 412593 241048
rect 367407 240990 367412 241046
rect 367468 240990 412532 241046
rect 412588 240990 412593 241046
rect 367407 240988 412593 240990
rect 367407 240985 367473 240988
rect 412527 240985 412593 240988
rect 241551 240900 241617 240903
rect 369135 240900 369201 240903
rect 241551 240898 369201 240900
rect 241551 240842 241556 240898
rect 241612 240842 369140 240898
rect 369196 240842 369201 240898
rect 241551 240840 369201 240842
rect 241551 240837 241617 240840
rect 369135 240837 369201 240840
rect 379311 240900 379377 240903
rect 413775 240900 413841 240903
rect 379311 240898 413841 240900
rect 379311 240842 379316 240898
rect 379372 240842 413780 240898
rect 413836 240842 413841 240898
rect 379311 240840 413841 240842
rect 379311 240837 379377 240840
rect 413775 240837 413841 240840
rect 240975 240752 241041 240755
rect 370191 240752 370257 240755
rect 240975 240750 370257 240752
rect 240975 240694 240980 240750
rect 241036 240694 370196 240750
rect 370252 240694 370257 240750
rect 240975 240692 370257 240694
rect 240975 240689 241041 240692
rect 370191 240689 370257 240692
rect 377103 240752 377169 240755
rect 409359 240752 409425 240755
rect 377103 240750 409425 240752
rect 377103 240694 377108 240750
rect 377164 240694 409364 240750
rect 409420 240694 409425 240750
rect 377103 240692 409425 240694
rect 377103 240689 377169 240692
rect 409359 240689 409425 240692
rect 146031 240604 146097 240607
rect 140802 240602 146097 240604
rect 140802 240546 146036 240602
rect 146092 240546 146097 240602
rect 140802 240544 146097 240546
rect 146031 240541 146097 240544
rect 215823 240604 215889 240607
rect 394767 240604 394833 240607
rect 215823 240602 394833 240604
rect 215823 240546 215828 240602
rect 215884 240546 394772 240602
rect 394828 240546 394833 240602
rect 215823 240544 394833 240546
rect 215823 240541 215889 240544
rect 394767 240541 394833 240544
rect 149583 240456 149649 240459
rect 208911 240456 208977 240459
rect 149583 240454 208977 240456
rect 149583 240398 149588 240454
rect 149644 240398 208916 240454
rect 208972 240398 208977 240454
rect 149583 240396 208977 240398
rect 149583 240393 149649 240396
rect 208911 240393 208977 240396
rect 215919 240456 215985 240459
rect 415311 240456 415377 240459
rect 215919 240454 415377 240456
rect 215919 240398 215924 240454
rect 215980 240398 415316 240454
rect 415372 240398 415377 240454
rect 215919 240396 415377 240398
rect 215919 240393 215985 240396
rect 415311 240393 415377 240396
rect 285711 240308 285777 240311
rect 299151 240308 299217 240311
rect 285711 240306 299217 240308
rect 285711 240250 285716 240306
rect 285772 240250 299156 240306
rect 299212 240250 299217 240306
rect 285711 240248 299217 240250
rect 285711 240245 285777 240248
rect 299151 240245 299217 240248
rect 342831 240308 342897 240311
rect 351375 240308 351441 240311
rect 342831 240306 351441 240308
rect 342831 240250 342836 240306
rect 342892 240250 351380 240306
rect 351436 240250 351441 240306
rect 342831 240248 351441 240250
rect 342831 240245 342897 240248
rect 351375 240245 351441 240248
rect 365199 240308 365265 240311
rect 408111 240308 408177 240311
rect 365199 240306 408177 240308
rect 365199 240250 365204 240306
rect 365260 240250 408116 240306
rect 408172 240250 408177 240306
rect 365199 240248 408177 240250
rect 365199 240245 365265 240248
rect 408111 240245 408177 240248
rect 241839 240160 241905 240163
rect 368463 240160 368529 240163
rect 241839 240158 368529 240160
rect 241839 240102 241844 240158
rect 241900 240102 368468 240158
rect 368524 240102 368529 240158
rect 241839 240100 368529 240102
rect 241839 240097 241905 240100
rect 368463 240097 368529 240100
rect 378447 240160 378513 240163
rect 412047 240160 412113 240163
rect 378447 240158 412113 240160
rect 378447 240102 378452 240158
rect 378508 240102 412052 240158
rect 412108 240102 412113 240158
rect 378447 240100 412113 240102
rect 378447 240097 378513 240100
rect 412047 240097 412113 240100
rect 342735 240012 342801 240015
rect 350607 240012 350673 240015
rect 342735 240010 350673 240012
rect 342735 239954 342740 240010
rect 342796 239954 350612 240010
rect 350668 239954 350673 240010
rect 342735 239952 350673 239954
rect 342735 239949 342801 239952
rect 350607 239949 350673 239952
rect 377487 240012 377553 240015
rect 410319 240012 410385 240015
rect 377487 240010 410385 240012
rect 377487 239954 377492 240010
rect 377548 239954 410324 240010
rect 410380 239954 410385 240010
rect 377487 239952 410385 239954
rect 377487 239949 377553 239952
rect 410319 239949 410385 239952
rect 144015 239864 144081 239867
rect 140832 239862 144081 239864
rect 140832 239806 144020 239862
rect 144076 239806 144081 239862
rect 140832 239804 144081 239806
rect 144015 239801 144081 239804
rect 208719 239864 208785 239867
rect 285423 239864 285489 239867
rect 293295 239864 293361 239867
rect 208719 239862 213054 239864
rect 208719 239806 208724 239862
rect 208780 239806 213054 239862
rect 208719 239804 213054 239806
rect 208719 239801 208785 239804
rect 208911 239716 208977 239719
rect 209871 239716 209937 239719
rect 208911 239714 212862 239716
rect 208911 239658 208916 239714
rect 208972 239658 209876 239714
rect 209932 239658 212862 239714
rect 208911 239656 212862 239658
rect 208911 239653 208977 239656
rect 209871 239653 209937 239656
rect 212802 239420 212862 239656
rect 212994 239568 213054 239804
rect 285423 239862 293361 239864
rect 285423 239806 285428 239862
rect 285484 239806 293300 239862
rect 293356 239806 293361 239862
rect 285423 239804 293361 239806
rect 285423 239801 285489 239804
rect 293295 239801 293361 239804
rect 377007 239864 377073 239867
rect 408303 239864 408369 239867
rect 377007 239862 408369 239864
rect 377007 239806 377012 239862
rect 377068 239806 408308 239862
rect 408364 239806 408369 239862
rect 377007 239804 408369 239806
rect 377007 239801 377073 239804
rect 408303 239801 408369 239804
rect 215439 239716 215505 239719
rect 325455 239716 325521 239719
rect 215439 239714 325521 239716
rect 215439 239658 215444 239714
rect 215500 239658 325460 239714
rect 325516 239658 325521 239714
rect 215439 239656 325521 239658
rect 215439 239653 215505 239656
rect 325455 239653 325521 239656
rect 377871 239716 377937 239719
rect 410895 239716 410961 239719
rect 377871 239714 410961 239716
rect 377871 239658 377876 239714
rect 377932 239658 410900 239714
rect 410956 239658 410961 239714
rect 377871 239656 410961 239658
rect 377871 239653 377937 239656
rect 410895 239653 410961 239656
rect 358863 239568 358929 239571
rect 212994 239566 358929 239568
rect 212994 239510 358868 239566
rect 358924 239510 358929 239566
rect 212994 239508 358929 239510
rect 358863 239505 358929 239508
rect 383055 239568 383121 239571
rect 395247 239568 395313 239571
rect 383055 239566 395313 239568
rect 383055 239510 383060 239566
rect 383116 239510 395252 239566
rect 395308 239510 395313 239566
rect 383055 239508 395313 239510
rect 383055 239505 383121 239508
rect 395247 239505 395313 239508
rect 359439 239420 359505 239423
rect 212802 239418 359505 239420
rect 212802 239362 359444 239418
rect 359500 239362 359505 239418
rect 212802 239360 359505 239362
rect 359439 239357 359505 239360
rect 140655 239272 140721 239275
rect 505551 239272 505617 239275
rect 674607 239274 674673 239275
rect 674554 239272 674560 239274
rect 140655 239270 505617 239272
rect 140655 239214 140660 239270
rect 140716 239214 505556 239270
rect 505612 239214 505617 239270
rect 140655 239212 505617 239214
rect 674516 239212 674560 239272
rect 674624 239270 674673 239274
rect 674668 239214 674673 239270
rect 140655 239209 140721 239212
rect 505551 239209 505617 239212
rect 674554 239210 674560 239212
rect 674624 239210 674673 239214
rect 674607 239209 674673 239210
rect 674991 239272 675057 239275
rect 675322 239272 675328 239274
rect 674991 239270 675328 239272
rect 674991 239214 674996 239270
rect 675052 239214 675328 239270
rect 674991 239212 675328 239214
rect 674991 239209 675057 239212
rect 675322 239210 675328 239212
rect 675392 239210 675398 239274
rect 140751 239124 140817 239127
rect 510351 239124 510417 239127
rect 140751 239122 510417 239124
rect 140751 239066 140756 239122
rect 140812 239066 510356 239122
rect 510412 239066 510417 239122
rect 140751 239064 510417 239066
rect 140751 239061 140817 239064
rect 510351 239061 510417 239064
rect 638415 239124 638481 239127
rect 639279 239124 639345 239127
rect 638415 239122 639345 239124
rect 638415 239066 638420 239122
rect 638476 239066 639284 239122
rect 639340 239066 639345 239122
rect 638415 239064 639345 239066
rect 638415 239061 638481 239064
rect 639279 239061 639345 239064
rect 232047 238976 232113 238979
rect 345615 238976 345681 238979
rect 675183 238978 675249 238979
rect 232047 238974 345681 238976
rect 232047 238918 232052 238974
rect 232108 238918 345620 238974
rect 345676 238918 345681 238974
rect 232047 238916 345681 238918
rect 232047 238913 232113 238916
rect 345615 238913 345681 238916
rect 675130 238914 675136 238978
rect 675200 238976 675249 238978
rect 675200 238974 675292 238976
rect 675244 238918 675292 238974
rect 675200 238916 675292 238918
rect 675200 238914 675249 238916
rect 675183 238913 675249 238914
rect 230223 238828 230289 238831
rect 344847 238828 344913 238831
rect 230223 238826 344913 238828
rect 230223 238770 230228 238826
rect 230284 238770 344852 238826
rect 344908 238770 344913 238826
rect 230223 238768 344913 238770
rect 230223 238765 230289 238768
rect 344847 238765 344913 238768
rect 144111 238680 144177 238683
rect 140832 238678 144177 238680
rect 140832 238622 144116 238678
rect 144172 238622 144177 238678
rect 140832 238620 144177 238622
rect 144111 238617 144177 238620
rect 227439 238680 227505 238683
rect 343407 238680 343473 238683
rect 227439 238678 343473 238680
rect 227439 238622 227444 238678
rect 227500 238622 343412 238678
rect 343468 238622 343473 238678
rect 227439 238620 343473 238622
rect 227439 238617 227505 238620
rect 343407 238617 343473 238620
rect 674362 238618 674368 238682
rect 674432 238680 674438 238682
rect 675471 238680 675537 238683
rect 674432 238678 675537 238680
rect 674432 238622 675476 238678
rect 675532 238622 675537 238678
rect 674432 238620 675537 238622
rect 674432 238618 674438 238620
rect 675471 238617 675537 238620
rect 222735 238532 222801 238535
rect 341199 238532 341265 238535
rect 222735 238530 341265 238532
rect 222735 238474 222740 238530
rect 222796 238474 341204 238530
rect 341260 238474 341265 238530
rect 222735 238472 341265 238474
rect 222735 238469 222801 238472
rect 341199 238469 341265 238472
rect 221007 238384 221073 238387
rect 338991 238384 339057 238387
rect 221007 238382 339057 238384
rect 221007 238326 221012 238382
rect 221068 238326 338996 238382
rect 339052 238326 339057 238382
rect 221007 238324 339057 238326
rect 221007 238321 221073 238324
rect 338991 238321 339057 238324
rect 225807 238236 225873 238239
rect 342735 238236 342801 238239
rect 225807 238234 342801 238236
rect 225807 238178 225812 238234
rect 225868 238178 342740 238234
rect 342796 238178 342801 238234
rect 225807 238176 342801 238178
rect 225807 238173 225873 238176
rect 342735 238173 342801 238176
rect 224175 238088 224241 238091
rect 342159 238088 342225 238091
rect 224175 238086 342225 238088
rect 224175 238030 224180 238086
rect 224236 238030 342164 238086
rect 342220 238030 342225 238086
rect 224175 238028 342225 238030
rect 224175 238025 224241 238028
rect 342159 238025 342225 238028
rect 42447 237942 42513 237943
rect 42447 237938 42496 237942
rect 42560 237940 42566 237942
rect 217071 237940 217137 237943
rect 344367 237940 344433 237943
rect 42447 237882 42452 237938
rect 42447 237878 42496 237882
rect 42560 237880 42604 237940
rect 217071 237938 344433 237940
rect 217071 237882 217076 237938
rect 217132 237882 344372 237938
rect 344428 237882 344433 237938
rect 217071 237880 344433 237882
rect 42560 237878 42566 237880
rect 42447 237877 42513 237878
rect 217071 237877 217137 237880
rect 344367 237877 344433 237880
rect 218799 237792 218865 237795
rect 352239 237792 352305 237795
rect 218799 237790 352305 237792
rect 218799 237734 218804 237790
rect 218860 237734 352244 237790
rect 352300 237734 352305 237790
rect 218799 237732 352305 237734
rect 218799 237729 218865 237732
rect 352239 237729 352305 237732
rect 218991 237644 219057 237647
rect 354447 237644 354513 237647
rect 218991 237642 354513 237644
rect 218991 237586 218996 237642
rect 219052 237586 354452 237642
rect 354508 237586 354513 237642
rect 218991 237584 354513 237586
rect 218991 237581 219057 237584
rect 354447 237581 354513 237584
rect 235119 237496 235185 237499
rect 347055 237496 347121 237499
rect 235119 237494 347121 237496
rect 235119 237438 235124 237494
rect 235180 237438 347060 237494
rect 347116 237438 347121 237494
rect 235119 237436 347121 237438
rect 235119 237433 235185 237436
rect 347055 237433 347121 237436
rect 140802 236904 140862 237392
rect 238191 237348 238257 237351
rect 348783 237348 348849 237351
rect 238191 237346 348849 237348
rect 238191 237290 238196 237346
rect 238252 237290 348788 237346
rect 348844 237290 348849 237346
rect 238191 237288 348849 237290
rect 238191 237285 238257 237288
rect 348783 237285 348849 237288
rect 210298 237138 210304 237202
rect 210368 237200 210374 237202
rect 211503 237200 211569 237203
rect 210368 237198 211569 237200
rect 210368 237142 211508 237198
rect 211564 237142 211569 237198
rect 210368 237140 211569 237142
rect 210368 237138 210374 237140
rect 211503 237137 211569 237140
rect 146223 236904 146289 236907
rect 140802 236902 146289 236904
rect 140802 236846 146228 236902
rect 146284 236846 146289 236902
rect 140802 236844 146289 236846
rect 146223 236841 146289 236844
rect 675759 236904 675825 236907
rect 676090 236904 676096 236906
rect 675759 236902 676096 236904
rect 675759 236846 675764 236902
rect 675820 236846 676096 236902
rect 675759 236844 676096 236846
rect 675759 236841 675825 236844
rect 676090 236842 676096 236844
rect 676160 236842 676166 236906
rect 144015 236312 144081 236315
rect 140802 236310 144081 236312
rect 140802 236254 144020 236310
rect 144076 236254 144081 236310
rect 140802 236252 144081 236254
rect 140802 236210 140862 236252
rect 144015 236249 144081 236252
rect 146415 235128 146481 235131
rect 140832 235126 146481 235128
rect 140832 235070 146420 235126
rect 146476 235070 146481 235126
rect 140832 235068 146481 235070
rect 146415 235065 146481 235068
rect 211450 234622 211456 234686
rect 211520 234684 211526 234686
rect 541455 234684 541521 234687
rect 211520 234682 541521 234684
rect 211520 234626 541460 234682
rect 541516 234626 541521 234682
rect 211520 234624 541521 234626
rect 211520 234622 211526 234624
rect 541455 234621 541521 234624
rect 211887 234092 211953 234095
rect 212794 234092 212800 234094
rect 211887 234090 212800 234092
rect 211887 234034 211892 234090
rect 211948 234034 212800 234090
rect 211887 234032 212800 234034
rect 211887 234029 211953 234032
rect 212794 234030 212800 234032
rect 212864 234030 212870 234094
rect 637498 234030 637504 234094
rect 637568 234092 637574 234094
rect 638031 234092 638097 234095
rect 637568 234090 638097 234092
rect 637568 234034 638036 234090
rect 638092 234034 638097 234090
rect 637568 234032 638097 234034
rect 637568 234030 637574 234032
rect 638031 234029 638097 234032
rect 211066 233882 211072 233946
rect 211136 233944 211142 233946
rect 212271 233944 212337 233947
rect 211136 233942 212337 233944
rect 211136 233886 212276 233942
rect 212332 233886 212337 233942
rect 211136 233884 212337 233886
rect 211136 233882 211142 233884
rect 212271 233881 212337 233884
rect 637647 233946 637713 233947
rect 637647 233942 637696 233946
rect 637760 233944 637766 233946
rect 637647 233886 637652 233942
rect 637647 233882 637696 233886
rect 637760 233884 637804 233944
rect 637760 233882 637766 233884
rect 637647 233881 637713 233882
rect 140802 233648 140862 233840
rect 210490 233734 210496 233798
rect 210560 233796 210566 233798
rect 211503 233796 211569 233799
rect 210560 233794 211569 233796
rect 210560 233738 211508 233794
rect 211564 233738 211569 233794
rect 210560 233736 211569 233738
rect 210560 233734 210566 233736
rect 211503 233733 211569 233736
rect 212410 233734 212416 233798
rect 212480 233796 212486 233798
rect 216687 233796 216753 233799
rect 212480 233794 216753 233796
rect 212480 233738 216692 233794
rect 216748 233738 216753 233794
rect 212480 233736 216753 233738
rect 212480 233734 212486 233736
rect 216687 233733 216753 233736
rect 272367 233796 272433 233799
rect 280335 233796 280401 233799
rect 272367 233794 280401 233796
rect 272367 233738 272372 233794
rect 272428 233738 280340 233794
rect 280396 233738 280401 233794
rect 272367 233736 280401 233738
rect 272367 233733 272433 233736
rect 280335 233733 280401 233736
rect 306543 233796 306609 233799
rect 637167 233798 637233 233799
rect 637114 233796 637120 233798
rect 306543 233794 306750 233796
rect 306543 233738 306548 233794
rect 306604 233738 306750 233794
rect 306543 233736 306750 233738
rect 637076 233736 637120 233796
rect 637184 233794 637233 233798
rect 637228 233738 637233 233794
rect 306543 233733 306609 233736
rect 144015 233648 144081 233651
rect 140802 233646 144081 233648
rect 140802 233590 144020 233646
rect 144076 233590 144081 233646
rect 140802 233588 144081 233590
rect 144015 233585 144081 233588
rect 210682 233586 210688 233650
rect 210752 233648 210758 233650
rect 211311 233648 211377 233651
rect 210752 233646 211377 233648
rect 210752 233590 211316 233646
rect 211372 233590 211377 233646
rect 210752 233588 211377 233590
rect 210752 233586 210758 233588
rect 211311 233585 211377 233588
rect 212026 233586 212032 233650
rect 212096 233648 212102 233650
rect 214191 233648 214257 233651
rect 212096 233646 214257 233648
rect 212096 233590 214196 233646
rect 214252 233590 214257 233646
rect 212096 233588 214257 233590
rect 306690 233648 306750 233736
rect 637114 233734 637120 233736
rect 637184 233734 637233 233738
rect 637306 233734 637312 233798
rect 637376 233796 637382 233798
rect 639279 233796 639345 233799
rect 637376 233794 639345 233796
rect 637376 233738 639284 233794
rect 639340 233738 639345 233794
rect 637376 233736 639345 233738
rect 637376 233734 637382 233736
rect 637167 233733 637233 233734
rect 639279 233733 639345 233736
rect 306927 233648 306993 233651
rect 306690 233646 306993 233648
rect 306690 233590 306932 233646
rect 306988 233590 306993 233646
rect 306690 233588 306993 233590
rect 212096 233586 212102 233588
rect 214191 233585 214257 233588
rect 306927 233585 306993 233588
rect 636730 233586 636736 233650
rect 636800 233648 636806 233650
rect 638127 233648 638193 233651
rect 638511 233648 638577 233651
rect 636800 233646 638193 233648
rect 636800 233590 638132 233646
rect 638188 233590 638193 233646
rect 636800 233588 638193 233590
rect 636800 233586 636806 233588
rect 638127 233585 638193 233588
rect 638274 233646 638577 233648
rect 638274 233590 638516 233646
rect 638572 233590 638577 233646
rect 638274 233588 638577 233590
rect 211314 233500 211374 233585
rect 212218 233500 212224 233502
rect 211314 233440 212224 233500
rect 212218 233438 212224 233440
rect 212288 233438 212294 233502
rect 636922 233438 636928 233502
rect 636992 233500 636998 233502
rect 638274 233500 638334 233588
rect 638511 233585 638577 233588
rect 636992 233440 638334 233500
rect 636992 233438 636998 233440
rect 41338 233290 41344 233354
rect 41408 233352 41414 233354
rect 41775 233352 41841 233355
rect 41408 233350 41841 233352
rect 41408 233294 41780 233350
rect 41836 233294 41841 233350
rect 41408 233292 41841 233294
rect 41408 233290 41414 233292
rect 41775 233289 41841 233292
rect 210298 232994 210304 233058
rect 210368 233056 210374 233058
rect 211450 233056 211456 233058
rect 210368 232996 211456 233056
rect 210368 232994 210374 232996
rect 211450 232994 211456 232996
rect 211520 232994 211526 233058
rect 212410 232846 212416 232910
rect 212480 232908 212486 232910
rect 212986 232908 212992 232910
rect 212480 232848 212992 232908
rect 212480 232846 212486 232848
rect 212986 232846 212992 232848
rect 213056 232846 213062 232910
rect 206799 232760 206865 232763
rect 645711 232760 645777 232763
rect 206799 232758 210528 232760
rect 206799 232702 206804 232758
rect 206860 232702 210528 232758
rect 206799 232700 210528 232702
rect 640224 232758 645777 232760
rect 640224 232702 645716 232758
rect 645772 232702 645777 232758
rect 640224 232700 645777 232702
rect 206799 232697 206865 232700
rect 645711 232697 645777 232700
rect 140802 232168 140862 232656
rect 645519 232316 645585 232319
rect 640194 232314 645585 232316
rect 640194 232258 645524 232314
rect 645580 232258 645585 232314
rect 640194 232256 645585 232258
rect 640194 232212 640254 232256
rect 645519 232253 645585 232256
rect 144111 232168 144177 232171
rect 140802 232166 144177 232168
rect 140802 232110 144116 232166
rect 144172 232110 144177 232166
rect 140802 232108 144177 232110
rect 144111 232105 144177 232108
rect 206895 232168 206961 232171
rect 210498 232168 210558 232212
rect 206895 232166 210558 232168
rect 206895 232110 206900 232166
rect 206956 232110 210558 232166
rect 206895 232108 210558 232110
rect 206895 232105 206961 232108
rect 41871 231726 41937 231727
rect 41871 231724 41920 231726
rect 41828 231722 41920 231724
rect 41828 231666 41876 231722
rect 41828 231664 41920 231666
rect 41871 231662 41920 231664
rect 41984 231662 41990 231726
rect 206703 231724 206769 231727
rect 645231 231724 645297 231727
rect 206703 231722 210528 231724
rect 206703 231666 206708 231722
rect 206764 231666 210528 231722
rect 206703 231664 210528 231666
rect 640224 231722 645297 231724
rect 640224 231666 645236 231722
rect 645292 231666 645297 231722
rect 640224 231664 645297 231666
rect 41871 231661 41937 231662
rect 206703 231661 206769 231664
rect 645231 231661 645297 231664
rect 144015 231428 144081 231431
rect 140832 231426 144081 231428
rect 140832 231370 144020 231426
rect 144076 231370 144081 231426
rect 140832 231368 144081 231370
rect 144015 231365 144081 231368
rect 41775 231134 41841 231135
rect 41722 231070 41728 231134
rect 41792 231132 41841 231134
rect 206607 231132 206673 231135
rect 645135 231132 645201 231135
rect 41792 231130 41884 231132
rect 41836 231074 41884 231130
rect 41792 231072 41884 231074
rect 206607 231130 210528 231132
rect 206607 231074 206612 231130
rect 206668 231074 210528 231130
rect 206607 231072 210528 231074
rect 640224 231130 645201 231132
rect 640224 231074 645140 231130
rect 645196 231074 645201 231130
rect 640224 231072 645201 231074
rect 41792 231070 41841 231072
rect 41775 231069 41841 231070
rect 206607 231069 206673 231072
rect 645135 231069 645201 231072
rect 42063 230542 42129 230543
rect 42063 230538 42112 230542
rect 42176 230540 42182 230542
rect 204783 230540 204849 230543
rect 206991 230540 207057 230543
rect 645327 230540 645393 230543
rect 42063 230482 42068 230538
rect 42063 230478 42112 230482
rect 42176 230480 42220 230540
rect 204783 230538 210528 230540
rect 204783 230482 204788 230538
rect 204844 230482 206996 230538
rect 207052 230482 210528 230538
rect 204783 230480 210528 230482
rect 640224 230538 645393 230540
rect 640224 230482 645332 230538
rect 645388 230482 645393 230538
rect 640224 230480 645393 230482
rect 42176 230478 42182 230480
rect 42063 230477 42129 230478
rect 204783 230477 204849 230480
rect 206991 230477 207057 230480
rect 645327 230477 645393 230480
rect 144207 230244 144273 230247
rect 140832 230242 144273 230244
rect 140832 230186 144212 230242
rect 144268 230186 144273 230242
rect 140832 230184 144273 230186
rect 144207 230181 144273 230184
rect 146895 230096 146961 230099
rect 166863 230096 166929 230099
rect 146895 230094 166929 230096
rect 146895 230038 146900 230094
rect 146956 230038 166868 230094
rect 166924 230038 166929 230094
rect 146895 230036 166929 230038
rect 146895 230033 146961 230036
rect 166863 230033 166929 230036
rect 204879 230096 204945 230099
rect 206511 230096 206577 230099
rect 204879 230094 210528 230096
rect 204879 230038 204884 230094
rect 204940 230038 206516 230094
rect 206572 230038 210528 230094
rect 204879 230036 210528 230038
rect 204879 230033 204945 230036
rect 206511 230033 206577 230036
rect 41146 229590 41152 229654
rect 41216 229652 41222 229654
rect 41775 229652 41841 229655
rect 41216 229650 41841 229652
rect 41216 229594 41780 229650
rect 41836 229594 41841 229650
rect 41216 229592 41841 229594
rect 41216 229590 41222 229592
rect 41775 229589 41841 229592
rect 201711 229504 201777 229507
rect 674415 229504 674481 229507
rect 201711 229502 210528 229504
rect 201711 229446 201716 229502
rect 201772 229446 210528 229502
rect 201711 229444 210528 229446
rect 674415 229502 674784 229504
rect 674415 229446 674420 229502
rect 674476 229446 674784 229502
rect 674415 229444 674784 229446
rect 201711 229441 201777 229444
rect 674415 229441 674481 229444
rect 40954 228998 40960 229062
rect 41024 229060 41030 229062
rect 41775 229060 41841 229063
rect 41024 229058 41841 229060
rect 41024 229002 41780 229058
rect 41836 229002 41841 229058
rect 41024 229000 41841 229002
rect 41024 228998 41030 229000
rect 41775 228997 41841 229000
rect 140802 228468 140862 228956
rect 210063 228912 210129 228915
rect 674703 228912 674769 228915
rect 210063 228910 210528 228912
rect 210063 228854 210068 228910
rect 210124 228854 210528 228910
rect 210063 228852 210528 228854
rect 674703 228910 674814 228912
rect 674703 228854 674708 228910
rect 674764 228854 674814 228910
rect 210063 228849 210129 228852
rect 674703 228849 674814 228854
rect 674754 228660 674814 228849
rect 144015 228468 144081 228471
rect 140802 228466 144081 228468
rect 140802 228410 144020 228466
rect 144076 228410 144081 228466
rect 140802 228408 144081 228410
rect 144015 228405 144081 228408
rect 201615 228468 201681 228471
rect 201615 228466 210528 228468
rect 201615 228410 201620 228466
rect 201676 228410 210528 228466
rect 201615 228408 210528 228410
rect 201615 228405 201681 228408
rect 140802 227728 140862 227914
rect 201807 227876 201873 227879
rect 674415 227876 674481 227879
rect 201807 227874 210528 227876
rect 201807 227818 201812 227874
rect 201868 227818 210528 227874
rect 201807 227816 210528 227818
rect 674415 227874 674784 227876
rect 674415 227818 674420 227874
rect 674476 227818 674784 227874
rect 674415 227816 674784 227818
rect 201807 227813 201873 227816
rect 674415 227813 674481 227816
rect 144111 227728 144177 227731
rect 140802 227726 144177 227728
rect 140802 227670 144116 227726
rect 144172 227670 144177 227726
rect 140802 227668 144177 227670
rect 144111 227665 144177 227668
rect 40570 227518 40576 227582
rect 40640 227580 40646 227582
rect 41530 227580 41536 227582
rect 40640 227520 41536 227580
rect 40640 227518 40646 227520
rect 41530 227518 41536 227520
rect 41600 227518 41606 227582
rect 40378 227222 40384 227286
rect 40448 227284 40454 227286
rect 41775 227284 41841 227287
rect 40448 227282 41841 227284
rect 40448 227226 41780 227282
rect 41836 227226 41841 227282
rect 40448 227224 41841 227226
rect 40448 227222 40454 227224
rect 41775 227221 41841 227224
rect 201711 227284 201777 227287
rect 201711 227282 210528 227284
rect 201711 227226 201716 227282
rect 201772 227226 210528 227282
rect 201711 227224 210528 227226
rect 201711 227221 201777 227224
rect 40762 226778 40768 226842
rect 40832 226840 40838 226842
rect 41775 226840 41841 226843
rect 40832 226838 41841 226840
rect 40832 226782 41780 226838
rect 41836 226782 41841 226838
rect 40832 226780 41841 226782
rect 40832 226778 40838 226780
rect 41775 226777 41841 226780
rect 201807 226840 201873 226843
rect 675714 226842 675774 227032
rect 201807 226838 210528 226840
rect 201807 226782 201812 226838
rect 201868 226782 210528 226838
rect 201807 226780 210528 226782
rect 201807 226777 201873 226780
rect 675706 226778 675712 226842
rect 675776 226778 675782 226842
rect 144015 226692 144081 226695
rect 140832 226690 144081 226692
rect 140832 226634 144020 226690
rect 144076 226634 144081 226690
rect 140832 226632 144081 226634
rect 144015 226629 144081 226632
rect 201615 226248 201681 226251
rect 201615 226246 210528 226248
rect 201615 226190 201620 226246
rect 201676 226190 210528 226246
rect 201615 226188 210528 226190
rect 201615 226185 201681 226188
rect 673978 226186 673984 226250
rect 674048 226248 674054 226250
rect 674048 226188 674784 226248
rect 674048 226186 674054 226188
rect 40570 225890 40576 225954
rect 40640 225952 40646 225954
rect 41775 225952 41841 225955
rect 40640 225950 41841 225952
rect 40640 225894 41780 225950
rect 41836 225894 41841 225950
rect 40640 225892 41841 225894
rect 40640 225890 40646 225892
rect 41775 225889 41841 225892
rect 679791 225804 679857 225807
rect 679746 225802 679857 225804
rect 679746 225746 679796 225802
rect 679852 225746 679857 225802
rect 679746 225741 679857 225746
rect 197583 225656 197649 225659
rect 197583 225654 210528 225656
rect 197583 225598 197588 225654
rect 197644 225598 210528 225654
rect 197583 225596 210528 225598
rect 197583 225593 197649 225596
rect 679746 225552 679806 225741
rect 140802 225064 140862 225466
rect 201519 225212 201585 225215
rect 201519 225210 210528 225212
rect 201519 225154 201524 225210
rect 201580 225154 210528 225210
rect 201519 225152 210528 225154
rect 201519 225149 201585 225152
rect 144015 225064 144081 225067
rect 140802 225062 144081 225064
rect 140802 225006 144020 225062
rect 144076 225006 144081 225062
rect 140802 225004 144081 225006
rect 144015 225001 144081 225004
rect 679983 224916 680049 224919
rect 679938 224914 680049 224916
rect 679938 224858 679988 224914
rect 680044 224858 680049 224914
rect 679938 224853 680049 224858
rect 679938 224738 679998 224853
rect 201711 224620 201777 224623
rect 201711 224618 210528 224620
rect 201711 224562 201716 224618
rect 201772 224562 210528 224618
rect 201711 224560 210528 224562
rect 201711 224557 201777 224560
rect 140802 223732 140862 224220
rect 201615 224028 201681 224031
rect 201615 224026 210528 224028
rect 201615 223970 201620 224026
rect 201676 223970 210528 224026
rect 201615 223968 210528 223970
rect 201615 223965 201681 223968
rect 677250 223735 677310 223850
rect 144111 223732 144177 223735
rect 140802 223730 144177 223732
rect 140802 223674 144116 223730
rect 144172 223674 144177 223730
rect 140802 223672 144177 223674
rect 144111 223669 144177 223672
rect 677199 223730 677310 223735
rect 677199 223674 677204 223730
rect 677260 223674 677310 223730
rect 677199 223672 677310 223674
rect 677199 223669 677265 223672
rect 201711 223584 201777 223587
rect 201711 223582 210528 223584
rect 201711 223526 201716 223582
rect 201772 223526 210528 223582
rect 201711 223524 210528 223526
rect 201711 223521 201777 223524
rect 674362 223078 674368 223142
rect 674432 223140 674438 223142
rect 674432 223080 674784 223140
rect 674432 223078 674438 223080
rect 144015 222992 144081 222995
rect 140832 222990 144081 222992
rect 140832 222934 144020 222990
rect 144076 222934 144081 222990
rect 140832 222932 144081 222934
rect 144015 222929 144081 222932
rect 201807 222992 201873 222995
rect 201807 222990 210528 222992
rect 201807 222934 201812 222990
rect 201868 222934 210528 222990
rect 201807 222932 210528 222934
rect 201807 222929 201873 222932
rect 201519 222400 201585 222403
rect 201519 222398 210528 222400
rect 201519 222342 201524 222398
rect 201580 222342 210528 222398
rect 201519 222340 210528 222342
rect 201519 222337 201585 222340
rect 674415 222252 674481 222255
rect 674415 222250 674784 222252
rect 674415 222194 674420 222250
rect 674476 222194 674784 222250
rect 674415 222192 674784 222194
rect 674415 222189 674481 222192
rect 209967 221882 210033 221885
rect 209967 221880 210528 221882
rect 209967 221824 209972 221880
rect 210028 221824 210528 221880
rect 209967 221822 210528 221824
rect 209967 221819 210033 221822
rect 145594 221808 145600 221810
rect 140832 221748 145600 221808
rect 145594 221746 145600 221748
rect 145664 221746 145670 221810
rect 198639 221364 198705 221367
rect 198639 221362 210528 221364
rect 198639 221306 198644 221362
rect 198700 221306 210528 221362
rect 198639 221304 210528 221306
rect 198639 221301 198705 221304
rect 674946 221219 675006 221482
rect 674946 221214 675057 221219
rect 674946 221158 674996 221214
rect 675052 221158 675057 221214
rect 674946 221156 675057 221158
rect 674991 221153 675057 221156
rect 42351 221068 42417 221071
rect 42306 221066 42417 221068
rect 42306 221010 42356 221066
rect 42412 221010 42417 221066
rect 42306 221005 42417 221010
rect 42306 220890 42366 221005
rect 201711 220772 201777 220775
rect 201711 220770 210528 220772
rect 201711 220714 201716 220770
rect 201772 220714 210528 220770
rect 201711 220712 210528 220714
rect 201711 220709 201777 220712
rect 42351 220328 42417 220331
rect 42306 220326 42417 220328
rect 42306 220270 42356 220326
rect 42412 220270 42417 220326
rect 42306 220265 42417 220270
rect 42306 220076 42366 220265
rect 140802 220180 140862 220668
rect 677058 220627 677118 220742
rect 677007 220622 677118 220627
rect 677007 220566 677012 220622
rect 677068 220566 677118 220622
rect 677007 220564 677118 220566
rect 677007 220561 677073 220564
rect 209967 220254 210033 220257
rect 209967 220252 210528 220254
rect 209967 220196 209972 220252
rect 210028 220196 210528 220252
rect 209967 220194 210528 220196
rect 209967 220191 210033 220194
rect 144015 220180 144081 220183
rect 140802 220178 144081 220180
rect 140802 220122 144020 220178
rect 144076 220122 144081 220178
rect 140802 220120 144081 220122
rect 144015 220117 144081 220120
rect 677058 219739 677118 220002
rect 201615 219736 201681 219739
rect 201615 219734 210528 219736
rect 201615 219678 201620 219734
rect 201676 219678 210528 219734
rect 201615 219676 210528 219678
rect 677058 219734 677169 219739
rect 677058 219678 677108 219734
rect 677164 219678 677169 219734
rect 677058 219676 677169 219678
rect 201615 219673 201681 219676
rect 677103 219673 677169 219676
rect 42351 219440 42417 219443
rect 42306 219438 42417 219440
rect 42306 219382 42356 219438
rect 42412 219382 42417 219438
rect 42306 219377 42417 219382
rect 42306 219262 42366 219377
rect 140802 218996 140862 219482
rect 201807 219144 201873 219147
rect 201807 219142 210528 219144
rect 201807 219086 201812 219142
rect 201868 219086 210528 219142
rect 201807 219084 210528 219086
rect 201807 219081 201873 219084
rect 145786 218996 145792 218998
rect 140802 218936 145792 218996
rect 145786 218934 145792 218936
rect 145856 218934 145862 218998
rect 209967 218626 210033 218629
rect 209967 218624 210528 218626
rect 209967 218568 209972 218624
rect 210028 218568 210528 218624
rect 209967 218566 210528 218568
rect 209967 218563 210033 218566
rect 675138 218555 675198 219114
rect 675138 218550 675249 218555
rect 675138 218494 675188 218550
rect 675244 218494 675249 218550
rect 675138 218492 675249 218494
rect 675183 218489 675249 218492
rect 144015 218256 144081 218259
rect 140832 218254 144081 218256
rect 140832 218198 144020 218254
rect 144076 218198 144081 218254
rect 140832 218196 144081 218198
rect 144015 218193 144081 218196
rect 675138 218111 675198 218374
rect 201711 218108 201777 218111
rect 201711 218106 210528 218108
rect 201711 218050 201716 218106
rect 201772 218050 210528 218106
rect 201711 218048 210528 218050
rect 675087 218106 675198 218111
rect 675087 218050 675092 218106
rect 675148 218050 675198 218106
rect 675087 218048 675198 218050
rect 201711 218045 201777 218048
rect 675087 218045 675153 218048
rect 675130 217750 675136 217814
rect 675200 217812 675206 217814
rect 675279 217812 675345 217815
rect 675200 217810 675345 217812
rect 675200 217754 675284 217810
rect 675340 217754 675345 217810
rect 675200 217752 675345 217754
rect 675200 217750 675206 217752
rect 675279 217749 675345 217752
rect 43215 217664 43281 217667
rect 42336 217662 43281 217664
rect 42336 217606 43220 217662
rect 43276 217606 43281 217662
rect 42336 217604 43281 217606
rect 43215 217601 43281 217604
rect 198159 217516 198225 217519
rect 674319 217516 674385 217519
rect 198159 217514 210528 217516
rect 198159 217458 198164 217514
rect 198220 217458 210528 217514
rect 198159 217456 210528 217458
rect 674319 217514 674784 217516
rect 674319 217458 674324 217514
rect 674380 217458 674784 217514
rect 674319 217456 674784 217458
rect 198159 217453 198225 217456
rect 674319 217453 674385 217456
rect 43503 216924 43569 216927
rect 42336 216922 43569 216924
rect 42336 216866 43508 216922
rect 43564 216866 43569 216922
rect 42336 216864 43569 216866
rect 43503 216861 43569 216864
rect 140802 216480 140862 217034
rect 210159 216998 210225 217001
rect 210159 216996 210528 216998
rect 210159 216940 210164 216996
rect 210220 216940 210528 216996
rect 210159 216938 210528 216940
rect 210159 216935 210225 216938
rect 676866 216483 676926 216746
rect 145978 216480 145984 216482
rect 140802 216420 145984 216480
rect 145978 216418 145984 216420
rect 146048 216418 146054 216482
rect 197583 216480 197649 216483
rect 197583 216478 210528 216480
rect 197583 216422 197588 216478
rect 197644 216422 210528 216478
rect 197583 216420 210528 216422
rect 676866 216478 676977 216483
rect 676866 216422 676916 216478
rect 676972 216422 676977 216478
rect 676866 216420 676977 216422
rect 197583 216417 197649 216420
rect 676911 216417 676977 216420
rect 43311 216184 43377 216187
rect 42336 216182 43377 216184
rect 42336 216126 43316 216182
rect 43372 216126 43377 216182
rect 42336 216124 43377 216126
rect 43311 216121 43377 216124
rect 676866 215891 676926 216006
rect 201711 215888 201777 215891
rect 201711 215886 210528 215888
rect 201711 215830 201716 215886
rect 201772 215830 210528 215886
rect 201711 215828 210528 215830
rect 676815 215886 676926 215891
rect 676815 215830 676820 215886
rect 676876 215830 676926 215886
rect 676815 215828 676926 215830
rect 201711 215825 201777 215828
rect 676815 215825 676881 215828
rect 140802 215296 140862 215784
rect 209967 215370 210033 215373
rect 209967 215368 210528 215370
rect 209967 215312 209972 215368
rect 210028 215312 210528 215368
rect 209967 215310 210528 215312
rect 209967 215307 210033 215310
rect 144111 215296 144177 215299
rect 140802 215294 144177 215296
rect 40386 214706 40446 215266
rect 140802 215238 144116 215294
rect 144172 215238 144177 215294
rect 140802 215236 144177 215238
rect 144111 215233 144177 215236
rect 674946 215003 675006 215192
rect 674895 214998 675006 215003
rect 674895 214942 674900 214998
rect 674956 214942 675006 214998
rect 674895 214940 675006 214942
rect 674895 214937 674961 214940
rect 201615 214852 201681 214855
rect 201615 214850 210528 214852
rect 201615 214794 201620 214850
rect 201676 214794 210528 214850
rect 201615 214792 210528 214794
rect 201615 214789 201681 214792
rect 40378 214642 40384 214706
rect 40448 214642 40454 214706
rect 145359 214556 145425 214559
rect 140832 214554 145425 214556
rect 41922 213967 41982 214526
rect 140832 214498 145364 214554
rect 145420 214498 145425 214554
rect 140832 214496 145425 214498
rect 145359 214493 145425 214496
rect 674754 214263 674814 214378
rect 201231 214260 201297 214263
rect 201231 214258 210528 214260
rect 201231 214202 201236 214258
rect 201292 214202 210528 214258
rect 201231 214200 210528 214202
rect 674754 214258 674865 214263
rect 674754 214202 674804 214258
rect 674860 214202 674865 214258
rect 674754 214200 674865 214202
rect 201231 214197 201297 214200
rect 674799 214197 674865 214200
rect 41922 213962 42033 213967
rect 41922 213906 41972 213962
rect 42028 213906 42033 213962
rect 41922 213904 42033 213906
rect 41967 213901 42033 213904
rect 210159 213742 210225 213745
rect 210159 213740 210528 213742
rect 210159 213684 210164 213740
rect 210220 213684 210528 213740
rect 210159 213682 210528 213684
rect 210159 213679 210225 213682
rect 40578 213226 40638 213638
rect 674754 213375 674814 213564
rect 144015 213372 144081 213375
rect 140832 213370 144081 213372
rect 140832 213314 144020 213370
rect 144076 213314 144081 213370
rect 140832 213312 144081 213314
rect 144015 213309 144081 213312
rect 674703 213370 674814 213375
rect 674703 213314 674708 213370
rect 674764 213314 674814 213370
rect 674703 213312 674814 213314
rect 674703 213309 674769 213312
rect 40570 213162 40576 213226
rect 40640 213162 40646 213226
rect 201807 213224 201873 213227
rect 201807 213222 210528 213224
rect 201807 213166 201812 213222
rect 201868 213166 210528 213222
rect 201807 213164 210528 213166
rect 201807 213161 201873 213164
rect 40962 212486 41022 212898
rect 201711 212632 201777 212635
rect 201711 212630 210528 212632
rect 201711 212574 201716 212630
rect 201772 212574 210528 212630
rect 201711 212572 210528 212574
rect 201711 212569 201777 212572
rect 40954 212422 40960 212486
rect 41024 212422 41030 212486
rect 41154 211598 41214 212158
rect 140802 211744 140862 212232
rect 679746 212191 679806 212750
rect 679695 212186 679806 212191
rect 679695 212130 679700 212186
rect 679756 212130 679806 212186
rect 679695 212128 679806 212130
rect 679695 212125 679761 212128
rect 209967 212114 210033 212117
rect 209967 212112 210528 212114
rect 209967 212056 209972 212112
rect 210028 212056 210528 212112
rect 209967 212054 210528 212056
rect 209967 212051 210033 212054
rect 144015 211744 144081 211747
rect 140802 211742 144081 211744
rect 140802 211686 144020 211742
rect 144076 211686 144081 211742
rect 140802 211684 144081 211686
rect 144015 211681 144081 211684
rect 675130 211682 675136 211746
rect 675200 211744 675206 211746
rect 675279 211744 675345 211747
rect 675200 211742 675345 211744
rect 675200 211686 675284 211742
rect 675340 211686 675345 211742
rect 675200 211684 675345 211686
rect 675200 211682 675206 211684
rect 675279 211681 675345 211684
rect 41146 211534 41152 211598
rect 41216 211534 41222 211598
rect 201615 211596 201681 211599
rect 201615 211594 210528 211596
rect 201615 211538 201620 211594
rect 201676 211538 210528 211594
rect 201615 211536 210528 211538
rect 201615 211533 201681 211536
rect 674746 211534 674752 211598
rect 674816 211596 674822 211598
rect 675514 211596 675520 211598
rect 674816 211536 675520 211596
rect 674816 211534 674822 211536
rect 675514 211534 675520 211536
rect 675584 211534 675590 211598
rect 679695 211448 679761 211451
rect 679695 211446 679806 211448
rect 41922 210859 41982 211418
rect 679695 211390 679700 211446
rect 679756 211390 679806 211446
rect 679695 211385 679806 211390
rect 679746 211270 679806 211385
rect 41871 210854 41982 210859
rect 41871 210798 41876 210854
rect 41932 210798 41982 210854
rect 41871 210796 41982 210798
rect 41871 210793 41937 210796
rect 140802 210560 140862 211048
rect 646095 211004 646161 211007
rect 640224 211002 646161 211004
rect 640224 210946 646100 211002
rect 646156 210946 646161 211002
rect 640224 210944 646161 210946
rect 646095 210941 646161 210944
rect 145455 210560 145521 210563
rect 140802 210558 145521 210560
rect 40770 210414 40830 210530
rect 140802 210502 145460 210558
rect 145516 210502 145521 210558
rect 140802 210500 145521 210502
rect 145455 210497 145521 210500
rect 40762 210350 40768 210414
rect 40832 210350 40838 210414
rect 676090 210202 676096 210266
rect 676160 210264 676166 210266
rect 676911 210264 676977 210267
rect 676160 210262 676977 210264
rect 676160 210206 676916 210262
rect 676972 210206 676977 210262
rect 676160 210204 676977 210206
rect 676160 210202 676166 210204
rect 676911 210201 676977 210204
rect 675514 210054 675520 210118
rect 675584 210116 675590 210118
rect 677007 210116 677073 210119
rect 675584 210114 677073 210116
rect 675584 210058 677012 210114
rect 677068 210058 677073 210114
rect 675584 210056 677073 210058
rect 675584 210054 675590 210056
rect 677007 210053 677073 210056
rect 676282 209906 676288 209970
rect 676352 209968 676358 209970
rect 677103 209968 677169 209971
rect 676352 209966 677169 209968
rect 676352 209910 677108 209966
rect 677164 209910 677169 209966
rect 676352 209908 677169 209910
rect 676352 209906 676358 209908
rect 677103 209905 677169 209908
rect 43119 209820 43185 209823
rect 144111 209820 144177 209823
rect 42336 209818 43185 209820
rect 42336 209762 43124 209818
rect 43180 209762 43185 209818
rect 42336 209760 43185 209762
rect 140832 209818 144177 209820
rect 140832 209762 144116 209818
rect 144172 209762 144177 209818
rect 140832 209760 144177 209762
rect 43119 209757 43185 209760
rect 144111 209757 144177 209760
rect 675898 209758 675904 209822
rect 675968 209820 675974 209822
rect 677199 209820 677265 209823
rect 675968 209818 677265 209820
rect 675968 209762 677204 209818
rect 677260 209762 677265 209818
rect 675968 209760 677265 209762
rect 675968 209758 675974 209760
rect 677199 209757 677265 209760
rect 675706 209610 675712 209674
rect 675776 209672 675782 209674
rect 679791 209672 679857 209675
rect 675776 209670 679857 209672
rect 675776 209614 679796 209670
rect 679852 209614 679857 209670
rect 675776 209612 679857 209614
rect 675776 209610 675782 209612
rect 679791 209609 679857 209612
rect 676474 209462 676480 209526
rect 676544 209524 676550 209526
rect 679983 209524 680049 209527
rect 676544 209522 680049 209524
rect 676544 209466 679988 209522
rect 680044 209466 680049 209522
rect 676544 209464 680049 209466
rect 676544 209462 676550 209464
rect 679983 209461 680049 209464
rect 42114 208343 42174 208902
rect 210490 208722 210496 208786
rect 210560 208784 210566 208786
rect 210874 208784 210880 208786
rect 210560 208724 210880 208784
rect 210560 208722 210566 208724
rect 210874 208722 210880 208724
rect 210944 208722 210950 208786
rect 42063 208338 42174 208343
rect 42063 208282 42068 208338
rect 42124 208282 42174 208338
rect 42063 208280 42174 208282
rect 42063 208277 42129 208280
rect 37314 207751 37374 208088
rect 140802 208044 140862 208602
rect 145551 208044 145617 208047
rect 140802 208042 145617 208044
rect 140802 207986 145556 208042
rect 145612 207986 145617 208042
rect 140802 207984 145617 207986
rect 145551 207981 145617 207984
rect 37263 207746 37374 207751
rect 37263 207690 37268 207746
rect 37324 207690 37374 207746
rect 37263 207688 37374 207690
rect 37263 207685 37329 207688
rect 144015 207452 144081 207455
rect 140832 207450 144081 207452
rect 40194 207159 40254 207422
rect 140832 207394 144020 207450
rect 144076 207394 144081 207450
rect 140832 207392 144081 207394
rect 144015 207389 144081 207392
rect 40143 207154 40254 207159
rect 40143 207098 40148 207154
rect 40204 207098 40254 207154
rect 40143 207096 40254 207098
rect 40143 207093 40209 207096
rect 37314 206123 37374 206608
rect 210874 206354 210880 206418
rect 210944 206354 210950 206418
rect 37314 206118 37425 206123
rect 37314 206062 37364 206118
rect 37420 206062 37425 206118
rect 37314 206060 37425 206062
rect 37359 206057 37425 206060
rect 42306 205531 42366 205794
rect 140802 205676 140862 206154
rect 210882 205974 210942 206354
rect 210874 205910 210880 205974
rect 210944 205910 210950 205974
rect 145647 205676 145713 205679
rect 140802 205674 145713 205676
rect 140802 205618 145652 205674
rect 145708 205618 145713 205674
rect 140802 205616 145713 205618
rect 145647 205613 145713 205616
rect 42306 205526 42417 205531
rect 42306 205470 42356 205526
rect 42412 205470 42417 205526
rect 42306 205468 42417 205470
rect 42351 205465 42417 205468
rect 145839 205084 145905 205087
rect 140832 205082 145905 205084
rect 140832 205026 145844 205082
rect 145900 205026 145905 205082
rect 140832 205024 145905 205026
rect 145839 205021 145905 205024
rect 40194 204643 40254 204980
rect 40194 204638 40305 204643
rect 40194 204582 40244 204638
rect 40300 204582 40305 204638
rect 40194 204580 40305 204582
rect 40239 204577 40305 204580
rect 42159 204344 42225 204347
rect 42114 204342 42225 204344
rect 42114 204286 42164 204342
rect 42220 204286 42225 204342
rect 42114 204281 42225 204286
rect 675759 204344 675825 204347
rect 675898 204344 675904 204346
rect 675759 204342 675904 204344
rect 675759 204286 675764 204342
rect 675820 204286 675904 204342
rect 675759 204284 675904 204286
rect 675759 204281 675825 204284
rect 675898 204282 675904 204284
rect 675968 204282 675974 204346
rect 42114 204166 42174 204281
rect 140802 203308 140862 203796
rect 144207 203308 144273 203311
rect 140802 203306 144273 203308
rect 140802 203250 144212 203306
rect 144268 203250 144273 203306
rect 140802 203248 144273 203250
rect 144207 203245 144273 203248
rect 42159 203012 42225 203015
rect 42114 203010 42225 203012
rect 42114 202954 42164 203010
rect 42220 202954 42225 203010
rect 42114 202949 42225 202954
rect 42114 202686 42174 202949
rect 206415 202864 206481 202867
rect 206415 202862 210528 202864
rect 206415 202806 206420 202862
rect 206476 202806 210528 202862
rect 206415 202804 210528 202806
rect 206415 202801 206481 202804
rect 140802 202124 140862 202612
rect 146799 202124 146865 202127
rect 140802 202122 146865 202124
rect 140802 202066 146804 202122
rect 146860 202066 146865 202122
rect 140802 202064 146865 202066
rect 146799 202061 146865 202064
rect 145743 201384 145809 201387
rect 140832 201382 145809 201384
rect 140832 201326 145748 201382
rect 145804 201326 145809 201382
rect 140832 201324 145809 201326
rect 145743 201321 145809 201324
rect 140802 199608 140862 200142
rect 674746 199694 674752 199758
rect 674816 199756 674822 199758
rect 675087 199756 675153 199759
rect 674816 199754 675153 199756
rect 674816 199698 675092 199754
rect 675148 199698 675153 199754
rect 674816 199696 675153 199698
rect 674816 199694 674822 199696
rect 675087 199693 675153 199696
rect 146703 199608 146769 199611
rect 140802 199606 146769 199608
rect 140802 199550 146708 199606
rect 146764 199550 146769 199606
rect 140802 199548 146769 199550
rect 146703 199545 146769 199548
rect 675183 199166 675249 199167
rect 675130 199164 675136 199166
rect 675092 199104 675136 199164
rect 675200 199162 675249 199166
rect 675244 199106 675249 199162
rect 675130 199102 675136 199104
rect 675200 199102 675249 199106
rect 675183 199101 675249 199102
rect 146799 199016 146865 199019
rect 140832 199014 146865 199016
rect 140832 198958 146804 199014
rect 146860 198958 146865 199014
rect 140832 198956 146865 198958
rect 146799 198953 146865 198956
rect 675471 198426 675537 198427
rect 675471 198422 675520 198426
rect 675584 198424 675590 198426
rect 675471 198366 675476 198422
rect 675471 198362 675520 198366
rect 675584 198364 675628 198424
rect 675584 198362 675590 198364
rect 675471 198361 675537 198362
rect 146799 197832 146865 197835
rect 140832 197830 146865 197832
rect 140832 197774 146804 197830
rect 146860 197774 146865 197830
rect 140832 197772 146865 197774
rect 146799 197769 146865 197772
rect 42159 197684 42225 197687
rect 42298 197684 42304 197686
rect 42159 197682 42304 197684
rect 42159 197626 42164 197682
rect 42220 197626 42304 197682
rect 42159 197624 42304 197626
rect 42159 197621 42225 197624
rect 42298 197622 42304 197624
rect 42368 197622 42374 197686
rect 42106 197326 42112 197390
rect 42176 197388 42182 197390
rect 42351 197388 42417 197391
rect 42176 197386 42417 197388
rect 42176 197330 42356 197386
rect 42412 197330 42417 197386
rect 42176 197328 42417 197330
rect 42176 197326 42182 197328
rect 42351 197325 42417 197328
rect 144783 196648 144849 196651
rect 140832 196646 144849 196648
rect 140832 196590 144788 196646
rect 144844 196590 144849 196646
rect 140832 196588 144849 196590
rect 144783 196585 144849 196588
rect 675183 195760 675249 195763
rect 675322 195760 675328 195762
rect 675183 195758 675328 195760
rect 675183 195702 675188 195758
rect 675244 195702 675328 195758
rect 675183 195700 675328 195702
rect 675183 195697 675249 195700
rect 675322 195698 675328 195700
rect 675392 195698 675398 195762
rect 675087 195612 675153 195615
rect 675514 195612 675520 195614
rect 675087 195610 675520 195612
rect 675087 195554 675092 195610
rect 675148 195554 675520 195610
rect 675087 195552 675520 195554
rect 675087 195549 675153 195552
rect 675514 195550 675520 195552
rect 675584 195550 675590 195614
rect 42351 195170 42417 195171
rect 42298 195168 42304 195170
rect 42260 195108 42304 195168
rect 42368 195166 42417 195170
rect 42412 195110 42417 195166
rect 42298 195106 42304 195108
rect 42368 195106 42417 195110
rect 42351 195105 42417 195106
rect 140802 194872 140862 195360
rect 675759 195316 675825 195319
rect 676090 195316 676096 195318
rect 675759 195314 676096 195316
rect 675759 195258 675764 195314
rect 675820 195258 676096 195314
rect 675759 195256 676096 195258
rect 675759 195253 675825 195256
rect 676090 195254 676096 195256
rect 676160 195254 676166 195318
rect 144591 194872 144657 194875
rect 140802 194870 144657 194872
rect 140802 194814 144596 194870
rect 144652 194814 144657 194870
rect 140802 194812 144657 194814
rect 144591 194809 144657 194812
rect 140802 193688 140862 194176
rect 146799 193688 146865 193691
rect 140802 193686 146865 193688
rect 140802 193630 146804 193686
rect 146860 193630 146865 193686
rect 140802 193628 146865 193630
rect 146799 193625 146865 193628
rect 674362 193478 674368 193542
rect 674432 193540 674438 193542
rect 675375 193540 675441 193543
rect 674432 193538 675441 193540
rect 674432 193482 675380 193538
rect 675436 193482 675441 193538
rect 674432 193480 675441 193482
rect 674432 193478 674438 193480
rect 675375 193477 675441 193480
rect 146799 192948 146865 192951
rect 140832 192946 146865 192948
rect 140832 192890 146804 192946
rect 146860 192890 146865 192946
rect 140832 192888 146865 192890
rect 146799 192885 146865 192888
rect 146703 191764 146769 191767
rect 140832 191762 146769 191764
rect 140832 191706 146708 191762
rect 146764 191706 146769 191762
rect 140832 191704 146769 191706
rect 146703 191701 146769 191704
rect 675759 191616 675825 191619
rect 676282 191616 676288 191618
rect 675759 191614 676288 191616
rect 675759 191558 675764 191614
rect 675820 191558 676288 191614
rect 675759 191556 676288 191558
rect 675759 191553 675825 191556
rect 676282 191554 676288 191556
rect 676352 191554 676358 191618
rect 42063 191026 42129 191027
rect 42063 191024 42112 191026
rect 42020 191022 42112 191024
rect 42020 190966 42068 191022
rect 42020 190964 42112 190966
rect 42063 190962 42112 190964
rect 42176 190962 42182 191026
rect 42063 190961 42129 190962
rect 41146 190074 41152 190138
rect 41216 190136 41222 190138
rect 41775 190136 41841 190139
rect 41216 190134 41841 190136
rect 41216 190078 41780 190134
rect 41836 190078 41841 190134
rect 41216 190076 41841 190078
rect 140802 190136 140862 190476
rect 145935 190136 146001 190139
rect 140802 190134 146001 190136
rect 140802 190078 145940 190134
rect 145996 190078 146001 190134
rect 140802 190076 146001 190078
rect 41216 190074 41222 190076
rect 41775 190073 41841 190076
rect 145935 190073 146001 190076
rect 146703 189396 146769 189399
rect 140832 189394 146769 189396
rect 140832 189338 146708 189394
rect 146764 189338 146769 189394
rect 140832 189336 146769 189338
rect 146703 189333 146769 189336
rect 41871 189102 41937 189103
rect 41871 189098 41920 189102
rect 41984 189100 41990 189102
rect 41871 189042 41876 189098
rect 41871 189038 41920 189042
rect 41984 189040 42028 189100
rect 41984 189038 41990 189040
rect 41871 189037 41937 189038
rect 41775 188362 41841 188363
rect 41722 188298 41728 188362
rect 41792 188360 41841 188362
rect 41792 188358 41884 188360
rect 41836 188302 41884 188358
rect 41792 188300 41884 188302
rect 41792 188298 41841 188300
rect 41775 188297 41841 188298
rect 146799 188212 146865 188215
rect 140832 188210 146865 188212
rect 140832 188154 146804 188210
rect 146860 188154 146865 188210
rect 140832 188152 146865 188154
rect 146799 188149 146865 188152
rect 140802 186436 140862 186924
rect 146127 186436 146193 186439
rect 140802 186434 146193 186436
rect 140802 186378 146132 186434
rect 146188 186378 146193 186434
rect 140802 186376 146193 186378
rect 146127 186373 146193 186376
rect 40954 185930 40960 185994
rect 41024 185992 41030 185994
rect 41775 185992 41841 185995
rect 41024 185990 41841 185992
rect 41024 185934 41780 185990
rect 41836 185934 41841 185990
rect 41024 185932 41841 185934
rect 41024 185930 41030 185932
rect 41775 185929 41841 185932
rect 140802 185252 140862 185740
rect 146319 185252 146385 185255
rect 140802 185250 146385 185252
rect 140802 185194 146324 185250
rect 146380 185194 146385 185250
rect 140802 185192 146385 185194
rect 146319 185189 146385 185192
rect 144015 184512 144081 184515
rect 140832 184510 144081 184512
rect 140832 184454 144020 184510
rect 144076 184454 144081 184510
rect 140832 184452 144081 184454
rect 144015 184449 144081 184452
rect 674415 184512 674481 184515
rect 674415 184510 674784 184512
rect 674415 184454 674420 184510
rect 674476 184454 674784 184510
rect 674415 184452 674784 184454
rect 674415 184449 674481 184452
rect 40378 184154 40384 184218
rect 40448 184216 40454 184218
rect 41775 184216 41841 184219
rect 40448 184214 41841 184216
rect 40448 184158 41780 184214
rect 41836 184158 41841 184214
rect 40448 184156 41841 184158
rect 40448 184154 40454 184156
rect 41775 184153 41841 184156
rect 674703 183920 674769 183923
rect 674703 183918 674814 183920
rect 674703 183862 674708 183918
rect 674764 183862 674814 183918
rect 674703 183857 674814 183862
rect 674754 183668 674814 183857
rect 40762 183562 40768 183626
rect 40832 183624 40838 183626
rect 41775 183624 41841 183627
rect 40832 183622 41841 183624
rect 40832 183566 41780 183622
rect 41836 183566 41841 183622
rect 40832 183564 41841 183566
rect 40832 183562 40838 183564
rect 41775 183561 41841 183564
rect 146415 183328 146481 183331
rect 140832 183326 146481 183328
rect 140832 183270 146420 183326
rect 146476 183270 146481 183326
rect 140832 183268 146481 183270
rect 146415 183265 146481 183268
rect 40570 182822 40576 182886
rect 40640 182884 40646 182886
rect 41775 182884 41841 182887
rect 40640 182882 41841 182884
rect 40640 182826 41780 182882
rect 41836 182826 41841 182882
rect 40640 182824 41841 182826
rect 40640 182822 40646 182824
rect 41775 182821 41841 182824
rect 674415 182884 674481 182887
rect 674415 182882 674784 182884
rect 674415 182826 674420 182882
rect 674476 182826 674784 182882
rect 674415 182824 674784 182826
rect 674415 182821 674481 182824
rect 210106 182674 210112 182738
rect 210176 182736 210182 182738
rect 210874 182736 210880 182738
rect 210176 182676 210880 182736
rect 210176 182674 210182 182676
rect 210874 182674 210880 182676
rect 210944 182674 210950 182738
rect 673978 182526 673984 182590
rect 674048 182588 674054 182590
rect 674048 182528 674814 182588
rect 674048 182526 674054 182528
rect 140802 181848 140862 182188
rect 674754 182040 674814 182528
rect 210298 181934 210304 181998
rect 210368 181996 210374 181998
rect 210874 181996 210880 181998
rect 210368 181936 210880 181996
rect 210368 181934 210374 181936
rect 210874 181934 210880 181936
rect 210944 181934 210950 181998
rect 144015 181848 144081 181851
rect 140802 181846 144081 181848
rect 140802 181790 144020 181846
rect 144076 181790 144081 181846
rect 140802 181788 144081 181790
rect 144015 181785 144081 181788
rect 673978 181194 673984 181258
rect 674048 181256 674054 181258
rect 674048 181196 674784 181256
rect 674048 181194 674054 181196
rect 140802 180516 140862 180994
rect 675706 180898 675712 180962
rect 675776 180898 675782 180962
rect 144111 180516 144177 180519
rect 140802 180514 144177 180516
rect 140802 180458 144116 180514
rect 144172 180458 144177 180514
rect 140802 180456 144177 180458
rect 144111 180453 144177 180456
rect 675714 179924 675774 180898
rect 679695 179924 679761 179927
rect 675714 179922 679761 179924
rect 675714 179866 679700 179922
rect 679756 179866 679761 179922
rect 675714 179864 679761 179866
rect 679695 179861 679761 179864
rect 146799 179776 146865 179779
rect 140832 179774 146865 179776
rect 140832 179718 146804 179774
rect 146860 179718 146865 179774
rect 140832 179716 146865 179718
rect 146799 179713 146865 179716
rect 676482 179482 676542 179746
rect 676474 179418 676480 179482
rect 676544 179480 676550 179482
rect 679791 179480 679857 179483
rect 676544 179478 679857 179480
rect 676544 179422 679796 179478
rect 679852 179422 679857 179478
rect 676544 179420 679857 179422
rect 676544 179418 676550 179420
rect 679791 179417 679857 179420
rect 674031 178888 674097 178891
rect 674031 178886 674784 178888
rect 674031 178830 674036 178886
rect 674092 178830 674784 178886
rect 674031 178828 674784 178830
rect 674031 178825 674097 178828
rect 144015 178592 144081 178595
rect 140832 178590 144081 178592
rect 140832 178534 144020 178590
rect 144076 178534 144081 178590
rect 140832 178532 144081 178534
rect 144015 178529 144081 178532
rect 674170 178086 674176 178150
rect 674240 178148 674246 178150
rect 674240 178088 674784 178148
rect 674240 178086 674246 178088
rect 31738 177050 31744 177114
rect 31808 177112 31814 177114
rect 42735 177112 42801 177115
rect 31808 177110 42801 177112
rect 31808 177054 42740 177110
rect 42796 177054 42801 177110
rect 31808 177052 42801 177054
rect 31808 177050 31814 177052
rect 42735 177049 42801 177052
rect 140802 176816 140862 177304
rect 674415 177260 674481 177263
rect 674415 177258 674784 177260
rect 674415 177202 674420 177258
rect 674476 177202 674784 177258
rect 674415 177200 674784 177202
rect 674415 177197 674481 177200
rect 144015 176816 144081 176819
rect 140802 176814 144081 176816
rect 140802 176758 144020 176814
rect 144076 176758 144081 176814
rect 140802 176756 144081 176758
rect 144015 176753 144081 176756
rect 677058 176227 677118 176490
rect 677007 176222 677118 176227
rect 677007 176166 677012 176222
rect 677068 176166 677118 176222
rect 677007 176164 677118 176166
rect 677007 176161 677073 176164
rect 146607 176076 146673 176079
rect 140832 176074 146673 176076
rect 140832 176018 146612 176074
rect 146668 176018 146673 176074
rect 140832 176016 146673 176018
rect 146607 176013 146673 176016
rect 676911 175632 676977 175635
rect 677058 175632 677118 175750
rect 676911 175630 677118 175632
rect 676911 175574 676916 175630
rect 676972 175574 677118 175630
rect 676911 175572 677118 175574
rect 676911 175569 676977 175572
rect 140802 174448 140862 174982
rect 677250 174747 677310 175010
rect 677199 174742 677310 174747
rect 677199 174686 677204 174742
rect 677260 174686 677310 174742
rect 677199 174684 677310 174686
rect 677199 174681 677265 174684
rect 144879 174448 144945 174451
rect 140802 174446 144945 174448
rect 140802 174390 144884 174446
rect 144940 174390 144945 174446
rect 140802 174388 144945 174390
rect 144879 174385 144945 174388
rect 675138 174007 675198 174122
rect 675138 174002 675249 174007
rect 675138 173946 675188 174002
rect 675244 173946 675249 174002
rect 675138 173944 675249 173946
rect 675183 173941 675249 173944
rect 140802 173412 140862 173752
rect 144015 173412 144081 173415
rect 140802 173410 144081 173412
rect 140802 173354 144020 173410
rect 144076 173354 144081 173410
rect 140802 173352 144081 173354
rect 144015 173349 144081 173352
rect 674946 173119 675006 173382
rect 674895 173114 675006 173119
rect 674895 173058 674900 173114
rect 674956 173058 675006 173114
rect 674895 173056 675006 173058
rect 674895 173053 674961 173056
rect 140802 172080 140862 172562
rect 674946 172379 675006 172494
rect 674946 172374 675057 172379
rect 674946 172318 674996 172374
rect 675052 172318 675057 172374
rect 674946 172316 675057 172318
rect 674991 172313 675057 172316
rect 145071 172080 145137 172083
rect 140802 172078 145137 172080
rect 140802 172022 145076 172078
rect 145132 172022 145137 172078
rect 140802 172020 145137 172022
rect 145071 172017 145137 172020
rect 677058 171491 677118 171754
rect 677058 171486 677169 171491
rect 677058 171430 677108 171486
rect 677164 171430 677169 171486
rect 677058 171428 677169 171430
rect 677103 171425 677169 171428
rect 144015 171340 144081 171343
rect 140832 171338 144081 171340
rect 140832 171282 144020 171338
rect 144076 171282 144081 171338
rect 140832 171280 144081 171282
rect 144015 171277 144081 171280
rect 676866 170899 676926 171014
rect 676815 170894 676926 170899
rect 676815 170838 676820 170894
rect 676876 170838 676926 170894
rect 676815 170836 676926 170838
rect 676815 170833 676881 170836
rect 145263 170156 145329 170159
rect 140832 170154 145329 170156
rect 140832 170098 145268 170154
rect 145324 170098 145329 170154
rect 140832 170096 145329 170098
rect 145263 170093 145329 170096
rect 675138 170011 675198 170200
rect 675087 170006 675198 170011
rect 675087 169950 675092 170006
rect 675148 169950 675198 170006
rect 675087 169948 675198 169950
rect 675087 169945 675153 169948
rect 674319 169416 674385 169419
rect 674319 169414 674784 169416
rect 674319 169358 674324 169414
rect 674380 169358 674784 169414
rect 674319 169356 674784 169358
rect 674319 169353 674385 169356
rect 140802 168380 140862 168868
rect 144111 168380 144177 168383
rect 140802 168378 144177 168380
rect 140802 168322 144116 168378
rect 144172 168322 144177 168378
rect 140802 168320 144177 168322
rect 144111 168317 144177 168320
rect 674511 168380 674577 168383
rect 674754 168380 674814 168572
rect 674511 168378 674814 168380
rect 674511 168322 674516 168378
rect 674572 168322 674814 168378
rect 674511 168320 674814 168322
rect 674511 168317 674577 168320
rect 144015 167640 144081 167643
rect 140832 167638 144081 167640
rect 140832 167582 144020 167638
rect 144076 167582 144081 167638
rect 140832 167580 144081 167582
rect 144015 167577 144081 167580
rect 674754 167347 674814 167758
rect 674703 167342 674814 167347
rect 674703 167286 674708 167342
rect 674764 167286 674814 167342
rect 674703 167284 674814 167286
rect 674703 167281 674769 167284
rect 646191 166900 646257 166903
rect 640224 166898 646257 166900
rect 640224 166842 646196 166898
rect 646252 166842 646257 166898
rect 640224 166840 646257 166842
rect 646191 166837 646257 166840
rect 144015 166604 144081 166607
rect 140832 166602 144081 166604
rect 140832 166546 144020 166602
rect 144076 166546 144081 166602
rect 140832 166544 144081 166546
rect 144015 166541 144081 166544
rect 674607 166604 674673 166607
rect 674754 166604 674814 166944
rect 679695 166604 679761 166607
rect 674607 166602 674814 166604
rect 674607 166546 674612 166602
rect 674668 166546 674814 166602
rect 674607 166544 674814 166546
rect 674946 166602 679761 166604
rect 674946 166546 679700 166602
rect 679756 166546 679761 166602
rect 674946 166544 679761 166546
rect 674607 166541 674673 166544
rect 645903 166456 645969 166459
rect 640224 166454 645969 166456
rect 640224 166398 645908 166454
rect 645964 166398 645969 166454
rect 640224 166396 645969 166398
rect 645903 166393 645969 166396
rect 674554 166394 674560 166458
rect 674624 166456 674630 166458
rect 674946 166456 675006 166544
rect 679695 166541 679761 166544
rect 674624 166396 675006 166456
rect 675279 166456 675345 166459
rect 679791 166456 679857 166459
rect 675279 166454 679857 166456
rect 675279 166398 675284 166454
rect 675340 166398 679796 166454
rect 679852 166398 679857 166454
rect 675279 166396 679857 166398
rect 674624 166394 674630 166396
rect 675279 166393 675345 166396
rect 679791 166393 679857 166396
rect 647919 165864 647985 165867
rect 640224 165862 647985 165864
rect 640224 165806 647924 165862
rect 647980 165806 647985 165862
rect 640224 165804 647985 165806
rect 647919 165801 647985 165804
rect 674754 165719 674814 166278
rect 674703 165714 674814 165719
rect 674703 165658 674708 165714
rect 674764 165658 674814 165714
rect 674703 165656 674814 165658
rect 674703 165653 674769 165656
rect 674362 165506 674368 165570
rect 674432 165568 674438 165570
rect 675279 165568 675345 165571
rect 674432 165566 675345 165568
rect 674432 165510 675284 165566
rect 675340 165510 675345 165566
rect 674432 165508 675345 165510
rect 674432 165506 674438 165508
rect 675279 165505 675345 165508
rect 140802 164828 140862 165316
rect 145167 164828 145233 164831
rect 140802 164826 145233 164828
rect 140802 164770 145172 164826
rect 145228 164770 145233 164826
rect 140802 164768 145233 164770
rect 145167 164765 145233 164768
rect 140802 163644 140862 164130
rect 676282 164026 676288 164090
rect 676352 164088 676358 164090
rect 676911 164088 676977 164091
rect 676352 164086 676977 164088
rect 676352 164030 676916 164086
rect 676972 164030 676977 164086
rect 676352 164028 676977 164030
rect 676352 164026 676358 164028
rect 676911 164025 676977 164028
rect 676666 163878 676672 163942
rect 676736 163940 676742 163942
rect 677199 163940 677265 163943
rect 676736 163938 677265 163940
rect 676736 163882 677204 163938
rect 677260 163882 677265 163938
rect 676736 163880 677265 163882
rect 676736 163878 676742 163880
rect 677199 163877 677265 163880
rect 144111 163644 144177 163647
rect 140802 163642 144177 163644
rect 140802 163586 144116 163642
rect 144172 163586 144177 163642
rect 140802 163584 144177 163586
rect 144111 163581 144177 163584
rect 676474 163582 676480 163646
rect 676544 163644 676550 163646
rect 677103 163644 677169 163647
rect 676544 163642 677169 163644
rect 676544 163586 677108 163642
rect 677164 163586 677169 163642
rect 676544 163584 677169 163586
rect 676544 163582 676550 163584
rect 677103 163581 677169 163584
rect 144015 162904 144081 162907
rect 140832 162902 144081 162904
rect 140832 162846 144020 162902
rect 144076 162846 144081 162902
rect 140832 162844 144081 162846
rect 144015 162841 144081 162844
rect 140802 161424 140862 161682
rect 144975 161424 145041 161427
rect 140802 161422 145041 161424
rect 140802 161366 144980 161422
rect 145036 161366 145041 161422
rect 140802 161364 145041 161366
rect 144975 161361 145041 161364
rect 210159 161276 210225 161279
rect 210682 161276 210688 161278
rect 210159 161274 210688 161276
rect 210159 161218 210164 161274
rect 210220 161218 210688 161274
rect 210159 161216 210688 161218
rect 210159 161213 210225 161216
rect 210682 161214 210688 161216
rect 210752 161214 210758 161278
rect 140802 159944 140862 160432
rect 144495 159944 144561 159947
rect 140802 159942 144561 159944
rect 140802 159886 144500 159942
rect 144556 159886 144561 159942
rect 140802 159884 144561 159886
rect 144495 159881 144561 159884
rect 144015 159352 144081 159355
rect 140832 159350 144081 159352
rect 140832 159294 144020 159350
rect 144076 159294 144081 159350
rect 140832 159292 144081 159294
rect 144015 159289 144081 159292
rect 144303 158168 144369 158171
rect 140832 158166 144369 158168
rect 140832 158110 144308 158166
rect 144364 158110 144369 158166
rect 140832 158108 144369 158110
rect 144303 158105 144369 158108
rect 146799 157280 146865 157283
rect 146754 157278 146865 157280
rect 146754 157222 146804 157278
rect 146860 157222 146865 157278
rect 146754 157217 146865 157222
rect 140802 156392 140862 156880
rect 146607 156836 146673 156839
rect 146754 156836 146814 157217
rect 146607 156834 146814 156836
rect 146607 156778 146612 156834
rect 146668 156778 146814 156834
rect 146607 156776 146814 156778
rect 146607 156773 146673 156776
rect 144207 156392 144273 156395
rect 140802 156390 144273 156392
rect 140802 156334 144212 156390
rect 144268 156334 144273 156390
rect 140802 156332 144273 156334
rect 144207 156329 144273 156332
rect 140802 155652 140862 155696
rect 144015 155652 144081 155655
rect 140802 155650 144081 155652
rect 140802 155594 144020 155650
rect 144076 155594 144081 155650
rect 140802 155592 144081 155594
rect 144015 155589 144081 155592
rect 675471 154618 675537 154619
rect 675471 154616 675520 154618
rect 675428 154614 675520 154616
rect 675428 154558 675476 154614
rect 675428 154556 675520 154558
rect 675471 154554 675520 154556
rect 675584 154554 675590 154618
rect 675471 154553 675537 154554
rect 144111 154468 144177 154471
rect 140832 154466 144177 154468
rect 140832 154410 144116 154466
rect 144172 154410 144177 154466
rect 140832 154408 144177 154410
rect 144111 154405 144177 154408
rect 210682 154258 210688 154322
rect 210752 154258 210758 154322
rect 675130 154258 675136 154322
rect 675200 154320 675206 154322
rect 675375 154320 675441 154323
rect 675200 154318 675441 154320
rect 675200 154262 675380 154318
rect 675436 154262 675441 154318
rect 675200 154260 675441 154262
rect 675200 154258 675206 154260
rect 210490 154110 210496 154174
rect 210560 154172 210566 154174
rect 210690 154172 210750 154258
rect 675375 154257 675441 154260
rect 210560 154112 210750 154172
rect 210560 154110 210566 154112
rect 675759 153432 675825 153435
rect 676282 153432 676288 153434
rect 675759 153430 676288 153432
rect 675759 153374 675764 153430
rect 675820 153374 676288 153430
rect 675759 153372 676288 153374
rect 675759 153369 675825 153372
rect 676282 153370 676288 153372
rect 676352 153370 676358 153434
rect 210159 153284 210225 153287
rect 210874 153284 210880 153286
rect 210159 153282 210880 153284
rect 140802 152988 140862 153250
rect 210159 153226 210164 153282
rect 210220 153226 210880 153282
rect 210159 153224 210880 153226
rect 210159 153221 210225 153224
rect 210874 153222 210880 153224
rect 210944 153222 210950 153286
rect 144015 152988 144081 152991
rect 140802 152986 144081 152988
rect 140802 152930 144020 152986
rect 144076 152930 144081 152986
rect 140802 152928 144081 152930
rect 144015 152925 144081 152928
rect 140802 151656 140862 152144
rect 144111 151656 144177 151659
rect 140802 151654 144177 151656
rect 140802 151598 144116 151654
rect 144172 151598 144177 151654
rect 140802 151596 144177 151598
rect 144111 151593 144177 151596
rect 144015 150916 144081 150919
rect 140832 150914 144081 150916
rect 140832 150858 144020 150914
rect 144076 150858 144081 150914
rect 140832 150856 144081 150858
rect 144015 150853 144081 150856
rect 675759 150324 675825 150327
rect 676474 150324 676480 150326
rect 675759 150322 676480 150324
rect 675759 150266 675764 150322
rect 675820 150266 676480 150322
rect 675759 150264 676480 150266
rect 675759 150261 675825 150264
rect 676474 150262 676480 150264
rect 676544 150262 676550 150326
rect 140802 149140 140862 149702
rect 144495 149140 144561 149143
rect 140802 149138 144561 149140
rect 140802 149082 144500 149138
rect 144556 149082 144561 149138
rect 140802 149080 144561 149082
rect 144495 149077 144561 149080
rect 674170 148486 674176 148550
rect 674240 148548 674246 148550
rect 675471 148548 675537 148551
rect 674240 148546 675537 148548
rect 674240 148490 675476 148546
rect 675532 148490 675537 148546
rect 674240 148488 675537 148490
rect 674240 148486 674246 148488
rect 675471 148485 675537 148488
rect 140802 147956 140862 148444
rect 144207 147956 144273 147959
rect 140802 147954 144273 147956
rect 140802 147898 144212 147954
rect 144268 147898 144273 147954
rect 140802 147896 144273 147898
rect 144207 147893 144273 147896
rect 140802 147216 140862 147260
rect 144015 147216 144081 147219
rect 140802 147214 144081 147216
rect 140802 147158 144020 147214
rect 144076 147158 144081 147214
rect 140802 147156 144081 147158
rect 144015 147153 144081 147156
rect 675759 146624 675825 146627
rect 676666 146624 676672 146626
rect 675759 146622 676672 146624
rect 675759 146566 675764 146622
rect 675820 146566 676672 146622
rect 675759 146564 676672 146566
rect 675759 146561 675825 146564
rect 676666 146562 676672 146564
rect 676736 146562 676742 146626
rect 144207 146032 144273 146035
rect 140832 146030 144273 146032
rect 140832 145974 144212 146030
rect 144268 145974 144273 146030
rect 140832 145972 144273 145974
rect 144207 145969 144273 145972
rect 140802 144256 140862 144790
rect 144879 144256 144945 144259
rect 140802 144254 144945 144256
rect 140802 144198 144884 144254
rect 144940 144198 144945 144254
rect 140802 144196 144945 144198
rect 144879 144193 144945 144196
rect 210682 144046 210688 144110
rect 210752 144046 210758 144110
rect 210490 143898 210496 143962
rect 210560 143960 210566 143962
rect 210690 143960 210750 144046
rect 210560 143900 210750 143960
rect 210560 143898 210566 143900
rect 140802 143220 140862 143708
rect 144399 143220 144465 143223
rect 140802 143218 144465 143220
rect 140802 143162 144404 143218
rect 144460 143162 144465 143218
rect 140802 143160 144465 143162
rect 144399 143157 144465 143160
rect 144207 142480 144273 142483
rect 140832 142478 144273 142480
rect 140832 142422 144212 142478
rect 144268 142422 144273 142478
rect 140832 142420 144273 142422
rect 144207 142417 144273 142420
rect 144687 141296 144753 141299
rect 140832 141294 144753 141296
rect 140832 141238 144692 141294
rect 144748 141238 144753 141294
rect 140832 141236 144753 141238
rect 144687 141233 144753 141236
rect 140802 139520 140862 140008
rect 144399 139520 144465 139523
rect 140802 139518 144465 139520
rect 140802 139462 144404 139518
rect 144460 139462 144465 139518
rect 140802 139460 144465 139462
rect 144399 139457 144465 139460
rect 674754 139079 674814 139342
rect 674703 139074 674814 139079
rect 674703 139018 674708 139074
rect 674764 139018 674814 139074
rect 674703 139016 674814 139018
rect 674703 139013 674769 139016
rect 140802 138484 140862 138824
rect 144207 138484 144273 138487
rect 140802 138482 144273 138484
rect 140802 138426 144212 138482
rect 144268 138426 144273 138482
rect 140802 138424 144273 138426
rect 144207 138421 144273 138424
rect 674415 138484 674481 138487
rect 674415 138482 674784 138484
rect 674415 138426 674420 138482
rect 674476 138426 674784 138482
rect 674415 138424 674784 138426
rect 674415 138421 674481 138424
rect 141519 137596 141585 137599
rect 140832 137594 141585 137596
rect 140832 137538 141524 137594
rect 141580 137538 141585 137594
rect 140832 137536 141585 137538
rect 141519 137533 141585 137536
rect 674607 137300 674673 137303
rect 674754 137300 674814 137640
rect 674607 137298 674814 137300
rect 674607 137242 674612 137298
rect 674668 137242 674814 137298
rect 674607 137240 674814 137242
rect 674607 137237 674673 137240
rect 673978 136794 673984 136858
rect 674048 136856 674054 136858
rect 674048 136796 674784 136856
rect 674048 136794 674054 136796
rect 140802 135968 140862 136522
rect 144687 135968 144753 135971
rect 140802 135966 144753 135968
rect 140802 135910 144692 135966
rect 144748 135910 144753 135966
rect 140802 135908 144753 135910
rect 144687 135905 144753 135908
rect 674754 135675 674814 136012
rect 674703 135670 674814 135675
rect 674703 135614 674708 135670
rect 674764 135614 674814 135670
rect 674703 135612 674814 135614
rect 674703 135609 674769 135612
rect 674554 135462 674560 135526
rect 674624 135462 674630 135526
rect 674562 135376 674622 135462
rect 674562 135316 674784 135376
rect 140802 135080 140862 135272
rect 144495 135080 144561 135083
rect 140802 135078 144561 135080
rect 140802 135022 144500 135078
rect 144556 135022 144561 135078
rect 140802 135020 144561 135022
rect 144495 135017 144561 135020
rect 673359 134932 673425 134935
rect 674554 134932 674560 134934
rect 673359 134930 674560 134932
rect 673359 134874 673364 134930
rect 673420 134874 674560 134930
rect 673359 134872 674560 134874
rect 673359 134869 673425 134872
rect 674554 134870 674560 134872
rect 674624 134870 674630 134934
rect 674362 134500 674368 134564
rect 674432 134562 674438 134564
rect 674432 134502 674784 134562
rect 674432 134500 674438 134502
rect 144399 134044 144465 134047
rect 140832 134042 144465 134044
rect 140832 133986 144404 134042
rect 144460 133986 144465 134042
rect 140832 133984 144465 133986
rect 144399 133981 144465 133984
rect 674415 133748 674481 133751
rect 674415 133746 674784 133748
rect 674415 133690 674420 133746
rect 674476 133690 674784 133746
rect 674415 133688 674784 133690
rect 674415 133685 674481 133688
rect 674170 132872 674176 132936
rect 674240 132934 674246 132936
rect 674240 132874 674784 132934
rect 674240 132872 674246 132874
rect 144207 132860 144273 132863
rect 140832 132858 144273 132860
rect 140832 132802 144212 132858
rect 144268 132802 144273 132858
rect 140832 132800 144273 132802
rect 144207 132797 144273 132800
rect 675138 131827 675198 132090
rect 675087 131822 675198 131827
rect 675087 131766 675092 131822
rect 675148 131766 675198 131822
rect 675087 131764 675198 131766
rect 675087 131761 675153 131764
rect 140802 131084 140862 131572
rect 674127 131232 674193 131235
rect 674127 131230 674784 131232
rect 674127 131174 674132 131230
rect 674188 131174 674784 131230
rect 674127 131172 674784 131174
rect 674127 131169 674193 131172
rect 144207 131084 144273 131087
rect 140802 131082 144273 131084
rect 140802 131026 144212 131082
rect 144268 131026 144273 131082
rect 140802 131024 144273 131026
rect 144207 131021 144273 131024
rect 140802 130048 140862 130388
rect 677058 130347 677118 130610
rect 677007 130342 677118 130347
rect 677007 130286 677012 130342
rect 677068 130286 677118 130342
rect 677007 130284 677118 130286
rect 677007 130281 677073 130284
rect 144207 130048 144273 130051
rect 140802 130046 144273 130048
rect 140802 129990 144212 130046
rect 144268 129990 144273 130046
rect 140802 129988 144273 129990
rect 144207 129985 144273 129988
rect 677058 129607 677118 129722
rect 677058 129602 677169 129607
rect 677058 129546 677108 129602
rect 677164 129546 677169 129602
rect 677058 129544 677169 129546
rect 677103 129541 677169 129544
rect 146511 129308 146577 129311
rect 140832 129306 146577 129308
rect 140832 129250 146516 129306
rect 146572 129250 146577 129306
rect 140832 129248 146577 129250
rect 146511 129245 146577 129248
rect 675138 128719 675198 128982
rect 675138 128714 675249 128719
rect 675138 128658 675188 128714
rect 675244 128658 675249 128714
rect 675138 128656 675249 128658
rect 675183 128653 675249 128656
rect 674223 128124 674289 128127
rect 674223 128122 674784 128124
rect 140802 127532 140862 128090
rect 674223 128066 674228 128122
rect 674284 128066 674784 128122
rect 674223 128064 674784 128066
rect 674223 128061 674289 128064
rect 146895 127532 146961 127535
rect 140802 127530 146961 127532
rect 140802 127474 146900 127530
rect 146956 127474 146961 127530
rect 140802 127472 146961 127474
rect 146895 127469 146961 127472
rect 674319 127384 674385 127387
rect 674319 127382 674784 127384
rect 674319 127326 674324 127382
rect 674380 127326 674784 127382
rect 674319 127324 674784 127326
rect 674319 127321 674385 127324
rect 146895 126940 146961 126943
rect 140832 126938 146961 126940
rect 140832 126882 146900 126938
rect 146956 126882 146961 126938
rect 140832 126880 146961 126882
rect 146895 126877 146961 126880
rect 210298 126730 210304 126794
rect 210368 126792 210374 126794
rect 210490 126792 210496 126794
rect 210368 126732 210496 126792
rect 210368 126730 210374 126732
rect 210490 126730 210496 126732
rect 210560 126730 210566 126794
rect 676866 126351 676926 126466
rect 676866 126346 676977 126351
rect 676866 126290 676916 126346
rect 676972 126290 676977 126346
rect 676866 126288 676977 126290
rect 676911 126285 676977 126288
rect 31738 125250 31744 125314
rect 31808 125312 31814 125314
rect 31808 125252 36222 125312
rect 31808 125250 31814 125252
rect 36162 124986 36222 125252
rect 140802 125164 140862 125642
rect 676866 125611 676926 125874
rect 676815 125606 676926 125611
rect 676815 125550 676820 125606
rect 676876 125550 676926 125606
rect 676815 125548 676926 125550
rect 676815 125545 676881 125548
rect 144783 125164 144849 125167
rect 140802 125162 144849 125164
rect 140802 125106 144788 125162
rect 144844 125106 144849 125162
rect 140802 125104 144849 125106
rect 144783 125101 144849 125104
rect 674946 124871 675006 124986
rect 674895 124866 675006 124871
rect 674895 124810 674900 124866
rect 674956 124810 675006 124866
rect 674895 124808 675006 124810
rect 674895 124805 674961 124808
rect 144591 124424 144657 124427
rect 140832 124422 144657 124424
rect 140832 124366 144596 124422
rect 144652 124366 144657 124422
rect 140832 124364 144657 124366
rect 144591 124361 144657 124364
rect 674511 123980 674577 123983
rect 674754 123980 674814 124246
rect 674511 123978 674814 123980
rect 674511 123922 674516 123978
rect 674572 123922 674814 123978
rect 674511 123920 674814 123922
rect 674511 123917 674577 123920
rect 674031 123388 674097 123391
rect 674031 123386 674784 123388
rect 674031 123330 674036 123386
rect 674092 123330 674784 123386
rect 674031 123328 674784 123330
rect 674031 123325 674097 123328
rect 140802 122648 140862 123136
rect 144783 122648 144849 122651
rect 140802 122646 144849 122648
rect 140802 122590 144788 122646
rect 144844 122590 144849 122646
rect 140802 122588 144849 122590
rect 144783 122585 144849 122588
rect 674754 122207 674814 122544
rect 674754 122202 674865 122207
rect 674754 122146 674804 122202
rect 674860 122146 674865 122202
rect 674754 122144 674865 122146
rect 674799 122141 674865 122144
rect 140802 121612 140862 121952
rect 647823 121760 647889 121763
rect 640224 121758 647889 121760
rect 640224 121702 647828 121758
rect 647884 121702 647889 121758
rect 640224 121700 647889 121702
rect 647823 121697 647889 121700
rect 144591 121612 144657 121615
rect 140802 121610 144657 121612
rect 140802 121554 144596 121610
rect 144652 121554 144657 121610
rect 140802 121552 144657 121554
rect 144591 121549 144657 121552
rect 674607 121612 674673 121615
rect 674754 121612 674814 121730
rect 674607 121610 674814 121612
rect 674607 121554 674612 121610
rect 674668 121554 674814 121610
rect 674607 121552 674814 121554
rect 674607 121549 674673 121552
rect 674703 121316 674769 121319
rect 674703 121314 674814 121316
rect 674703 121258 674708 121314
rect 674764 121258 674814 121314
rect 674703 121253 674814 121258
rect 640194 121168 640254 121212
rect 647919 121168 647985 121171
rect 640194 121166 647985 121168
rect 640194 121110 647924 121166
rect 647980 121110 647985 121166
rect 640194 121108 647985 121110
rect 647919 121105 647985 121108
rect 674754 121064 674814 121253
rect 141519 121020 141585 121023
rect 144399 121020 144465 121023
rect 141519 121018 144465 121020
rect 141519 120962 141524 121018
rect 141580 120962 144404 121018
rect 144460 120962 144465 121018
rect 141519 120960 144465 120962
rect 141519 120957 141585 120960
rect 144399 120957 144465 120960
rect 144591 120872 144657 120875
rect 140832 120870 144657 120872
rect 140832 120814 144596 120870
rect 144652 120814 144657 120870
rect 140832 120812 144657 120814
rect 144591 120809 144657 120812
rect 647823 120724 647889 120727
rect 640224 120722 647889 120724
rect 640224 120666 647828 120722
rect 647884 120666 647889 120722
rect 640224 120664 647889 120666
rect 647823 120661 647889 120664
rect 675706 120366 675712 120430
rect 675776 120428 675782 120430
rect 677007 120428 677073 120431
rect 675776 120426 677073 120428
rect 675776 120370 677012 120426
rect 677068 120370 677073 120426
rect 675776 120368 677073 120370
rect 675776 120366 675782 120368
rect 677007 120365 677073 120368
rect 646479 120132 646545 120135
rect 640224 120130 646545 120132
rect 640224 120074 646484 120130
rect 646540 120074 646545 120130
rect 640224 120072 646545 120074
rect 646479 120069 646545 120072
rect 140802 119096 140862 119630
rect 144783 119096 144849 119099
rect 140802 119094 144849 119096
rect 140802 119038 144788 119094
rect 144844 119038 144849 119094
rect 140802 119036 144849 119038
rect 144783 119033 144849 119036
rect 141039 118652 141105 118655
rect 140610 118650 141105 118652
rect 140610 118594 141044 118650
rect 141100 118594 141105 118650
rect 140610 118592 141105 118594
rect 140610 118474 140670 118592
rect 141039 118589 141105 118592
rect 141039 118356 141105 118359
rect 144591 118356 144657 118359
rect 141039 118354 144657 118356
rect 141039 118298 141044 118354
rect 141100 118298 144596 118354
rect 144652 118298 144657 118354
rect 141039 118296 144657 118298
rect 141039 118293 141105 118296
rect 144591 118293 144657 118296
rect 676666 117998 676672 118062
rect 676736 118060 676742 118062
rect 677103 118060 677169 118063
rect 676736 118058 677169 118060
rect 676736 118002 677108 118058
rect 677164 118002 677169 118058
rect 676736 118000 677169 118002
rect 676736 117998 676742 118000
rect 677103 117997 677169 118000
rect 140802 116728 140862 117210
rect 144591 116728 144657 116731
rect 140802 116726 144657 116728
rect 140802 116670 144596 116726
rect 144652 116670 144657 116726
rect 140802 116668 144657 116670
rect 144591 116665 144657 116668
rect 140802 115396 140862 115958
rect 146703 115396 146769 115399
rect 140802 115394 146769 115396
rect 140802 115338 146708 115394
rect 146764 115338 146769 115394
rect 140802 115336 146769 115338
rect 146703 115333 146769 115336
rect 146703 115248 146769 115251
rect 147087 115248 147153 115251
rect 146703 115246 147153 115248
rect 146703 115190 146708 115246
rect 146764 115190 147092 115246
rect 147148 115190 147153 115246
rect 146703 115188 147153 115190
rect 146703 115185 146769 115188
rect 147087 115185 147153 115188
rect 140802 114212 140862 114762
rect 144591 114212 144657 114215
rect 140802 114210 144657 114212
rect 140802 114154 144596 114210
rect 144652 114154 144657 114210
rect 140802 114152 144657 114154
rect 144591 114149 144657 114152
rect 140802 113176 140862 113664
rect 144783 113176 144849 113179
rect 140802 113174 144849 113176
rect 140802 113118 144788 113174
rect 144844 113118 144849 113174
rect 140802 113116 144849 113118
rect 144783 113113 144849 113116
rect 665199 112880 665265 112883
rect 665154 112878 665265 112880
rect 665154 112822 665204 112878
rect 665260 112822 665265 112878
rect 665154 112817 665265 112822
rect 144591 112436 144657 112439
rect 140832 112434 144657 112436
rect 140832 112378 144596 112434
rect 144652 112378 144657 112434
rect 665154 112424 665214 112817
rect 140832 112376 144657 112378
rect 144591 112373 144657 112376
rect 665154 111551 665214 112059
rect 665154 111546 665265 111551
rect 665154 111490 665204 111546
rect 665260 111490 665265 111546
rect 665154 111488 665265 111490
rect 665199 111485 665265 111488
rect 674746 111400 674752 111402
rect 665442 111340 674752 111400
rect 665442 111337 665502 111340
rect 674746 111338 674752 111340
rect 674816 111338 674822 111402
rect 144783 111252 144849 111255
rect 140832 111250 144849 111252
rect 140832 111194 144788 111250
rect 144844 111194 144849 111250
rect 140832 111192 144849 111194
rect 144783 111189 144849 111192
rect 675471 110070 675537 110071
rect 675471 110066 675520 110070
rect 675584 110068 675590 110070
rect 675471 110010 675476 110066
rect 675471 110006 675520 110010
rect 675584 110008 675628 110068
rect 675584 110006 675590 110008
rect 675471 110005 675537 110006
rect 140802 109772 140862 109964
rect 144591 109772 144657 109775
rect 140802 109770 144657 109772
rect 140802 109714 144596 109770
rect 144652 109714 144657 109770
rect 140802 109712 144657 109714
rect 144591 109709 144657 109712
rect 674746 109414 674752 109478
rect 674816 109476 674822 109478
rect 675375 109476 675441 109479
rect 674816 109474 675441 109476
rect 674816 109418 675380 109474
rect 675436 109418 675441 109474
rect 674816 109416 675441 109418
rect 674816 109414 674822 109416
rect 675375 109413 675441 109416
rect 140802 108292 140862 108778
rect 146031 108292 146097 108295
rect 140802 108290 146097 108292
rect 140802 108234 146036 108290
rect 146092 108234 146097 108290
rect 140802 108232 146097 108234
rect 146031 108229 146097 108232
rect 675663 108146 675729 108147
rect 675663 108142 675712 108146
rect 675776 108144 675782 108146
rect 675663 108086 675668 108142
rect 675663 108082 675712 108086
rect 675776 108084 675820 108144
rect 675776 108082 675782 108084
rect 675663 108081 675729 108082
rect 144591 107552 144657 107555
rect 140832 107550 144657 107552
rect 140832 107494 144596 107550
rect 144652 107494 144657 107550
rect 140832 107492 144657 107494
rect 144591 107489 144657 107492
rect 144687 106664 144753 106667
rect 144826 106664 144832 106666
rect 144687 106662 144832 106664
rect 144687 106606 144692 106662
rect 144748 106606 144832 106662
rect 144687 106604 144832 106606
rect 144687 106601 144753 106604
rect 144826 106602 144832 106604
rect 144896 106602 144902 106666
rect 144303 106516 144369 106519
rect 144303 106514 144510 106516
rect 144303 106458 144308 106514
rect 144364 106458 144510 106514
rect 144303 106456 144510 106458
rect 144303 106453 144369 106456
rect 140802 105924 140862 106412
rect 144450 106368 144510 106456
rect 144591 106368 144657 106371
rect 144450 106366 144657 106368
rect 144450 106310 144596 106366
rect 144652 106310 144657 106366
rect 144450 106308 144657 106310
rect 144591 106305 144657 106308
rect 144111 105924 144177 105927
rect 140802 105922 144177 105924
rect 140802 105866 144116 105922
rect 144172 105866 144177 105922
rect 140802 105864 144177 105866
rect 144111 105861 144177 105864
rect 140802 104888 140862 105228
rect 209914 105122 209920 105186
rect 209984 105184 209990 105186
rect 210298 105184 210304 105186
rect 209984 105124 210304 105184
rect 209984 105122 209990 105124
rect 210298 105122 210304 105124
rect 210368 105122 210374 105186
rect 144015 104888 144081 104891
rect 140802 104886 144081 104888
rect 140802 104830 144020 104886
rect 144076 104830 144081 104886
rect 140802 104828 144081 104830
rect 144015 104825 144081 104828
rect 647919 104444 647985 104447
rect 640224 104442 647985 104444
rect 640224 104386 647924 104442
rect 647980 104386 647985 104442
rect 640224 104384 647985 104386
rect 647919 104381 647985 104384
rect 144015 104000 144081 104003
rect 140832 103998 144081 104000
rect 140832 103942 144020 103998
rect 144076 103942 144081 103998
rect 140832 103940 144081 103942
rect 144015 103937 144081 103940
rect 210106 103494 210112 103558
rect 210176 103556 210182 103558
rect 210874 103556 210880 103558
rect 210176 103496 210880 103556
rect 210176 103494 210182 103496
rect 210874 103494 210880 103496
rect 210944 103494 210950 103558
rect 674170 103198 674176 103262
rect 674240 103260 674246 103262
rect 675375 103260 675441 103263
rect 674240 103258 675441 103260
rect 674240 103202 675380 103258
rect 675436 103202 675441 103258
rect 674240 103200 675441 103202
rect 674240 103198 674246 103200
rect 675375 103197 675441 103200
rect 144111 102816 144177 102819
rect 140832 102814 144177 102816
rect 140832 102758 144116 102814
rect 144172 102758 144177 102814
rect 140832 102756 144177 102758
rect 144111 102753 144177 102756
rect 210490 102310 210496 102374
rect 210560 102372 210566 102374
rect 210874 102372 210880 102374
rect 210560 102312 210880 102372
rect 210560 102310 210566 102312
rect 210874 102310 210880 102312
rect 210944 102310 210950 102374
rect 199983 102224 200049 102227
rect 199983 102222 210528 102224
rect 199983 102166 199988 102222
rect 200044 102166 210528 102222
rect 199983 102164 210528 102166
rect 199983 102161 200049 102164
rect 201711 101632 201777 101635
rect 201711 101630 210528 101632
rect 201711 101574 201716 101630
rect 201772 101574 210528 101630
rect 201711 101572 210528 101574
rect 201711 101569 201777 101572
rect 140802 101336 140862 101528
rect 675759 101484 675825 101487
rect 676666 101484 676672 101486
rect 675759 101482 676672 101484
rect 675759 101426 675764 101482
rect 675820 101426 676672 101482
rect 675759 101424 676672 101426
rect 675759 101421 675825 101424
rect 676666 101422 676672 101424
rect 676736 101422 676742 101486
rect 144015 101336 144081 101339
rect 140802 101334 144081 101336
rect 140802 101278 144020 101334
rect 144076 101278 144081 101334
rect 140802 101276 144081 101278
rect 144015 101273 144081 101276
rect 210159 101114 210225 101117
rect 210159 101112 210528 101114
rect 210159 101056 210164 101112
rect 210220 101056 210528 101112
rect 210159 101054 210528 101056
rect 210159 101051 210225 101054
rect 144687 100892 144753 100895
rect 144826 100892 144832 100894
rect 144687 100890 144832 100892
rect 144687 100834 144692 100890
rect 144748 100834 144832 100890
rect 144687 100832 144832 100834
rect 144687 100829 144753 100832
rect 144826 100830 144832 100832
rect 144896 100830 144902 100894
rect 201711 100596 201777 100599
rect 201711 100594 210528 100596
rect 201711 100538 201716 100594
rect 201772 100538 210528 100594
rect 201711 100536 210528 100538
rect 201711 100533 201777 100536
rect 140802 99856 140862 100344
rect 201711 100004 201777 100007
rect 201711 100002 210528 100004
rect 201711 99946 201716 100002
rect 201772 99946 210528 100002
rect 201711 99944 210528 99946
rect 201711 99941 201777 99944
rect 144015 99856 144081 99859
rect 140802 99854 144081 99856
rect 140802 99798 144020 99854
rect 144076 99798 144081 99854
rect 140802 99796 144081 99798
rect 144015 99793 144081 99796
rect 210159 99486 210225 99489
rect 210159 99484 210528 99486
rect 210159 99428 210164 99484
rect 210220 99428 210528 99484
rect 210159 99426 210528 99428
rect 210159 99423 210225 99426
rect 144111 99116 144177 99119
rect 140832 99114 144177 99116
rect 140832 99058 144116 99114
rect 144172 99058 144177 99114
rect 140832 99056 144177 99058
rect 144111 99053 144177 99056
rect 201615 98968 201681 98971
rect 201615 98966 210528 98968
rect 201615 98910 201620 98966
rect 201676 98910 210528 98966
rect 201615 98908 210528 98910
rect 201615 98905 201681 98908
rect 201807 98376 201873 98379
rect 201807 98374 210528 98376
rect 201807 98318 201812 98374
rect 201868 98318 210528 98374
rect 201807 98316 210528 98318
rect 201807 98313 201873 98316
rect 144015 98080 144081 98083
rect 140832 98078 144081 98080
rect 140832 98022 144020 98078
rect 144076 98022 144081 98078
rect 140832 98020 144081 98022
rect 144015 98017 144081 98020
rect 210159 97858 210225 97861
rect 210159 97856 210528 97858
rect 210159 97800 210164 97856
rect 210220 97800 210528 97856
rect 210159 97798 210528 97800
rect 210159 97795 210225 97798
rect 202959 97340 203025 97343
rect 202959 97338 210528 97340
rect 202959 97282 202964 97338
rect 203020 97282 210528 97338
rect 202959 97280 210528 97282
rect 202959 97277 203025 97280
rect 140802 96304 140862 96792
rect 201711 96748 201777 96751
rect 201711 96746 210528 96748
rect 201711 96690 201716 96746
rect 201772 96690 210528 96746
rect 201711 96688 210528 96690
rect 201711 96685 201777 96688
rect 144015 96304 144081 96307
rect 140802 96302 144081 96304
rect 140802 96246 144020 96302
rect 144076 96246 144081 96302
rect 140802 96244 144081 96246
rect 144015 96241 144081 96244
rect 210159 96230 210225 96233
rect 210159 96228 210528 96230
rect 210159 96172 210164 96228
rect 210220 96172 210528 96228
rect 210159 96170 210528 96172
rect 210159 96167 210225 96170
rect 201615 95712 201681 95715
rect 201615 95710 210528 95712
rect 201615 95654 201620 95710
rect 201676 95654 210528 95710
rect 201615 95652 210528 95654
rect 201615 95649 201681 95652
rect 146511 95564 146577 95567
rect 140832 95562 146577 95564
rect 140832 95506 146516 95562
rect 146572 95506 146577 95562
rect 140832 95504 146577 95506
rect 146511 95501 146577 95504
rect 201807 95120 201873 95123
rect 201807 95118 210528 95120
rect 201807 95062 201812 95118
rect 201868 95062 210528 95118
rect 201807 95060 210528 95062
rect 201807 95057 201873 95060
rect 209722 94762 209728 94826
rect 209792 94824 209798 94826
rect 210874 94824 210880 94826
rect 209792 94764 210880 94824
rect 209792 94762 209798 94764
rect 210874 94762 210880 94764
rect 210944 94762 210950 94826
rect 210159 94602 210225 94605
rect 210159 94600 210528 94602
rect 210159 94544 210164 94600
rect 210220 94544 210528 94600
rect 210159 94542 210528 94544
rect 210159 94539 210225 94542
rect 144111 94380 144177 94383
rect 140832 94378 144177 94380
rect 140832 94322 144116 94378
rect 144172 94322 144177 94378
rect 140832 94320 144177 94322
rect 144111 94317 144177 94320
rect 201711 94084 201777 94087
rect 201711 94082 210528 94084
rect 201711 94026 201716 94082
rect 201772 94026 210528 94082
rect 201711 94024 210528 94026
rect 201711 94021 201777 94024
rect 210490 93726 210496 93790
rect 210560 93788 210566 93790
rect 210874 93788 210880 93790
rect 210560 93728 210880 93788
rect 210560 93726 210566 93728
rect 210874 93726 210880 93728
rect 210944 93726 210950 93790
rect 200175 93492 200241 93495
rect 200175 93490 210528 93492
rect 200175 93434 200180 93490
rect 200236 93434 210528 93490
rect 200175 93432 210528 93434
rect 200175 93429 200241 93432
rect 197295 93344 197361 93347
rect 197295 93342 210558 93344
rect 197295 93286 197300 93342
rect 197356 93286 210558 93342
rect 197295 93284 210558 93286
rect 197295 93281 197361 93284
rect 140802 92752 140862 93092
rect 210498 92944 210558 93284
rect 144015 92752 144081 92755
rect 140802 92750 144081 92752
rect 140802 92694 144020 92750
rect 144076 92694 144081 92750
rect 140802 92692 144081 92694
rect 144015 92689 144081 92692
rect 201615 92456 201681 92459
rect 201615 92454 210528 92456
rect 201615 92398 201620 92454
rect 201676 92398 210528 92454
rect 201615 92396 210528 92398
rect 201615 92393 201681 92396
rect 140802 91420 140862 91908
rect 201711 91864 201777 91867
rect 201711 91862 210528 91864
rect 201711 91806 201716 91862
rect 201772 91806 210528 91862
rect 201711 91804 210528 91806
rect 201711 91801 201777 91804
rect 197679 91716 197745 91719
rect 197679 91714 210558 91716
rect 197679 91658 197684 91714
rect 197740 91658 210558 91714
rect 197679 91656 210558 91658
rect 197679 91653 197745 91656
rect 146223 91420 146289 91423
rect 140802 91418 146289 91420
rect 140802 91362 146228 91418
rect 146284 91362 146289 91418
rect 140802 91360 146289 91362
rect 146223 91357 146289 91360
rect 210498 91316 210558 91656
rect 144111 90828 144177 90831
rect 140832 90826 144177 90828
rect 140832 90770 144116 90826
rect 144172 90770 144177 90826
rect 140832 90768 144177 90770
rect 144111 90765 144177 90768
rect 194415 90828 194481 90831
rect 194415 90826 210528 90828
rect 194415 90770 194420 90826
rect 194476 90770 210528 90826
rect 194415 90768 210528 90770
rect 194415 90765 194481 90768
rect 201615 90236 201681 90239
rect 201615 90234 210528 90236
rect 201615 90178 201620 90234
rect 201676 90178 210528 90234
rect 201615 90176 210528 90178
rect 201615 90173 201681 90176
rect 144015 89644 144081 89647
rect 140832 89642 144081 89644
rect 140832 89586 144020 89642
rect 144076 89586 144081 89642
rect 140832 89584 144081 89586
rect 144015 89581 144081 89584
rect 201807 89644 201873 89647
rect 201807 89642 210528 89644
rect 201807 89586 201812 89642
rect 201868 89586 210528 89642
rect 201807 89584 210528 89586
rect 201807 89581 201873 89584
rect 201711 89200 201777 89203
rect 647631 89200 647697 89203
rect 201711 89198 210528 89200
rect 201711 89142 201716 89198
rect 201772 89142 210528 89198
rect 201711 89140 210528 89142
rect 640224 89198 647697 89200
rect 640224 89142 647636 89198
rect 647692 89142 647697 89198
rect 640224 89140 647697 89142
rect 201711 89137 201777 89140
rect 647631 89137 647697 89140
rect 198735 88608 198801 88611
rect 646287 88608 646353 88611
rect 198735 88606 210528 88608
rect 198735 88550 198740 88606
rect 198796 88550 210528 88606
rect 198735 88548 210528 88550
rect 640224 88606 646353 88608
rect 640224 88550 646292 88606
rect 646348 88550 646353 88606
rect 640224 88548 646353 88550
rect 198735 88545 198801 88548
rect 646287 88545 646353 88548
rect 140802 87868 140862 88356
rect 201519 88016 201585 88019
rect 647919 88016 647985 88019
rect 201519 88014 210528 88016
rect 201519 87958 201524 88014
rect 201580 87958 210528 88014
rect 201519 87956 210528 87958
rect 640224 88014 647985 88016
rect 640224 87958 647924 88014
rect 647980 87958 647985 88014
rect 640224 87956 647985 87958
rect 201519 87953 201585 87956
rect 647919 87953 647985 87956
rect 144015 87868 144081 87871
rect 140802 87866 144081 87868
rect 140802 87810 144020 87866
rect 144076 87810 144081 87866
rect 140802 87808 144081 87810
rect 144015 87805 144081 87808
rect 210106 87806 210112 87870
rect 210176 87868 210182 87870
rect 210874 87868 210880 87870
rect 210176 87808 210880 87868
rect 210176 87806 210182 87808
rect 210874 87806 210880 87808
rect 210944 87806 210950 87870
rect 210159 87720 210225 87723
rect 210682 87720 210688 87722
rect 210159 87718 210688 87720
rect 210159 87662 210164 87718
rect 210220 87662 210688 87718
rect 210159 87660 210688 87662
rect 210159 87657 210225 87660
rect 210682 87658 210688 87660
rect 210752 87658 210758 87722
rect 201615 87572 201681 87575
rect 647439 87572 647505 87575
rect 201615 87570 210528 87572
rect 201615 87514 201620 87570
rect 201676 87514 210528 87570
rect 201615 87512 210528 87514
rect 640224 87570 647505 87572
rect 640224 87514 647444 87570
rect 647500 87514 647505 87570
rect 640224 87512 647505 87514
rect 201615 87509 201681 87512
rect 647439 87509 647505 87512
rect 144783 87128 144849 87131
rect 140832 87126 144849 87128
rect 140832 87070 144788 87126
rect 144844 87070 144849 87126
rect 140832 87068 144849 87070
rect 144783 87065 144849 87068
rect 201807 86980 201873 86983
rect 646383 86980 646449 86983
rect 201807 86978 210528 86980
rect 201807 86922 201812 86978
rect 201868 86922 210528 86978
rect 201807 86920 210528 86922
rect 640224 86978 646449 86980
rect 640224 86922 646388 86978
rect 646444 86922 646449 86978
rect 640224 86920 646449 86922
rect 201807 86917 201873 86920
rect 646383 86917 646449 86920
rect 650895 86980 650961 86983
rect 650895 86978 656736 86980
rect 650895 86922 650900 86978
rect 650956 86922 656736 86978
rect 650895 86920 656736 86922
rect 650895 86917 650961 86920
rect 201711 86388 201777 86391
rect 646095 86388 646161 86391
rect 201711 86386 210528 86388
rect 201711 86330 201716 86386
rect 201772 86330 210528 86386
rect 201711 86328 210528 86330
rect 640224 86386 646161 86388
rect 640224 86330 646100 86386
rect 646156 86330 646161 86386
rect 640224 86328 646161 86330
rect 201711 86325 201777 86328
rect 646095 86325 646161 86328
rect 651183 86240 651249 86243
rect 651183 86238 656736 86240
rect 651183 86182 651188 86238
rect 651244 86182 656736 86238
rect 651183 86180 656736 86182
rect 651183 86177 651249 86180
rect 209914 86030 209920 86094
rect 209984 86092 209990 86094
rect 210874 86092 210880 86094
rect 209984 86032 210880 86092
rect 209984 86030 209990 86032
rect 210874 86030 210880 86032
rect 210944 86030 210950 86094
rect 144015 85944 144081 85947
rect 140832 85942 144081 85944
rect 140832 85886 144020 85942
rect 144076 85886 144081 85942
rect 140832 85884 144081 85886
rect 144015 85881 144081 85884
rect 201711 85944 201777 85947
rect 647247 85944 647313 85947
rect 201711 85942 210528 85944
rect 201711 85886 201716 85942
rect 201772 85886 210528 85942
rect 201711 85884 210528 85886
rect 640224 85942 647313 85944
rect 640224 85886 647252 85942
rect 647308 85886 647313 85942
rect 640224 85884 647313 85886
rect 201711 85881 201777 85884
rect 647247 85881 647313 85884
rect 663618 85651 663678 86210
rect 663567 85646 663678 85651
rect 663567 85590 663572 85646
rect 663628 85590 663678 85646
rect 663567 85588 663678 85590
rect 663567 85585 663633 85588
rect 201615 85352 201681 85355
rect 647823 85352 647889 85355
rect 201615 85350 210528 85352
rect 201615 85294 201620 85350
rect 201676 85294 210528 85350
rect 201615 85292 210528 85294
rect 640224 85350 647889 85352
rect 640224 85294 647828 85350
rect 647884 85294 647889 85350
rect 640224 85292 647889 85294
rect 201615 85289 201681 85292
rect 647823 85289 647889 85292
rect 650991 85352 651057 85355
rect 650991 85350 656736 85352
rect 650991 85294 650996 85350
rect 651052 85294 656736 85350
rect 650991 85292 656736 85294
rect 650991 85289 651057 85292
rect 663279 85204 663345 85207
rect 663234 85202 663345 85204
rect 663234 85146 663284 85202
rect 663340 85146 663345 85202
rect 663234 85141 663345 85146
rect 201807 84760 201873 84763
rect 646479 84760 646545 84763
rect 201807 84758 210528 84760
rect 201807 84702 201812 84758
rect 201868 84702 210528 84758
rect 201807 84700 210528 84702
rect 640224 84758 646545 84760
rect 640224 84702 646484 84758
rect 646540 84702 646545 84758
rect 640224 84700 646545 84702
rect 201807 84697 201873 84700
rect 646479 84697 646545 84700
rect 140802 84168 140862 84656
rect 210106 84550 210112 84614
rect 210176 84612 210182 84614
rect 210682 84612 210688 84614
rect 210176 84552 210688 84612
rect 210176 84550 210182 84552
rect 210682 84550 210688 84552
rect 210752 84550 210758 84614
rect 663234 84582 663294 85141
rect 663426 84763 663486 85322
rect 663426 84758 663537 84763
rect 663426 84702 663476 84758
rect 663532 84702 663537 84758
rect 663426 84700 663537 84702
rect 663471 84697 663537 84700
rect 201519 84316 201585 84319
rect 645999 84316 646065 84319
rect 201519 84314 210528 84316
rect 201519 84258 201524 84314
rect 201580 84258 210528 84314
rect 201519 84256 210528 84258
rect 640224 84314 646065 84316
rect 640224 84258 646004 84314
rect 646060 84258 646065 84314
rect 640224 84256 646065 84258
rect 201519 84253 201585 84256
rect 645999 84253 646065 84256
rect 650991 84316 651057 84319
rect 650991 84314 656736 84316
rect 650991 84258 650996 84314
rect 651052 84258 656736 84314
rect 650991 84256 656736 84258
rect 650991 84253 651057 84256
rect 146511 84168 146577 84171
rect 140802 84166 146577 84168
rect 140802 84110 146516 84166
rect 146572 84110 146577 84166
rect 140802 84108 146577 84110
rect 146511 84105 146577 84108
rect 201903 83724 201969 83727
rect 652335 83724 652401 83727
rect 201903 83722 210528 83724
rect 201903 83666 201908 83722
rect 201964 83666 210528 83722
rect 201903 83664 210528 83666
rect 640224 83722 652401 83724
rect 640224 83666 652340 83722
rect 652396 83666 652401 83722
rect 640224 83664 652401 83666
rect 201903 83661 201969 83664
rect 652335 83661 652401 83664
rect 140802 83576 140862 83618
rect 145935 83576 146001 83579
rect 140802 83574 146001 83576
rect 140802 83518 145940 83574
rect 145996 83518 146001 83574
rect 140802 83516 146001 83518
rect 145935 83513 146001 83516
rect 210255 83430 210321 83431
rect 210255 83428 210304 83430
rect 210212 83426 210304 83428
rect 210212 83370 210260 83426
rect 210212 83368 210304 83370
rect 210255 83366 210304 83368
rect 210368 83366 210374 83430
rect 651087 83428 651153 83431
rect 651087 83426 656736 83428
rect 651087 83370 651092 83426
rect 651148 83370 656736 83426
rect 651087 83368 656736 83370
rect 210255 83365 210321 83366
rect 651087 83365 651153 83368
rect 201039 83132 201105 83135
rect 646287 83132 646353 83135
rect 201039 83130 210528 83132
rect 201039 83074 201044 83130
rect 201100 83074 210528 83130
rect 201039 83072 210528 83074
rect 640224 83130 646353 83132
rect 640224 83074 646292 83130
rect 646348 83074 646353 83130
rect 640224 83072 646353 83074
rect 201039 83069 201105 83072
rect 646287 83069 646353 83072
rect 663426 82839 663486 83398
rect 663375 82834 663486 82839
rect 663375 82778 663380 82834
rect 663436 82778 663486 82834
rect 663375 82776 663486 82778
rect 663375 82773 663441 82776
rect 201711 82688 201777 82691
rect 646095 82688 646161 82691
rect 201711 82686 210528 82688
rect 201711 82630 201716 82686
rect 201772 82630 210528 82686
rect 201711 82628 210528 82630
rect 640224 82686 646161 82688
rect 640224 82630 646100 82686
rect 646156 82630 646161 82686
rect 640224 82628 646161 82630
rect 201711 82625 201777 82628
rect 646095 82625 646161 82628
rect 650895 82688 650961 82691
rect 650895 82686 656736 82688
rect 650895 82630 650900 82686
rect 650956 82630 656736 82686
rect 650895 82628 656736 82630
rect 650895 82625 650961 82628
rect 144015 82392 144081 82395
rect 140832 82390 144081 82392
rect 140832 82334 144020 82390
rect 144076 82334 144081 82390
rect 140832 82332 144081 82334
rect 144015 82329 144081 82332
rect 209722 82330 209728 82394
rect 209792 82392 209798 82394
rect 210874 82392 210880 82394
rect 209792 82332 210880 82392
rect 209792 82330 209798 82332
rect 210874 82330 210880 82332
rect 210944 82330 210950 82394
rect 663234 82099 663294 82658
rect 197775 82096 197841 82099
rect 647535 82096 647601 82099
rect 197775 82094 210528 82096
rect 197775 82038 197780 82094
rect 197836 82038 210528 82094
rect 197775 82036 210528 82038
rect 640224 82094 647601 82096
rect 640224 82038 647540 82094
rect 647596 82038 647601 82094
rect 640224 82036 647601 82038
rect 663234 82094 663345 82099
rect 663234 82038 663284 82094
rect 663340 82038 663345 82094
rect 663234 82036 663345 82038
rect 197775 82033 197841 82036
rect 647535 82033 647601 82036
rect 663279 82033 663345 82036
rect 201615 81504 201681 81507
rect 647919 81504 647985 81507
rect 201615 81502 210528 81504
rect 201615 81446 201620 81502
rect 201676 81446 210528 81502
rect 201615 81444 210528 81446
rect 640224 81502 647985 81504
rect 640224 81446 647924 81502
rect 647980 81446 647985 81502
rect 640224 81444 647985 81446
rect 201615 81441 201681 81444
rect 647919 81441 647985 81444
rect 194607 81356 194673 81359
rect 647343 81356 647409 81359
rect 194607 81354 210558 81356
rect 194607 81298 194612 81354
rect 194668 81298 210558 81354
rect 194607 81296 210558 81298
rect 194607 81293 194673 81296
rect 144015 81208 144081 81211
rect 140832 81206 144081 81208
rect 140832 81150 144020 81206
rect 144076 81150 144081 81206
rect 140832 81148 144081 81150
rect 144015 81145 144081 81148
rect 210498 80956 210558 81296
rect 640194 81354 647409 81356
rect 640194 81298 647348 81354
rect 647404 81298 647409 81354
rect 640194 81296 647409 81298
rect 640194 80956 640254 81296
rect 647343 81293 647409 81296
rect 662895 81208 662961 81211
rect 663042 81208 663102 81770
rect 662895 81206 663102 81208
rect 662895 81150 662900 81206
rect 662956 81150 663102 81206
rect 662895 81148 663102 81150
rect 662895 81145 662961 81148
rect 200271 80468 200337 80471
rect 647919 80468 647985 80471
rect 200271 80466 210528 80468
rect 200271 80410 200276 80466
rect 200332 80410 210528 80466
rect 200271 80408 210528 80410
rect 640224 80466 647985 80468
rect 640224 80410 647924 80466
rect 647980 80410 647985 80466
rect 640224 80408 647985 80410
rect 200271 80405 200337 80408
rect 647919 80405 647985 80408
rect 140802 79432 140862 79920
rect 197391 79876 197457 79879
rect 646863 79876 646929 79879
rect 197391 79874 210528 79876
rect 197391 79818 197396 79874
rect 197452 79818 210528 79874
rect 197391 79816 210528 79818
rect 640224 79874 646929 79876
rect 640224 79818 646868 79874
rect 646924 79818 646929 79874
rect 640224 79816 646929 79818
rect 197391 79813 197457 79816
rect 646863 79813 646929 79816
rect 194511 79728 194577 79731
rect 194511 79726 210558 79728
rect 194511 79670 194516 79726
rect 194572 79670 210558 79726
rect 194511 79668 210558 79670
rect 194511 79665 194577 79668
rect 144111 79432 144177 79435
rect 140802 79430 144177 79432
rect 140802 79374 144116 79430
rect 144172 79374 144177 79430
rect 140802 79372 144177 79374
rect 144111 79369 144177 79372
rect 210498 79328 210558 79668
rect 640194 78988 640254 79328
rect 646479 78988 646545 78991
rect 640194 78986 646545 78988
rect 640194 78930 646484 78986
rect 646540 78930 646545 78986
rect 640194 78928 646545 78930
rect 646479 78925 646545 78928
rect 200367 78840 200433 78843
rect 646863 78840 646929 78843
rect 200367 78838 210528 78840
rect 200367 78782 200372 78838
rect 200428 78782 210528 78838
rect 200367 78780 210528 78782
rect 640224 78838 646929 78840
rect 640224 78782 646868 78838
rect 646924 78782 646929 78838
rect 640224 78780 646929 78782
rect 200367 78777 200433 78780
rect 646863 78777 646929 78780
rect 144015 78692 144081 78695
rect 140832 78690 144081 78692
rect 140832 78634 144020 78690
rect 144076 78634 144081 78690
rect 140832 78632 144081 78634
rect 144015 78629 144081 78632
rect 201711 78248 201777 78251
rect 646863 78248 646929 78251
rect 201711 78246 210528 78248
rect 201711 78190 201716 78246
rect 201772 78190 210528 78246
rect 201711 78188 210528 78190
rect 640224 78246 646929 78248
rect 640224 78190 646868 78246
rect 646924 78190 646929 78246
rect 640224 78188 646929 78190
rect 201711 78185 201777 78188
rect 646863 78185 646929 78188
rect 210255 77730 210321 77733
rect 210255 77728 210528 77730
rect 210255 77672 210260 77728
rect 210316 77672 210528 77728
rect 210255 77670 210528 77672
rect 210255 77667 210321 77670
rect 640194 77656 640254 77700
rect 647823 77656 647889 77659
rect 640194 77654 647889 77656
rect 640194 77598 647828 77654
rect 647884 77598 647889 77654
rect 640194 77596 647889 77598
rect 647823 77593 647889 77596
rect 146895 77508 146961 77511
rect 140832 77506 146961 77508
rect 140832 77450 146900 77506
rect 146956 77450 146961 77506
rect 140832 77448 146961 77450
rect 146895 77445 146961 77448
rect 201711 77212 201777 77215
rect 647919 77212 647985 77215
rect 201711 77210 210528 77212
rect 201711 77154 201716 77210
rect 201772 77154 210528 77210
rect 201711 77152 210528 77154
rect 640224 77210 647985 77212
rect 640224 77154 647924 77210
rect 647980 77154 647985 77210
rect 640224 77152 647985 77154
rect 201711 77149 201777 77152
rect 647919 77149 647985 77152
rect 201615 76620 201681 76623
rect 646671 76620 646737 76623
rect 201615 76618 210528 76620
rect 201615 76562 201620 76618
rect 201676 76562 210528 76618
rect 201615 76560 210528 76562
rect 640224 76618 646737 76620
rect 640224 76562 646676 76618
rect 646732 76562 646737 76618
rect 640224 76560 646737 76562
rect 201615 76557 201681 76560
rect 646671 76557 646737 76560
rect 195567 76472 195633 76475
rect 646287 76472 646353 76475
rect 195567 76470 210558 76472
rect 195567 76414 195572 76470
rect 195628 76414 210558 76470
rect 195567 76412 210558 76414
rect 195567 76409 195633 76412
rect 140802 75732 140862 76220
rect 210498 76072 210558 76412
rect 640194 76470 646353 76472
rect 640194 76414 646292 76470
rect 646348 76414 646353 76470
rect 640194 76412 646353 76414
rect 640194 76072 640254 76412
rect 646287 76409 646353 76412
rect 144111 75732 144177 75735
rect 140802 75730 144177 75732
rect 140802 75674 144116 75730
rect 144172 75674 144177 75730
rect 140802 75672 144177 75674
rect 144111 75669 144177 75672
rect 201807 75584 201873 75587
rect 646479 75584 646545 75587
rect 201807 75582 210528 75584
rect 201807 75526 201812 75582
rect 201868 75526 210528 75582
rect 201807 75524 210528 75526
rect 640224 75582 646545 75584
rect 640224 75526 646484 75582
rect 646540 75526 646545 75582
rect 640224 75524 646545 75526
rect 201807 75521 201873 75524
rect 646479 75521 646545 75524
rect 140802 75140 140862 75184
rect 144015 75140 144081 75143
rect 140802 75138 144081 75140
rect 140802 75082 144020 75138
rect 144076 75082 144081 75138
rect 140802 75080 144081 75082
rect 144015 75077 144081 75080
rect 201519 74992 201585 74995
rect 647919 74992 647985 74995
rect 201519 74990 210528 74992
rect 201519 74934 201524 74990
rect 201580 74934 210528 74990
rect 201519 74932 210528 74934
rect 640224 74990 647985 74992
rect 640224 74934 647924 74990
rect 647980 74934 647985 74990
rect 640224 74932 647985 74934
rect 201519 74929 201585 74932
rect 647919 74929 647985 74932
rect 210255 74474 210321 74477
rect 210255 74472 210528 74474
rect 210255 74416 210260 74472
rect 210316 74416 210528 74472
rect 210255 74414 210528 74416
rect 210255 74411 210321 74414
rect 640194 74104 640254 74444
rect 646095 74104 646161 74107
rect 640194 74102 646161 74104
rect 640194 74046 646100 74102
rect 646156 74046 646161 74102
rect 640194 74044 646161 74046
rect 646095 74041 646161 74044
rect 144015 73956 144081 73959
rect 140832 73954 144081 73956
rect 140832 73898 144020 73954
rect 144076 73898 144081 73954
rect 140832 73896 144081 73898
rect 144015 73893 144081 73896
rect 201039 73956 201105 73959
rect 647151 73956 647217 73959
rect 201039 73954 210528 73956
rect 201039 73898 201044 73954
rect 201100 73898 210528 73954
rect 201039 73896 210528 73898
rect 640224 73954 647217 73956
rect 640224 73898 647156 73954
rect 647212 73898 647217 73954
rect 640224 73896 647217 73898
rect 201039 73893 201105 73896
rect 647151 73893 647217 73896
rect 198351 73364 198417 73367
rect 646287 73364 646353 73367
rect 198351 73362 210528 73364
rect 198351 73306 198356 73362
rect 198412 73306 210528 73362
rect 198351 73304 210528 73306
rect 640224 73362 646353 73364
rect 640224 73306 646292 73362
rect 646348 73306 646353 73362
rect 640224 73304 646353 73306
rect 198351 73301 198417 73304
rect 646287 73301 646353 73304
rect 200943 73216 201009 73219
rect 646383 73216 646449 73219
rect 200943 73214 210558 73216
rect 200943 73158 200948 73214
rect 201004 73158 210558 73214
rect 200943 73156 210558 73158
rect 200943 73153 201009 73156
rect 210498 72816 210558 73156
rect 640194 73214 646449 73216
rect 640194 73158 646388 73214
rect 646444 73158 646449 73214
rect 640194 73156 646449 73158
rect 640194 72816 640254 73156
rect 646383 73153 646449 73156
rect 144111 72772 144177 72775
rect 140832 72770 144177 72772
rect 140832 72714 144116 72770
rect 144172 72714 144177 72770
rect 140832 72712 144177 72714
rect 144111 72709 144177 72712
rect 201711 72328 201777 72331
rect 646671 72328 646737 72331
rect 201711 72326 210528 72328
rect 201711 72270 201716 72326
rect 201772 72270 210528 72326
rect 201711 72268 210528 72270
rect 640224 72326 646737 72328
rect 640224 72270 646676 72326
rect 646732 72270 646737 72326
rect 640224 72268 646737 72270
rect 201711 72265 201777 72268
rect 646671 72265 646737 72268
rect 209967 71886 210033 71887
rect 209914 71822 209920 71886
rect 209984 71884 210033 71886
rect 209984 71882 210076 71884
rect 210028 71826 210076 71882
rect 209984 71824 210076 71826
rect 209984 71822 210033 71824
rect 209967 71821 210033 71822
rect 201711 71736 201777 71739
rect 201711 71734 210528 71736
rect 201711 71678 201716 71734
rect 201772 71678 210528 71734
rect 201711 71676 210528 71678
rect 201711 71673 201777 71676
rect 140802 70996 140862 71484
rect 209967 71218 210033 71221
rect 209967 71216 210528 71218
rect 209967 71160 209972 71216
rect 210028 71160 210528 71216
rect 209967 71158 210528 71160
rect 209967 71155 210033 71158
rect 144015 70996 144081 70999
rect 140802 70994 144081 70996
rect 140802 70938 144020 70994
rect 144076 70938 144081 70994
rect 140802 70936 144081 70938
rect 144015 70933 144081 70936
rect 201615 70700 201681 70703
rect 201615 70698 210528 70700
rect 201615 70642 201620 70698
rect 201676 70642 210528 70698
rect 201615 70640 210528 70642
rect 201615 70637 201681 70640
rect 140802 69812 140862 70290
rect 201807 70108 201873 70111
rect 201807 70106 210528 70108
rect 201807 70050 201812 70106
rect 201868 70050 210528 70106
rect 201807 70048 210528 70050
rect 201807 70045 201873 70048
rect 144015 69812 144081 69815
rect 140802 69810 144081 69812
rect 140802 69754 144020 69810
rect 144076 69754 144081 69810
rect 140802 69752 144081 69754
rect 144015 69749 144081 69752
rect 200463 69516 200529 69519
rect 200463 69514 210528 69516
rect 200463 69458 200468 69514
rect 200524 69458 210528 69514
rect 200463 69456 210528 69458
rect 200463 69453 200529 69456
rect 144207 69072 144273 69075
rect 140832 69070 144273 69072
rect 140832 69014 144212 69070
rect 144268 69014 144273 69070
rect 140832 69012 144273 69014
rect 144207 69009 144273 69012
rect 194703 69072 194769 69075
rect 194703 69070 210528 69072
rect 194703 69014 194708 69070
rect 194764 69014 210528 69070
rect 194703 69012 210528 69014
rect 194703 69009 194769 69012
rect 201711 68480 201777 68483
rect 201711 68478 210528 68480
rect 201711 68422 201716 68478
rect 201772 68422 210528 68478
rect 201711 68420 210528 68422
rect 201711 68417 201777 68420
rect 140802 67592 140862 67932
rect 201615 67888 201681 67891
rect 201615 67886 210528 67888
rect 201615 67830 201620 67886
rect 201676 67830 210528 67886
rect 201615 67828 210528 67830
rect 201615 67825 201681 67828
rect 144015 67592 144081 67595
rect 140802 67590 144081 67592
rect 140802 67534 144020 67590
rect 144076 67534 144081 67590
rect 140802 67532 144081 67534
rect 144015 67529 144081 67532
rect 201807 67444 201873 67447
rect 201807 67442 210528 67444
rect 201807 67386 201812 67442
rect 201868 67386 210528 67442
rect 201807 67384 210528 67386
rect 201807 67381 201873 67384
rect 201519 66852 201585 66855
rect 201519 66850 210528 66852
rect 201519 66794 201524 66850
rect 201580 66794 210528 66850
rect 201519 66792 210528 66794
rect 201519 66789 201585 66792
rect 140802 66408 140862 66748
rect 144015 66408 144081 66411
rect 140802 66406 144081 66408
rect 140802 66350 144020 66406
rect 144076 66350 144081 66406
rect 140802 66348 144081 66350
rect 144015 66345 144081 66348
rect 201615 66260 201681 66263
rect 201615 66258 210528 66260
rect 201615 66202 201620 66258
rect 201676 66202 210528 66258
rect 201615 66200 210528 66202
rect 201615 66197 201681 66200
rect 201711 65816 201777 65819
rect 201711 65814 210528 65816
rect 201711 65758 201716 65814
rect 201772 65758 210528 65814
rect 201711 65756 210528 65758
rect 201711 65753 201777 65756
rect 146223 65520 146289 65523
rect 140832 65518 146289 65520
rect 140832 65462 146228 65518
rect 146284 65462 146289 65518
rect 140832 65460 146289 65462
rect 146223 65457 146289 65460
rect 200175 65224 200241 65227
rect 200175 65222 210528 65224
rect 200175 65166 200180 65222
rect 200236 65166 210528 65222
rect 200175 65164 210528 65166
rect 200175 65161 200241 65164
rect 144015 64780 144081 64783
rect 140802 64778 144081 64780
rect 140802 64722 144020 64778
rect 144076 64722 144081 64778
rect 140802 64720 144081 64722
rect 140802 64334 140862 64720
rect 144015 64717 144081 64720
rect 201711 64632 201777 64635
rect 201711 64630 210528 64632
rect 201711 64574 201716 64630
rect 201772 64574 210528 64630
rect 201711 64572 210528 64574
rect 201711 64569 201777 64572
rect 193743 64188 193809 64191
rect 193743 64186 210528 64188
rect 193743 64130 193748 64186
rect 193804 64130 210528 64186
rect 193743 64128 210528 64130
rect 193743 64125 193809 64128
rect 201711 63596 201777 63599
rect 201711 63594 210528 63596
rect 201711 63538 201716 63594
rect 201772 63538 210528 63594
rect 201711 63536 210528 63538
rect 201711 63533 201777 63536
rect 140802 62708 140862 63048
rect 201711 63004 201777 63007
rect 201711 63002 210528 63004
rect 201711 62946 201716 63002
rect 201772 62946 210528 63002
rect 201711 62944 210528 62946
rect 201711 62941 201777 62944
rect 144015 62708 144081 62711
rect 140802 62706 144081 62708
rect 140802 62650 144020 62706
rect 144076 62650 144081 62706
rect 140802 62648 144081 62650
rect 144015 62645 144081 62648
rect 194127 62560 194193 62563
rect 194127 62558 210528 62560
rect 194127 62502 194132 62558
rect 194188 62502 210528 62558
rect 194127 62500 210528 62502
rect 194127 62497 194193 62500
rect 146895 62412 146961 62415
rect 140802 62410 146961 62412
rect 140802 62354 146900 62410
rect 146956 62354 146961 62410
rect 140802 62352 146961 62354
rect 140802 61864 140862 62352
rect 146895 62349 146961 62352
rect 201615 61968 201681 61971
rect 201615 61966 210528 61968
rect 201615 61910 201620 61966
rect 201676 61910 210528 61966
rect 201615 61908 210528 61910
rect 201615 61905 201681 61908
rect 199311 61376 199377 61379
rect 199311 61374 210528 61376
rect 199311 61318 199316 61374
rect 199372 61318 210528 61374
rect 199311 61316 210528 61318
rect 199311 61313 199377 61316
rect 209967 60858 210033 60861
rect 209967 60856 210528 60858
rect 209967 60800 209972 60856
rect 210028 60800 210528 60856
rect 209967 60798 210528 60800
rect 209967 60795 210033 60798
rect 146895 60784 146961 60787
rect 140832 60782 146961 60784
rect 140832 60726 146900 60782
rect 146956 60726 146961 60782
rect 140832 60724 146961 60726
rect 146895 60721 146961 60724
rect 201615 60340 201681 60343
rect 201615 60338 210528 60340
rect 201615 60282 201620 60338
rect 201676 60282 210528 60338
rect 201615 60280 210528 60282
rect 201615 60277 201681 60280
rect 201711 59748 201777 59751
rect 201711 59746 210528 59748
rect 201711 59690 201716 59746
rect 201772 59690 210528 59746
rect 201711 59688 210528 59690
rect 201711 59685 201777 59688
rect 146511 59600 146577 59603
rect 140832 59598 146577 59600
rect 140832 59542 146516 59598
rect 146572 59542 146577 59598
rect 140832 59540 146577 59542
rect 146511 59537 146577 59540
rect 209967 59230 210033 59233
rect 209967 59228 210528 59230
rect 209967 59172 209972 59228
rect 210028 59172 210528 59228
rect 209967 59170 210528 59172
rect 209967 59167 210033 59170
rect 144015 58712 144081 58715
rect 140802 58710 144081 58712
rect 140802 58654 144020 58710
rect 144076 58654 144081 58710
rect 140802 58652 144081 58654
rect 140802 58322 140862 58652
rect 144015 58649 144081 58652
rect 210882 58418 210942 58682
rect 210874 58354 210880 58418
rect 210944 58354 210950 58418
rect 209967 58120 210033 58123
rect 209967 58118 210528 58120
rect 209967 58062 209972 58118
rect 210028 58062 210528 58118
rect 209967 58060 210528 58062
rect 209967 58057 210033 58060
rect 144015 57380 144081 57383
rect 140802 57378 144081 57380
rect 140802 57322 144020 57378
rect 144076 57322 144081 57378
rect 140802 57320 144081 57322
rect 140802 57128 140862 57320
rect 144015 57317 144081 57320
rect 210498 57234 210558 57572
rect 210490 57170 210496 57234
rect 210560 57170 210566 57234
rect 210159 57084 210225 57087
rect 210159 57082 210528 57084
rect 210159 57026 210164 57082
rect 210220 57026 210528 57082
rect 210159 57024 210528 57026
rect 210159 57021 210225 57024
rect 144111 56492 144177 56495
rect 140802 56490 144177 56492
rect 140802 56434 144116 56490
rect 144172 56434 144177 56490
rect 140802 56432 144177 56434
rect 140802 55874 140862 56432
rect 144111 56429 144177 56432
rect 210255 56492 210321 56495
rect 210255 56490 210528 56492
rect 210255 56434 210260 56490
rect 210316 56434 210528 56490
rect 210255 56432 210528 56434
rect 210255 56429 210321 56432
rect 207279 55604 207345 55607
rect 210498 55604 210558 55944
rect 207279 55602 210558 55604
rect 207279 55546 207284 55602
rect 207340 55546 210558 55602
rect 207279 55544 210558 55546
rect 207279 55541 207345 55544
rect 210882 55162 210942 55426
rect 210874 55098 210880 55162
rect 210944 55098 210950 55162
rect 144015 54716 144081 54719
rect 140832 54714 144081 54716
rect 140832 54658 144020 54714
rect 144076 54658 144081 54714
rect 140832 54656 144081 54658
rect 144015 54653 144081 54656
rect 210690 54423 210750 54834
rect 210351 54422 210417 54423
rect 210298 54420 210304 54422
rect 210260 54360 210304 54420
rect 210368 54418 210417 54422
rect 210412 54362 210417 54418
rect 210298 54358 210304 54360
rect 210368 54358 210417 54362
rect 210351 54357 210417 54358
rect 210639 54418 210750 54423
rect 210639 54362 210644 54418
rect 210700 54362 210750 54418
rect 210639 54360 210750 54362
rect 210639 54357 210705 54360
rect 210874 54358 210880 54422
rect 210944 54420 210950 54422
rect 220623 54420 220689 54423
rect 210944 54418 220689 54420
rect 210944 54362 220628 54418
rect 220684 54362 220689 54418
rect 210944 54360 220689 54362
rect 210944 54358 210950 54360
rect 220623 54357 220689 54360
rect 203151 54272 203217 54275
rect 218607 54272 218673 54275
rect 203151 54270 218673 54272
rect 203151 54214 203156 54270
rect 203212 54214 218612 54270
rect 218668 54214 218673 54270
rect 203151 54212 218673 54214
rect 203151 54209 203217 54212
rect 218607 54209 218673 54212
rect 209914 54062 209920 54126
rect 209984 54124 209990 54126
rect 210063 54124 210129 54127
rect 209984 54122 210129 54124
rect 209984 54066 210068 54122
rect 210124 54066 210129 54122
rect 209984 54064 210129 54066
rect 209984 54062 209990 54064
rect 210063 54061 210129 54064
rect 210682 54062 210688 54126
rect 210752 54124 210758 54126
rect 214191 54124 214257 54127
rect 210752 54122 214257 54124
rect 210752 54066 214196 54122
rect 214252 54066 214257 54122
rect 210752 54064 214257 54066
rect 210752 54062 210758 54064
rect 214191 54061 214257 54064
rect 210490 53914 210496 53978
rect 210560 53976 210566 53978
rect 229647 53976 229713 53979
rect 210560 53974 229713 53976
rect 210560 53918 229652 53974
rect 229708 53918 229713 53974
rect 210560 53916 229713 53918
rect 210560 53914 210566 53916
rect 229647 53913 229713 53916
rect 144015 53828 144081 53831
rect 140802 53826 144081 53828
rect 140802 53770 144020 53826
rect 144076 53770 144081 53826
rect 140802 53768 144081 53770
rect 140802 53576 140862 53768
rect 144015 53765 144081 53768
rect 212602 53766 212608 53830
rect 212672 53828 212678 53830
rect 212672 53768 217038 53828
rect 212672 53766 212678 53768
rect 211450 53618 211456 53682
rect 211520 53680 211526 53682
rect 216978 53680 217038 53768
rect 211520 53646 215262 53680
rect 216978 53646 217086 53680
rect 211520 53641 215265 53646
rect 211520 53620 215204 53641
rect 211520 53618 211526 53620
rect 215199 53585 215204 53620
rect 215260 53585 215265 53641
rect 216978 53641 217089 53646
rect 216978 53620 217028 53641
rect 215199 53580 215265 53585
rect 217023 53585 217028 53620
rect 217084 53585 217089 53641
rect 217023 53580 217089 53585
rect 211066 53470 211072 53534
rect 211136 53532 211142 53534
rect 211791 53532 211857 53535
rect 211136 53530 211857 53532
rect 211136 53474 211796 53530
rect 211852 53474 211857 53530
rect 211136 53472 211857 53474
rect 211136 53470 211142 53472
rect 211791 53469 211857 53472
rect 212986 53470 212992 53534
rect 213056 53532 213062 53534
rect 214863 53532 214929 53535
rect 213056 53530 214929 53532
rect 213056 53474 214868 53530
rect 214924 53474 214929 53530
rect 213056 53472 214929 53474
rect 213056 53470 213062 53472
rect 214863 53469 214929 53472
rect 246978 53472 249726 53532
rect 209679 53384 209745 53387
rect 212943 53384 213009 53387
rect 209679 53382 213009 53384
rect 209679 53326 209684 53382
rect 209740 53326 212948 53382
rect 213004 53326 213009 53382
rect 209679 53324 213009 53326
rect 209679 53321 209745 53324
rect 212943 53321 213009 53324
rect 229647 53384 229713 53387
rect 246978 53384 247038 53472
rect 229647 53382 247038 53384
rect 229647 53326 229652 53382
rect 229708 53326 247038 53382
rect 229647 53324 247038 53326
rect 229647 53321 229713 53324
rect 210106 53174 210112 53238
rect 210176 53236 210182 53238
rect 221103 53236 221169 53239
rect 210176 53234 221169 53236
rect 210176 53178 221108 53234
rect 221164 53178 221169 53234
rect 210176 53176 221169 53178
rect 249666 53236 249726 53472
rect 423279 53384 423345 53387
rect 443439 53384 443505 53387
rect 465658 53384 465664 53386
rect 423279 53382 443505 53384
rect 423279 53326 423284 53382
rect 423340 53326 443444 53382
rect 443500 53326 443505 53382
rect 423279 53324 443505 53326
rect 423279 53321 423345 53324
rect 443439 53321 443505 53324
rect 453570 53324 465664 53384
rect 354255 53236 354321 53239
rect 453570 53236 453630 53324
rect 465658 53322 465664 53324
rect 465728 53322 465734 53386
rect 249666 53176 282366 53236
rect 210176 53174 210182 53176
rect 221103 53173 221169 53176
rect 211834 53026 211840 53090
rect 211904 53088 211910 53090
rect 216687 53088 216753 53091
rect 211904 53086 216753 53088
rect 211904 53030 216692 53086
rect 216748 53030 216753 53086
rect 211904 53028 216753 53030
rect 211904 53026 211910 53028
rect 216687 53025 216753 53028
rect 282306 52940 282366 53176
rect 306498 53234 354321 53236
rect 306498 53178 354260 53234
rect 354316 53178 354321 53234
rect 306498 53176 354321 53178
rect 306498 52940 306558 53176
rect 354255 53173 354321 53176
rect 383106 53176 413118 53236
rect 377530 53026 377536 53090
rect 377600 53088 377606 53090
rect 383106 53088 383166 53176
rect 377600 53028 383166 53088
rect 377600 53026 377606 53028
rect 282306 52880 306558 52940
rect 374319 52940 374385 52943
rect 377338 52940 377344 52942
rect 374319 52938 377344 52940
rect 374319 52882 374324 52938
rect 374380 52882 377344 52938
rect 374319 52880 377344 52882
rect 374319 52877 374385 52880
rect 377338 52878 377344 52880
rect 377408 52878 377414 52942
rect 413058 52940 413118 53176
rect 433410 53176 453630 53236
rect 433410 52940 433470 53176
rect 413058 52880 433470 52940
rect 221871 52644 221937 52647
rect 636730 52644 636736 52646
rect 221871 52642 636736 52644
rect 221871 52586 221876 52642
rect 221932 52586 636736 52642
rect 221871 52584 636736 52586
rect 221871 52581 221937 52584
rect 636730 52582 636736 52584
rect 636800 52582 636806 52646
rect 222543 52496 222609 52499
rect 637498 52496 637504 52498
rect 222543 52494 637504 52496
rect 222543 52438 222548 52494
rect 222604 52438 637504 52494
rect 222543 52436 637504 52438
rect 222543 52433 222609 52436
rect 637498 52434 637504 52436
rect 637568 52434 637574 52498
rect 223695 52348 223761 52351
rect 637114 52348 637120 52350
rect 223695 52346 637120 52348
rect 223695 52290 223700 52346
rect 223756 52290 637120 52346
rect 223695 52288 637120 52290
rect 223695 52285 223761 52288
rect 637114 52286 637120 52288
rect 637184 52286 637190 52350
rect 223311 52200 223377 52203
rect 637690 52200 637696 52202
rect 223311 52198 637696 52200
rect 223311 52142 223316 52198
rect 223372 52142 637696 52198
rect 223311 52140 637696 52142
rect 223311 52137 223377 52140
rect 637690 52138 637696 52140
rect 637760 52138 637766 52202
rect 212655 52052 212721 52055
rect 636922 52052 636928 52054
rect 212655 52050 636928 52052
rect 212655 51994 212660 52050
rect 212716 51994 636928 52050
rect 212655 51992 636928 51994
rect 212655 51989 212721 51992
rect 636922 51990 636928 51992
rect 636992 51990 636998 52054
rect 211887 51904 211953 51907
rect 637306 51904 637312 51906
rect 211887 51902 637312 51904
rect 211887 51846 211892 51902
rect 211948 51846 637312 51902
rect 211887 51844 637312 51846
rect 211887 51841 211953 51844
rect 637306 51842 637312 51844
rect 637376 51842 637382 51906
rect 434895 51756 434961 51759
rect 459279 51756 459345 51759
rect 434895 51754 459345 51756
rect 434895 51698 434900 51754
rect 434956 51698 459284 51754
rect 459340 51698 459345 51754
rect 434895 51696 459345 51698
rect 434895 51693 434961 51696
rect 459279 51693 459345 51696
rect 601935 51756 602001 51759
rect 621999 51756 622065 51759
rect 601935 51754 622065 51756
rect 601935 51698 601940 51754
rect 601996 51698 622004 51754
rect 622060 51698 622065 51754
rect 601935 51696 622065 51698
rect 601935 51693 602001 51696
rect 621999 51693 622065 51696
rect 362895 51608 362961 51611
rect 382959 51608 383025 51611
rect 362895 51606 383025 51608
rect 362895 51550 362900 51606
rect 362956 51550 382964 51606
rect 383020 51550 383025 51606
rect 362895 51548 383025 51550
rect 362895 51545 362961 51548
rect 382959 51545 383025 51548
rect 403215 51608 403281 51611
rect 423279 51608 423345 51611
rect 403215 51606 423345 51608
rect 403215 51550 403220 51606
rect 403276 51550 423284 51606
rect 423340 51550 423345 51606
rect 403215 51548 423345 51550
rect 403215 51545 403281 51548
rect 423279 51545 423345 51548
rect 489615 51608 489681 51611
rect 509583 51608 509649 51611
rect 489615 51606 509649 51608
rect 489615 51550 489620 51606
rect 489676 51550 509588 51606
rect 509644 51550 509649 51606
rect 489615 51548 509649 51550
rect 489615 51545 489681 51548
rect 509583 51545 509649 51548
rect 145978 51250 145984 51314
rect 146048 51312 146054 51314
rect 237231 51312 237297 51315
rect 146048 51310 237297 51312
rect 146048 51254 237236 51310
rect 237292 51254 237297 51310
rect 146048 51252 237297 51254
rect 146048 51250 146054 51252
rect 237231 51249 237297 51252
rect 145786 51102 145792 51166
rect 145856 51164 145862 51166
rect 237807 51164 237873 51167
rect 145856 51162 237873 51164
rect 145856 51106 237812 51162
rect 237868 51106 237873 51162
rect 145856 51104 237873 51106
rect 145856 51102 145862 51104
rect 237807 51101 237873 51104
rect 145402 50954 145408 51018
rect 145472 51016 145478 51018
rect 243471 51016 243537 51019
rect 145472 51014 243537 51016
rect 145472 50958 243476 51014
rect 243532 50958 243537 51014
rect 145472 50956 243537 50958
rect 145472 50954 145478 50956
rect 243471 50953 243537 50956
rect 145594 50806 145600 50870
rect 145664 50868 145670 50870
rect 238191 50868 238257 50871
rect 145664 50866 238257 50868
rect 145664 50810 238196 50866
rect 238252 50810 238257 50866
rect 145664 50808 238257 50810
rect 145664 50806 145670 50808
rect 238191 50805 238257 50808
rect 302415 48944 302481 48947
rect 306682 48944 306688 48946
rect 302415 48942 306688 48944
rect 302415 48886 302420 48942
rect 302476 48886 306688 48942
rect 302415 48884 306688 48886
rect 302415 48881 302481 48884
rect 306682 48882 306688 48884
rect 306752 48882 306758 48946
rect 207183 48796 207249 48799
rect 219951 48796 220017 48799
rect 207183 48794 220017 48796
rect 207183 48738 207188 48794
rect 207244 48738 219956 48794
rect 220012 48738 220017 48794
rect 207183 48736 220017 48738
rect 207183 48733 207249 48736
rect 219951 48733 220017 48736
rect 168399 48648 168465 48651
rect 242991 48648 243057 48651
rect 168399 48646 243057 48648
rect 168399 48590 168404 48646
rect 168460 48590 242996 48646
rect 243052 48590 243057 48646
rect 168399 48588 243057 48590
rect 168399 48585 168465 48588
rect 242991 48585 243057 48588
rect 171279 48500 171345 48503
rect 242223 48500 242289 48503
rect 171279 48498 242289 48500
rect 171279 48442 171284 48498
rect 171340 48442 242228 48498
rect 242284 48442 242289 48498
rect 171279 48440 242289 48442
rect 171279 48437 171345 48440
rect 242223 48437 242289 48440
rect 174159 48352 174225 48355
rect 243375 48352 243441 48355
rect 174159 48350 243441 48352
rect 174159 48294 174164 48350
rect 174220 48294 243380 48350
rect 243436 48294 243441 48350
rect 174159 48292 243441 48294
rect 174159 48289 174225 48292
rect 243375 48289 243441 48292
rect 188559 48204 188625 48207
rect 239439 48204 239505 48207
rect 188559 48202 239505 48204
rect 188559 48146 188564 48202
rect 188620 48146 239444 48202
rect 239500 48146 239505 48202
rect 188559 48144 239505 48146
rect 188559 48141 188625 48144
rect 239439 48141 239505 48144
rect 194319 48056 194385 48059
rect 240015 48056 240081 48059
rect 194319 48054 240081 48056
rect 194319 47998 194324 48054
rect 194380 47998 240020 48054
rect 240076 47998 240081 48054
rect 194319 47996 240081 47998
rect 194319 47993 194385 47996
rect 240015 47993 240081 47996
rect 162639 47908 162705 47911
rect 241647 47908 241713 47911
rect 162639 47906 241713 47908
rect 162639 47850 162644 47906
rect 162700 47850 241652 47906
rect 241708 47850 241713 47906
rect 162639 47848 241713 47850
rect 162639 47845 162705 47848
rect 241647 47845 241713 47848
rect 205167 47760 205233 47763
rect 220719 47760 220785 47763
rect 205167 47758 220785 47760
rect 205167 47702 205172 47758
rect 205228 47702 220724 47758
rect 220780 47702 220785 47758
rect 205167 47700 220785 47702
rect 205167 47697 205233 47700
rect 220719 47697 220785 47700
rect 165519 47612 165585 47615
rect 242607 47612 242673 47615
rect 165519 47610 242673 47612
rect 165519 47554 165524 47610
rect 165580 47554 242612 47610
rect 242668 47554 242673 47610
rect 165519 47552 242673 47554
rect 165519 47549 165585 47552
rect 242607 47549 242673 47552
rect 353583 46132 353649 46135
rect 356986 46132 356992 46134
rect 353583 46130 356992 46132
rect 353583 46074 353588 46130
rect 353644 46074 356992 46130
rect 353583 46072 356992 46074
rect 353583 46069 353649 46072
rect 356986 46070 356992 46072
rect 357056 46070 357062 46134
rect 212079 45392 212145 45395
rect 302458 45392 302464 45394
rect 212079 45390 302464 45392
rect 212079 45334 212084 45390
rect 212140 45334 302464 45390
rect 212079 45332 302464 45334
rect 212079 45329 212145 45332
rect 302458 45330 302464 45332
rect 302528 45330 302534 45394
rect 211311 45244 211377 45247
rect 360058 45244 360064 45246
rect 211311 45242 360064 45244
rect 211311 45186 211316 45242
rect 211372 45186 360064 45242
rect 211311 45184 360064 45186
rect 211311 45181 211377 45184
rect 360058 45182 360064 45184
rect 360128 45182 360134 45246
rect 211695 45096 211761 45099
rect 362938 45096 362944 45098
rect 211695 45094 362944 45096
rect 211695 45038 211700 45094
rect 211756 45038 362944 45094
rect 211695 45036 362944 45038
rect 211695 45033 211761 45036
rect 362938 45034 362944 45036
rect 363008 45034 363014 45098
rect 213135 44948 213201 44951
rect 409018 44948 409024 44950
rect 213135 44946 409024 44948
rect 213135 44890 213140 44946
rect 213196 44890 409024 44946
rect 213135 44888 409024 44890
rect 213135 44885 213201 44888
rect 409018 44886 409024 44888
rect 409088 44886 409094 44950
rect 215055 44800 215121 44803
rect 518799 44800 518865 44803
rect 215055 44798 518865 44800
rect 215055 44742 215060 44798
rect 215116 44742 518804 44798
rect 518860 44742 518865 44798
rect 215055 44740 518865 44742
rect 215055 44737 215121 44740
rect 518799 44737 518865 44740
rect 215343 44652 215409 44655
rect 529263 44652 529329 44655
rect 215343 44650 529329 44652
rect 215343 44594 215348 44650
rect 215404 44594 529268 44650
rect 529324 44594 529329 44650
rect 215343 44592 529329 44594
rect 215343 44589 215409 44592
rect 529263 44589 529329 44592
rect 302511 43322 302577 43323
rect 302458 43320 302464 43322
rect 302420 43260 302464 43320
rect 302528 43318 302577 43322
rect 302572 43262 302577 43318
rect 302458 43258 302464 43260
rect 302528 43258 302577 43262
rect 360058 43258 360064 43322
rect 360128 43320 360134 43322
rect 361743 43320 361809 43323
rect 360128 43318 361809 43320
rect 360128 43262 361748 43318
rect 361804 43262 361809 43318
rect 360128 43260 361809 43262
rect 360128 43258 360134 43260
rect 302511 43257 302577 43258
rect 361743 43257 361809 43260
rect 362938 43258 362944 43322
rect 363008 43320 363014 43322
rect 364911 43320 364977 43323
rect 363008 43318 364977 43320
rect 363008 43262 364916 43318
rect 364972 43262 364977 43318
rect 363008 43260 364977 43262
rect 363008 43258 363014 43260
rect 364911 43257 364977 43260
rect 409018 43258 409024 43322
rect 409088 43320 409094 43322
rect 410799 43320 410865 43323
rect 409088 43318 410865 43320
rect 409088 43262 410804 43318
rect 410860 43262 410865 43318
rect 409088 43260 410865 43262
rect 409088 43258 409094 43260
rect 410799 43257 410865 43260
rect 306735 42138 306801 42139
rect 306682 42074 306688 42138
rect 306752 42136 306801 42138
rect 306752 42134 306844 42136
rect 306796 42078 306844 42134
rect 306752 42076 306844 42078
rect 306752 42074 306801 42076
rect 356986 42074 356992 42138
rect 357056 42136 357062 42138
rect 357135 42136 357201 42139
rect 357056 42134 357201 42136
rect 357056 42078 357140 42134
rect 357196 42078 357201 42134
rect 357056 42076 357201 42078
rect 357056 42074 357062 42076
rect 306735 42073 306801 42074
rect 357135 42073 357201 42076
rect 408879 42136 408945 42139
rect 416271 42136 416337 42139
rect 408879 42134 416337 42136
rect 408879 42078 408884 42134
rect 408940 42078 416276 42134
rect 416332 42078 416337 42134
rect 408879 42076 416337 42078
rect 408879 42073 408945 42076
rect 416271 42073 416337 42076
rect 187599 41840 187665 41843
rect 189946 41840 189952 41842
rect 187599 41838 189952 41840
rect 187599 41782 187604 41838
rect 187660 41782 189952 41838
rect 187599 41780 189952 41782
rect 187599 41777 187665 41780
rect 189946 41778 189952 41780
rect 190016 41778 190022 41842
rect 194319 41840 194385 41843
rect 194938 41840 194944 41842
rect 194319 41838 194944 41840
rect 194319 41782 194324 41838
rect 194380 41782 194944 41838
rect 194319 41780 194944 41782
rect 194319 41777 194385 41780
rect 194938 41778 194944 41780
rect 195008 41778 195014 41842
rect 458170 41778 458176 41842
rect 458240 41840 458246 41842
rect 463695 41840 463761 41843
rect 465711 41842 465777 41843
rect 465658 41840 465664 41842
rect 458240 41838 463761 41840
rect 458240 41782 463700 41838
rect 463756 41782 463761 41838
rect 458240 41780 463761 41782
rect 465620 41780 465664 41840
rect 465728 41838 465777 41842
rect 465772 41782 465777 41838
rect 458240 41778 458246 41780
rect 463695 41777 463761 41780
rect 465658 41778 465664 41780
rect 465728 41778 465777 41782
rect 465711 41777 465777 41778
rect 189946 40742 189952 40806
rect 190016 40804 190022 40806
rect 210735 40804 210801 40807
rect 190016 40802 210801 40804
rect 190016 40746 210740 40802
rect 210796 40746 210801 40802
rect 190016 40744 210801 40746
rect 190016 40742 190022 40744
rect 210735 40741 210801 40744
rect 194938 40594 194944 40658
rect 195008 40656 195014 40658
rect 625071 40656 625137 40659
rect 195008 40654 625137 40656
rect 195008 40598 625076 40654
rect 625132 40598 625137 40654
rect 195008 40596 625137 40598
rect 195008 40594 195014 40596
rect 625071 40593 625137 40596
rect 141807 40360 141873 40363
rect 457743 40362 457809 40363
rect 457743 40360 457792 40362
rect 141762 40358 141873 40360
rect 141762 40302 141812 40358
rect 141868 40302 141873 40358
rect 141762 40297 141873 40302
rect 457700 40358 457792 40360
rect 457700 40302 457748 40358
rect 457700 40300 457792 40302
rect 457743 40298 457792 40300
rect 457856 40298 457862 40362
rect 457743 40297 457809 40298
rect 141762 39886 141822 40297
<< via3 >>
rect 42112 968762 42176 968766
rect 42112 968706 42124 968762
rect 42124 968706 42176 968762
rect 42112 968702 42176 968706
rect 40384 967074 40448 967138
rect 674368 966334 674432 966398
rect 676480 965742 676544 965806
rect 40960 965002 41024 965066
rect 675904 965002 675968 965066
rect 42496 963966 42560 964030
rect 41344 963374 41408 963438
rect 675328 963286 675392 963290
rect 675328 963230 675380 963286
rect 675380 963230 675392 963286
rect 675328 963226 675392 963230
rect 42304 962782 42368 962846
rect 674752 962634 674816 962698
rect 674560 962190 674624 962254
rect 41728 962042 41792 962106
rect 676096 961302 676160 961366
rect 675712 960770 675776 960774
rect 675712 960714 675724 960770
rect 675724 960714 675776 960770
rect 675712 960710 675776 960714
rect 675520 960178 675584 960182
rect 675520 960122 675532 960178
rect 675532 960122 675584 960178
rect 675520 960118 675584 960122
rect 41152 959674 41216 959738
rect 41536 959082 41600 959146
rect 41920 958402 41984 958406
rect 41920 958346 41972 958402
rect 41972 958346 41984 958402
rect 41920 958342 41984 958346
rect 40768 957750 40832 957814
rect 674944 957602 675008 957666
rect 40576 956122 40640 956186
rect 675136 955974 675200 956038
rect 677056 953458 677120 953522
rect 676864 953310 676928 953374
rect 42880 953162 42944 953226
rect 42688 947598 42752 947602
rect 42688 947542 42700 947598
rect 42700 947542 42752 947598
rect 42688 947538 42752 947542
rect 42688 947390 42752 947454
rect 42880 947390 42944 947454
rect 43072 947242 43136 947306
rect 42688 944726 42752 944790
rect 40576 944430 40640 944494
rect 40384 943690 40448 943754
rect 40768 941618 40832 941682
rect 41728 941174 41792 941238
rect 675904 940878 675968 940942
rect 42112 940582 42176 940646
rect 41920 938806 41984 938870
rect 674368 938658 674432 938722
rect 675328 938362 675392 938426
rect 41536 938066 41600 938130
rect 40960 937326 41024 937390
rect 41344 936438 41408 936502
rect 41152 935846 41216 935910
rect 676480 935846 676544 935910
rect 674752 935254 674816 935318
rect 42304 934958 42368 935022
rect 674560 934514 674624 934578
rect 42496 934070 42560 934134
rect 675136 933330 675200 933394
rect 43072 933094 43136 933098
rect 43072 933038 43084 933094
rect 43084 933038 43136 933094
rect 43072 933034 43136 933038
rect 674944 932886 675008 932950
rect 676096 932146 676160 932210
rect 677056 931406 677120 931470
rect 676864 930222 676928 930286
rect 42496 912906 42560 912970
rect 43072 912906 43136 912970
rect 42496 907134 42560 907198
rect 43072 887214 43136 887218
rect 43072 887158 43124 887214
rect 43124 887158 43136 887214
rect 43072 887154 43136 887158
rect 674560 876350 674624 876414
rect 676096 876350 676160 876414
rect 674944 876202 675008 876266
rect 675520 875758 675584 875822
rect 675712 875610 675776 875674
rect 674752 873982 674816 874046
rect 674368 873390 674432 873454
rect 674176 872798 674240 872862
rect 42496 872502 42560 872566
rect 43072 872502 43136 872566
rect 675328 869898 675392 869902
rect 675328 869842 675380 869898
rect 675380 869842 675392 869898
rect 675328 869838 675392 869842
rect 675136 866878 675200 866942
rect 675712 864718 675776 864722
rect 675712 864662 675724 864718
rect 675724 864662 675776 864718
rect 675712 864658 675776 864662
rect 675520 862942 675584 862946
rect 675520 862886 675532 862942
rect 675532 862886 675584 862942
rect 675520 862882 675584 862886
rect 42496 846750 42560 846814
rect 43072 846750 43136 846814
rect 41920 832246 41984 832310
rect 43072 832246 43136 832310
rect 42112 819518 42176 819582
rect 40768 818630 40832 818694
rect 41920 816262 41984 816326
rect 42688 816262 42752 816326
rect 42496 811970 42560 812034
rect 42880 811970 42944 812034
rect 42496 803594 42560 803598
rect 42496 803538 42508 803594
rect 42508 803538 42560 803594
rect 42496 803534 42560 803538
rect 41344 802202 41408 802266
rect 40384 802054 40448 802118
rect 41536 801906 41600 801970
rect 41728 800338 41792 800342
rect 41728 800282 41780 800338
rect 41780 800282 41792 800338
rect 41728 800278 41792 800282
rect 42496 800278 42560 800342
rect 42304 800042 42368 800046
rect 42304 799986 42316 800042
rect 42316 799986 42368 800042
rect 42304 799982 42368 799986
rect 42304 797910 42368 797974
rect 42496 794802 42560 794866
rect 41728 794270 41792 794274
rect 41728 794214 41780 794270
rect 41780 794214 41792 794270
rect 41728 794210 41792 794214
rect 41536 791842 41600 791906
rect 41344 791694 41408 791758
rect 41728 791310 41792 791314
rect 41728 791254 41780 791310
rect 41780 791254 41792 791310
rect 41728 791250 41792 791254
rect 41920 790954 41984 791018
rect 42496 790954 42560 791018
rect 676288 787846 676352 787910
rect 673984 787402 674048 787466
rect 676480 786662 676544 786726
rect 675904 784146 675968 784210
rect 676672 781926 676736 781990
rect 677056 780446 677120 780510
rect 677056 777486 677120 777550
rect 676864 777338 676928 777402
rect 40384 776746 40448 776810
rect 41344 775858 41408 775922
rect 40768 775118 40832 775182
rect 676864 773046 676928 773110
rect 677824 773046 677888 773110
rect 676864 772898 676928 772962
rect 677248 772898 677312 772962
rect 677248 772602 677312 772666
rect 42112 765942 42176 766006
rect 41536 764018 41600 764082
rect 674944 762390 675008 762454
rect 675712 761650 675776 761714
rect 674560 760466 674624 760530
rect 40960 760170 41024 760234
rect 674752 760022 674816 760086
rect 675328 759134 675392 759198
rect 40384 758542 40448 758606
rect 675520 758542 675584 758606
rect 676096 757358 676160 757422
rect 674368 756322 674432 756386
rect 674176 755434 674240 755498
rect 675136 755286 675200 755350
rect 676864 754398 676928 754462
rect 677824 753806 677888 753870
rect 677248 752918 677312 752982
rect 42880 751942 42944 751946
rect 42880 751886 42892 751942
rect 42892 751886 42944 751942
rect 42880 751882 42944 751886
rect 41536 751734 41600 751798
rect 42880 751646 42944 751650
rect 42880 751590 42892 751646
rect 42892 751590 42944 751646
rect 42880 751586 42944 751590
rect 41728 748686 41792 748690
rect 41728 748630 41780 748686
rect 41780 748630 41792 748686
rect 41728 748626 41792 748630
rect 42112 747502 42176 747506
rect 42112 747446 42164 747502
rect 42164 747446 42176 747502
rect 42112 747442 42176 747446
rect 41920 747354 41984 747358
rect 41920 747298 41972 747354
rect 41972 747298 41984 747354
rect 41920 747294 41984 747298
rect 40384 747146 40448 747210
rect 40960 746850 41024 746914
rect 41920 745814 41984 745878
rect 42112 745370 42176 745434
rect 674560 743298 674624 743362
rect 674176 742114 674240 742178
rect 674752 740190 674816 740254
rect 674368 740042 674432 740106
rect 675520 739214 675584 739218
rect 675520 739158 675532 739214
rect 675532 739158 675584 739214
rect 675520 739154 675584 739158
rect 676096 738710 676160 738774
rect 674944 737674 675008 737738
rect 676672 737674 676736 737738
rect 42112 735958 42176 735962
rect 42112 735902 42124 735958
rect 42124 735902 42176 735958
rect 42112 735898 42176 735902
rect 676864 734862 676928 734926
rect 675136 734122 675200 734186
rect 41344 733826 41408 733890
rect 40576 733086 40640 733150
rect 40768 733086 40832 733150
rect 40960 732198 41024 732262
rect 42112 725894 42176 725898
rect 42112 725838 42124 725894
rect 42124 725838 42176 725894
rect 42112 725834 42176 725838
rect 42688 723762 42752 723826
rect 42304 722578 42368 722642
rect 41344 720802 41408 720866
rect 676480 717102 676544 717166
rect 40384 716954 40448 717018
rect 41152 716658 41216 716722
rect 41536 716066 41600 716130
rect 676288 715770 676352 715834
rect 41920 713906 41984 713910
rect 41920 713850 41932 713906
rect 41932 713850 41984 713906
rect 41920 713846 41984 713850
rect 42496 713846 42560 713910
rect 673984 712070 674048 712134
rect 675904 711922 675968 711986
rect 41920 711686 41984 711690
rect 41920 711630 41932 711686
rect 41932 711630 41984 711686
rect 41920 711626 41984 711630
rect 42496 710738 42560 710802
rect 41344 708518 41408 708582
rect 677056 708370 677120 708434
rect 42688 707778 42752 707842
rect 41536 706742 41600 706806
rect 42304 706150 42368 706214
rect 41344 704670 41408 704734
rect 41728 704730 41792 704734
rect 41728 704674 41780 704730
rect 41780 704674 41792 704730
rect 41728 704670 41792 704674
rect 41536 704078 41600 704142
rect 42112 704078 42176 704142
rect 41152 703634 41216 703698
rect 40384 703486 40448 703550
rect 675904 703042 675968 703106
rect 676288 703042 676352 703106
rect 676096 702450 676160 702514
rect 675328 697922 675392 697926
rect 675328 697866 675380 697922
rect 675380 697866 675392 697922
rect 675328 697862 675392 697866
rect 673984 697270 674048 697334
rect 675904 697122 675968 697186
rect 675520 694814 675584 694818
rect 675520 694758 675532 694814
rect 675532 694758 675584 694814
rect 675520 694754 675584 694758
rect 674944 694310 675008 694374
rect 676672 694310 676736 694374
rect 674944 693422 675008 693486
rect 41344 692742 41408 692746
rect 41344 692686 41396 692742
rect 41396 692686 41408 692742
rect 41344 692682 41408 692686
rect 676288 691942 676352 692006
rect 40576 690314 40640 690378
rect 40960 689574 41024 689638
rect 42304 689574 42368 689638
rect 674176 689426 674240 689490
rect 675712 689426 675776 689490
rect 42112 688686 42176 688750
rect 677056 688242 677120 688306
rect 40576 686318 40640 686382
rect 677056 685578 677120 685642
rect 40960 683210 41024 683274
rect 41728 680842 41792 680906
rect 674176 679658 674240 679722
rect 676480 679658 676544 679722
rect 674176 679510 674240 679574
rect 674944 679570 675008 679574
rect 674944 679514 674996 679570
rect 674996 679514 675008 679570
rect 674944 679510 675008 679514
rect 675904 679570 675968 679574
rect 675904 679514 675916 679570
rect 675916 679514 675968 679570
rect 675904 679510 675968 679514
rect 42496 678326 42560 678390
rect 674944 675366 675008 675430
rect 675328 675366 675392 675430
rect 674752 672258 674816 672322
rect 674752 671518 674816 671582
rect 675136 671282 675200 671286
rect 675136 671226 675148 671282
rect 675148 671226 675200 671282
rect 675136 671222 675200 671226
rect 41344 670986 41408 670990
rect 41344 670930 41396 670986
rect 41396 670930 41408 670986
rect 41344 670926 41408 670930
rect 42880 670926 42944 670990
rect 41920 670778 41984 670842
rect 42688 670778 42752 670842
rect 42688 670630 42752 670694
rect 675136 670690 675200 670694
rect 675136 670634 675148 670690
rect 675148 670634 675200 670690
rect 675136 670630 675200 670634
rect 675328 670630 675392 670694
rect 674560 670482 674624 670546
rect 674560 670334 674624 670398
rect 674368 669224 674432 669288
rect 42496 668766 42560 668770
rect 42496 668710 42548 668766
rect 42548 668710 42560 668766
rect 42496 668706 42560 668710
rect 675712 667522 675776 667586
rect 41728 666694 41792 666698
rect 41728 666638 41780 666694
rect 41780 666638 41792 666694
rect 41728 666634 41792 666638
rect 676096 666634 676160 666698
rect 42688 666486 42752 666550
rect 676480 665894 676544 665958
rect 41344 665450 41408 665514
rect 41536 665302 41600 665366
rect 41536 665006 41600 665070
rect 42688 665006 42752 665070
rect 42880 664710 42944 664774
rect 675136 664266 675200 664330
rect 677248 663526 677312 663590
rect 676864 662342 676928 662406
rect 42688 661454 42752 661518
rect 41920 660774 41984 660778
rect 41920 660718 41932 660774
rect 41932 660718 41984 660774
rect 41920 660714 41984 660718
rect 674752 658346 674816 658410
rect 676480 658346 676544 658410
rect 40960 656718 41024 656782
rect 40576 656126 40640 656190
rect 675904 652574 675968 652638
rect 674176 652130 674240 652194
rect 675136 651390 675200 651454
rect 676288 650946 676352 651010
rect 676096 649614 676160 649678
rect 674944 647986 675008 648050
rect 42304 647394 42368 647458
rect 42112 646654 42176 646718
rect 674368 645322 674432 645386
rect 40576 643102 40640 643166
rect 675520 642510 675584 642574
rect 676288 642510 676352 642574
rect 674752 641178 674816 641242
rect 675328 640882 675392 640946
rect 675904 640882 675968 640946
rect 675520 640734 675584 640798
rect 674560 640586 674624 640650
rect 674944 640586 675008 640650
rect 676480 640438 676544 640502
rect 676480 640290 676544 640354
rect 674944 640142 675008 640206
rect 40768 639994 40832 640058
rect 675328 638574 675392 638578
rect 675328 638518 675380 638574
rect 675380 638518 675392 638574
rect 675328 638514 675392 638518
rect 42304 637626 42368 637690
rect 43072 627918 43136 627922
rect 43072 627862 43124 627918
rect 43124 627862 43136 627918
rect 43072 627858 43136 627862
rect 41920 627474 41984 627478
rect 41920 627418 41932 627474
rect 41932 627418 41984 627474
rect 41920 627414 41984 627418
rect 42112 627474 42176 627478
rect 42112 627418 42164 627474
rect 42164 627418 42176 627474
rect 42112 627414 42176 627418
rect 675904 627266 675968 627330
rect 675520 625638 675584 625702
rect 676288 624750 676352 624814
rect 42688 623862 42752 623926
rect 42304 623418 42368 623482
rect 41920 623270 41984 623334
rect 673984 621938 674048 622002
rect 676672 621642 676736 621706
rect 674944 620902 675008 620966
rect 43072 620754 43136 620818
rect 42112 620222 42176 620226
rect 42112 620166 42124 620222
rect 42124 620166 42176 620222
rect 42112 620162 42176 620166
rect 674752 619126 674816 619190
rect 41920 618446 41984 618450
rect 41920 618390 41972 618446
rect 41972 618390 41984 618446
rect 41920 618386 41984 618390
rect 40768 618238 40832 618302
rect 40576 618090 40640 618154
rect 41728 617854 41792 617858
rect 41728 617798 41780 617854
rect 41780 617798 41792 617854
rect 41728 617794 41792 617798
rect 677056 617794 677120 617858
rect 674752 607730 674816 607794
rect 673984 607434 674048 607498
rect 675520 606458 675584 606462
rect 675520 606402 675532 606458
rect 675532 606402 675584 606458
rect 675520 606398 675584 606402
rect 674944 604770 675008 604834
rect 675904 600182 675968 600246
rect 40576 599886 40640 599950
rect 40960 596778 41024 596842
rect 676672 595298 676736 595362
rect 676288 593374 676352 593438
rect 42880 585382 42944 585446
rect 42496 584702 42560 584706
rect 42496 584646 42548 584702
rect 42548 584646 42560 584702
rect 42496 584642 42560 584646
rect 41536 584198 41600 584262
rect 42304 584198 42368 584262
rect 675136 581682 675200 581746
rect 676480 581238 676544 581302
rect 675712 580350 675776 580414
rect 42304 580054 42368 580118
rect 676096 579610 676160 579674
rect 676096 578870 676160 578934
rect 674368 578352 674432 578416
rect 42880 578338 42944 578342
rect 42880 578282 42932 578338
rect 42932 578282 42944 578338
rect 42880 578278 42944 578282
rect 675328 578130 675392 578194
rect 41536 577094 41600 577158
rect 674176 576724 674240 576788
rect 674560 576058 674624 576122
rect 42496 575910 42560 575974
rect 41920 575230 41984 575234
rect 41920 575174 41972 575230
rect 41972 575174 41984 575230
rect 41920 575170 41984 575174
rect 41728 574638 41792 574642
rect 41728 574582 41780 574638
rect 41780 574582 41792 574638
rect 41728 574578 41792 574582
rect 40960 573986 41024 574050
rect 40576 573838 40640 573902
rect 675328 562946 675392 562950
rect 675328 562890 675340 562946
rect 675340 562890 675392 562946
rect 675328 562886 675392 562890
rect 674176 561702 674240 561766
rect 674560 561554 674624 561618
rect 675136 558890 675200 558954
rect 674368 557706 674432 557770
rect 675712 550158 675776 550222
rect 676096 547050 676160 547114
rect 675712 546902 675776 546966
rect 41152 544238 41216 544302
rect 40960 542906 41024 542970
rect 42112 541278 42176 541342
rect 42880 541130 42944 541194
rect 43072 540982 43136 541046
rect 42112 538762 42176 538826
rect 675520 536986 675584 537050
rect 42880 536898 42944 536902
rect 42880 536842 42932 536898
rect 42932 536842 42944 536898
rect 42880 536838 42944 536842
rect 676672 536246 676736 536310
rect 43072 535654 43136 535718
rect 674752 535358 674816 535422
rect 674944 534618 675008 534682
rect 675904 533730 675968 533794
rect 676288 532694 676352 532758
rect 40960 532546 41024 532610
rect 41152 532250 41216 532314
rect 41920 532014 41984 532018
rect 41920 531958 41932 532014
rect 41932 531958 41984 532014
rect 41920 531954 41984 531958
rect 673984 531658 674048 531722
rect 41728 531274 41792 531278
rect 41728 531218 41780 531274
rect 41780 531218 41792 531274
rect 41728 531214 41792 531218
rect 674560 492290 674624 492354
rect 675328 491402 675392 491466
rect 674176 487702 674240 487766
rect 675136 487406 675200 487470
rect 674368 483780 674432 483844
rect 40576 432646 40640 432710
rect 40384 431906 40448 431970
rect 40768 430722 40832 430786
rect 40960 429390 41024 429454
rect 41344 428354 41408 428418
rect 41536 427614 41600 427678
rect 41152 426282 41216 426346
rect 42112 425098 42176 425162
rect 676480 412134 676544 412138
rect 676480 412078 676532 412134
rect 676532 412078 676544 412134
rect 676480 412074 676544 412078
rect 676672 411986 676736 411990
rect 676672 411930 676684 411986
rect 676684 411930 676736 411986
rect 676672 411926 676736 411930
rect 676480 406154 676544 406218
rect 41536 406006 41600 406070
rect 674176 405858 674240 405922
rect 675520 405266 675584 405330
rect 676672 405266 676736 405330
rect 41920 404882 41984 404886
rect 41920 404826 41972 404882
rect 41972 404826 41984 404882
rect 41920 404822 41984 404826
rect 41728 403846 41792 403850
rect 41728 403790 41780 403846
rect 41780 403790 41792 403846
rect 41728 403786 41792 403790
rect 674944 403194 675008 403258
rect 42112 402662 42176 402666
rect 42112 402606 42164 402662
rect 42164 402606 42176 402662
rect 42112 402602 42176 402606
rect 41344 401862 41408 401926
rect 674560 400530 674624 400594
rect 674368 400382 674432 400446
rect 40768 400086 40832 400150
rect 41920 399938 41984 400002
rect 41152 399494 41216 399558
rect 40960 398754 41024 398818
rect 40576 390170 40640 390234
rect 40384 389134 40448 389198
rect 40768 387506 40832 387570
rect 40960 386026 41024 386090
rect 41344 385138 41408 385202
rect 41152 383066 41216 383130
rect 41536 381882 41600 381946
rect 674560 378774 674624 378838
rect 675328 374482 675392 374546
rect 674944 373890 675008 373954
rect 674368 371966 674432 372030
rect 675712 371670 675776 371734
rect 42112 371522 42176 371586
rect 42112 362850 42176 362854
rect 42112 362794 42124 362850
rect 42124 362794 42176 362850
rect 42112 362790 42176 362794
rect 41920 361962 41984 361966
rect 41920 361906 41932 361962
rect 41932 361906 41984 361962
rect 41920 361902 41984 361906
rect 674368 361384 674432 361448
rect 41728 361370 41792 361374
rect 41728 361314 41780 361370
rect 41780 361314 41792 361370
rect 41728 361310 41792 361314
rect 674176 360718 674240 360782
rect 675520 360126 675584 360190
rect 673984 359978 674048 360042
rect 41536 359386 41600 359450
rect 41344 358646 41408 358710
rect 40768 356870 40832 356934
rect 41152 356426 41216 356490
rect 40960 355538 41024 355602
rect 40576 346806 40640 346870
rect 42112 346214 42176 346278
rect 40384 345918 40448 345982
rect 42304 345918 42368 345982
rect 676672 345474 676736 345538
rect 676096 345326 676160 345390
rect 676480 345178 676544 345242
rect 676288 344438 676352 344502
rect 40960 344290 41024 344354
rect 40768 342810 40832 342874
rect 41344 341922 41408 341986
rect 40384 341182 40448 341246
rect 41152 339850 41216 339914
rect 41536 338666 41600 338730
rect 42688 336150 42752 336214
rect 675328 335026 675392 335030
rect 675328 334970 675340 335026
rect 675340 334970 675392 335026
rect 675328 334966 675392 334970
rect 675520 333842 675584 333846
rect 675520 333786 675572 333842
rect 675572 333786 675584 333842
rect 675520 333782 675584 333786
rect 676096 333486 676160 333550
rect 676288 330526 676352 330590
rect 675328 329490 675392 329554
rect 676672 328010 676736 328074
rect 42496 327418 42560 327482
rect 676480 326826 676544 326890
rect 42496 322978 42560 323042
rect 40384 319722 40448 319786
rect 41920 318746 41984 318750
rect 41920 318690 41932 318746
rect 41932 318690 41984 318746
rect 41920 318686 41984 318690
rect 41728 318006 41792 318010
rect 41728 317950 41780 318006
rect 41780 317950 41792 318006
rect 41728 317946 41792 317950
rect 42688 317354 42752 317418
rect 674368 317206 674432 317270
rect 674368 316392 674432 316456
rect 41536 316170 41600 316234
rect 674176 315726 674240 315790
rect 41344 315430 41408 315494
rect 673984 314838 674048 314902
rect 40960 313654 41024 313718
rect 41152 313210 41216 313274
rect 674560 312618 674624 312682
rect 40768 312322 40832 312386
rect 42112 303738 42176 303802
rect 42304 302998 42368 303062
rect 40768 302258 40832 302322
rect 40960 301074 41024 301138
rect 41152 299594 41216 299658
rect 675712 299446 675776 299510
rect 676672 299298 676736 299362
rect 40576 298706 40640 298770
rect 40384 297966 40448 298030
rect 40576 296634 40640 296698
rect 41344 296634 41408 296698
rect 41536 296634 41600 296698
rect 40576 295450 40640 295514
rect 675328 290034 675392 290038
rect 675328 289978 675340 290034
rect 675340 289978 675392 290034
rect 675328 289974 675392 289978
rect 675520 289590 675584 289594
rect 675520 289534 675532 289590
rect 675532 289534 675584 289590
rect 675520 289530 675584 289534
rect 675712 285298 675776 285302
rect 675712 285242 675724 285298
rect 675724 285242 675776 285298
rect 675712 285238 675776 285242
rect 675136 284942 675200 285006
rect 42304 283670 42368 283674
rect 42304 283614 42316 283670
rect 42316 283614 42368 283670
rect 42304 283610 42368 283614
rect 674560 283610 674624 283674
rect 676672 281834 676736 281898
rect 42304 281538 42368 281602
rect 40384 276506 40448 276570
rect 674944 275322 675008 275386
rect 41920 275234 41984 275238
rect 41920 275178 41972 275234
rect 41972 275178 41984 275234
rect 41920 275174 41984 275178
rect 41728 274642 41792 274646
rect 41728 274586 41780 274642
rect 41780 274586 41792 274642
rect 41728 274582 41792 274586
rect 41920 273990 41984 274054
rect 40576 272806 40640 272870
rect 41536 272362 41600 272426
rect 674368 272214 674432 272278
rect 675712 270882 675776 270946
rect 40960 270586 41024 270650
rect 41920 270438 41984 270502
rect 674176 270142 674240 270206
rect 674560 270142 674624 270206
rect 41344 269994 41408 270058
rect 673984 269846 674048 269910
rect 675328 269698 675392 269762
rect 41152 269106 41216 269170
rect 674752 268514 674816 268578
rect 674368 268218 674432 268282
rect 42112 260374 42176 260438
rect 40768 259486 40832 259550
rect 40384 257858 40448 257922
rect 40576 256378 40640 256442
rect 675136 256230 675200 256294
rect 676288 256230 676352 256294
rect 40960 255638 41024 255702
rect 41344 254750 41408 254814
rect 676096 253566 676160 253630
rect 40768 253418 40832 253482
rect 675904 253418 675968 253482
rect 41152 252382 41216 252446
rect 674752 250458 674816 250522
rect 40576 247794 40640 247858
rect 41536 247646 41600 247710
rect 210688 246314 210752 246378
rect 210304 246166 210368 246230
rect 337024 245130 337088 245194
rect 337024 244982 337088 245046
rect 676288 245130 676352 245194
rect 675136 244302 675200 244306
rect 675136 244246 675188 244302
rect 675188 244246 675200 244302
rect 675136 244242 675200 244246
rect 675904 243502 675968 243566
rect 41728 243354 41792 243418
rect 145408 242022 145472 242086
rect 675520 241282 675584 241346
rect 42112 240750 42176 240754
rect 42112 240694 42124 240750
rect 42124 240694 42176 240750
rect 42112 240690 42176 240694
rect 42496 240690 42560 240754
rect 674560 239270 674624 239274
rect 674560 239214 674612 239270
rect 674612 239214 674624 239270
rect 674560 239210 674624 239214
rect 675328 239210 675392 239274
rect 675136 238974 675200 238978
rect 675136 238918 675188 238974
rect 675188 238918 675200 238974
rect 675136 238914 675200 238918
rect 674368 238618 674432 238682
rect 42496 237938 42560 237942
rect 42496 237882 42508 237938
rect 42508 237882 42560 237938
rect 42496 237878 42560 237882
rect 210304 237138 210368 237202
rect 676096 236842 676160 236906
rect 211456 234622 211520 234686
rect 212800 234030 212864 234094
rect 637504 234030 637568 234094
rect 211072 233882 211136 233946
rect 637696 233942 637760 233946
rect 637696 233886 637708 233942
rect 637708 233886 637760 233942
rect 637696 233882 637760 233886
rect 210496 233734 210560 233798
rect 212416 233734 212480 233798
rect 637120 233794 637184 233798
rect 637120 233738 637172 233794
rect 637172 233738 637184 233794
rect 210688 233586 210752 233650
rect 212032 233586 212096 233650
rect 637120 233734 637184 233738
rect 637312 233734 637376 233798
rect 636736 233586 636800 233650
rect 212224 233438 212288 233502
rect 636928 233438 636992 233502
rect 41344 233290 41408 233354
rect 210304 232994 210368 233058
rect 211456 232994 211520 233058
rect 212416 232846 212480 232910
rect 212992 232846 213056 232910
rect 41920 231722 41984 231726
rect 41920 231666 41932 231722
rect 41932 231666 41984 231722
rect 41920 231662 41984 231666
rect 41728 231130 41792 231134
rect 41728 231074 41780 231130
rect 41780 231074 41792 231130
rect 41728 231070 41792 231074
rect 42112 230538 42176 230542
rect 42112 230482 42124 230538
rect 42124 230482 42176 230538
rect 42112 230478 42176 230482
rect 41152 229590 41216 229654
rect 40960 228998 41024 229062
rect 40576 227518 40640 227582
rect 41536 227518 41600 227582
rect 40384 227222 40448 227286
rect 40768 226778 40832 226842
rect 675712 226778 675776 226842
rect 673984 226186 674048 226250
rect 40576 225890 40640 225954
rect 674368 223078 674432 223142
rect 145600 221746 145664 221810
rect 145792 218934 145856 218998
rect 675136 217750 675200 217814
rect 145984 216418 146048 216482
rect 40384 214642 40448 214706
rect 40576 213162 40640 213226
rect 40960 212422 41024 212486
rect 675136 211682 675200 211746
rect 41152 211534 41216 211598
rect 674752 211534 674816 211598
rect 675520 211534 675584 211598
rect 40768 210350 40832 210414
rect 676096 210202 676160 210266
rect 675520 210054 675584 210118
rect 676288 209906 676352 209970
rect 675904 209758 675968 209822
rect 675712 209610 675776 209674
rect 676480 209462 676544 209526
rect 210496 208722 210560 208786
rect 210880 208722 210944 208786
rect 210880 206354 210944 206418
rect 210880 205910 210944 205974
rect 675904 204282 675968 204346
rect 674752 199694 674816 199758
rect 675136 199162 675200 199166
rect 675136 199106 675188 199162
rect 675188 199106 675200 199162
rect 675136 199102 675200 199106
rect 675520 198422 675584 198426
rect 675520 198366 675532 198422
rect 675532 198366 675584 198422
rect 675520 198362 675584 198366
rect 42304 197622 42368 197686
rect 42112 197326 42176 197390
rect 675328 195698 675392 195762
rect 675520 195550 675584 195614
rect 42304 195166 42368 195170
rect 42304 195110 42356 195166
rect 42356 195110 42368 195166
rect 42304 195106 42368 195110
rect 676096 195254 676160 195318
rect 674368 193478 674432 193542
rect 676288 191554 676352 191618
rect 42112 191022 42176 191026
rect 42112 190966 42124 191022
rect 42124 190966 42176 191022
rect 42112 190962 42176 190966
rect 41152 190074 41216 190138
rect 41920 189098 41984 189102
rect 41920 189042 41932 189098
rect 41932 189042 41984 189098
rect 41920 189038 41984 189042
rect 41728 188358 41792 188362
rect 41728 188302 41780 188358
rect 41780 188302 41792 188358
rect 41728 188298 41792 188302
rect 40960 185930 41024 185994
rect 40384 184154 40448 184218
rect 40768 183562 40832 183626
rect 40576 182822 40640 182886
rect 210112 182674 210176 182738
rect 210880 182674 210944 182738
rect 673984 182526 674048 182590
rect 210304 181934 210368 181998
rect 210880 181934 210944 181998
rect 673984 181194 674048 181258
rect 675712 180898 675776 180962
rect 676480 179418 676544 179482
rect 674176 178086 674240 178150
rect 31744 177050 31808 177114
rect 674560 166394 674624 166458
rect 674368 165506 674432 165570
rect 676288 164026 676352 164090
rect 676672 163878 676736 163942
rect 676480 163582 676544 163646
rect 210688 161214 210752 161278
rect 675520 154614 675584 154618
rect 675520 154558 675532 154614
rect 675532 154558 675584 154614
rect 675520 154554 675584 154558
rect 210688 154258 210752 154322
rect 675136 154258 675200 154322
rect 210496 154110 210560 154174
rect 676288 153370 676352 153434
rect 210880 153222 210944 153286
rect 676480 150262 676544 150326
rect 674176 148486 674240 148550
rect 676672 146562 676736 146626
rect 210688 144046 210752 144110
rect 210496 143898 210560 143962
rect 673984 136794 674048 136858
rect 674560 135462 674624 135526
rect 674560 134870 674624 134934
rect 674368 134500 674432 134564
rect 674176 132872 674240 132936
rect 210304 126730 210368 126794
rect 210496 126730 210560 126794
rect 31744 125250 31808 125314
rect 675712 120366 675776 120430
rect 676672 117998 676736 118062
rect 674752 111338 674816 111402
rect 675520 110066 675584 110070
rect 675520 110010 675532 110066
rect 675532 110010 675584 110066
rect 675520 110006 675584 110010
rect 674752 109414 674816 109478
rect 675712 108142 675776 108146
rect 675712 108086 675724 108142
rect 675724 108086 675776 108142
rect 675712 108082 675776 108086
rect 144832 106602 144896 106666
rect 209920 105122 209984 105186
rect 210304 105122 210368 105186
rect 210112 103494 210176 103558
rect 210880 103494 210944 103558
rect 674176 103198 674240 103262
rect 210496 102310 210560 102374
rect 210880 102310 210944 102374
rect 676672 101422 676736 101486
rect 144832 100830 144896 100894
rect 209728 94762 209792 94826
rect 210880 94762 210944 94826
rect 210496 93726 210560 93790
rect 210880 93726 210944 93790
rect 210112 87806 210176 87870
rect 210880 87806 210944 87870
rect 210688 87658 210752 87722
rect 209920 86030 209984 86094
rect 210880 86030 210944 86094
rect 210112 84550 210176 84614
rect 210688 84550 210752 84614
rect 210304 83426 210368 83430
rect 210304 83370 210316 83426
rect 210316 83370 210368 83426
rect 210304 83366 210368 83370
rect 209728 82330 209792 82394
rect 210880 82330 210944 82394
rect 209920 71882 209984 71886
rect 209920 71826 209972 71882
rect 209972 71826 209984 71882
rect 209920 71822 209984 71826
rect 210880 58354 210944 58418
rect 210496 57170 210560 57234
rect 210880 55098 210944 55162
rect 210304 54418 210368 54422
rect 210304 54362 210356 54418
rect 210356 54362 210368 54418
rect 210304 54358 210368 54362
rect 210880 54358 210944 54422
rect 209920 54062 209984 54126
rect 210688 54062 210752 54126
rect 210496 53914 210560 53978
rect 212608 53766 212672 53830
rect 211456 53618 211520 53682
rect 211072 53470 211136 53534
rect 212992 53470 213056 53534
rect 210112 53174 210176 53238
rect 465664 53322 465728 53386
rect 211840 53026 211904 53090
rect 377536 53026 377600 53090
rect 377344 52878 377408 52942
rect 636736 52582 636800 52646
rect 637504 52434 637568 52498
rect 637120 52286 637184 52350
rect 637696 52138 637760 52202
rect 636928 51990 636992 52054
rect 637312 51842 637376 51906
rect 145984 51250 146048 51314
rect 145792 51102 145856 51166
rect 145408 50954 145472 51018
rect 145600 50806 145664 50870
rect 306688 48882 306752 48946
rect 356992 46070 357056 46134
rect 302464 45330 302528 45394
rect 360064 45182 360128 45246
rect 362944 45034 363008 45098
rect 409024 44886 409088 44950
rect 302464 43318 302528 43322
rect 302464 43262 302516 43318
rect 302516 43262 302528 43318
rect 302464 43258 302528 43262
rect 360064 43258 360128 43322
rect 362944 43258 363008 43322
rect 409024 43258 409088 43322
rect 306688 42134 306752 42138
rect 306688 42078 306740 42134
rect 306740 42078 306752 42134
rect 306688 42074 306752 42078
rect 356992 42074 357056 42138
rect 189952 41778 190016 41842
rect 194944 41778 195008 41842
rect 458176 41778 458240 41842
rect 465664 41838 465728 41842
rect 465664 41782 465716 41838
rect 465716 41782 465728 41838
rect 465664 41778 465728 41782
rect 189952 40742 190016 40806
rect 194944 40594 195008 40658
rect 457792 40358 457856 40362
rect 457792 40302 457804 40358
rect 457804 40302 457856 40358
rect 457792 40298 457856 40302
<< metal4 >>
rect 42111 968766 42177 968767
rect 42111 968702 42112 968766
rect 42176 968702 42177 968766
rect 42111 968701 42177 968702
rect 40383 967138 40449 967139
rect 40383 967074 40384 967138
rect 40448 967074 40449 967138
rect 40383 967073 40449 967074
rect 40386 943755 40446 967073
rect 40959 965066 41025 965067
rect 40959 965002 40960 965066
rect 41024 965002 41025 965066
rect 40959 965001 41025 965002
rect 40767 957814 40833 957815
rect 40767 957750 40768 957814
rect 40832 957750 40833 957814
rect 40767 957749 40833 957750
rect 40575 956186 40641 956187
rect 40575 956122 40576 956186
rect 40640 956122 40641 956186
rect 40575 956121 40641 956122
rect 40578 944495 40638 956121
rect 40575 944494 40641 944495
rect 40575 944430 40576 944494
rect 40640 944430 40641 944494
rect 40575 944429 40641 944430
rect 40383 943754 40449 943755
rect 40383 943690 40384 943754
rect 40448 943690 40449 943754
rect 40383 943689 40449 943690
rect 40770 941683 40830 957749
rect 40767 941682 40833 941683
rect 40767 941618 40768 941682
rect 40832 941618 40833 941682
rect 40767 941617 40833 941618
rect 40962 937391 41022 965001
rect 41343 963438 41409 963439
rect 41343 963374 41344 963438
rect 41408 963374 41409 963438
rect 41343 963373 41409 963374
rect 41151 959738 41217 959739
rect 41151 959674 41152 959738
rect 41216 959674 41217 959738
rect 41151 959673 41217 959674
rect 40959 937390 41025 937391
rect 40959 937326 40960 937390
rect 41024 937326 41025 937390
rect 40959 937325 41025 937326
rect 41154 935911 41214 959673
rect 41346 936503 41406 963373
rect 41727 962106 41793 962107
rect 41727 962042 41728 962106
rect 41792 962042 41793 962106
rect 41727 962041 41793 962042
rect 41535 959146 41601 959147
rect 41535 959082 41536 959146
rect 41600 959082 41601 959146
rect 41535 959081 41601 959082
rect 41538 938131 41598 959081
rect 41730 941239 41790 962041
rect 41919 958406 41985 958407
rect 41919 958342 41920 958406
rect 41984 958342 41985 958406
rect 41919 958341 41985 958342
rect 41727 941238 41793 941239
rect 41727 941174 41728 941238
rect 41792 941174 41793 941238
rect 41727 941173 41793 941174
rect 41922 938871 41982 958341
rect 42114 940647 42174 968701
rect 674367 966398 674433 966399
rect 674367 966334 674368 966398
rect 674432 966334 674433 966398
rect 674367 966333 674433 966334
rect 42495 964030 42561 964031
rect 42495 963966 42496 964030
rect 42560 963966 42561 964030
rect 42495 963965 42561 963966
rect 42303 962846 42369 962847
rect 42303 962782 42304 962846
rect 42368 962782 42369 962846
rect 42303 962781 42369 962782
rect 42111 940646 42177 940647
rect 42111 940582 42112 940646
rect 42176 940582 42177 940646
rect 42111 940581 42177 940582
rect 41919 938870 41985 938871
rect 41919 938806 41920 938870
rect 41984 938806 41985 938870
rect 41919 938805 41985 938806
rect 41535 938130 41601 938131
rect 41535 938066 41536 938130
rect 41600 938066 41601 938130
rect 41535 938065 41601 938066
rect 41343 936502 41409 936503
rect 41343 936438 41344 936502
rect 41408 936438 41409 936502
rect 41343 936437 41409 936438
rect 41151 935910 41217 935911
rect 41151 935846 41152 935910
rect 41216 935846 41217 935910
rect 41151 935845 41217 935846
rect 42306 935023 42366 962781
rect 42303 935022 42369 935023
rect 42303 934958 42304 935022
rect 42368 934958 42369 935022
rect 42303 934957 42369 934958
rect 42498 934135 42558 963965
rect 42879 953226 42945 953227
rect 42879 953162 42880 953226
rect 42944 953162 42945 953226
rect 42879 953161 42945 953162
rect 42687 947602 42753 947603
rect 42687 947538 42688 947602
rect 42752 947538 42753 947602
rect 42687 947537 42753 947538
rect 42690 947455 42750 947537
rect 42882 947455 42942 953161
rect 42687 947454 42753 947455
rect 42687 947390 42688 947454
rect 42752 947390 42753 947454
rect 42687 947389 42753 947390
rect 42879 947454 42945 947455
rect 42879 947390 42880 947454
rect 42944 947390 42945 947454
rect 42879 947389 42945 947390
rect 43071 947306 43137 947307
rect 43071 947242 43072 947306
rect 43136 947242 43137 947306
rect 43071 947241 43137 947242
rect 42687 944790 42753 944791
rect 42687 944726 42688 944790
rect 42752 944726 42753 944790
rect 42687 944725 42753 944726
rect 42495 934134 42561 934135
rect 42495 934070 42496 934134
rect 42560 934070 42561 934134
rect 42495 934069 42561 934070
rect 42495 912970 42561 912971
rect 42495 912906 42496 912970
rect 42560 912906 42561 912970
rect 42495 912905 42561 912906
rect 42498 907199 42558 912905
rect 42495 907198 42561 907199
rect 42495 907134 42496 907198
rect 42560 907134 42561 907198
rect 42495 907133 42561 907134
rect 42495 872566 42561 872567
rect 42495 872502 42496 872566
rect 42560 872502 42561 872566
rect 42495 872501 42561 872502
rect 42498 846815 42558 872501
rect 42495 846814 42561 846815
rect 42495 846750 42496 846814
rect 42560 846750 42561 846814
rect 42495 846749 42561 846750
rect 41919 832310 41985 832311
rect 41919 832246 41920 832310
rect 41984 832246 41985 832310
rect 41919 832245 41985 832246
rect 40767 818694 40833 818695
rect 40767 818630 40768 818694
rect 40832 818630 40833 818694
rect 40767 818629 40833 818630
rect 40383 802118 40449 802119
rect 40383 802054 40384 802118
rect 40448 802054 40449 802118
rect 40383 802053 40449 802054
rect 40386 776811 40446 802053
rect 40383 776810 40449 776811
rect 40383 776746 40384 776810
rect 40448 776746 40449 776810
rect 40383 776745 40449 776746
rect 40770 775183 40830 818629
rect 41922 816327 41982 832245
rect 42690 822873 42750 944725
rect 43074 937425 43134 947241
rect 674370 938723 674430 966333
rect 676479 965806 676545 965807
rect 676479 965742 676480 965806
rect 676544 965742 676545 965806
rect 676479 965741 676545 965742
rect 675903 965066 675969 965067
rect 675903 965002 675904 965066
rect 675968 965002 675969 965066
rect 675903 965001 675969 965002
rect 675327 963290 675393 963291
rect 675327 963226 675328 963290
rect 675392 963226 675393 963290
rect 675327 963225 675393 963226
rect 674751 962698 674817 962699
rect 674751 962634 674752 962698
rect 674816 962634 674817 962698
rect 674751 962633 674817 962634
rect 674559 962254 674625 962255
rect 674559 962190 674560 962254
rect 674624 962190 674625 962254
rect 674559 962189 674625 962190
rect 674367 938722 674433 938723
rect 674367 938658 674368 938722
rect 674432 938658 674433 938722
rect 674367 938657 674433 938658
rect 42114 822813 42750 822873
rect 42882 937365 43134 937425
rect 42114 819583 42174 822813
rect 42111 819582 42177 819583
rect 42111 819518 42112 819582
rect 42176 819518 42177 819582
rect 42111 819517 42177 819518
rect 41919 816326 41985 816327
rect 41919 816262 41920 816326
rect 41984 816262 41985 816326
rect 41919 816261 41985 816262
rect 42687 816326 42753 816327
rect 42687 816262 42688 816326
rect 42752 816262 42753 816326
rect 42687 816261 42753 816262
rect 42495 812034 42561 812035
rect 42495 811970 42496 812034
rect 42560 811970 42561 812034
rect 42495 811969 42561 811970
rect 42498 803599 42558 811969
rect 42495 803598 42561 803599
rect 42495 803534 42496 803598
rect 42560 803534 42561 803598
rect 42495 803533 42561 803534
rect 41343 802266 41409 802267
rect 41343 802202 41344 802266
rect 41408 802202 41409 802266
rect 41343 802201 41409 802202
rect 41346 791759 41406 802201
rect 41535 801970 41601 801971
rect 41535 801906 41536 801970
rect 41600 801906 41601 801970
rect 41535 801905 41601 801906
rect 41538 791907 41598 801905
rect 41727 800342 41793 800343
rect 41727 800278 41728 800342
rect 41792 800278 41793 800342
rect 41727 800277 41793 800278
rect 42495 800342 42561 800343
rect 42495 800278 42496 800342
rect 42560 800278 42561 800342
rect 42495 800277 42561 800278
rect 41730 794275 41790 800277
rect 42303 800046 42369 800047
rect 42303 799982 42304 800046
rect 42368 799982 42369 800046
rect 42303 799981 42369 799982
rect 42306 797975 42366 799981
rect 42303 797974 42369 797975
rect 42303 797910 42304 797974
rect 42368 797910 42369 797974
rect 42303 797909 42369 797910
rect 42498 794867 42558 800277
rect 42495 794866 42561 794867
rect 42495 794802 42496 794866
rect 42560 794802 42561 794866
rect 42495 794801 42561 794802
rect 41727 794274 41793 794275
rect 41727 794210 41728 794274
rect 41792 794210 41793 794274
rect 42690 794235 42750 816261
rect 42882 812035 42942 937365
rect 674562 934579 674622 962189
rect 674754 935319 674814 962633
rect 674943 957666 675009 957667
rect 674943 957602 674944 957666
rect 675008 957602 675009 957666
rect 674943 957601 675009 957602
rect 674751 935318 674817 935319
rect 674751 935254 674752 935318
rect 674816 935254 674817 935318
rect 674751 935253 674817 935254
rect 674559 934578 674625 934579
rect 674559 934514 674560 934578
rect 674624 934514 674625 934578
rect 674559 934513 674625 934514
rect 43071 933098 43137 933099
rect 43071 933034 43072 933098
rect 43136 933034 43137 933098
rect 43071 933033 43137 933034
rect 43074 912971 43134 933033
rect 674946 932951 675006 957601
rect 675135 956038 675201 956039
rect 675135 955974 675136 956038
rect 675200 955974 675201 956038
rect 675135 955973 675201 955974
rect 675138 933395 675198 955973
rect 675330 938427 675390 963225
rect 675711 960774 675777 960775
rect 675711 960710 675712 960774
rect 675776 960710 675777 960774
rect 675711 960709 675777 960710
rect 675519 960182 675585 960183
rect 675519 960118 675520 960182
rect 675584 960118 675585 960182
rect 675519 960117 675585 960118
rect 675327 938426 675393 938427
rect 675327 938362 675328 938426
rect 675392 938362 675393 938426
rect 675327 938361 675393 938362
rect 675135 933394 675201 933395
rect 675135 933330 675136 933394
rect 675200 933330 675201 933394
rect 675135 933329 675201 933330
rect 674943 932950 675009 932951
rect 674943 932886 674944 932950
rect 675008 932886 675009 932950
rect 674943 932885 675009 932886
rect 43071 912970 43137 912971
rect 43071 912906 43072 912970
rect 43136 912906 43137 912970
rect 43071 912905 43137 912906
rect 43071 887218 43137 887219
rect 43071 887154 43072 887218
rect 43136 887154 43137 887218
rect 43071 887153 43137 887154
rect 43074 872567 43134 887153
rect 674559 876414 674625 876415
rect 674559 876350 674560 876414
rect 674624 876350 674625 876414
rect 674559 876349 674625 876350
rect 674367 873454 674433 873455
rect 674367 873390 674368 873454
rect 674432 873390 674433 873454
rect 674367 873389 674433 873390
rect 674175 872862 674241 872863
rect 674175 872798 674176 872862
rect 674240 872798 674241 872862
rect 674175 872797 674241 872798
rect 43071 872566 43137 872567
rect 43071 872502 43072 872566
rect 43136 872502 43137 872566
rect 43071 872501 43137 872502
rect 43071 846814 43137 846815
rect 43071 846750 43072 846814
rect 43136 846750 43137 846814
rect 43071 846749 43137 846750
rect 43074 832311 43134 846749
rect 43071 832310 43137 832311
rect 43071 832246 43072 832310
rect 43136 832246 43137 832310
rect 43071 832245 43137 832246
rect 42879 812034 42945 812035
rect 42879 811970 42880 812034
rect 42944 811970 42945 812034
rect 42879 811969 42945 811970
rect 41727 794209 41793 794210
rect 42498 794175 42750 794235
rect 41535 791906 41601 791907
rect 41535 791842 41536 791906
rect 41600 791842 41601 791906
rect 41535 791841 41601 791842
rect 41343 791758 41409 791759
rect 41343 791694 41344 791758
rect 41408 791694 41409 791758
rect 41343 791693 41409 791694
rect 41727 791314 41793 791315
rect 41727 791250 41728 791314
rect 41792 791250 41793 791314
rect 41727 791249 41793 791250
rect 41343 775922 41409 775923
rect 41343 775858 41344 775922
rect 41408 775858 41409 775922
rect 41343 775857 41409 775858
rect 40767 775182 40833 775183
rect 40767 775118 40768 775182
rect 40832 775118 40833 775182
rect 40767 775117 40833 775118
rect 40383 758606 40449 758607
rect 40383 758542 40384 758606
rect 40448 758542 40449 758606
rect 40383 758541 40449 758542
rect 40386 747211 40446 758541
rect 40383 747210 40449 747211
rect 40383 747146 40384 747210
rect 40448 747146 40449 747210
rect 40383 747145 40449 747146
rect 40770 733151 40830 775117
rect 40959 760234 41025 760235
rect 40959 760170 40960 760234
rect 41024 760170 41025 760234
rect 40959 760169 41025 760170
rect 40962 746915 41022 760169
rect 40959 746914 41025 746915
rect 40959 746850 40960 746914
rect 41024 746850 41025 746914
rect 40959 746849 41025 746850
rect 41346 733891 41406 775857
rect 41535 764082 41601 764083
rect 41535 764018 41536 764082
rect 41600 764018 41601 764082
rect 41535 764017 41601 764018
rect 41538 751799 41598 764017
rect 41535 751798 41601 751799
rect 41535 751734 41536 751798
rect 41600 751734 41601 751798
rect 41535 751733 41601 751734
rect 41730 748691 41790 791249
rect 42498 791019 42558 794175
rect 41919 791018 41985 791019
rect 41919 790954 41920 791018
rect 41984 790954 41985 791018
rect 41919 790953 41985 790954
rect 42495 791018 42561 791019
rect 42495 790954 42496 791018
rect 42560 790954 42561 791018
rect 42495 790953 42561 790954
rect 41727 748690 41793 748691
rect 41727 748626 41728 748690
rect 41792 748626 41793 748690
rect 41727 748625 41793 748626
rect 41343 733890 41409 733891
rect 41343 733826 41344 733890
rect 41408 733826 41409 733890
rect 41343 733825 41409 733826
rect 40575 733150 40641 733151
rect 40575 733086 40576 733150
rect 40640 733086 40641 733150
rect 40575 733085 40641 733086
rect 40767 733150 40833 733151
rect 40767 733086 40768 733150
rect 40832 733086 40833 733150
rect 40767 733085 40833 733086
rect 40383 717018 40449 717019
rect 40383 716954 40384 717018
rect 40448 716954 40449 717018
rect 40383 716953 40449 716954
rect 40386 703551 40446 716953
rect 40383 703550 40449 703551
rect 40383 703486 40384 703550
rect 40448 703486 40449 703550
rect 40383 703485 40449 703486
rect 40578 690379 40638 733085
rect 40959 732262 41025 732263
rect 40959 732198 40960 732262
rect 41024 732198 41025 732262
rect 40959 732197 41025 732198
rect 40575 690378 40641 690379
rect 40575 690314 40576 690378
rect 40640 690314 40641 690378
rect 40575 690313 40641 690314
rect 40962 689639 41022 732197
rect 41343 720866 41409 720867
rect 41343 720802 41344 720866
rect 41408 720802 41409 720866
rect 41343 720801 41409 720802
rect 41151 716722 41217 716723
rect 41151 716658 41152 716722
rect 41216 716658 41217 716722
rect 41151 716657 41217 716658
rect 41154 703699 41214 716657
rect 41346 708583 41406 720801
rect 41535 716130 41601 716131
rect 41535 716066 41536 716130
rect 41600 716066 41601 716130
rect 41535 716065 41601 716066
rect 41343 708582 41409 708583
rect 41343 708518 41344 708582
rect 41408 708518 41409 708582
rect 41343 708517 41409 708518
rect 41538 706807 41598 716065
rect 41535 706806 41601 706807
rect 41535 706742 41536 706806
rect 41600 706742 41601 706806
rect 41535 706741 41601 706742
rect 41730 704735 41790 748625
rect 41922 747359 41982 790953
rect 673983 787466 674049 787467
rect 673983 787402 673984 787466
rect 674048 787402 674049 787466
rect 673983 787401 674049 787402
rect 42111 766006 42177 766007
rect 42111 765942 42112 766006
rect 42176 765942 42177 766006
rect 42111 765941 42177 765942
rect 42114 747507 42174 765941
rect 42879 751946 42945 751947
rect 42879 751882 42880 751946
rect 42944 751882 42945 751946
rect 42879 751881 42945 751882
rect 42882 751651 42942 751881
rect 42879 751650 42945 751651
rect 42879 751586 42880 751650
rect 42944 751586 42945 751650
rect 42879 751585 42945 751586
rect 42111 747506 42177 747507
rect 42111 747442 42112 747506
rect 42176 747442 42177 747506
rect 42111 747441 42177 747442
rect 41919 747358 41985 747359
rect 41919 747294 41920 747358
rect 41984 747294 41985 747358
rect 41919 747293 41985 747294
rect 41922 745879 41982 747293
rect 41919 745878 41985 745879
rect 41919 745814 41920 745878
rect 41984 745814 41985 745878
rect 41919 745813 41985 745814
rect 42111 745434 42177 745435
rect 42111 745370 42112 745434
rect 42176 745370 42177 745434
rect 42111 745369 42177 745370
rect 42114 735963 42174 745369
rect 42111 735962 42177 735963
rect 42111 735898 42112 735962
rect 42176 735898 42177 735962
rect 42111 735897 42177 735898
rect 42111 725898 42177 725899
rect 42111 725834 42112 725898
rect 42176 725834 42177 725898
rect 42111 725833 42177 725834
rect 41919 713910 41985 713911
rect 41919 713846 41920 713910
rect 41984 713846 41985 713910
rect 41919 713845 41985 713846
rect 41922 711691 41982 713845
rect 41919 711690 41985 711691
rect 41919 711626 41920 711690
rect 41984 711626 41985 711690
rect 41919 711625 41985 711626
rect 41343 704734 41409 704735
rect 41343 704670 41344 704734
rect 41408 704670 41409 704734
rect 41343 704669 41409 704670
rect 41727 704734 41793 704735
rect 41727 704670 41728 704734
rect 41792 704670 41793 704734
rect 41727 704669 41793 704670
rect 41151 703698 41217 703699
rect 41151 703634 41152 703698
rect 41216 703634 41217 703698
rect 41151 703633 41217 703634
rect 41346 692747 41406 704669
rect 42114 704143 42174 725833
rect 42687 723826 42753 723827
rect 42687 723762 42688 723826
rect 42752 723762 42753 723826
rect 42687 723761 42753 723762
rect 42303 722642 42369 722643
rect 42303 722578 42304 722642
rect 42368 722578 42369 722642
rect 42303 722577 42369 722578
rect 42306 706215 42366 722577
rect 42495 713910 42561 713911
rect 42495 713846 42496 713910
rect 42560 713846 42561 713910
rect 42495 713845 42561 713846
rect 42498 710803 42558 713845
rect 42495 710802 42561 710803
rect 42495 710738 42496 710802
rect 42560 710738 42561 710802
rect 42495 710737 42561 710738
rect 42690 707843 42750 723761
rect 673986 712135 674046 787401
rect 674178 755499 674238 872797
rect 674370 756387 674430 873389
rect 674562 760531 674622 876349
rect 674943 876266 675009 876267
rect 674943 876202 674944 876266
rect 675008 876202 675009 876266
rect 674943 876201 675009 876202
rect 674751 874046 674817 874047
rect 674751 873982 674752 874046
rect 674816 873982 674817 874046
rect 674751 873981 674817 873982
rect 674559 760530 674625 760531
rect 674559 760466 674560 760530
rect 674624 760466 674625 760530
rect 674559 760465 674625 760466
rect 674754 760087 674814 873981
rect 674946 762455 675006 876201
rect 675522 875823 675582 960117
rect 675519 875822 675585 875823
rect 675519 875758 675520 875822
rect 675584 875758 675585 875822
rect 675519 875757 675585 875758
rect 675714 875675 675774 960709
rect 675906 940943 675966 965001
rect 676095 961366 676161 961367
rect 676095 961302 676096 961366
rect 676160 961302 676161 961366
rect 676095 961301 676161 961302
rect 675903 940942 675969 940943
rect 675903 940878 675904 940942
rect 675968 940878 675969 940942
rect 675903 940877 675969 940878
rect 676098 932211 676158 961301
rect 676482 935911 676542 965741
rect 677055 953522 677121 953523
rect 677055 953458 677056 953522
rect 677120 953458 677121 953522
rect 677055 953457 677121 953458
rect 676863 953374 676929 953375
rect 676863 953310 676864 953374
rect 676928 953310 676929 953374
rect 676863 953309 676929 953310
rect 676479 935910 676545 935911
rect 676479 935846 676480 935910
rect 676544 935846 676545 935910
rect 676479 935845 676545 935846
rect 676095 932210 676161 932211
rect 676095 932146 676096 932210
rect 676160 932146 676161 932210
rect 676095 932145 676161 932146
rect 676866 930287 676926 953309
rect 677058 931471 677118 953457
rect 677055 931470 677121 931471
rect 677055 931406 677056 931470
rect 677120 931406 677121 931470
rect 677055 931405 677121 931406
rect 676863 930286 676929 930287
rect 676863 930222 676864 930286
rect 676928 930222 676929 930286
rect 676863 930221 676929 930222
rect 676095 876414 676161 876415
rect 676095 876350 676096 876414
rect 676160 876350 676161 876414
rect 676095 876349 676161 876350
rect 675711 875674 675777 875675
rect 675711 875610 675712 875674
rect 675776 875610 675777 875674
rect 675711 875609 675777 875610
rect 675327 869902 675393 869903
rect 675327 869838 675328 869902
rect 675392 869838 675393 869902
rect 675327 869837 675393 869838
rect 675135 866942 675201 866943
rect 675135 866878 675136 866942
rect 675200 866878 675201 866942
rect 675135 866877 675201 866878
rect 674943 762454 675009 762455
rect 674943 762390 674944 762454
rect 675008 762390 675009 762454
rect 674943 762389 675009 762390
rect 674751 760086 674817 760087
rect 674751 760022 674752 760086
rect 674816 760022 674817 760086
rect 674751 760021 674817 760022
rect 674367 756386 674433 756387
rect 674367 756322 674368 756386
rect 674432 756322 674433 756386
rect 674367 756321 674433 756322
rect 674175 755498 674241 755499
rect 674175 755434 674176 755498
rect 674240 755434 674241 755498
rect 674175 755433 674241 755434
rect 675138 755351 675198 866877
rect 675330 759199 675390 869837
rect 675711 864722 675777 864723
rect 675711 864658 675712 864722
rect 675776 864658 675777 864722
rect 675711 864657 675777 864658
rect 675519 862946 675585 862947
rect 675519 862882 675520 862946
rect 675584 862882 675585 862946
rect 675519 862881 675585 862882
rect 675327 759198 675393 759199
rect 675327 759134 675328 759198
rect 675392 759134 675393 759198
rect 675327 759133 675393 759134
rect 675522 758607 675582 862881
rect 675714 761715 675774 864657
rect 675903 784210 675969 784211
rect 675903 784146 675904 784210
rect 675968 784146 675969 784210
rect 675903 784145 675969 784146
rect 675711 761714 675777 761715
rect 675711 761650 675712 761714
rect 675776 761650 675777 761714
rect 675711 761649 675777 761650
rect 675519 758606 675585 758607
rect 675519 758542 675520 758606
rect 675584 758542 675585 758606
rect 675519 758541 675585 758542
rect 675135 755350 675201 755351
rect 675135 755286 675136 755350
rect 675200 755286 675201 755350
rect 675135 755285 675201 755286
rect 674559 743362 674625 743363
rect 674559 743298 674560 743362
rect 674624 743298 674625 743362
rect 674559 743297 674625 743298
rect 674175 742178 674241 742179
rect 674175 742114 674176 742178
rect 674240 742114 674241 742178
rect 674175 742113 674241 742114
rect 673983 712134 674049 712135
rect 673983 712070 673984 712134
rect 674048 712070 674049 712134
rect 673983 712069 674049 712070
rect 42687 707842 42753 707843
rect 42687 707778 42688 707842
rect 42752 707778 42753 707842
rect 42687 707777 42753 707778
rect 42303 706214 42369 706215
rect 42303 706150 42304 706214
rect 42368 706150 42369 706214
rect 42303 706149 42369 706150
rect 41535 704142 41601 704143
rect 41535 704078 41536 704142
rect 41600 704078 41601 704142
rect 41535 704077 41601 704078
rect 42111 704142 42177 704143
rect 42111 704078 42112 704142
rect 42176 704078 42177 704142
rect 42111 704077 42177 704078
rect 41343 692746 41409 692747
rect 41343 692682 41344 692746
rect 41408 692682 41409 692746
rect 41343 692681 41409 692682
rect 41538 690339 41598 704077
rect 673983 697334 674049 697335
rect 673983 697270 673984 697334
rect 674048 697270 674049 697334
rect 673983 697269 674049 697270
rect 41538 690279 42750 690339
rect 40959 689638 41025 689639
rect 40959 689574 40960 689638
rect 41024 689574 41025 689638
rect 40959 689573 41025 689574
rect 42303 689638 42369 689639
rect 42303 689574 42304 689638
rect 42368 689574 42369 689638
rect 42303 689573 42369 689574
rect 42111 688750 42177 688751
rect 42111 688686 42112 688750
rect 42176 688686 42177 688750
rect 42111 688685 42177 688686
rect 40575 686382 40641 686383
rect 40575 686318 40576 686382
rect 40640 686318 40641 686382
rect 40575 686317 40641 686318
rect 40578 656191 40638 686317
rect 40959 683274 41025 683275
rect 40959 683210 40960 683274
rect 41024 683210 41025 683274
rect 40959 683209 41025 683210
rect 40962 656783 41022 683209
rect 41727 680906 41793 680907
rect 41727 680842 41728 680906
rect 41792 680842 41793 680906
rect 41727 680841 41793 680842
rect 41343 670990 41409 670991
rect 41343 670926 41344 670990
rect 41408 670926 41409 670990
rect 41343 670925 41409 670926
rect 41346 665515 41406 670925
rect 41730 666699 41790 680841
rect 41919 670842 41985 670843
rect 41919 670778 41920 670842
rect 41984 670778 41985 670842
rect 41919 670777 41985 670778
rect 41727 666698 41793 666699
rect 41727 666634 41728 666698
rect 41792 666634 41793 666698
rect 41727 666633 41793 666634
rect 41343 665514 41409 665515
rect 41343 665450 41344 665514
rect 41408 665450 41409 665514
rect 41343 665449 41409 665450
rect 41535 665366 41601 665367
rect 41535 665302 41536 665366
rect 41600 665302 41601 665366
rect 41535 665301 41601 665302
rect 41538 665071 41598 665301
rect 41535 665070 41601 665071
rect 41535 665006 41536 665070
rect 41600 665006 41601 665070
rect 41535 665005 41601 665006
rect 41922 660779 41982 670777
rect 41919 660778 41985 660779
rect 41919 660714 41920 660778
rect 41984 660714 41985 660778
rect 41919 660713 41985 660714
rect 40959 656782 41025 656783
rect 40959 656718 40960 656782
rect 41024 656718 41025 656782
rect 40959 656717 41025 656718
rect 40575 656190 40641 656191
rect 40575 656126 40576 656190
rect 40640 656126 40641 656190
rect 40575 656125 40641 656126
rect 40575 643166 40641 643167
rect 40575 643102 40576 643166
rect 40640 643102 40641 643166
rect 40575 643101 40641 643102
rect 40578 618155 40638 643101
rect 40767 640058 40833 640059
rect 40767 639994 40768 640058
rect 40832 639994 40833 640058
rect 40767 639993 40833 639994
rect 40770 618303 40830 639993
rect 41922 627735 41982 660713
rect 42114 646719 42174 688685
rect 42306 647459 42366 689573
rect 42495 678390 42561 678391
rect 42495 678326 42496 678390
rect 42560 678326 42561 678390
rect 42495 678325 42561 678326
rect 42498 668771 42558 678325
rect 42690 670843 42750 690279
rect 42879 670990 42945 670991
rect 42879 670926 42880 670990
rect 42944 670926 42945 670990
rect 42879 670925 42945 670926
rect 42687 670842 42753 670843
rect 42687 670778 42688 670842
rect 42752 670778 42753 670842
rect 42687 670777 42753 670778
rect 42687 670694 42753 670695
rect 42687 670630 42688 670694
rect 42752 670630 42753 670694
rect 42687 670629 42753 670630
rect 42495 668770 42561 668771
rect 42495 668706 42496 668770
rect 42560 668706 42561 668770
rect 42495 668705 42561 668706
rect 42690 666551 42750 670629
rect 42687 666550 42753 666551
rect 42687 666486 42688 666550
rect 42752 666486 42753 666550
rect 42687 666485 42753 666486
rect 42687 665070 42753 665071
rect 42687 665006 42688 665070
rect 42752 665006 42753 665070
rect 42687 665005 42753 665006
rect 42690 661519 42750 665005
rect 42882 664775 42942 670925
rect 42879 664774 42945 664775
rect 42879 664710 42880 664774
rect 42944 664710 42945 664774
rect 42879 664709 42945 664710
rect 42687 661518 42753 661519
rect 42687 661454 42688 661518
rect 42752 661454 42753 661518
rect 42687 661453 42753 661454
rect 42303 647458 42369 647459
rect 42303 647394 42304 647458
rect 42368 647394 42369 647458
rect 42303 647393 42369 647394
rect 42111 646718 42177 646719
rect 42111 646654 42112 646718
rect 42176 646654 42177 646718
rect 42111 646653 42177 646654
rect 42303 637690 42369 637691
rect 42303 637626 42304 637690
rect 42368 637626 42369 637690
rect 42303 637625 42369 637626
rect 41730 627675 41982 627735
rect 40767 618302 40833 618303
rect 40767 618238 40768 618302
rect 40832 618238 40833 618302
rect 40767 618237 40833 618238
rect 40575 618154 40641 618155
rect 40575 618090 40576 618154
rect 40640 618090 40641 618154
rect 40575 618089 40641 618090
rect 41730 617859 41790 627675
rect 41919 627478 41985 627479
rect 41919 627414 41920 627478
rect 41984 627414 41985 627478
rect 41919 627413 41985 627414
rect 42111 627478 42177 627479
rect 42111 627414 42112 627478
rect 42176 627414 42177 627478
rect 42111 627413 42177 627414
rect 41922 623335 41982 627413
rect 41919 623334 41985 623335
rect 41919 623270 41920 623334
rect 41984 623270 41985 623334
rect 41919 623269 41985 623270
rect 42114 620227 42174 627413
rect 42306 623483 42366 637625
rect 42690 623927 42750 661453
rect 43071 627922 43137 627923
rect 43071 627858 43072 627922
rect 43136 627858 43137 627922
rect 43071 627857 43137 627858
rect 42687 623926 42753 623927
rect 42687 623862 42688 623926
rect 42752 623862 42753 623926
rect 42687 623861 42753 623862
rect 42303 623482 42369 623483
rect 42303 623418 42304 623482
rect 42368 623418 42369 623482
rect 42303 623417 42369 623418
rect 43074 620819 43134 627857
rect 673986 622003 674046 697269
rect 674178 689491 674238 742113
rect 674367 740106 674433 740107
rect 674367 740042 674368 740106
rect 674432 740042 674433 740106
rect 674367 740041 674433 740042
rect 674175 689490 674241 689491
rect 674175 689426 674176 689490
rect 674240 689426 674241 689490
rect 674175 689425 674241 689426
rect 674175 679722 674241 679723
rect 674175 679658 674176 679722
rect 674240 679658 674241 679722
rect 674175 679657 674241 679658
rect 674178 679575 674238 679657
rect 674175 679574 674241 679575
rect 674175 679510 674176 679574
rect 674240 679510 674241 679574
rect 674175 679509 674241 679510
rect 674370 669289 674430 740041
rect 674562 670547 674622 743297
rect 674751 740254 674817 740255
rect 674751 740190 674752 740254
rect 674816 740190 674817 740254
rect 674751 740189 674817 740190
rect 674754 672323 674814 740189
rect 675519 739218 675585 739219
rect 675519 739154 675520 739218
rect 675584 739154 675585 739218
rect 675519 739153 675585 739154
rect 674943 737738 675009 737739
rect 674943 737674 674944 737738
rect 675008 737674 675009 737738
rect 674943 737673 675009 737674
rect 674946 694375 675006 737673
rect 675135 734186 675201 734187
rect 675135 734122 675136 734186
rect 675200 734122 675201 734186
rect 675135 734121 675201 734122
rect 674943 694374 675009 694375
rect 674943 694310 674944 694374
rect 675008 694310 675009 694374
rect 674943 694309 675009 694310
rect 674943 693486 675009 693487
rect 674943 693422 674944 693486
rect 675008 693422 675009 693486
rect 674943 693421 675009 693422
rect 674946 679575 675006 693421
rect 674943 679574 675009 679575
rect 674943 679510 674944 679574
rect 675008 679510 675009 679574
rect 674943 679509 675009 679510
rect 674943 675430 675009 675431
rect 674943 675366 674944 675430
rect 675008 675366 675009 675430
rect 674943 675365 675009 675366
rect 674751 672322 674817 672323
rect 674751 672258 674752 672322
rect 674816 672258 674817 672322
rect 674751 672257 674817 672258
rect 674751 671582 674817 671583
rect 674751 671518 674752 671582
rect 674816 671518 674817 671582
rect 674751 671517 674817 671518
rect 674559 670546 674625 670547
rect 674559 670482 674560 670546
rect 674624 670482 674625 670546
rect 674559 670481 674625 670482
rect 674559 670398 674625 670399
rect 674559 670334 674560 670398
rect 674624 670334 674625 670398
rect 674559 670333 674625 670334
rect 674367 669288 674433 669289
rect 674367 669224 674368 669288
rect 674432 669224 674433 669288
rect 674367 669223 674433 669224
rect 674175 652194 674241 652195
rect 674175 652130 674176 652194
rect 674240 652130 674241 652194
rect 674175 652129 674241 652130
rect 673983 622002 674049 622003
rect 673983 621938 673984 622002
rect 674048 621938 674049 622002
rect 673983 621937 674049 621938
rect 43071 620818 43137 620819
rect 43071 620754 43072 620818
rect 43136 620754 43137 620818
rect 43071 620753 43137 620754
rect 42111 620226 42177 620227
rect 42111 620162 42112 620226
rect 42176 620162 42177 620226
rect 42111 620161 42177 620162
rect 41919 618450 41985 618451
rect 41919 618386 41920 618450
rect 41984 618386 41985 618450
rect 41919 618385 41985 618386
rect 41727 617858 41793 617859
rect 41727 617794 41728 617858
rect 41792 617794 41793 617858
rect 41727 617793 41793 617794
rect 40575 599950 40641 599951
rect 40575 599886 40576 599950
rect 40640 599886 40641 599950
rect 40575 599885 40641 599886
rect 40578 573903 40638 599885
rect 40959 596842 41025 596843
rect 40959 596778 40960 596842
rect 41024 596778 41025 596842
rect 40959 596777 41025 596778
rect 40962 574051 41022 596777
rect 41535 584262 41601 584263
rect 41535 584198 41536 584262
rect 41600 584198 41601 584262
rect 41535 584197 41601 584198
rect 41538 577159 41598 584197
rect 41535 577158 41601 577159
rect 41535 577094 41536 577158
rect 41600 577094 41601 577158
rect 41535 577093 41601 577094
rect 41730 574643 41790 617793
rect 41922 575235 41982 618385
rect 673983 607498 674049 607499
rect 673983 607434 673984 607498
rect 674048 607434 674049 607498
rect 673983 607433 674049 607434
rect 42879 585446 42945 585447
rect 42879 585382 42880 585446
rect 42944 585382 42945 585446
rect 42879 585381 42945 585382
rect 42495 584706 42561 584707
rect 42495 584642 42496 584706
rect 42560 584642 42561 584706
rect 42495 584641 42561 584642
rect 42303 584262 42369 584263
rect 42303 584198 42304 584262
rect 42368 584198 42369 584262
rect 42303 584197 42369 584198
rect 42306 580119 42366 584197
rect 42303 580118 42369 580119
rect 42303 580054 42304 580118
rect 42368 580054 42369 580118
rect 42303 580053 42369 580054
rect 42498 575975 42558 584641
rect 42882 578343 42942 585381
rect 42879 578342 42945 578343
rect 42879 578278 42880 578342
rect 42944 578278 42945 578342
rect 42879 578277 42945 578278
rect 42495 575974 42561 575975
rect 42495 575910 42496 575974
rect 42560 575910 42561 575974
rect 42495 575909 42561 575910
rect 41919 575234 41985 575235
rect 41919 575170 41920 575234
rect 41984 575170 41985 575234
rect 41919 575169 41985 575170
rect 41727 574642 41793 574643
rect 41727 574578 41728 574642
rect 41792 574578 41793 574642
rect 41727 574577 41793 574578
rect 40959 574050 41025 574051
rect 40959 573986 40960 574050
rect 41024 573986 41025 574050
rect 40959 573985 41025 573986
rect 40575 573902 40641 573903
rect 40575 573838 40576 573902
rect 40640 573838 40641 573902
rect 40575 573837 40641 573838
rect 41151 544302 41217 544303
rect 41151 544238 41152 544302
rect 41216 544238 41217 544302
rect 41151 544237 41217 544238
rect 40959 542970 41025 542971
rect 40959 542906 40960 542970
rect 41024 542906 41025 542970
rect 40959 542905 41025 542906
rect 40962 532611 41022 542905
rect 40959 532610 41025 532611
rect 40959 532546 40960 532610
rect 41024 532546 41025 532610
rect 40959 532545 41025 532546
rect 41154 532315 41214 544237
rect 41151 532314 41217 532315
rect 41151 532250 41152 532314
rect 41216 532250 41217 532314
rect 41151 532249 41217 532250
rect 41730 531279 41790 574577
rect 41922 532019 41982 575169
rect 42111 541342 42177 541343
rect 42111 541278 42112 541342
rect 42176 541278 42177 541342
rect 42111 541277 42177 541278
rect 42114 538827 42174 541277
rect 42879 541194 42945 541195
rect 42879 541130 42880 541194
rect 42944 541130 42945 541194
rect 42879 541129 42945 541130
rect 42111 538826 42177 538827
rect 42111 538762 42112 538826
rect 42176 538762 42177 538826
rect 42111 538761 42177 538762
rect 42882 536903 42942 541129
rect 43071 541046 43137 541047
rect 43071 540982 43072 541046
rect 43136 540982 43137 541046
rect 43071 540981 43137 540982
rect 42879 536902 42945 536903
rect 42879 536838 42880 536902
rect 42944 536838 42945 536902
rect 42879 536837 42945 536838
rect 43074 535719 43134 540981
rect 43071 535718 43137 535719
rect 43071 535654 43072 535718
rect 43136 535654 43137 535718
rect 43071 535653 43137 535654
rect 41919 532018 41985 532019
rect 41919 531954 41920 532018
rect 41984 531954 41985 532018
rect 41919 531953 41985 531954
rect 41727 531278 41793 531279
rect 41727 531214 41728 531278
rect 41792 531214 41793 531278
rect 41727 531213 41793 531214
rect 40575 432710 40641 432711
rect 40575 432646 40576 432710
rect 40640 432646 40641 432710
rect 40575 432645 40641 432646
rect 40383 431970 40449 431971
rect 40383 431906 40384 431970
rect 40448 431906 40449 431970
rect 40383 431905 40449 431906
rect 40386 389199 40446 431905
rect 40578 390235 40638 432645
rect 40767 430786 40833 430787
rect 40767 430722 40768 430786
rect 40832 430722 40833 430786
rect 40767 430721 40833 430722
rect 40770 400151 40830 430721
rect 40959 429454 41025 429455
rect 40959 429390 40960 429454
rect 41024 429390 41025 429454
rect 40959 429389 41025 429390
rect 40767 400150 40833 400151
rect 40767 400086 40768 400150
rect 40832 400086 40833 400150
rect 40767 400085 40833 400086
rect 40962 398819 41022 429389
rect 41343 428418 41409 428419
rect 41343 428354 41344 428418
rect 41408 428354 41409 428418
rect 41343 428353 41409 428354
rect 41151 426346 41217 426347
rect 41151 426282 41152 426346
rect 41216 426282 41217 426346
rect 41151 426281 41217 426282
rect 41154 399559 41214 426281
rect 41346 401927 41406 428353
rect 41535 427678 41601 427679
rect 41535 427614 41536 427678
rect 41600 427614 41601 427678
rect 41535 427613 41601 427614
rect 41538 406071 41598 427613
rect 41535 406070 41601 406071
rect 41535 406006 41536 406070
rect 41600 406006 41601 406070
rect 41535 406005 41601 406006
rect 41730 403851 41790 531213
rect 41922 404887 41982 531953
rect 673986 531723 674046 607433
rect 674178 576789 674238 652129
rect 674367 645386 674433 645387
rect 674367 645322 674368 645386
rect 674432 645322 674433 645386
rect 674367 645321 674433 645322
rect 674370 578417 674430 645321
rect 674562 641055 674622 670333
rect 674754 658411 674814 671517
rect 674751 658410 674817 658411
rect 674751 658346 674752 658410
rect 674816 658346 674817 658410
rect 674751 658345 674817 658346
rect 674946 657705 675006 675365
rect 675138 671287 675198 734121
rect 675522 711651 675582 739153
rect 675906 711987 675966 784145
rect 676098 757423 676158 876349
rect 676287 787910 676353 787911
rect 676287 787846 676288 787910
rect 676352 787846 676353 787910
rect 676287 787845 676353 787846
rect 676095 757422 676161 757423
rect 676095 757358 676096 757422
rect 676160 757358 676161 757422
rect 676095 757357 676161 757358
rect 676095 738774 676161 738775
rect 676095 738710 676096 738774
rect 676160 738710 676161 738774
rect 676095 738709 676161 738710
rect 675903 711986 675969 711987
rect 675903 711922 675904 711986
rect 675968 711922 675969 711986
rect 675903 711921 675969 711922
rect 675522 711591 675966 711651
rect 675906 703107 675966 711591
rect 675903 703106 675969 703107
rect 675903 703042 675904 703106
rect 675968 703042 675969 703106
rect 675903 703041 675969 703042
rect 676098 702515 676158 738709
rect 676290 715835 676350 787845
rect 676479 786726 676545 786727
rect 676479 786662 676480 786726
rect 676544 786662 676545 786726
rect 676479 786661 676545 786662
rect 676482 717167 676542 786661
rect 676671 781990 676737 781991
rect 676671 781926 676672 781990
rect 676736 781926 676737 781990
rect 676671 781925 676737 781926
rect 676674 737739 676734 781925
rect 677055 780510 677121 780511
rect 677055 780446 677056 780510
rect 677120 780446 677121 780510
rect 677055 780445 677121 780446
rect 677058 780249 677118 780445
rect 677058 780189 677310 780249
rect 677055 777550 677121 777551
rect 677055 777486 677056 777550
rect 677120 777486 677121 777550
rect 677055 777485 677121 777486
rect 676863 777402 676929 777403
rect 676863 777338 676864 777402
rect 676928 777338 676929 777402
rect 676863 777337 676929 777338
rect 676866 773111 676926 777337
rect 676863 773110 676929 773111
rect 676863 773046 676864 773110
rect 676928 773046 676929 773110
rect 676863 773045 676929 773046
rect 676863 772962 676929 772963
rect 676863 772898 676864 772962
rect 676928 772898 676929 772962
rect 676863 772897 676929 772898
rect 676866 754463 676926 772897
rect 676863 754462 676929 754463
rect 676863 754398 676864 754462
rect 676928 754398 676929 754462
rect 676863 754397 676929 754398
rect 676671 737738 676737 737739
rect 676671 737674 676672 737738
rect 676736 737674 676737 737738
rect 676671 737673 676737 737674
rect 676863 734926 676929 734927
rect 676863 734862 676864 734926
rect 676928 734862 676929 734926
rect 676863 734861 676929 734862
rect 676479 717166 676545 717167
rect 676479 717102 676480 717166
rect 676544 717102 676545 717166
rect 676479 717101 676545 717102
rect 676287 715834 676353 715835
rect 676287 715770 676288 715834
rect 676352 715770 676353 715834
rect 676287 715769 676353 715770
rect 676287 703106 676353 703107
rect 676287 703042 676288 703106
rect 676352 703042 676353 703106
rect 676287 703041 676353 703042
rect 676095 702514 676161 702515
rect 676095 702450 676096 702514
rect 676160 702450 676161 702514
rect 676095 702449 676161 702450
rect 676290 702327 676350 703041
rect 676098 702267 676350 702327
rect 675327 697926 675393 697927
rect 675327 697862 675328 697926
rect 675392 697862 675393 697926
rect 675327 697861 675393 697862
rect 675330 675431 675390 697861
rect 675903 697186 675969 697187
rect 675903 697122 675904 697186
rect 675968 697122 675969 697186
rect 675903 697121 675969 697122
rect 675519 694818 675585 694819
rect 675519 694754 675520 694818
rect 675584 694754 675585 694818
rect 675519 694753 675585 694754
rect 675327 675430 675393 675431
rect 675327 675366 675328 675430
rect 675392 675366 675393 675430
rect 675327 675365 675393 675366
rect 675135 671286 675201 671287
rect 675135 671222 675136 671286
rect 675200 671222 675201 671286
rect 675135 671221 675201 671222
rect 675135 670694 675201 670695
rect 675135 670630 675136 670694
rect 675200 670630 675201 670694
rect 675135 670629 675201 670630
rect 675327 670694 675393 670695
rect 675327 670630 675328 670694
rect 675392 670630 675393 670694
rect 675327 670629 675393 670630
rect 675138 664331 675198 670629
rect 675135 664330 675201 664331
rect 675135 664266 675136 664330
rect 675200 664266 675201 664330
rect 675135 664265 675201 664266
rect 674754 657645 675006 657705
rect 674754 641243 674814 657645
rect 675135 651454 675201 651455
rect 675135 651390 675136 651454
rect 675200 651390 675201 651454
rect 675135 651389 675201 651390
rect 674943 648050 675009 648051
rect 674943 647986 674944 648050
rect 675008 647986 675009 648050
rect 674943 647985 675009 647986
rect 674751 641242 674817 641243
rect 674751 641178 674752 641242
rect 674816 641178 674817 641242
rect 674751 641177 674817 641178
rect 674562 640995 674814 641055
rect 674559 640650 674625 640651
rect 674559 640586 674560 640650
rect 674624 640586 674625 640650
rect 674559 640585 674625 640586
rect 674367 578416 674433 578417
rect 674367 578352 674368 578416
rect 674432 578352 674433 578416
rect 674367 578351 674433 578352
rect 674175 576788 674241 576789
rect 674175 576724 674176 576788
rect 674240 576724 674241 576788
rect 674175 576723 674241 576724
rect 674562 576123 674622 640585
rect 674754 619191 674814 640995
rect 674946 640651 675006 647985
rect 674943 640650 675009 640651
rect 674943 640586 674944 640650
rect 675008 640586 675009 640650
rect 674943 640585 675009 640586
rect 674943 640206 675009 640207
rect 674943 640142 674944 640206
rect 675008 640142 675009 640206
rect 674943 640141 675009 640142
rect 674946 620967 675006 640141
rect 674943 620966 675009 620967
rect 674943 620902 674944 620966
rect 675008 620902 675009 620966
rect 674943 620901 675009 620902
rect 674751 619190 674817 619191
rect 674751 619126 674752 619190
rect 674816 619126 674817 619190
rect 674751 619125 674817 619126
rect 674751 607794 674817 607795
rect 674751 607730 674752 607794
rect 674816 607730 674817 607794
rect 674751 607729 674817 607730
rect 674559 576122 674625 576123
rect 674559 576058 674560 576122
rect 674624 576058 674625 576122
rect 674559 576057 674625 576058
rect 674175 561766 674241 561767
rect 674175 561702 674176 561766
rect 674240 561702 674241 561766
rect 674175 561701 674241 561702
rect 673983 531722 674049 531723
rect 673983 531658 673984 531722
rect 674048 531658 674049 531722
rect 673983 531657 674049 531658
rect 674178 487767 674238 561701
rect 674559 561618 674625 561619
rect 674559 561554 674560 561618
rect 674624 561554 674625 561618
rect 674559 561553 674625 561554
rect 674367 557770 674433 557771
rect 674367 557706 674368 557770
rect 674432 557706 674433 557770
rect 674367 557705 674433 557706
rect 674175 487766 674241 487767
rect 674175 487702 674176 487766
rect 674240 487702 674241 487766
rect 674175 487701 674241 487702
rect 674370 483845 674430 557705
rect 674562 492355 674622 561553
rect 674754 535423 674814 607729
rect 674943 604834 675009 604835
rect 674943 604770 674944 604834
rect 675008 604770 675009 604834
rect 674943 604769 675009 604770
rect 674751 535422 674817 535423
rect 674751 535358 674752 535422
rect 674816 535358 674817 535422
rect 674751 535357 674817 535358
rect 674946 534683 675006 604769
rect 675138 581747 675198 651389
rect 675330 640947 675390 670629
rect 675522 642575 675582 694753
rect 675711 689490 675777 689491
rect 675711 689426 675712 689490
rect 675776 689426 675777 689490
rect 675711 689425 675777 689426
rect 675714 667587 675774 689425
rect 675906 679575 675966 697121
rect 675903 679574 675969 679575
rect 675903 679510 675904 679574
rect 675968 679510 675969 679574
rect 675903 679509 675969 679510
rect 675711 667586 675777 667587
rect 675711 667522 675712 667586
rect 675776 667522 675777 667586
rect 675711 667521 675777 667522
rect 676098 666699 676158 702267
rect 676671 694374 676737 694375
rect 676671 694310 676672 694374
rect 676736 694310 676737 694374
rect 676671 694309 676737 694310
rect 676287 692006 676353 692007
rect 676287 691942 676288 692006
rect 676352 691942 676353 692006
rect 676287 691941 676353 691942
rect 676095 666698 676161 666699
rect 676095 666634 676096 666698
rect 676160 666634 676161 666698
rect 676095 666633 676161 666634
rect 675903 652638 675969 652639
rect 675903 652574 675904 652638
rect 675968 652574 675969 652638
rect 675903 652573 675969 652574
rect 675519 642574 675585 642575
rect 675519 642510 675520 642574
rect 675584 642510 675585 642574
rect 675519 642509 675585 642510
rect 675906 642387 675966 652573
rect 676290 651011 676350 691941
rect 676479 679722 676545 679723
rect 676479 679658 676480 679722
rect 676544 679658 676545 679722
rect 676479 679657 676545 679658
rect 676482 665959 676542 679657
rect 676479 665958 676545 665959
rect 676479 665894 676480 665958
rect 676544 665894 676545 665958
rect 676479 665893 676545 665894
rect 676479 658410 676545 658411
rect 676479 658346 676480 658410
rect 676544 658346 676545 658410
rect 676479 658345 676545 658346
rect 676287 651010 676353 651011
rect 676287 650946 676288 651010
rect 676352 650946 676353 651010
rect 676287 650945 676353 650946
rect 676095 649678 676161 649679
rect 676095 649614 676096 649678
rect 676160 649614 676161 649678
rect 676095 649613 676161 649614
rect 675522 642327 675966 642387
rect 675522 641055 675582 642327
rect 675522 640995 675774 641055
rect 675327 640946 675393 640947
rect 675327 640882 675328 640946
rect 675392 640882 675393 640946
rect 675327 640881 675393 640882
rect 675519 640798 675585 640799
rect 675519 640734 675520 640798
rect 675584 640734 675585 640798
rect 675519 640733 675585 640734
rect 675327 638578 675393 638579
rect 675327 638514 675328 638578
rect 675392 638514 675393 638578
rect 675327 638513 675393 638514
rect 675135 581746 675201 581747
rect 675135 581682 675136 581746
rect 675200 581682 675201 581746
rect 675135 581681 675201 581682
rect 675330 578195 675390 638513
rect 675522 625703 675582 640733
rect 675519 625702 675585 625703
rect 675519 625638 675520 625702
rect 675584 625638 675585 625702
rect 675519 625637 675585 625638
rect 675519 606462 675585 606463
rect 675519 606398 675520 606462
rect 675584 606398 675585 606462
rect 675519 606397 675585 606398
rect 675327 578194 675393 578195
rect 675327 578130 675328 578194
rect 675392 578130 675393 578194
rect 675327 578129 675393 578130
rect 675327 562950 675393 562951
rect 675327 562886 675328 562950
rect 675392 562886 675393 562950
rect 675327 562885 675393 562886
rect 675135 558954 675201 558955
rect 675135 558890 675136 558954
rect 675200 558890 675201 558954
rect 675135 558889 675201 558890
rect 674943 534682 675009 534683
rect 674943 534618 674944 534682
rect 675008 534618 675009 534682
rect 674943 534617 675009 534618
rect 674559 492354 674625 492355
rect 674559 492290 674560 492354
rect 674624 492290 674625 492354
rect 674559 492289 674625 492290
rect 675138 487471 675198 558889
rect 675330 491467 675390 562885
rect 675522 537051 675582 606397
rect 675714 580415 675774 640995
rect 675903 640946 675969 640947
rect 675903 640882 675904 640946
rect 675968 640882 675969 640946
rect 675903 640881 675969 640882
rect 675906 627331 675966 640881
rect 675903 627330 675969 627331
rect 675903 627266 675904 627330
rect 675968 627266 675969 627330
rect 675903 627265 675969 627266
rect 675903 600246 675969 600247
rect 675903 600182 675904 600246
rect 675968 600182 675969 600246
rect 675903 600181 675969 600182
rect 675711 580414 675777 580415
rect 675711 580350 675712 580414
rect 675776 580350 675777 580414
rect 675711 580349 675777 580350
rect 675711 550222 675777 550223
rect 675711 550158 675712 550222
rect 675776 550158 675777 550222
rect 675711 550157 675777 550158
rect 675714 546967 675774 550157
rect 675711 546966 675777 546967
rect 675711 546902 675712 546966
rect 675776 546902 675777 546966
rect 675711 546901 675777 546902
rect 675519 537050 675585 537051
rect 675519 536986 675520 537050
rect 675584 536986 675585 537050
rect 675519 536985 675585 536986
rect 675906 533795 675966 600181
rect 676098 579675 676158 649613
rect 676287 642574 676353 642575
rect 676287 642510 676288 642574
rect 676352 642510 676353 642574
rect 676287 642509 676353 642510
rect 676290 624815 676350 642509
rect 676482 640503 676542 658345
rect 676479 640502 676545 640503
rect 676479 640438 676480 640502
rect 676544 640438 676545 640502
rect 676479 640437 676545 640438
rect 676479 640354 676545 640355
rect 676479 640290 676480 640354
rect 676544 640290 676545 640354
rect 676479 640289 676545 640290
rect 676287 624814 676353 624815
rect 676287 624750 676288 624814
rect 676352 624750 676353 624814
rect 676287 624749 676353 624750
rect 676287 593438 676353 593439
rect 676287 593374 676288 593438
rect 676352 593374 676353 593438
rect 676287 593373 676353 593374
rect 676095 579674 676161 579675
rect 676095 579610 676096 579674
rect 676160 579610 676161 579674
rect 676095 579609 676161 579610
rect 676095 578934 676161 578935
rect 676095 578870 676096 578934
rect 676160 578870 676161 578934
rect 676095 578869 676161 578870
rect 676098 547115 676158 578869
rect 676095 547114 676161 547115
rect 676095 547050 676096 547114
rect 676160 547050 676161 547114
rect 676095 547049 676161 547050
rect 675903 533794 675969 533795
rect 675903 533730 675904 533794
rect 675968 533730 675969 533794
rect 675903 533729 675969 533730
rect 676290 532759 676350 593373
rect 676482 581303 676542 640289
rect 676674 621707 676734 694309
rect 676866 662407 676926 734861
rect 677058 708435 677118 777485
rect 677250 772963 677310 780189
rect 677823 773110 677889 773111
rect 677823 773046 677824 773110
rect 677888 773046 677889 773110
rect 677823 773045 677889 773046
rect 677247 772962 677313 772963
rect 677247 772898 677248 772962
rect 677312 772898 677313 772962
rect 677247 772897 677313 772898
rect 677247 772666 677313 772667
rect 677247 772602 677248 772666
rect 677312 772602 677313 772666
rect 677247 772601 677313 772602
rect 677250 752983 677310 772601
rect 677826 753871 677886 773045
rect 677823 753870 677889 753871
rect 677823 753806 677824 753870
rect 677888 753806 677889 753870
rect 677823 753805 677889 753806
rect 677247 752982 677313 752983
rect 677247 752918 677248 752982
rect 677312 752918 677313 752982
rect 677247 752917 677313 752918
rect 677055 708434 677121 708435
rect 677055 708370 677056 708434
rect 677120 708370 677121 708434
rect 677055 708369 677121 708370
rect 677055 688306 677121 688307
rect 677055 688242 677056 688306
rect 677120 688242 677121 688306
rect 677055 688241 677121 688242
rect 677058 687675 677118 688241
rect 677058 687615 677310 687675
rect 677055 685642 677121 685643
rect 677055 685578 677056 685642
rect 677120 685578 677121 685642
rect 677055 685577 677121 685578
rect 676863 662406 676929 662407
rect 676863 662342 676864 662406
rect 676928 662342 676929 662406
rect 676863 662341 676929 662342
rect 676671 621706 676737 621707
rect 676671 621642 676672 621706
rect 676736 621642 676737 621706
rect 676671 621641 676737 621642
rect 677058 617859 677118 685577
rect 677250 663591 677310 687615
rect 677247 663590 677313 663591
rect 677247 663526 677248 663590
rect 677312 663526 677313 663590
rect 677247 663525 677313 663526
rect 677055 617858 677121 617859
rect 677055 617794 677056 617858
rect 677120 617794 677121 617858
rect 677055 617793 677121 617794
rect 676671 595362 676737 595363
rect 676671 595298 676672 595362
rect 676736 595298 676737 595362
rect 676671 595297 676737 595298
rect 676479 581302 676545 581303
rect 676479 581238 676480 581302
rect 676544 581238 676545 581302
rect 676479 581237 676545 581238
rect 676674 536311 676734 595297
rect 676671 536310 676737 536311
rect 676671 536246 676672 536310
rect 676736 536246 676737 536310
rect 676671 536245 676737 536246
rect 676287 532758 676353 532759
rect 676287 532694 676288 532758
rect 676352 532694 676353 532758
rect 676287 532693 676353 532694
rect 675327 491466 675393 491467
rect 675327 491402 675328 491466
rect 675392 491402 675393 491466
rect 675327 491401 675393 491402
rect 675135 487470 675201 487471
rect 675135 487406 675136 487470
rect 675200 487406 675201 487470
rect 675135 487405 675201 487406
rect 674367 483844 674433 483845
rect 674367 483780 674368 483844
rect 674432 483780 674433 483844
rect 674367 483779 674433 483780
rect 42111 425162 42177 425163
rect 42111 425098 42112 425162
rect 42176 425098 42177 425162
rect 42111 425097 42177 425098
rect 41919 404886 41985 404887
rect 41919 404822 41920 404886
rect 41984 404822 41985 404886
rect 41919 404821 41985 404822
rect 41727 403850 41793 403851
rect 41727 403786 41728 403850
rect 41792 403786 41793 403850
rect 41727 403785 41793 403786
rect 41343 401926 41409 401927
rect 41343 401862 41344 401926
rect 41408 401862 41409 401926
rect 41343 401861 41409 401862
rect 41151 399558 41217 399559
rect 41151 399494 41152 399558
rect 41216 399494 41217 399558
rect 41151 399493 41217 399494
rect 40959 398818 41025 398819
rect 40959 398754 40960 398818
rect 41024 398754 41025 398818
rect 40959 398753 41025 398754
rect 40575 390234 40641 390235
rect 40575 390170 40576 390234
rect 40640 390170 40641 390234
rect 40575 390169 40641 390170
rect 40383 389198 40449 389199
rect 40383 389134 40384 389198
rect 40448 389134 40449 389198
rect 40383 389133 40449 389134
rect 40386 345983 40446 389133
rect 40578 346871 40638 390169
rect 40767 387570 40833 387571
rect 40767 387506 40768 387570
rect 40832 387506 40833 387570
rect 40767 387505 40833 387506
rect 40770 356935 40830 387505
rect 40959 386090 41025 386091
rect 40959 386026 40960 386090
rect 41024 386026 41025 386090
rect 40959 386025 41025 386026
rect 40767 356934 40833 356935
rect 40767 356870 40768 356934
rect 40832 356870 40833 356934
rect 40767 356869 40833 356870
rect 40962 355603 41022 386025
rect 41343 385202 41409 385203
rect 41343 385138 41344 385202
rect 41408 385138 41409 385202
rect 41343 385137 41409 385138
rect 41151 383130 41217 383131
rect 41151 383066 41152 383130
rect 41216 383066 41217 383130
rect 41151 383065 41217 383066
rect 41154 356491 41214 383065
rect 41346 358711 41406 385137
rect 41535 381946 41601 381947
rect 41535 381882 41536 381946
rect 41600 381882 41601 381946
rect 41535 381881 41601 381882
rect 41538 359451 41598 381881
rect 41730 361375 41790 403785
rect 42114 402667 42174 425097
rect 676479 412138 676545 412139
rect 676479 412074 676480 412138
rect 676544 412074 676545 412138
rect 676479 412073 676545 412074
rect 676482 406219 676542 412073
rect 676671 411990 676737 411991
rect 676671 411926 676672 411990
rect 676736 411926 676737 411990
rect 676671 411925 676737 411926
rect 676479 406218 676545 406219
rect 676479 406154 676480 406218
rect 676544 406154 676545 406218
rect 676479 406153 676545 406154
rect 674175 405922 674241 405923
rect 674175 405858 674176 405922
rect 674240 405858 674241 405922
rect 674175 405857 674241 405858
rect 42111 402666 42177 402667
rect 42111 402602 42112 402666
rect 42176 402602 42177 402666
rect 42111 402601 42177 402602
rect 41919 400002 41985 400003
rect 41919 399938 41920 400002
rect 41984 399938 41985 400002
rect 41919 399937 41985 399938
rect 41922 361967 41982 399937
rect 42111 371586 42177 371587
rect 42111 371522 42112 371586
rect 42176 371522 42177 371586
rect 42111 371521 42177 371522
rect 42114 362855 42174 371521
rect 42111 362854 42177 362855
rect 42111 362790 42112 362854
rect 42176 362790 42177 362854
rect 42111 362789 42177 362790
rect 41919 361966 41985 361967
rect 41919 361902 41920 361966
rect 41984 361902 41985 361966
rect 41919 361901 41985 361902
rect 41727 361374 41793 361375
rect 41727 361310 41728 361374
rect 41792 361310 41793 361374
rect 41727 361309 41793 361310
rect 41535 359450 41601 359451
rect 41535 359386 41536 359450
rect 41600 359386 41601 359450
rect 41535 359385 41601 359386
rect 41343 358710 41409 358711
rect 41343 358646 41344 358710
rect 41408 358646 41409 358710
rect 41343 358645 41409 358646
rect 41151 356490 41217 356491
rect 41151 356426 41152 356490
rect 41216 356426 41217 356490
rect 41151 356425 41217 356426
rect 40959 355602 41025 355603
rect 40959 355538 40960 355602
rect 41024 355538 41025 355602
rect 40959 355537 41025 355538
rect 40575 346870 40641 346871
rect 40575 346806 40576 346870
rect 40640 346806 40641 346870
rect 40575 346805 40641 346806
rect 40383 345982 40449 345983
rect 40383 345918 40384 345982
rect 40448 345918 40449 345982
rect 40383 345917 40449 345918
rect 40959 344354 41025 344355
rect 40959 344290 40960 344354
rect 41024 344290 41025 344354
rect 40959 344289 41025 344290
rect 40767 342874 40833 342875
rect 40767 342810 40768 342874
rect 40832 342810 40833 342874
rect 40767 342809 40833 342810
rect 40383 341246 40449 341247
rect 40383 341182 40384 341246
rect 40448 341182 40449 341246
rect 40383 341181 40449 341182
rect 40386 319787 40446 341181
rect 40383 319786 40449 319787
rect 40383 319722 40384 319786
rect 40448 319722 40449 319786
rect 40383 319721 40449 319722
rect 40770 312387 40830 342809
rect 40962 313719 41022 344289
rect 41343 341986 41409 341987
rect 41343 341922 41344 341986
rect 41408 341922 41409 341986
rect 41343 341921 41409 341922
rect 41151 339914 41217 339915
rect 41151 339850 41152 339914
rect 41216 339850 41217 339914
rect 41151 339849 41217 339850
rect 40959 313718 41025 313719
rect 40959 313654 40960 313718
rect 41024 313654 41025 313718
rect 40959 313653 41025 313654
rect 41154 313275 41214 339849
rect 41346 315495 41406 341921
rect 41535 338730 41601 338731
rect 41535 338666 41536 338730
rect 41600 338666 41601 338730
rect 41535 338665 41601 338666
rect 41538 316235 41598 338665
rect 41730 318011 41790 361309
rect 41922 318751 41982 361901
rect 674178 360783 674238 405857
rect 676674 405331 676734 411925
rect 675519 405330 675585 405331
rect 675519 405266 675520 405330
rect 675584 405266 675585 405330
rect 675519 405265 675585 405266
rect 676671 405330 676737 405331
rect 676671 405266 676672 405330
rect 676736 405266 676737 405330
rect 676671 405265 676737 405266
rect 674943 403258 675009 403259
rect 674943 403194 674944 403258
rect 675008 403194 675009 403258
rect 674943 403193 675009 403194
rect 674559 400594 674625 400595
rect 674559 400530 674560 400594
rect 674624 400530 674625 400594
rect 674559 400529 674625 400530
rect 674367 400446 674433 400447
rect 674367 400382 674368 400446
rect 674432 400382 674433 400446
rect 674367 400381 674433 400382
rect 674370 372031 674430 400381
rect 674562 378839 674622 400529
rect 674559 378838 674625 378839
rect 674559 378774 674560 378838
rect 674624 378774 674625 378838
rect 674559 378773 674625 378774
rect 674946 373955 675006 403193
rect 675327 374546 675393 374547
rect 675327 374482 675328 374546
rect 675392 374482 675393 374546
rect 675327 374481 675393 374482
rect 674943 373954 675009 373955
rect 674943 373890 674944 373954
rect 675008 373890 675009 373954
rect 674943 373889 675009 373890
rect 674367 372030 674433 372031
rect 674367 371966 674368 372030
rect 674432 371966 674433 372030
rect 674367 371965 674433 371966
rect 674367 361448 674433 361449
rect 674367 361384 674368 361448
rect 674432 361384 674433 361448
rect 674367 361383 674433 361384
rect 674175 360782 674241 360783
rect 674175 360718 674176 360782
rect 674240 360718 674241 360782
rect 674175 360717 674241 360718
rect 673983 360042 674049 360043
rect 673983 359978 673984 360042
rect 674048 359978 674049 360042
rect 673983 359977 674049 359978
rect 42111 346278 42177 346279
rect 42111 346214 42112 346278
rect 42176 346214 42177 346278
rect 42111 346213 42177 346214
rect 41919 318750 41985 318751
rect 41919 318686 41920 318750
rect 41984 318686 41985 318750
rect 41919 318685 41985 318686
rect 41727 318010 41793 318011
rect 41727 317946 41728 318010
rect 41792 317946 41793 318010
rect 41727 317945 41793 317946
rect 41535 316234 41601 316235
rect 41535 316170 41536 316234
rect 41600 316170 41601 316234
rect 41535 316169 41601 316170
rect 41343 315494 41409 315495
rect 41343 315430 41344 315494
rect 41408 315430 41409 315494
rect 41343 315429 41409 315430
rect 41151 313274 41217 313275
rect 41151 313210 41152 313274
rect 41216 313210 41217 313274
rect 41151 313209 41217 313210
rect 40767 312386 40833 312387
rect 40767 312322 40768 312386
rect 40832 312322 40833 312386
rect 40767 312321 40833 312322
rect 40767 302322 40833 302323
rect 40767 302258 40768 302322
rect 40832 302258 40833 302322
rect 40767 302257 40833 302258
rect 40575 298770 40641 298771
rect 40575 298706 40576 298770
rect 40640 298706 40641 298770
rect 40575 298705 40641 298706
rect 40383 298030 40449 298031
rect 40383 297966 40384 298030
rect 40448 297966 40449 298030
rect 40383 297965 40449 297966
rect 40386 276571 40446 297965
rect 40578 296699 40638 298705
rect 40575 296698 40641 296699
rect 40575 296634 40576 296698
rect 40640 296634 40641 296698
rect 40575 296633 40641 296634
rect 40575 295514 40641 295515
rect 40575 295450 40576 295514
rect 40640 295450 40641 295514
rect 40575 295449 40641 295450
rect 40383 276570 40449 276571
rect 40383 276506 40384 276570
rect 40448 276506 40449 276570
rect 40383 276505 40449 276506
rect 40578 272871 40638 295449
rect 40575 272870 40641 272871
rect 40575 272806 40576 272870
rect 40640 272806 40641 272870
rect 40575 272805 40641 272806
rect 40770 259551 40830 302257
rect 40959 301138 41025 301139
rect 40959 301074 40960 301138
rect 41024 301074 41025 301138
rect 40959 301073 41025 301074
rect 40962 270651 41022 301073
rect 41151 299658 41217 299659
rect 41151 299594 41152 299658
rect 41216 299594 41217 299658
rect 41151 299593 41217 299594
rect 40959 270650 41025 270651
rect 40959 270586 40960 270650
rect 41024 270586 41025 270650
rect 40959 270585 41025 270586
rect 41154 269171 41214 299593
rect 41343 296698 41409 296699
rect 41343 296634 41344 296698
rect 41408 296634 41409 296698
rect 41343 296633 41409 296634
rect 41535 296698 41601 296699
rect 41535 296634 41536 296698
rect 41600 296634 41601 296698
rect 41535 296633 41601 296634
rect 41346 270059 41406 296633
rect 41538 272427 41598 296633
rect 41730 274647 41790 317945
rect 41922 275239 41982 318685
rect 42114 303803 42174 346213
rect 42303 345982 42369 345983
rect 42303 345918 42304 345982
rect 42368 345918 42369 345982
rect 42303 345917 42369 345918
rect 42111 303802 42177 303803
rect 42111 303738 42112 303802
rect 42176 303738 42177 303802
rect 42111 303737 42177 303738
rect 41919 275238 41985 275239
rect 41919 275174 41920 275238
rect 41984 275174 41985 275238
rect 41919 275173 41985 275174
rect 41727 274646 41793 274647
rect 41727 274582 41728 274646
rect 41792 274582 41793 274646
rect 41727 274581 41793 274582
rect 41922 274055 41982 275173
rect 41919 274054 41985 274055
rect 41919 273990 41920 274054
rect 41984 273990 41985 274054
rect 41919 273989 41985 273990
rect 41535 272426 41601 272427
rect 41535 272362 41536 272426
rect 41600 272362 41601 272426
rect 41535 272361 41601 272362
rect 41919 270502 41985 270503
rect 41919 270438 41920 270502
rect 41984 270438 41985 270502
rect 41919 270437 41985 270438
rect 41343 270058 41409 270059
rect 41343 269994 41344 270058
rect 41408 269994 41409 270058
rect 41343 269993 41409 269994
rect 41151 269170 41217 269171
rect 41151 269106 41152 269170
rect 41216 269106 41217 269170
rect 41151 269105 41217 269106
rect 40767 259550 40833 259551
rect 40767 259486 40768 259550
rect 40832 259486 40833 259550
rect 40767 259485 40833 259486
rect 40383 257922 40449 257923
rect 40383 257858 40384 257922
rect 40448 257858 40449 257922
rect 40383 257857 40449 257858
rect 40386 227287 40446 257857
rect 40575 256442 40641 256443
rect 40575 256378 40576 256442
rect 40640 256378 40641 256442
rect 40575 256377 40641 256378
rect 40578 247859 40638 256377
rect 40959 255702 41025 255703
rect 40959 255638 40960 255702
rect 41024 255638 41025 255702
rect 40959 255637 41025 255638
rect 40767 253482 40833 253483
rect 40767 253418 40768 253482
rect 40832 253418 40833 253482
rect 40767 253417 40833 253418
rect 40575 247858 40641 247859
rect 40575 247794 40576 247858
rect 40640 247794 40641 247858
rect 40575 247793 40641 247794
rect 40575 227582 40641 227583
rect 40575 227518 40576 227582
rect 40640 227518 40641 227582
rect 40575 227517 40641 227518
rect 40383 227286 40449 227287
rect 40383 227222 40384 227286
rect 40448 227222 40449 227286
rect 40383 227221 40449 227222
rect 40578 225955 40638 227517
rect 40770 226843 40830 253417
rect 40962 229063 41022 255637
rect 41343 254814 41409 254815
rect 41343 254750 41344 254814
rect 41408 254750 41409 254814
rect 41343 254749 41409 254750
rect 41151 252446 41217 252447
rect 41151 252382 41152 252446
rect 41216 252382 41217 252446
rect 41151 252381 41217 252382
rect 41154 229655 41214 252381
rect 41346 233355 41406 254749
rect 41535 247710 41601 247711
rect 41535 247646 41536 247710
rect 41600 247646 41601 247710
rect 41535 247645 41601 247646
rect 41343 233354 41409 233355
rect 41343 233290 41344 233354
rect 41408 233290 41409 233354
rect 41343 233289 41409 233290
rect 41151 229654 41217 229655
rect 41151 229590 41152 229654
rect 41216 229590 41217 229654
rect 41151 229589 41217 229590
rect 40959 229062 41025 229063
rect 40959 228998 40960 229062
rect 41024 228998 41025 229062
rect 40959 228997 41025 228998
rect 41538 227583 41598 247645
rect 41727 243418 41793 243419
rect 41727 243354 41728 243418
rect 41792 243354 41793 243418
rect 41727 243353 41793 243354
rect 41730 231135 41790 243353
rect 41922 231727 41982 270437
rect 42114 260439 42174 303737
rect 42306 303063 42366 345917
rect 42687 336214 42753 336215
rect 42687 336150 42688 336214
rect 42752 336150 42753 336214
rect 42687 336149 42753 336150
rect 42495 327482 42561 327483
rect 42495 327418 42496 327482
rect 42560 327418 42561 327482
rect 42495 327417 42561 327418
rect 42498 323043 42558 327417
rect 42495 323042 42561 323043
rect 42495 322978 42496 323042
rect 42560 322978 42561 323042
rect 42495 322977 42561 322978
rect 42690 317419 42750 336149
rect 42687 317418 42753 317419
rect 42687 317354 42688 317418
rect 42752 317354 42753 317418
rect 42687 317353 42753 317354
rect 673986 314903 674046 359977
rect 674178 315791 674238 360717
rect 674370 317271 674430 361383
rect 675330 335031 675390 374481
rect 675522 360191 675582 405265
rect 675711 371734 675777 371735
rect 675711 371670 675712 371734
rect 675776 371670 675777 371734
rect 675711 371669 675777 371670
rect 675519 360190 675585 360191
rect 675519 360126 675520 360190
rect 675584 360126 675585 360190
rect 675519 360125 675585 360126
rect 675327 335030 675393 335031
rect 675327 334966 675328 335030
rect 675392 334966 675393 335030
rect 675327 334965 675393 334966
rect 675714 334029 675774 371669
rect 676671 345538 676737 345539
rect 676671 345474 676672 345538
rect 676736 345474 676737 345538
rect 676671 345473 676737 345474
rect 676095 345390 676161 345391
rect 676095 345326 676096 345390
rect 676160 345326 676161 345390
rect 676095 345325 676161 345326
rect 675522 333969 675774 334029
rect 675522 333847 675582 333969
rect 675519 333846 675585 333847
rect 675519 333782 675520 333846
rect 675584 333782 675585 333846
rect 675519 333781 675585 333782
rect 675327 329554 675393 329555
rect 675327 329490 675328 329554
rect 675392 329490 675393 329554
rect 675327 329489 675393 329490
rect 674367 317270 674433 317271
rect 674367 317206 674368 317270
rect 674432 317206 674433 317270
rect 674367 317205 674433 317206
rect 674367 316456 674433 316457
rect 674367 316392 674368 316456
rect 674432 316392 674433 316456
rect 674367 316391 674433 316392
rect 674175 315790 674241 315791
rect 674175 315726 674176 315790
rect 674240 315726 674241 315790
rect 674175 315725 674241 315726
rect 673983 314902 674049 314903
rect 673983 314838 673984 314902
rect 674048 314838 674049 314902
rect 673983 314837 674049 314838
rect 42303 303062 42369 303063
rect 42303 302998 42304 303062
rect 42368 302998 42369 303062
rect 42303 302997 42369 302998
rect 42303 283674 42369 283675
rect 42303 283610 42304 283674
rect 42368 283610 42369 283674
rect 42303 283609 42369 283610
rect 42306 281603 42366 283609
rect 42303 281602 42369 281603
rect 42303 281538 42304 281602
rect 42368 281538 42369 281602
rect 42303 281537 42369 281538
rect 673986 269911 674046 314837
rect 674178 270207 674238 315725
rect 674370 272279 674430 316391
rect 674559 312682 674625 312683
rect 674559 312618 674560 312682
rect 674624 312618 674625 312682
rect 674559 312617 674625 312618
rect 674562 283675 674622 312617
rect 675330 290039 675390 329489
rect 675327 290038 675393 290039
rect 675327 289974 675328 290038
rect 675392 289974 675393 290038
rect 675327 289973 675393 289974
rect 675522 289595 675582 333781
rect 676098 333551 676158 345325
rect 676479 345242 676545 345243
rect 676479 345178 676480 345242
rect 676544 345178 676545 345242
rect 676479 345177 676545 345178
rect 676287 344502 676353 344503
rect 676287 344438 676288 344502
rect 676352 344438 676353 344502
rect 676287 344437 676353 344438
rect 676095 333550 676161 333551
rect 676095 333486 676096 333550
rect 676160 333486 676161 333550
rect 676095 333485 676161 333486
rect 676290 330591 676350 344437
rect 676287 330590 676353 330591
rect 676287 330526 676288 330590
rect 676352 330526 676353 330590
rect 676287 330525 676353 330526
rect 676482 326891 676542 345177
rect 676674 328075 676734 345473
rect 676671 328074 676737 328075
rect 676671 328010 676672 328074
rect 676736 328010 676737 328074
rect 676671 328009 676737 328010
rect 676479 326890 676545 326891
rect 676479 326826 676480 326890
rect 676544 326826 676545 326890
rect 676479 326825 676545 326826
rect 675711 299510 675777 299511
rect 675711 299446 675712 299510
rect 675776 299446 675777 299510
rect 675711 299445 675777 299446
rect 675519 289594 675585 289595
rect 675519 289530 675520 289594
rect 675584 289530 675585 289594
rect 675519 289529 675585 289530
rect 675714 285303 675774 299445
rect 676671 299362 676737 299363
rect 676671 299298 676672 299362
rect 676736 299298 676737 299362
rect 676671 299297 676737 299298
rect 675711 285302 675777 285303
rect 675711 285238 675712 285302
rect 675776 285238 675777 285302
rect 675711 285237 675777 285238
rect 675135 285006 675201 285007
rect 675135 284942 675136 285006
rect 675200 284942 675201 285006
rect 675135 284941 675201 284942
rect 674559 283674 674625 283675
rect 674559 283610 674560 283674
rect 674624 283610 674625 283674
rect 674559 283609 674625 283610
rect 674943 275386 675009 275387
rect 674943 275322 674944 275386
rect 675008 275322 675009 275386
rect 674943 275321 675009 275322
rect 674367 272278 674433 272279
rect 674367 272214 674368 272278
rect 674432 272214 674433 272278
rect 674367 272213 674433 272214
rect 674175 270206 674241 270207
rect 674175 270142 674176 270206
rect 674240 270142 674241 270206
rect 674175 270141 674241 270142
rect 674559 270206 674625 270207
rect 674559 270142 674560 270206
rect 674624 270142 674625 270206
rect 674559 270141 674625 270142
rect 673983 269910 674049 269911
rect 673983 269846 673984 269910
rect 674048 269846 674049 269910
rect 673983 269845 674049 269846
rect 674367 268282 674433 268283
rect 674367 268218 674368 268282
rect 674432 268218 674433 268282
rect 674367 268217 674433 268218
rect 42111 260438 42177 260439
rect 42111 260374 42112 260438
rect 42176 260374 42177 260438
rect 42111 260373 42177 260374
rect 210687 246378 210753 246379
rect 210687 246314 210688 246378
rect 210752 246314 210753 246378
rect 210687 246313 210753 246314
rect 210303 246230 210369 246231
rect 210303 246166 210304 246230
rect 210368 246166 210369 246230
rect 210303 246165 210369 246166
rect 145407 242086 145473 242087
rect 145407 242022 145408 242086
rect 145472 242022 145473 242086
rect 145407 242021 145473 242022
rect 42111 240754 42177 240755
rect 42111 240690 42112 240754
rect 42176 240690 42177 240754
rect 42111 240689 42177 240690
rect 42495 240754 42561 240755
rect 42495 240690 42496 240754
rect 42560 240690 42561 240754
rect 42495 240689 42561 240690
rect 41919 231726 41985 231727
rect 41919 231662 41920 231726
rect 41984 231662 41985 231726
rect 41919 231661 41985 231662
rect 41727 231134 41793 231135
rect 41727 231070 41728 231134
rect 41792 231070 41793 231134
rect 41727 231069 41793 231070
rect 41535 227582 41601 227583
rect 41535 227518 41536 227582
rect 41600 227518 41601 227582
rect 41535 227517 41601 227518
rect 40767 226842 40833 226843
rect 40767 226778 40768 226842
rect 40832 226778 40833 226842
rect 40767 226777 40833 226778
rect 40575 225954 40641 225955
rect 40575 225890 40576 225954
rect 40640 225890 40641 225954
rect 40575 225889 40641 225890
rect 40383 214706 40449 214707
rect 40383 214642 40384 214706
rect 40448 214642 40449 214706
rect 40383 214641 40449 214642
rect 40386 184219 40446 214641
rect 40575 213226 40641 213227
rect 40575 213162 40576 213226
rect 40640 213162 40641 213226
rect 40575 213161 40641 213162
rect 40383 184218 40449 184219
rect 40383 184154 40384 184218
rect 40448 184154 40449 184218
rect 40383 184153 40449 184154
rect 40578 182887 40638 213161
rect 40959 212486 41025 212487
rect 40959 212422 40960 212486
rect 41024 212422 41025 212486
rect 40959 212421 41025 212422
rect 40767 210414 40833 210415
rect 40767 210350 40768 210414
rect 40832 210350 40833 210414
rect 40767 210349 40833 210350
rect 40770 183627 40830 210349
rect 40962 185995 41022 212421
rect 41151 211598 41217 211599
rect 41151 211534 41152 211598
rect 41216 211534 41217 211598
rect 41151 211533 41217 211534
rect 41154 190139 41214 211533
rect 41151 190138 41217 190139
rect 41151 190074 41152 190138
rect 41216 190074 41217 190138
rect 41151 190073 41217 190074
rect 41730 188363 41790 231069
rect 41922 189103 41982 231661
rect 42114 230543 42174 240689
rect 42498 237943 42558 240689
rect 42495 237942 42561 237943
rect 42495 237878 42496 237942
rect 42560 237878 42561 237942
rect 42495 237877 42561 237878
rect 42111 230542 42177 230543
rect 42111 230478 42112 230542
rect 42176 230478 42177 230542
rect 42111 230477 42177 230478
rect 42303 197686 42369 197687
rect 42303 197622 42304 197686
rect 42368 197622 42369 197686
rect 42303 197621 42369 197622
rect 42111 197390 42177 197391
rect 42111 197326 42112 197390
rect 42176 197326 42177 197390
rect 42111 197325 42177 197326
rect 42114 191027 42174 197325
rect 42306 195171 42366 197621
rect 42303 195170 42369 195171
rect 42303 195106 42304 195170
rect 42368 195106 42369 195170
rect 42303 195105 42369 195106
rect 42111 191026 42177 191027
rect 42111 190962 42112 191026
rect 42176 190962 42177 191026
rect 42111 190961 42177 190962
rect 41919 189102 41985 189103
rect 41919 189038 41920 189102
rect 41984 189038 41985 189102
rect 41919 189037 41985 189038
rect 41727 188362 41793 188363
rect 41727 188298 41728 188362
rect 41792 188298 41793 188362
rect 41727 188297 41793 188298
rect 40959 185994 41025 185995
rect 40959 185930 40960 185994
rect 41024 185930 41025 185994
rect 40959 185929 41025 185930
rect 40767 183626 40833 183627
rect 40767 183562 40768 183626
rect 40832 183562 40833 183626
rect 40767 183561 40833 183562
rect 40575 182886 40641 182887
rect 40575 182822 40576 182886
rect 40640 182822 40641 182886
rect 40575 182821 40641 182822
rect 31743 177114 31809 177115
rect 31743 177050 31744 177114
rect 31808 177050 31809 177114
rect 31743 177049 31809 177050
rect 31746 125315 31806 177049
rect 31743 125314 31809 125315
rect 31743 125250 31744 125314
rect 31808 125250 31809 125314
rect 31743 125249 31809 125250
rect 144831 106666 144897 106667
rect 144831 106602 144832 106666
rect 144896 106602 144897 106666
rect 144831 106601 144897 106602
rect 144834 100895 144894 106601
rect 144831 100894 144897 100895
rect 144831 100830 144832 100894
rect 144896 100830 144897 100894
rect 144831 100829 144897 100830
rect 145410 51019 145470 242021
rect 210306 237203 210366 246165
rect 210303 237202 210369 237203
rect 210303 237138 210304 237202
rect 210368 237138 210369 237202
rect 210303 237137 210369 237138
rect 210495 233798 210561 233799
rect 210495 233734 210496 233798
rect 210560 233734 210561 233798
rect 210495 233733 210561 233734
rect 210303 233058 210369 233059
rect 210303 232994 210304 233058
rect 210368 232994 210369 233058
rect 210303 232993 210369 232994
rect 145599 221810 145665 221811
rect 145599 221746 145600 221810
rect 145664 221746 145665 221810
rect 145599 221745 145665 221746
rect 145407 51018 145473 51019
rect 145407 50954 145408 51018
rect 145472 50954 145473 51018
rect 145407 50953 145473 50954
rect 145602 50871 145662 221745
rect 145791 218998 145857 218999
rect 145791 218934 145792 218998
rect 145856 218934 145857 218998
rect 145791 218933 145857 218934
rect 145794 51167 145854 218933
rect 145983 216482 146049 216483
rect 145983 216418 145984 216482
rect 146048 216418 146049 216482
rect 145983 216417 146049 216418
rect 145986 51315 146046 216417
rect 210306 202161 210366 232993
rect 210498 223473 210558 233733
rect 210690 233651 210750 246313
rect 337023 245194 337089 245195
rect 337023 245130 337024 245194
rect 337088 245130 337089 245194
rect 337023 245129 337089 245130
rect 337026 245047 337086 245129
rect 337023 245046 337089 245047
rect 337023 244982 337024 245046
rect 337088 244982 337089 245046
rect 337023 244981 337089 244982
rect 674370 238683 674430 268217
rect 674562 239275 674622 270141
rect 674751 268578 674817 268579
rect 674751 268514 674752 268578
rect 674816 268514 674817 268578
rect 674751 268513 674817 268514
rect 674754 250523 674814 268513
rect 674946 256107 675006 275321
rect 675138 256295 675198 284941
rect 676674 281899 676734 299297
rect 676671 281898 676737 281899
rect 676671 281834 676672 281898
rect 676736 281834 676737 281898
rect 676671 281833 676737 281834
rect 675711 270946 675777 270947
rect 675711 270882 675712 270946
rect 675776 270882 675777 270946
rect 675711 270881 675777 270882
rect 675327 269762 675393 269763
rect 675327 269698 675328 269762
rect 675392 269698 675393 269762
rect 675327 269697 675393 269698
rect 675135 256294 675201 256295
rect 675135 256230 675136 256294
rect 675200 256230 675201 256294
rect 675135 256229 675201 256230
rect 674946 256047 675198 256107
rect 674751 250522 674817 250523
rect 674751 250458 674752 250522
rect 674816 250458 674817 250522
rect 674751 250457 674817 250458
rect 675138 244307 675198 256047
rect 675135 244306 675201 244307
rect 675135 244242 675136 244306
rect 675200 244242 675201 244306
rect 675135 244241 675201 244242
rect 675330 239275 675390 269697
rect 675519 241346 675585 241347
rect 675519 241282 675520 241346
rect 675584 241282 675585 241346
rect 675519 241281 675585 241282
rect 674559 239274 674625 239275
rect 674559 239210 674560 239274
rect 674624 239210 674625 239274
rect 674559 239209 674625 239210
rect 675327 239274 675393 239275
rect 675327 239210 675328 239274
rect 675392 239210 675393 239274
rect 675327 239209 675393 239210
rect 675135 238978 675201 238979
rect 675135 238914 675136 238978
rect 675200 238914 675201 238978
rect 675135 238913 675201 238914
rect 674367 238682 674433 238683
rect 674367 238618 674368 238682
rect 674432 238618 674433 238682
rect 674367 238617 674433 238618
rect 211455 234686 211521 234687
rect 211455 234622 211456 234686
rect 211520 234622 211521 234686
rect 211455 234621 211521 234622
rect 211071 233946 211137 233947
rect 211071 233882 211072 233946
rect 211136 233882 211137 233946
rect 211071 233881 211137 233882
rect 210687 233650 210753 233651
rect 210687 233586 210688 233650
rect 210752 233586 210753 233650
rect 210687 233585 210753 233586
rect 211074 223473 211134 233881
rect 211458 233059 211518 234621
rect 212799 234094 212865 234095
rect 212799 234030 212800 234094
rect 212864 234030 212865 234094
rect 212799 234029 212865 234030
rect 637503 234094 637569 234095
rect 637503 234030 637504 234094
rect 637568 234030 637569 234094
rect 637503 234029 637569 234030
rect 212415 233798 212481 233799
rect 212415 233734 212416 233798
rect 212480 233734 212481 233798
rect 212415 233733 212481 233734
rect 212031 233650 212097 233651
rect 212031 233648 212032 233650
rect 211842 233588 212032 233648
rect 211455 233058 211521 233059
rect 211455 232994 211456 233058
rect 211520 232994 211521 233058
rect 211455 232993 211521 232994
rect 210498 223413 210750 223473
rect 211074 223413 211710 223473
rect 210495 208786 210561 208787
rect 210495 208722 210496 208786
rect 210560 208722 210561 208786
rect 210495 208721 210561 208722
rect 210162 202101 210366 202161
rect 210498 202161 210558 208721
rect 210690 206157 210750 223413
rect 211650 208821 211710 223413
rect 210882 208787 211710 208821
rect 210879 208786 211710 208787
rect 210879 208722 210880 208786
rect 210944 208761 211710 208786
rect 210944 208722 210945 208761
rect 210879 208721 210945 208722
rect 211842 206823 211902 233588
rect 212031 233586 212032 233588
rect 212096 233586 212097 233650
rect 212031 233585 212097 233586
rect 212223 233502 212289 233503
rect 212223 233438 212224 233502
rect 212288 233438 212289 233502
rect 212223 233437 212289 233438
rect 212226 223473 212286 233437
rect 212418 232911 212478 233733
rect 212415 232910 212481 232911
rect 212415 232846 212416 232910
rect 212480 232846 212481 232910
rect 212415 232845 212481 232846
rect 212226 223413 212478 223473
rect 210882 206763 211902 206823
rect 210882 206419 210942 206763
rect 210879 206418 210945 206419
rect 210879 206354 210880 206418
rect 210944 206354 210945 206418
rect 210879 206353 210945 206354
rect 210690 206097 212094 206157
rect 210879 205974 210945 205975
rect 210879 205910 210880 205974
rect 210944 205910 210945 205974
rect 210879 205909 210945 205910
rect 210882 205676 210942 205909
rect 210882 205616 211902 205676
rect 210498 202101 211518 202161
rect 210162 201495 210222 202101
rect 210114 201435 210222 201495
rect 210114 182739 210174 201435
rect 211458 198165 211518 202101
rect 210306 198105 211518 198165
rect 210111 182738 210177 182739
rect 210111 182674 210112 182738
rect 210176 182674 210177 182738
rect 210111 182673 210177 182674
rect 210306 181999 210366 198105
rect 211842 195501 211902 205616
rect 210690 195441 211902 195501
rect 210303 181998 210369 181999
rect 210303 181934 210304 181998
rect 210368 181934 210369 181998
rect 210303 181933 210369 181934
rect 210690 161279 210750 195441
rect 212034 194835 212094 206097
rect 211842 194775 212094 194835
rect 211842 184179 211902 194775
rect 211458 184119 211902 184179
rect 210879 182738 210945 182739
rect 210879 182674 210880 182738
rect 210944 182736 210945 182738
rect 210944 182676 211134 182736
rect 210944 182674 210945 182676
rect 210879 182673 210945 182674
rect 210879 181998 210945 181999
rect 210879 181934 210880 181998
rect 210944 181934 210945 181998
rect 210879 181933 210945 181934
rect 210687 161278 210753 161279
rect 210687 161214 210688 161278
rect 210752 161214 210753 161278
rect 210687 161213 210753 161214
rect 210882 155541 210942 181933
rect 210690 155481 210942 155541
rect 210690 154323 210750 155481
rect 210687 154322 210753 154323
rect 210687 154258 210688 154322
rect 210752 154258 210753 154322
rect 210687 154257 210753 154258
rect 210495 154174 210561 154175
rect 210495 154110 210496 154174
rect 210560 154110 210561 154174
rect 211074 154172 211134 182676
rect 210495 154109 210561 154110
rect 210690 154112 211134 154172
rect 210498 146883 210558 154109
rect 210690 151545 210750 154112
rect 210879 153286 210945 153287
rect 210879 153222 210880 153286
rect 210944 153222 210945 153286
rect 210879 153221 210945 153222
rect 210882 152211 210942 153221
rect 211458 152877 211518 184119
rect 212418 183513 212478 223413
rect 212802 221475 212862 234029
rect 637119 233798 637185 233799
rect 637119 233734 637120 233798
rect 637184 233734 637185 233798
rect 637119 233733 637185 233734
rect 637311 233798 637377 233799
rect 637311 233734 637312 233798
rect 637376 233734 637377 233798
rect 637311 233733 637377 233734
rect 636735 233650 636801 233651
rect 636735 233586 636736 233650
rect 636800 233586 636801 233650
rect 636735 233585 636801 233586
rect 212991 232910 213057 232911
rect 212991 232846 212992 232910
rect 213056 232846 213057 232910
rect 212991 232845 213057 232846
rect 212226 183453 212478 183513
rect 212610 221415 212862 221475
rect 212226 182736 212286 183453
rect 212610 182736 212670 221415
rect 212994 220809 213054 232845
rect 212802 220749 213054 220809
rect 212802 200829 212862 220749
rect 212802 200769 213054 200829
rect 211842 182676 212286 182736
rect 212418 182676 212670 182736
rect 211842 167529 211902 182676
rect 212418 168861 212478 182676
rect 212994 181996 213054 200769
rect 212802 181936 213054 181996
rect 212418 168801 212670 168861
rect 212610 167529 212670 168801
rect 211842 167469 212286 167529
rect 212226 164199 212286 167469
rect 211650 164139 212286 164199
rect 212418 167469 212670 167529
rect 211650 161276 211710 164139
rect 211650 161216 212286 161276
rect 211458 152817 212094 152877
rect 210882 152151 211710 152211
rect 210690 151485 211134 151545
rect 210498 146823 210750 146883
rect 210690 144111 210750 146823
rect 210687 144110 210753 144111
rect 210687 144046 210688 144110
rect 210752 144046 210753 144110
rect 210687 144045 210753 144046
rect 210495 143962 210561 143963
rect 210495 143898 210496 143962
rect 210560 143898 210561 143962
rect 210495 143897 210561 143898
rect 210498 126795 210558 143897
rect 211074 135561 211134 151485
rect 211650 136893 211710 152151
rect 211650 136833 211902 136893
rect 211074 135501 211710 135561
rect 210303 126794 210369 126795
rect 210303 126730 210304 126794
rect 210368 126730 210369 126794
rect 210303 126729 210369 126730
rect 210495 126794 210561 126795
rect 210495 126730 210496 126794
rect 210560 126730 210561 126794
rect 210495 126729 210561 126730
rect 210306 105187 210366 126729
rect 211650 120909 211710 135501
rect 210690 120849 211710 120909
rect 209919 105186 209985 105187
rect 209919 105122 209920 105186
rect 209984 105122 209985 105186
rect 209919 105121 209985 105122
rect 210303 105186 210369 105187
rect 210303 105122 210304 105186
rect 210368 105122 210369 105186
rect 210303 105121 210369 105122
rect 209727 94826 209793 94827
rect 209727 94762 209728 94826
rect 209792 94762 209793 94826
rect 209727 94761 209793 94762
rect 209730 82395 209790 94761
rect 209922 86095 209982 105121
rect 210111 103558 210177 103559
rect 210111 103494 210112 103558
rect 210176 103494 210177 103558
rect 210111 103493 210177 103494
rect 210114 93603 210174 103493
rect 210495 102374 210561 102375
rect 210495 102310 210496 102374
rect 210560 102310 210561 102374
rect 210495 102309 210561 102310
rect 210498 93791 210558 102309
rect 210690 100929 210750 120849
rect 211842 112917 211902 136833
rect 210882 112857 211902 112917
rect 210882 103559 210942 112857
rect 212034 112251 212094 152817
rect 211266 112191 212094 112251
rect 210879 103558 210945 103559
rect 210879 103494 210880 103558
rect 210944 103494 210945 103558
rect 210879 103493 210945 103494
rect 211266 102927 211326 112191
rect 212226 102927 212286 161216
rect 212418 146883 212478 167469
rect 212418 146823 212670 146883
rect 212610 137559 212670 146823
rect 212418 137499 212670 137559
rect 212418 118245 212478 137499
rect 212802 134895 212862 181936
rect 212802 134835 213054 134895
rect 212418 118185 212862 118245
rect 210882 102867 211326 102927
rect 211458 102867 212286 102927
rect 210882 102375 210942 102867
rect 210879 102374 210945 102375
rect 210879 102310 210880 102374
rect 210944 102310 210945 102374
rect 210879 102309 210945 102310
rect 210690 100869 210942 100929
rect 210882 100263 210942 100869
rect 210690 100203 210942 100263
rect 210495 93790 210561 93791
rect 210495 93726 210496 93790
rect 210560 93726 210561 93790
rect 210495 93725 210561 93726
rect 210114 93543 210366 93603
rect 210111 87870 210177 87871
rect 210111 87806 210112 87870
rect 210176 87806 210177 87870
rect 210111 87805 210177 87806
rect 209919 86094 209985 86095
rect 209919 86030 209920 86094
rect 209984 86030 209985 86094
rect 209919 86029 209985 86030
rect 210114 84615 210174 87805
rect 210111 84614 210177 84615
rect 210111 84550 210112 84614
rect 210176 84550 210177 84614
rect 210111 84549 210177 84550
rect 210306 83613 210366 93543
rect 210690 87723 210750 100203
rect 210879 94826 210945 94827
rect 210879 94762 210880 94826
rect 210944 94824 210945 94826
rect 211458 94824 211518 102867
rect 212802 101595 212862 118185
rect 210944 94764 211518 94824
rect 211650 101535 212862 101595
rect 210944 94762 210945 94764
rect 210879 94761 210945 94762
rect 210879 93790 210945 93791
rect 210879 93726 210880 93790
rect 210944 93726 210945 93790
rect 210879 93725 210945 93726
rect 210882 87871 210942 93725
rect 210879 87870 210945 87871
rect 210879 87806 210880 87870
rect 210944 87806 210945 87870
rect 210879 87805 210945 87806
rect 210687 87722 210753 87723
rect 210687 87658 210688 87722
rect 210752 87658 210753 87722
rect 211650 87720 211710 101535
rect 210687 87657 210753 87658
rect 210882 87660 211710 87720
rect 210882 86277 210942 87660
rect 210690 86217 210942 86277
rect 210690 84945 210750 86217
rect 210879 86094 210945 86095
rect 210879 86030 210880 86094
rect 210944 86092 210945 86094
rect 210944 86032 212094 86092
rect 210944 86030 210945 86032
rect 210879 86029 210945 86030
rect 212034 85611 212094 86032
rect 212034 85551 212670 85611
rect 210690 84885 211902 84945
rect 210687 84614 210753 84615
rect 210687 84550 210688 84614
rect 210752 84550 210753 84614
rect 210687 84549 210753 84550
rect 210114 83553 210366 83613
rect 209727 82394 209793 82395
rect 209727 82330 209728 82394
rect 209792 82330 209793 82394
rect 209727 82329 209793 82330
rect 209919 71886 209985 71887
rect 209919 71822 209920 71886
rect 209984 71822 209985 71886
rect 209919 71821 209985 71822
rect 209922 54127 209982 71821
rect 209919 54126 209985 54127
rect 209919 54062 209920 54126
rect 209984 54062 209985 54126
rect 209919 54061 209985 54062
rect 210114 53239 210174 83553
rect 210303 83430 210369 83431
rect 210303 83366 210304 83430
rect 210368 83366 210369 83430
rect 210303 83365 210369 83366
rect 210306 54423 210366 83365
rect 210495 57234 210561 57235
rect 210495 57170 210496 57234
rect 210560 57170 210561 57234
rect 210495 57169 210561 57170
rect 210303 54422 210369 54423
rect 210303 54358 210304 54422
rect 210368 54358 210369 54422
rect 210303 54357 210369 54358
rect 210498 53979 210558 57169
rect 210690 54127 210750 84549
rect 210879 82394 210945 82395
rect 210879 82330 210880 82394
rect 210944 82392 210945 82394
rect 210944 82332 211134 82392
rect 210944 82330 210945 82332
rect 210879 82329 210945 82330
rect 211074 80283 211134 82332
rect 211074 80223 211518 80283
rect 210879 58418 210945 58419
rect 210879 58354 210880 58418
rect 210944 58354 210945 58418
rect 210879 58353 210945 58354
rect 210882 55641 210942 58353
rect 210882 55581 211134 55641
rect 210879 55162 210945 55163
rect 210879 55098 210880 55162
rect 210944 55098 210945 55162
rect 210879 55097 210945 55098
rect 210882 54423 210942 55097
rect 210879 54422 210945 54423
rect 210879 54358 210880 54422
rect 210944 54358 210945 54422
rect 210879 54357 210945 54358
rect 210687 54126 210753 54127
rect 210687 54062 210688 54126
rect 210752 54062 210753 54126
rect 210687 54061 210753 54062
rect 210495 53978 210561 53979
rect 210495 53914 210496 53978
rect 210560 53914 210561 53978
rect 210495 53913 210561 53914
rect 211074 53535 211134 55581
rect 211458 53683 211518 80223
rect 211455 53682 211521 53683
rect 211455 53618 211456 53682
rect 211520 53618 211521 53682
rect 211455 53617 211521 53618
rect 211071 53534 211137 53535
rect 211071 53470 211072 53534
rect 211136 53470 211137 53534
rect 211071 53469 211137 53470
rect 210111 53238 210177 53239
rect 210111 53174 210112 53238
rect 210176 53174 210177 53238
rect 210111 53173 210177 53174
rect 211842 53091 211902 84885
rect 212610 53831 212670 85551
rect 212607 53830 212673 53831
rect 212607 53766 212608 53830
rect 212672 53766 212673 53830
rect 212607 53765 212673 53766
rect 212994 53535 213054 134835
rect 212991 53534 213057 53535
rect 212991 53470 212992 53534
rect 213056 53470 213057 53534
rect 212991 53469 213057 53470
rect 465663 53386 465729 53387
rect 465663 53322 465664 53386
rect 465728 53322 465729 53386
rect 465663 53321 465729 53322
rect 211839 53090 211905 53091
rect 211839 53026 211840 53090
rect 211904 53026 211905 53090
rect 211839 53025 211905 53026
rect 377535 53090 377601 53091
rect 377535 53026 377536 53090
rect 377600 53026 377601 53090
rect 377535 53025 377601 53026
rect 377343 52942 377409 52943
rect 377343 52878 377344 52942
rect 377408 52878 377409 52942
rect 377343 52877 377409 52878
rect 377346 52311 377406 52877
rect 377538 52311 377598 53025
rect 377346 52251 377598 52311
rect 145983 51314 146049 51315
rect 145983 51250 145984 51314
rect 146048 51250 146049 51314
rect 145983 51249 146049 51250
rect 145791 51166 145857 51167
rect 145791 51102 145792 51166
rect 145856 51102 145857 51166
rect 145791 51101 145857 51102
rect 145599 50870 145665 50871
rect 145599 50806 145600 50870
rect 145664 50806 145665 50870
rect 145599 50805 145665 50806
rect 306687 48946 306753 48947
rect 306687 48882 306688 48946
rect 306752 48882 306753 48946
rect 306687 48881 306753 48882
rect 302463 45394 302529 45395
rect 302463 45330 302464 45394
rect 302528 45330 302529 45394
rect 302463 45329 302529 45330
rect 302466 43323 302526 45329
rect 302463 43322 302529 43323
rect 302463 43258 302464 43322
rect 302528 43258 302529 43322
rect 302463 43257 302529 43258
rect 306690 42139 306750 48881
rect 356991 46134 357057 46135
rect 356991 46070 356992 46134
rect 357056 46070 357057 46134
rect 356991 46069 357057 46070
rect 356994 42139 357054 46069
rect 360063 45246 360129 45247
rect 360063 45182 360064 45246
rect 360128 45182 360129 45246
rect 360063 45181 360129 45182
rect 360066 43323 360126 45181
rect 362943 45098 363009 45099
rect 362943 45034 362944 45098
rect 363008 45034 363009 45098
rect 362943 45033 363009 45034
rect 362946 43323 363006 45033
rect 409023 44950 409089 44951
rect 409023 44886 409024 44950
rect 409088 44886 409089 44950
rect 409023 44885 409089 44886
rect 409026 43323 409086 44885
rect 360063 43322 360129 43323
rect 360063 43258 360064 43322
rect 360128 43258 360129 43322
rect 360063 43257 360129 43258
rect 362943 43322 363009 43323
rect 362943 43258 362944 43322
rect 363008 43258 363009 43322
rect 362943 43257 363009 43258
rect 409023 43322 409089 43323
rect 409023 43258 409024 43322
rect 409088 43258 409089 43322
rect 409023 43257 409089 43258
rect 306687 42138 306753 42139
rect 306687 42074 306688 42138
rect 306752 42074 306753 42138
rect 306687 42073 306753 42074
rect 356991 42138 357057 42139
rect 356991 42074 356992 42138
rect 357056 42074 357057 42138
rect 356991 42073 357057 42074
rect 465666 41843 465726 53321
rect 636738 52647 636798 233585
rect 636927 233502 636993 233503
rect 636927 233438 636928 233502
rect 636992 233438 636993 233502
rect 636927 233437 636993 233438
rect 636735 52646 636801 52647
rect 636735 52582 636736 52646
rect 636800 52582 636801 52646
rect 636735 52581 636801 52582
rect 636930 52055 636990 233437
rect 637122 52351 637182 233733
rect 637119 52350 637185 52351
rect 637119 52286 637120 52350
rect 637184 52286 637185 52350
rect 637119 52285 637185 52286
rect 636927 52054 636993 52055
rect 636927 51990 636928 52054
rect 636992 51990 636993 52054
rect 636927 51989 636993 51990
rect 637314 51907 637374 233733
rect 637506 52499 637566 234029
rect 637695 233946 637761 233947
rect 637695 233882 637696 233946
rect 637760 233882 637761 233946
rect 637695 233881 637761 233882
rect 637503 52498 637569 52499
rect 637503 52434 637504 52498
rect 637568 52434 637569 52498
rect 637503 52433 637569 52434
rect 637698 52203 637758 233881
rect 673983 226250 674049 226251
rect 673983 226186 673984 226250
rect 674048 226186 674049 226250
rect 673983 226185 674049 226186
rect 673986 182591 674046 226185
rect 674367 223142 674433 223143
rect 674367 223078 674368 223142
rect 674432 223078 674433 223142
rect 674367 223077 674433 223078
rect 674370 193543 674430 223077
rect 675138 217815 675198 238913
rect 675135 217814 675201 217815
rect 675135 217750 675136 217814
rect 675200 217750 675201 217814
rect 675135 217749 675201 217750
rect 675135 211746 675201 211747
rect 675135 211682 675136 211746
rect 675200 211682 675201 211746
rect 675135 211681 675201 211682
rect 674751 211598 674817 211599
rect 674751 211534 674752 211598
rect 674816 211534 674817 211598
rect 674751 211533 674817 211534
rect 674754 199759 674814 211533
rect 674751 199758 674817 199759
rect 674751 199694 674752 199758
rect 674816 199694 674817 199758
rect 674751 199693 674817 199694
rect 675138 199167 675198 211681
rect 675522 211599 675582 241281
rect 675714 226843 675774 270881
rect 676287 256294 676353 256295
rect 676287 256230 676288 256294
rect 676352 256230 676353 256294
rect 676287 256229 676353 256230
rect 676095 253630 676161 253631
rect 676095 253566 676096 253630
rect 676160 253566 676161 253630
rect 676095 253565 676161 253566
rect 675903 253482 675969 253483
rect 675903 253418 675904 253482
rect 675968 253418 675969 253482
rect 675903 253417 675969 253418
rect 675906 243567 675966 253417
rect 675903 243566 675969 243567
rect 675903 243502 675904 243566
rect 675968 243502 675969 243566
rect 675903 243501 675969 243502
rect 676098 236907 676158 253565
rect 676290 245195 676350 256229
rect 676287 245194 676353 245195
rect 676287 245130 676288 245194
rect 676352 245130 676353 245194
rect 676287 245129 676353 245130
rect 676095 236906 676161 236907
rect 676095 236842 676096 236906
rect 676160 236842 676161 236906
rect 676095 236841 676161 236842
rect 675711 226842 675777 226843
rect 675711 226778 675712 226842
rect 675776 226778 675777 226842
rect 675711 226777 675777 226778
rect 675519 211598 675585 211599
rect 675519 211534 675520 211598
rect 675584 211534 675585 211598
rect 675519 211533 675585 211534
rect 676095 210266 676161 210267
rect 676095 210202 676096 210266
rect 676160 210202 676161 210266
rect 676095 210201 676161 210202
rect 675519 210118 675585 210119
rect 675519 210054 675520 210118
rect 675584 210054 675585 210118
rect 675519 210053 675585 210054
rect 675135 199166 675201 199167
rect 675135 199102 675136 199166
rect 675200 199102 675201 199166
rect 675135 199101 675201 199102
rect 675522 198427 675582 210053
rect 675903 209822 675969 209823
rect 675903 209758 675904 209822
rect 675968 209758 675969 209822
rect 675903 209757 675969 209758
rect 675711 209674 675777 209675
rect 675711 209610 675712 209674
rect 675776 209610 675777 209674
rect 675711 209609 675777 209610
rect 675519 198426 675585 198427
rect 675519 198362 675520 198426
rect 675584 198362 675585 198426
rect 675519 198361 675585 198362
rect 675327 195762 675393 195763
rect 675327 195698 675328 195762
rect 675392 195698 675393 195762
rect 675327 195697 675393 195698
rect 674367 193542 674433 193543
rect 674367 193478 674368 193542
rect 674432 193478 674433 193542
rect 674367 193477 674433 193478
rect 673983 182590 674049 182591
rect 673983 182526 673984 182590
rect 674048 182526 674049 182590
rect 673983 182525 674049 182526
rect 673983 181258 674049 181259
rect 673983 181194 673984 181258
rect 674048 181194 674049 181258
rect 673983 181193 674049 181194
rect 673986 136859 674046 181193
rect 674175 178150 674241 178151
rect 674175 178086 674176 178150
rect 674240 178086 674241 178150
rect 674175 178085 674241 178086
rect 674178 148551 674238 178085
rect 674559 166458 674625 166459
rect 674559 166394 674560 166458
rect 674624 166394 674625 166458
rect 674559 166393 674625 166394
rect 674367 165570 674433 165571
rect 674367 165506 674368 165570
rect 674432 165506 674433 165570
rect 674367 165505 674433 165506
rect 674175 148550 674241 148551
rect 674175 148486 674176 148550
rect 674240 148486 674241 148550
rect 674175 148485 674241 148486
rect 673983 136858 674049 136859
rect 673983 136794 673984 136858
rect 674048 136794 674049 136858
rect 673983 136793 674049 136794
rect 674370 134565 674430 165505
rect 674562 135527 674622 166393
rect 675330 155541 675390 195697
rect 675519 195614 675585 195615
rect 675519 195550 675520 195614
rect 675584 195550 675585 195614
rect 675519 195549 675585 195550
rect 675138 155481 675390 155541
rect 675138 154323 675198 155481
rect 675522 154619 675582 195549
rect 675714 180963 675774 209609
rect 675906 204347 675966 209757
rect 675903 204346 675969 204347
rect 675903 204282 675904 204346
rect 675968 204282 675969 204346
rect 675903 204281 675969 204282
rect 676098 195319 676158 210201
rect 676287 209970 676353 209971
rect 676287 209906 676288 209970
rect 676352 209906 676353 209970
rect 676287 209905 676353 209906
rect 676095 195318 676161 195319
rect 676095 195254 676096 195318
rect 676160 195254 676161 195318
rect 676095 195253 676161 195254
rect 676290 191619 676350 209905
rect 676479 209526 676545 209527
rect 676479 209462 676480 209526
rect 676544 209462 676545 209526
rect 676479 209461 676545 209462
rect 676287 191618 676353 191619
rect 676287 191554 676288 191618
rect 676352 191554 676353 191618
rect 676287 191553 676353 191554
rect 675711 180962 675777 180963
rect 675711 180898 675712 180962
rect 675776 180898 675777 180962
rect 675711 180897 675777 180898
rect 676482 179483 676542 209461
rect 676479 179482 676545 179483
rect 676479 179418 676480 179482
rect 676544 179418 676545 179482
rect 676479 179417 676545 179418
rect 676287 164090 676353 164091
rect 676287 164026 676288 164090
rect 676352 164026 676353 164090
rect 676287 164025 676353 164026
rect 675519 154618 675585 154619
rect 675519 154554 675520 154618
rect 675584 154554 675585 154618
rect 675519 154553 675585 154554
rect 675135 154322 675201 154323
rect 675135 154258 675136 154322
rect 675200 154258 675201 154322
rect 675135 154257 675201 154258
rect 675138 135561 675198 154257
rect 674559 135526 674625 135527
rect 674559 135462 674560 135526
rect 674624 135462 674625 135526
rect 674559 135461 674625 135462
rect 674754 135501 675198 135561
rect 674559 134934 674625 134935
rect 674559 134870 674560 134934
rect 674624 134895 674625 134934
rect 674754 134895 674814 135501
rect 674624 134870 674814 134895
rect 674559 134869 674814 134870
rect 674562 134835 674814 134869
rect 674367 134564 674433 134565
rect 674367 134500 674368 134564
rect 674432 134500 674433 134564
rect 674367 134499 674433 134500
rect 674175 132936 674241 132937
rect 674175 132872 674176 132936
rect 674240 132872 674241 132936
rect 674175 132871 674241 132872
rect 674178 103263 674238 132871
rect 674754 111403 674814 134835
rect 674751 111402 674817 111403
rect 674751 111338 674752 111402
rect 674816 111338 674817 111402
rect 674751 111337 674817 111338
rect 674754 109479 674814 111337
rect 675522 110071 675582 154553
rect 676290 153435 676350 164025
rect 676671 163942 676737 163943
rect 676671 163878 676672 163942
rect 676736 163878 676737 163942
rect 676671 163877 676737 163878
rect 676479 163646 676545 163647
rect 676479 163582 676480 163646
rect 676544 163582 676545 163646
rect 676479 163581 676545 163582
rect 676287 153434 676353 153435
rect 676287 153370 676288 153434
rect 676352 153370 676353 153434
rect 676287 153369 676353 153370
rect 676482 150327 676542 163581
rect 676479 150326 676545 150327
rect 676479 150262 676480 150326
rect 676544 150262 676545 150326
rect 676479 150261 676545 150262
rect 676674 146627 676734 163877
rect 676671 146626 676737 146627
rect 676671 146562 676672 146626
rect 676736 146562 676737 146626
rect 676671 146561 676737 146562
rect 675711 120430 675777 120431
rect 675711 120366 675712 120430
rect 675776 120366 675777 120430
rect 675711 120365 675777 120366
rect 675519 110070 675585 110071
rect 675519 110006 675520 110070
rect 675584 110006 675585 110070
rect 675519 110005 675585 110006
rect 674751 109478 674817 109479
rect 674751 109414 674752 109478
rect 674816 109414 674817 109478
rect 674751 109413 674817 109414
rect 675714 108147 675774 120365
rect 676671 118062 676737 118063
rect 676671 117998 676672 118062
rect 676736 117998 676737 118062
rect 676671 117997 676737 117998
rect 675711 108146 675777 108147
rect 675711 108082 675712 108146
rect 675776 108082 675777 108146
rect 675711 108081 675777 108082
rect 674175 103262 674241 103263
rect 674175 103198 674176 103262
rect 674240 103198 674241 103262
rect 674175 103197 674241 103198
rect 676674 101487 676734 117997
rect 676671 101486 676737 101487
rect 676671 101422 676672 101486
rect 676736 101422 676737 101486
rect 676671 101421 676737 101422
rect 637695 52202 637761 52203
rect 637695 52138 637696 52202
rect 637760 52138 637761 52202
rect 637695 52137 637761 52138
rect 637311 51906 637377 51907
rect 637311 51842 637312 51906
rect 637376 51842 637377 51906
rect 637311 51841 637377 51842
rect 189951 41842 190017 41843
rect 189951 41778 189952 41842
rect 190016 41778 190017 41842
rect 189951 41777 190017 41778
rect 194943 41842 195009 41843
rect 194943 41778 194944 41842
rect 195008 41778 195009 41842
rect 194943 41777 195009 41778
rect 458175 41842 458241 41843
rect 458175 41778 458176 41842
rect 458240 41778 458241 41842
rect 458175 41777 458241 41778
rect 465663 41842 465729 41843
rect 465663 41778 465664 41842
rect 465728 41778 465729 41842
rect 465663 41777 465729 41778
rect 189954 40807 190014 41777
rect 189951 40806 190017 40807
rect 189951 40742 189952 40806
rect 190016 40742 190017 40806
rect 189951 40741 190017 40742
rect 194946 40659 195006 41777
rect 194943 40658 195009 40659
rect 194943 40594 194944 40658
rect 195008 40594 195009 40658
rect 194943 40593 195009 40594
rect 458178 40411 458238 41777
<< via4 >>
rect 457706 40362 457942 40411
rect 457706 40298 457792 40362
rect 457792 40298 457856 40362
rect 457856 40298 457942 40362
rect 457706 40175 457942 40298
rect 458090 40175 458326 40411
<< metal5 >>
rect 457664 40411 458368 40453
rect 457664 40175 457706 40411
rect 457942 40175 458090 40411
rect 458326 40175 458368 40411
rect 457664 40133 458368 40175
use user_id_programming  user_id_value
timestamp 1607580681
transform 1 0 656624 0 1 80926
box 0 0 7109 7077
use storage  storage
timestamp 1607580681
transform 1 0 52032 0 1 53156
box 38 0 88934 189234
use mgmt_core  soc
timestamp 1607580681
transform 1 0 210400 0 1 53700
box 0 0 430000 180000
use sky130_fd_sc_hvl__lsbufhv2lv_1_wrapped  rstb_level
timestamp 1607580681
transform -1 0 159876 0 -1 56488
box 66 33 5058 5084
use simple_por  por
timestamp 1607580681
transform 1 0 654176 0 1 104538
box 25 11 11344 8291
use gpio_control_block  gpio_control_bidir\[1\]
timestamp 1607580681
transform -1 0 708537 0 1 166200
box 38 0 33934 18344
use gpio_control_block  gpio_control_bidir\[0\]
timestamp 1607580681
transform -1 0 708537 0 1 121000
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[36\]
timestamp 1607580681
transform 1 0 8567 0 1 245800
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[37\]
timestamp 1607580681
transform 1 0 8567 0 1 202600
box 38 0 33934 18344
use mgmt_protect  mgmt_buffers
timestamp 1607580681
transform 1 0 215796 0 1 247292
box -1586 -1602 201502 12482
use gpio_control_block  gpio_control_in\[2\]
timestamp 1607580681
transform -1 0 708537 0 1 211200
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[3\]
timestamp 1607580681
transform -1 0 708537 0 1 256400
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[33\]
timestamp 1607580681
transform 1 0 8567 0 1 375400
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[34\]
timestamp 1607580681
transform 1 0 8567 0 1 332200
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[35\]
timestamp 1607580681
transform 1 0 8567 0 1 289000
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[4\]
timestamp 1607580681
transform -1 0 708537 0 1 301400
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[5\]
timestamp 1607580681
transform -1 0 708537 0 1 346400
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[7\]
timestamp 1607580681
transform -1 0 708537 0 1 479800
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[6\]
timestamp 1607580681
transform -1 0 708537 0 1 391600
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[32\]
timestamp 1607580681
transform 1 0 8567 0 1 418600
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[31\]
timestamp 1607580681
transform 1 0 8567 0 1 546200
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[30\]
timestamp 1607580681
transform 1 0 8567 0 1 589400
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[29\]
timestamp 1607580681
transform 1 0 8567 0 1 632600
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[9\]
timestamp 1607580681
transform -1 0 708537 0 1 568800
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[8\]
timestamp 1607580681
transform -1 0 708537 0 1 523800
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[10\]
timestamp 1607580681
transform -1 0 708537 0 1 614000
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[28\]
timestamp 1607580681
transform 1 0 8567 0 1 675800
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[27\]
timestamp 1607580681
transform 1 0 8567 0 1 719000
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[26\]
timestamp 1607580681
transform 1 0 8567 0 1 762200
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[13\]
timestamp 1607580681
transform -1 0 708537 0 1 749200
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[12\]
timestamp 1607580681
transform -1 0 708537 0 1 704200
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[11\]
timestamp 1607580681
transform -1 0 708537 0 1 659000
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[25\]
timestamp 1607580681
transform 1 0 8567 0 1 805400
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[24\]
timestamp 1607580681
transform 1 0 8567 0 1 931224
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[23\]
timestamp 1607580681
transform 0 1 97200 -1 0 1029747
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[22\]
timestamp 1607580681
transform 0 1 148600 -1 0 1029747
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[21\]
timestamp 1607580681
transform 0 1 200000 -1 0 1029747
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[20\]
timestamp 1607580681
transform 0 1 251400 -1 0 1029747
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[19\]
timestamp 1607580681
transform 0 1 303000 -1 0 1029747
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[18\]
timestamp 1607580681
transform 0 1 353400 -1 0 1029747
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[17\]
timestamp 1607580681
transform 0 1 420800 -1 0 1029747
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[16\]
timestamp 1607580681
transform 0 1 497800 -1 0 1029747
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[15\]
timestamp 1607580681
transform 0 1 549200 -1 0 1029747
box 38 0 33934 18344
use gpio_control_block  gpio_control_in\[14\]
timestamp 1607580681
transform -1 0 708537 0 1 927600
box 38 0 33934 18344
use user_project_wrapper  mprj
timestamp 1607580681
transform 1 0 65308 0 1 276608
box -8576 -7506 592500 711442
use chip_io  padframe
timestamp 1607580681
transform 1 0 0 0 1 0
box 0 0 717600 1037600
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
