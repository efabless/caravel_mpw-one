magic
tech sky130A
magscale 12 1
timestamp 1598787010
<< metal5 >>
rect 15 90 30 105
rect 0 75 30 90
rect 15 15 30 75
rect 0 0 45 15
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
