// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

/* Generated by Yosys 0.9+3621 (git sha1 84e9fa7, gcc 8.3.1 -fPIC -Os) */

module mgmt_protect(caravel_clk, caravel_clk2, caravel_rstn, mprj_cyc_o_core, mprj_cyc_o_user, mprj_stb_o_core, mprj_stb_o_user, mprj_we_o_core, mprj_we_o_user, user1_vcc_powergood, user1_vdd_powergood, user2_vcc_powergood, user2_vdd_powergood, user_clock, user_clock2, user_reset, user_resetn, vccd1, vssd1, vccd, vssd, vccd2, vssd2, vdda1, vssa1, vdda2, vssa2, la_data_in_core, la_data_in_mprj, la_data_out_core, la_data_out_mprj, la_oen_core, la_oen_mprj, mprj_adr_o_core, mprj_adr_o_user, mprj_dat_o_core, mprj_dat_o_user, mprj_sel_o_core, mprj_sel_o_user);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire _283_;
  wire _284_;
  wire _285_;
  wire _286_;
  wire _287_;
  wire _288_;
  wire _289_;
  wire _290_;
  wire _291_;
  wire _292_;
  wire _293_;
  wire _294_;
  wire _295_;
  wire _296_;
  wire _297_;
  wire _298_;
  wire _299_;
  wire _300_;
  wire _301_;
  wire _302_;
  wire _303_;
  wire _304_;
  wire _305_;
  wire _306_;
  wire _307_;
  wire _308_;
  wire _309_;
  wire _310_;
  wire _311_;
  wire _312_;
  wire _313_;
  wire _314_;
  wire _315_;
  wire _316_;
  wire _317_;
  wire _318_;
  wire _319_;
  wire _320_;
  wire _321_;
  wire _322_;
  wire _323_;
  wire _324_;
  wire _325_;
  wire _326_;
  wire _327_;
  wire _328_;
  wire _329_;
  input caravel_clk;
  input caravel_clk2;
  input caravel_rstn;
  output [127:0] la_data_in_core;
  output [127:0] la_data_in_mprj;
  wire \la_data_in_mprj_bar[0] ;
  wire \la_data_in_mprj_bar[100] ;
  wire \la_data_in_mprj_bar[101] ;
  wire \la_data_in_mprj_bar[102] ;
  wire \la_data_in_mprj_bar[103] ;
  wire \la_data_in_mprj_bar[104] ;
  wire \la_data_in_mprj_bar[105] ;
  wire \la_data_in_mprj_bar[106] ;
  wire \la_data_in_mprj_bar[107] ;
  wire \la_data_in_mprj_bar[108] ;
  wire \la_data_in_mprj_bar[109] ;
  wire \la_data_in_mprj_bar[10] ;
  wire \la_data_in_mprj_bar[110] ;
  wire \la_data_in_mprj_bar[111] ;
  wire \la_data_in_mprj_bar[112] ;
  wire \la_data_in_mprj_bar[113] ;
  wire \la_data_in_mprj_bar[114] ;
  wire \la_data_in_mprj_bar[115] ;
  wire \la_data_in_mprj_bar[116] ;
  wire \la_data_in_mprj_bar[117] ;
  wire \la_data_in_mprj_bar[118] ;
  wire \la_data_in_mprj_bar[119] ;
  wire \la_data_in_mprj_bar[11] ;
  wire \la_data_in_mprj_bar[120] ;
  wire \la_data_in_mprj_bar[121] ;
  wire \la_data_in_mprj_bar[122] ;
  wire \la_data_in_mprj_bar[123] ;
  wire \la_data_in_mprj_bar[124] ;
  wire \la_data_in_mprj_bar[125] ;
  wire \la_data_in_mprj_bar[126] ;
  wire \la_data_in_mprj_bar[127] ;
  wire \la_data_in_mprj_bar[12] ;
  wire \la_data_in_mprj_bar[13] ;
  wire \la_data_in_mprj_bar[14] ;
  wire \la_data_in_mprj_bar[15] ;
  wire \la_data_in_mprj_bar[16] ;
  wire \la_data_in_mprj_bar[17] ;
  wire \la_data_in_mprj_bar[18] ;
  wire \la_data_in_mprj_bar[19] ;
  wire \la_data_in_mprj_bar[1] ;
  wire \la_data_in_mprj_bar[20] ;
  wire \la_data_in_mprj_bar[21] ;
  wire \la_data_in_mprj_bar[22] ;
  wire \la_data_in_mprj_bar[23] ;
  wire \la_data_in_mprj_bar[24] ;
  wire \la_data_in_mprj_bar[25] ;
  wire \la_data_in_mprj_bar[26] ;
  wire \la_data_in_mprj_bar[27] ;
  wire \la_data_in_mprj_bar[28] ;
  wire \la_data_in_mprj_bar[29] ;
  wire \la_data_in_mprj_bar[2] ;
  wire \la_data_in_mprj_bar[30] ;
  wire \la_data_in_mprj_bar[31] ;
  wire \la_data_in_mprj_bar[32] ;
  wire \la_data_in_mprj_bar[33] ;
  wire \la_data_in_mprj_bar[34] ;
  wire \la_data_in_mprj_bar[35] ;
  wire \la_data_in_mprj_bar[36] ;
  wire \la_data_in_mprj_bar[37] ;
  wire \la_data_in_mprj_bar[38] ;
  wire \la_data_in_mprj_bar[39] ;
  wire \la_data_in_mprj_bar[3] ;
  wire \la_data_in_mprj_bar[40] ;
  wire \la_data_in_mprj_bar[41] ;
  wire \la_data_in_mprj_bar[42] ;
  wire \la_data_in_mprj_bar[43] ;
  wire \la_data_in_mprj_bar[44] ;
  wire \la_data_in_mprj_bar[45] ;
  wire \la_data_in_mprj_bar[46] ;
  wire \la_data_in_mprj_bar[47] ;
  wire \la_data_in_mprj_bar[48] ;
  wire \la_data_in_mprj_bar[49] ;
  wire \la_data_in_mprj_bar[4] ;
  wire \la_data_in_mprj_bar[50] ;
  wire \la_data_in_mprj_bar[51] ;
  wire \la_data_in_mprj_bar[52] ;
  wire \la_data_in_mprj_bar[53] ;
  wire \la_data_in_mprj_bar[54] ;
  wire \la_data_in_mprj_bar[55] ;
  wire \la_data_in_mprj_bar[56] ;
  wire \la_data_in_mprj_bar[57] ;
  wire \la_data_in_mprj_bar[58] ;
  wire \la_data_in_mprj_bar[59] ;
  wire \la_data_in_mprj_bar[5] ;
  wire \la_data_in_mprj_bar[60] ;
  wire \la_data_in_mprj_bar[61] ;
  wire \la_data_in_mprj_bar[62] ;
  wire \la_data_in_mprj_bar[63] ;
  wire \la_data_in_mprj_bar[64] ;
  wire \la_data_in_mprj_bar[65] ;
  wire \la_data_in_mprj_bar[66] ;
  wire \la_data_in_mprj_bar[67] ;
  wire \la_data_in_mprj_bar[68] ;
  wire \la_data_in_mprj_bar[69] ;
  wire \la_data_in_mprj_bar[6] ;
  wire \la_data_in_mprj_bar[70] ;
  wire \la_data_in_mprj_bar[71] ;
  wire \la_data_in_mprj_bar[72] ;
  wire \la_data_in_mprj_bar[73] ;
  wire \la_data_in_mprj_bar[74] ;
  wire \la_data_in_mprj_bar[75] ;
  wire \la_data_in_mprj_bar[76] ;
  wire \la_data_in_mprj_bar[77] ;
  wire \la_data_in_mprj_bar[78] ;
  wire \la_data_in_mprj_bar[79] ;
  wire \la_data_in_mprj_bar[7] ;
  wire \la_data_in_mprj_bar[80] ;
  wire \la_data_in_mprj_bar[81] ;
  wire \la_data_in_mprj_bar[82] ;
  wire \la_data_in_mprj_bar[83] ;
  wire \la_data_in_mprj_bar[84] ;
  wire \la_data_in_mprj_bar[85] ;
  wire \la_data_in_mprj_bar[86] ;
  wire \la_data_in_mprj_bar[87] ;
  wire \la_data_in_mprj_bar[88] ;
  wire \la_data_in_mprj_bar[89] ;
  wire \la_data_in_mprj_bar[8] ;
  wire \la_data_in_mprj_bar[90] ;
  wire \la_data_in_mprj_bar[91] ;
  wire \la_data_in_mprj_bar[92] ;
  wire \la_data_in_mprj_bar[93] ;
  wire \la_data_in_mprj_bar[94] ;
  wire \la_data_in_mprj_bar[95] ;
  wire \la_data_in_mprj_bar[96] ;
  wire \la_data_in_mprj_bar[97] ;
  wire \la_data_in_mprj_bar[98] ;
  wire \la_data_in_mprj_bar[99] ;
  wire \la_data_in_mprj_bar[9] ;
  input [127:0] la_data_out_core;
  input [127:0] la_data_out_mprj;
  output [127:0] la_oen_core;
  input [127:0] la_oen_mprj;
  wire mprj2_vdd_logic1;
  input [31:0] mprj_adr_o_core;
  output [31:0] mprj_adr_o_user;
  input mprj_cyc_o_core;
  output mprj_cyc_o_user;
  input [31:0] mprj_dat_o_core;
  output [31:0] mprj_dat_o_user;
  wire \mprj_logic1[0] ;
  wire \mprj_logic1[100] ;
  wire \mprj_logic1[101] ;
  wire \mprj_logic1[102] ;
  wire \mprj_logic1[103] ;
  wire \mprj_logic1[104] ;
  wire \mprj_logic1[105] ;
  wire \mprj_logic1[106] ;
  wire \mprj_logic1[107] ;
  wire \mprj_logic1[108] ;
  wire \mprj_logic1[109] ;
  wire \mprj_logic1[10] ;
  wire \mprj_logic1[110] ;
  wire \mprj_logic1[111] ;
  wire \mprj_logic1[112] ;
  wire \mprj_logic1[113] ;
  wire \mprj_logic1[114] ;
  wire \mprj_logic1[115] ;
  wire \mprj_logic1[116] ;
  wire \mprj_logic1[117] ;
  wire \mprj_logic1[118] ;
  wire \mprj_logic1[119] ;
  wire \mprj_logic1[11] ;
  wire \mprj_logic1[120] ;
  wire \mprj_logic1[121] ;
  wire \mprj_logic1[122] ;
  wire \mprj_logic1[123] ;
  wire \mprj_logic1[124] ;
  wire \mprj_logic1[125] ;
  wire \mprj_logic1[126] ;
  wire \mprj_logic1[127] ;
  wire \mprj_logic1[128] ;
  wire \mprj_logic1[129] ;
  wire \mprj_logic1[12] ;
  wire \mprj_logic1[130] ;
  wire \mprj_logic1[131] ;
  wire \mprj_logic1[132] ;
  wire \mprj_logic1[133] ;
  wire \mprj_logic1[134] ;
  wire \mprj_logic1[135] ;
  wire \mprj_logic1[136] ;
  wire \mprj_logic1[137] ;
  wire \mprj_logic1[138] ;
  wire \mprj_logic1[139] ;
  wire \mprj_logic1[13] ;
  wire \mprj_logic1[140] ;
  wire \mprj_logic1[141] ;
  wire \mprj_logic1[142] ;
  wire \mprj_logic1[143] ;
  wire \mprj_logic1[144] ;
  wire \mprj_logic1[145] ;
  wire \mprj_logic1[146] ;
  wire \mprj_logic1[147] ;
  wire \mprj_logic1[148] ;
  wire \mprj_logic1[149] ;
  wire \mprj_logic1[14] ;
  wire \mprj_logic1[150] ;
  wire \mprj_logic1[151] ;
  wire \mprj_logic1[152] ;
  wire \mprj_logic1[153] ;
  wire \mprj_logic1[154] ;
  wire \mprj_logic1[155] ;
  wire \mprj_logic1[156] ;
  wire \mprj_logic1[157] ;
  wire \mprj_logic1[158] ;
  wire \mprj_logic1[159] ;
  wire \mprj_logic1[15] ;
  wire \mprj_logic1[160] ;
  wire \mprj_logic1[161] ;
  wire \mprj_logic1[162] ;
  wire \mprj_logic1[163] ;
  wire \mprj_logic1[164] ;
  wire \mprj_logic1[165] ;
  wire \mprj_logic1[166] ;
  wire \mprj_logic1[167] ;
  wire \mprj_logic1[168] ;
  wire \mprj_logic1[169] ;
  wire \mprj_logic1[16] ;
  wire \mprj_logic1[170] ;
  wire \mprj_logic1[171] ;
  wire \mprj_logic1[172] ;
  wire \mprj_logic1[173] ;
  wire \mprj_logic1[174] ;
  wire \mprj_logic1[175] ;
  wire \mprj_logic1[176] ;
  wire \mprj_logic1[177] ;
  wire \mprj_logic1[178] ;
  wire \mprj_logic1[179] ;
  wire \mprj_logic1[17] ;
  wire \mprj_logic1[180] ;
  wire \mprj_logic1[181] ;
  wire \mprj_logic1[182] ;
  wire \mprj_logic1[183] ;
  wire \mprj_logic1[184] ;
  wire \mprj_logic1[185] ;
  wire \mprj_logic1[186] ;
  wire \mprj_logic1[187] ;
  wire \mprj_logic1[188] ;
  wire \mprj_logic1[189] ;
  wire \mprj_logic1[18] ;
  wire \mprj_logic1[190] ;
  wire \mprj_logic1[191] ;
  wire \mprj_logic1[192] ;
  wire \mprj_logic1[193] ;
  wire \mprj_logic1[194] ;
  wire \mprj_logic1[195] ;
  wire \mprj_logic1[196] ;
  wire \mprj_logic1[197] ;
  wire \mprj_logic1[198] ;
  wire \mprj_logic1[199] ;
  wire \mprj_logic1[19] ;
  wire \mprj_logic1[1] ;
  wire \mprj_logic1[200] ;
  wire \mprj_logic1[201] ;
  wire \mprj_logic1[202] ;
  wire \mprj_logic1[203] ;
  wire \mprj_logic1[204] ;
  wire \mprj_logic1[205] ;
  wire \mprj_logic1[206] ;
  wire \mprj_logic1[207] ;
  wire \mprj_logic1[208] ;
  wire \mprj_logic1[209] ;
  wire \mprj_logic1[20] ;
  wire \mprj_logic1[210] ;
  wire \mprj_logic1[211] ;
  wire \mprj_logic1[212] ;
  wire \mprj_logic1[213] ;
  wire \mprj_logic1[214] ;
  wire \mprj_logic1[215] ;
  wire \mprj_logic1[216] ;
  wire \mprj_logic1[217] ;
  wire \mprj_logic1[218] ;
  wire \mprj_logic1[219] ;
  wire \mprj_logic1[21] ;
  wire \mprj_logic1[220] ;
  wire \mprj_logic1[221] ;
  wire \mprj_logic1[222] ;
  wire \mprj_logic1[223] ;
  wire \mprj_logic1[224] ;
  wire \mprj_logic1[225] ;
  wire \mprj_logic1[226] ;
  wire \mprj_logic1[227] ;
  wire \mprj_logic1[228] ;
  wire \mprj_logic1[229] ;
  wire \mprj_logic1[22] ;
  wire \mprj_logic1[230] ;
  wire \mprj_logic1[231] ;
  wire \mprj_logic1[232] ;
  wire \mprj_logic1[233] ;
  wire \mprj_logic1[234] ;
  wire \mprj_logic1[235] ;
  wire \mprj_logic1[236] ;
  wire \mprj_logic1[237] ;
  wire \mprj_logic1[238] ;
  wire \mprj_logic1[239] ;
  wire \mprj_logic1[23] ;
  wire \mprj_logic1[240] ;
  wire \mprj_logic1[241] ;
  wire \mprj_logic1[242] ;
  wire \mprj_logic1[243] ;
  wire \mprj_logic1[244] ;
  wire \mprj_logic1[245] ;
  wire \mprj_logic1[246] ;
  wire \mprj_logic1[247] ;
  wire \mprj_logic1[248] ;
  wire \mprj_logic1[249] ;
  wire \mprj_logic1[24] ;
  wire \mprj_logic1[250] ;
  wire \mprj_logic1[251] ;
  wire \mprj_logic1[252] ;
  wire \mprj_logic1[253] ;
  wire \mprj_logic1[254] ;
  wire \mprj_logic1[255] ;
  wire \mprj_logic1[256] ;
  wire \mprj_logic1[257] ;
  wire \mprj_logic1[258] ;
  wire \mprj_logic1[259] ;
  wire \mprj_logic1[25] ;
  wire \mprj_logic1[260] ;
  wire \mprj_logic1[261] ;
  wire \mprj_logic1[262] ;
  wire \mprj_logic1[263] ;
  wire \mprj_logic1[264] ;
  wire \mprj_logic1[265] ;
  wire \mprj_logic1[266] ;
  wire \mprj_logic1[267] ;
  wire \mprj_logic1[268] ;
  wire \mprj_logic1[269] ;
  wire \mprj_logic1[26] ;
  wire \mprj_logic1[270] ;
  wire \mprj_logic1[271] ;
  wire \mprj_logic1[272] ;
  wire \mprj_logic1[273] ;
  wire \mprj_logic1[274] ;
  wire \mprj_logic1[275] ;
  wire \mprj_logic1[276] ;
  wire \mprj_logic1[277] ;
  wire \mprj_logic1[278] ;
  wire \mprj_logic1[279] ;
  wire \mprj_logic1[27] ;
  wire \mprj_logic1[280] ;
  wire \mprj_logic1[281] ;
  wire \mprj_logic1[282] ;
  wire \mprj_logic1[283] ;
  wire \mprj_logic1[284] ;
  wire \mprj_logic1[285] ;
  wire \mprj_logic1[286] ;
  wire \mprj_logic1[287] ;
  wire \mprj_logic1[288] ;
  wire \mprj_logic1[289] ;
  wire \mprj_logic1[28] ;
  wire \mprj_logic1[290] ;
  wire \mprj_logic1[291] ;
  wire \mprj_logic1[292] ;
  wire \mprj_logic1[293] ;
  wire \mprj_logic1[294] ;
  wire \mprj_logic1[295] ;
  wire \mprj_logic1[296] ;
  wire \mprj_logic1[297] ;
  wire \mprj_logic1[298] ;
  wire \mprj_logic1[299] ;
  wire \mprj_logic1[29] ;
  wire \mprj_logic1[2] ;
  wire \mprj_logic1[300] ;
  wire \mprj_logic1[301] ;
  wire \mprj_logic1[302] ;
  wire \mprj_logic1[303] ;
  wire \mprj_logic1[304] ;
  wire \mprj_logic1[305] ;
  wire \mprj_logic1[306] ;
  wire \mprj_logic1[307] ;
  wire \mprj_logic1[308] ;
  wire \mprj_logic1[309] ;
  wire \mprj_logic1[30] ;
  wire \mprj_logic1[310] ;
  wire \mprj_logic1[311] ;
  wire \mprj_logic1[312] ;
  wire \mprj_logic1[313] ;
  wire \mprj_logic1[314] ;
  wire \mprj_logic1[315] ;
  wire \mprj_logic1[316] ;
  wire \mprj_logic1[317] ;
  wire \mprj_logic1[318] ;
  wire \mprj_logic1[319] ;
  wire \mprj_logic1[31] ;
  wire \mprj_logic1[320] ;
  wire \mprj_logic1[321] ;
  wire \mprj_logic1[322] ;
  wire \mprj_logic1[323] ;
  wire \mprj_logic1[324] ;
  wire \mprj_logic1[325] ;
  wire \mprj_logic1[326] ;
  wire \mprj_logic1[327] ;
  wire \mprj_logic1[328] ;
  wire \mprj_logic1[329] ;
  wire \mprj_logic1[32] ;
  wire \mprj_logic1[330] ;
  wire \mprj_logic1[331] ;
  wire \mprj_logic1[332] ;
  wire \mprj_logic1[333] ;
  wire \mprj_logic1[334] ;
  wire \mprj_logic1[335] ;
  wire \mprj_logic1[336] ;
  wire \mprj_logic1[337] ;
  wire \mprj_logic1[338] ;
  wire \mprj_logic1[339] ;
  wire \mprj_logic1[33] ;
  wire \mprj_logic1[340] ;
  wire \mprj_logic1[341] ;
  wire \mprj_logic1[342] ;
  wire \mprj_logic1[343] ;
  wire \mprj_logic1[344] ;
  wire \mprj_logic1[345] ;
  wire \mprj_logic1[346] ;
  wire \mprj_logic1[347] ;
  wire \mprj_logic1[348] ;
  wire \mprj_logic1[349] ;
  wire \mprj_logic1[34] ;
  wire \mprj_logic1[350] ;
  wire \mprj_logic1[351] ;
  wire \mprj_logic1[352] ;
  wire \mprj_logic1[353] ;
  wire \mprj_logic1[354] ;
  wire \mprj_logic1[355] ;
  wire \mprj_logic1[356] ;
  wire \mprj_logic1[357] ;
  wire \mprj_logic1[358] ;
  wire \mprj_logic1[359] ;
  wire \mprj_logic1[35] ;
  wire \mprj_logic1[360] ;
  wire \mprj_logic1[361] ;
  wire \mprj_logic1[362] ;
  wire \mprj_logic1[363] ;
  wire \mprj_logic1[364] ;
  wire \mprj_logic1[365] ;
  wire \mprj_logic1[366] ;
  wire \mprj_logic1[367] ;
  wire \mprj_logic1[368] ;
  wire \mprj_logic1[369] ;
  wire \mprj_logic1[36] ;
  wire \mprj_logic1[370] ;
  wire \mprj_logic1[371] ;
  wire \mprj_logic1[372] ;
  wire \mprj_logic1[373] ;
  wire \mprj_logic1[374] ;
  wire \mprj_logic1[375] ;
  wire \mprj_logic1[376] ;
  wire \mprj_logic1[377] ;
  wire \mprj_logic1[378] ;
  wire \mprj_logic1[379] ;
  wire \mprj_logic1[37] ;
  wire \mprj_logic1[380] ;
  wire \mprj_logic1[381] ;
  wire \mprj_logic1[382] ;
  wire \mprj_logic1[383] ;
  wire \mprj_logic1[384] ;
  wire \mprj_logic1[385] ;
  wire \mprj_logic1[386] ;
  wire \mprj_logic1[387] ;
  wire \mprj_logic1[388] ;
  wire \mprj_logic1[389] ;
  wire \mprj_logic1[38] ;
  wire \mprj_logic1[390] ;
  wire \mprj_logic1[391] ;
  wire \mprj_logic1[392] ;
  wire \mprj_logic1[393] ;
  wire \mprj_logic1[394] ;
  wire \mprj_logic1[395] ;
  wire \mprj_logic1[396] ;
  wire \mprj_logic1[397] ;
  wire \mprj_logic1[398] ;
  wire \mprj_logic1[399] ;
  wire \mprj_logic1[39] ;
  wire \mprj_logic1[3] ;
  wire \mprj_logic1[400] ;
  wire \mprj_logic1[401] ;
  wire \mprj_logic1[402] ;
  wire \mprj_logic1[403] ;
  wire \mprj_logic1[404] ;
  wire \mprj_logic1[405] ;
  wire \mprj_logic1[406] ;
  wire \mprj_logic1[407] ;
  wire \mprj_logic1[408] ;
  wire \mprj_logic1[409] ;
  wire \mprj_logic1[40] ;
  wire \mprj_logic1[410] ;
  wire \mprj_logic1[411] ;
  wire \mprj_logic1[412] ;
  wire \mprj_logic1[413] ;
  wire \mprj_logic1[414] ;
  wire \mprj_logic1[415] ;
  wire \mprj_logic1[416] ;
  wire \mprj_logic1[417] ;
  wire \mprj_logic1[418] ;
  wire \mprj_logic1[419] ;
  wire \mprj_logic1[41] ;
  wire \mprj_logic1[420] ;
  wire \mprj_logic1[421] ;
  wire \mprj_logic1[422] ;
  wire \mprj_logic1[423] ;
  wire \mprj_logic1[424] ;
  wire \mprj_logic1[425] ;
  wire \mprj_logic1[426] ;
  wire \mprj_logic1[427] ;
  wire \mprj_logic1[428] ;
  wire \mprj_logic1[429] ;
  wire \mprj_logic1[42] ;
  wire \mprj_logic1[430] ;
  wire \mprj_logic1[431] ;
  wire \mprj_logic1[432] ;
  wire \mprj_logic1[433] ;
  wire \mprj_logic1[434] ;
  wire \mprj_logic1[435] ;
  wire \mprj_logic1[436] ;
  wire \mprj_logic1[437] ;
  wire \mprj_logic1[438] ;
  wire \mprj_logic1[439] ;
  wire \mprj_logic1[43] ;
  wire \mprj_logic1[440] ;
  wire \mprj_logic1[441] ;
  wire \mprj_logic1[442] ;
  wire \mprj_logic1[443] ;
  wire \mprj_logic1[444] ;
  wire \mprj_logic1[445] ;
  wire \mprj_logic1[446] ;
  wire \mprj_logic1[447] ;
  wire \mprj_logic1[448] ;
  wire \mprj_logic1[449] ;
  wire \mprj_logic1[44] ;
  wire \mprj_logic1[450] ;
  wire \mprj_logic1[451] ;
  wire \mprj_logic1[452] ;
  wire \mprj_logic1[453] ;
  wire \mprj_logic1[454] ;
  wire \mprj_logic1[455] ;
  wire \mprj_logic1[456] ;
  wire \mprj_logic1[457] ;
  wire \mprj_logic1[458] ;
  wire \mprj_logic1[45] ;
  wire \mprj_logic1[46] ;
  wire \mprj_logic1[47] ;
  wire \mprj_logic1[48] ;
  wire \mprj_logic1[49] ;
  wire \mprj_logic1[4] ;
  wire \mprj_logic1[50] ;
  wire \mprj_logic1[51] ;
  wire \mprj_logic1[52] ;
  wire \mprj_logic1[53] ;
  wire \mprj_logic1[54] ;
  wire \mprj_logic1[55] ;
  wire \mprj_logic1[56] ;
  wire \mprj_logic1[57] ;
  wire \mprj_logic1[58] ;
  wire \mprj_logic1[59] ;
  wire \mprj_logic1[5] ;
  wire \mprj_logic1[60] ;
  wire \mprj_logic1[61] ;
  wire \mprj_logic1[62] ;
  wire \mprj_logic1[63] ;
  wire \mprj_logic1[64] ;
  wire \mprj_logic1[65] ;
  wire \mprj_logic1[66] ;
  wire \mprj_logic1[67] ;
  wire \mprj_logic1[68] ;
  wire \mprj_logic1[69] ;
  wire \mprj_logic1[6] ;
  wire \mprj_logic1[70] ;
  wire \mprj_logic1[71] ;
  wire \mprj_logic1[72] ;
  wire \mprj_logic1[73] ;
  wire \mprj_logic1[74] ;
  wire \mprj_logic1[75] ;
  wire \mprj_logic1[76] ;
  wire \mprj_logic1[77] ;
  wire \mprj_logic1[78] ;
  wire \mprj_logic1[79] ;
  wire \mprj_logic1[7] ;
  wire \mprj_logic1[80] ;
  wire \mprj_logic1[81] ;
  wire \mprj_logic1[82] ;
  wire \mprj_logic1[83] ;
  wire \mprj_logic1[84] ;
  wire \mprj_logic1[85] ;
  wire \mprj_logic1[86] ;
  wire \mprj_logic1[87] ;
  wire \mprj_logic1[88] ;
  wire \mprj_logic1[89] ;
  wire \mprj_logic1[8] ;
  wire \mprj_logic1[90] ;
  wire \mprj_logic1[91] ;
  wire \mprj_logic1[92] ;
  wire \mprj_logic1[93] ;
  wire \mprj_logic1[94] ;
  wire \mprj_logic1[95] ;
  wire \mprj_logic1[96] ;
  wire \mprj_logic1[97] ;
  wire \mprj_logic1[98] ;
  wire \mprj_logic1[99] ;
  wire \mprj_logic1[9] ;
  input [3:0] mprj_sel_o_core;
  output [3:0] mprj_sel_o_user;
  input mprj_stb_o_core;
  output mprj_stb_o_user;
  wire mprj_vdd_logic1;
  input mprj_we_o_core;
  output mprj_we_o_user;
  output user1_vcc_powergood;
  output user1_vdd_powergood;
  output user2_vcc_powergood;
  output user2_vdd_powergood;
  output user_clock;
  output user_clock2;
  output user_reset;
  output user_resetn;
  input vccd;
  input vccd1;
  input vccd2;
  input vdda1;
  input vdda2;
  input vssa1;
  input vssa2;
  input vssd;
  input vssd1;
  input vssd2;
  sky130_fd_sc_hd__diode_2 ANTENNA_0 (
    .DIODE(la_oen_mprj[106]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_1 (
    .DIODE(la_oen_mprj[111]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_10 (
    .DIODE(la_oen_mprj[92]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_11 (
    .DIODE(la_oen_mprj[93]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_12 (
    .DIODE(la_oen_mprj[96]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_13 (
    .DIODE(la_oen_mprj[97]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_14 (
    .DIODE(la_oen_mprj[99]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_15 (
    .DIODE(mprj_sel_o_core[2]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_16 (
    .DIODE(mprj_we_o_core),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_2 (
    .DIODE(la_oen_mprj[121]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_3 (
    .DIODE(la_oen_mprj[125]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_4 (
    .DIODE(la_oen_mprj[68]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_5 (
    .DIODE(la_oen_mprj[78]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_6 (
    .DIODE(la_oen_mprj[80]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_7 (
    .DIODE(la_oen_mprj[82]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_8 (
    .DIODE(la_oen_mprj[89]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_9 (
    .DIODE(la_oen_mprj[91]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1002 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1013 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_1021 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1033 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1044 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_1052 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1055 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_106 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_1063 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1068 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_1080 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_1084 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_1086 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1099 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_1111 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_1115 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1117 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1128 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1139 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1157 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_1165 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1170 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_118 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1182 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1193 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_1205 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1213 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_1225 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1232 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1244 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_125 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1255 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_1267 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1275 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1286 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_1298 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_1303 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1310 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1325 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1337 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1348 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_1360 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1365 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_137 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1376 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1387 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1399 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1410 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_1422 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1430 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1441 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_1453 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1461 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1472 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_1484 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1489 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_149 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_1497 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_15 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1501 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1513 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_1520 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1525 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1537 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_1549 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_1551 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1556 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_0_156 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1567 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_1579 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1585 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1597 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_0_1609 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1613 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_162 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1624 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1636 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_1642 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1647 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_1659 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1666 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1678 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1690 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_0_1702 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1706 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_1714 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1728 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_173 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1740 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_1752 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1759 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1768 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1779 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1790 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1799 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1810 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1821 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_0_1830 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1836 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_1848 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_185 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1852 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1864 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_187 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1875 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_1887 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1895 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1906 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_1918 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_1923 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1927 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1938 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_0_1950 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_1954 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1961 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1972 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1985 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_199 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_1993 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1997 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_2009 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_2016 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_2022 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_2026 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_2037 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_2045 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_205 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_2050 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_2062 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_2069 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_2078 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_2086 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_209 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_2100 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_2121 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_2133 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_2140 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_218 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_223 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_234 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_246 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_249 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_253 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_264 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_27 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_0_276 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_280 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_292 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_296 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_3 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_300 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_308 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_311 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_32 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_323 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_335 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_0_342 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_348 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_359 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_371 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_376 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_388 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_0_400 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_404 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_415 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_427 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_433 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_435 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_44 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_447 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_453 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_457 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_466 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_473 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_48 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_484 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_497 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_509 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_521 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_531 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_542 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_554 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_562 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_574 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_578 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_0_586 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_590 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_598 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_60 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_608 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_621 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_629 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_639 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_66 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_661 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_673 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_681 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_683 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_695 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_707 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_714 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_726 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_738 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_754 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_766 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_77 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_774 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_785 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_796 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_804 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_816 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_824 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_829 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_847 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_855 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_860 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_869 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_880 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_89 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_891 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_909 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_917 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_921 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_929 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_94 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_940 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_948 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_953 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_971 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_982 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_990 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_1005 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_10_1008 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_101 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_1014 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1024 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_1032 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1042 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1059 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_1067 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1072 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_1080 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1086 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_1098 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1119 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_1127 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_1130 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1150 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1176 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_1188 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1200 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_1208 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_121 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1213 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_1221 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1240 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_1248 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1270 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1296 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_1308 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_1313 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_132 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1332 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_1340 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1360 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_1372 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_1374 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1396 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1422 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_143 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1438 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1464 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1475 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1486 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_1494 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1499 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_15 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_151 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1510 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_1522 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1542 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_1554 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1560 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1571 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_1583 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1602 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_1614 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1618 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1629 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1655 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_1663 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_172 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_183 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_19 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_194 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_206 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_215 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_23 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_237 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_263 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_294 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_3 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_305 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_317 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_10_32 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_328 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_355 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_366 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_378 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_38 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_389 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_398 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_405 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_417 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_429 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_10_441 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_450 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_10_459 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_465 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_484 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_510 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_518 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_538 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_550 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_569 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_57 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_577 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_584 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_596 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_616 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_633 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_651 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_663 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_673 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_690 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_703 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_714 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_731 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_748 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_760 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_773 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_790 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_802 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_815 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_823 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_825 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_83 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_837 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_848 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_859 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_876 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_884 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_895 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_10_907 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_91 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_922 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_93 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_933 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_945 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_950 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_962 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_966 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_976 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_993 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1003 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1024 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_1036 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_1038 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1060 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1077 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1088 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1096 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_11_1099 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1114 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1131 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_114 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1148 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_1156 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1169 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_1177 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1198 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1209 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_1217 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_1221 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1242 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_1254 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1273 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_1282 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_1286 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1290 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_1298 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1317 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1329 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1334 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_11_1343 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1352 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1378 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1389 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1401 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1407 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_141 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1433 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1444 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1455 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_1463 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1483 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_1495 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_15 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1517 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1526 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1552 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1563 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_1571 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1577 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_1585 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_11_1587 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1611 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1619 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1639 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1648 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1653 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_167 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_179 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_202 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_228 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_23 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_240 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_248 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_256 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_27 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_276 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_287 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_11_299 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_3 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_306 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_326 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_352 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_364 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_367 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_379 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_387 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_406 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_418 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_426 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_428 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_440 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_446 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_472 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_484 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_507 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_519 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_53 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_541 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_568 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_594 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_606 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_611 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_62 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_628 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_645 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_66 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_662 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_670 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_681 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_698 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_709 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_720 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_742 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_759 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_771 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_775 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_785 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_794 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_807 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_818 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_830 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_840 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_85 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_852 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_858 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_870 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_880 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_897 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_11_909 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_925 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_93 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_942 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_954 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_958 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_968 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_986 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1017 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1034 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1060 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1072 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1083 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_12_1095 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1119 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1127 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1139 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_1151 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1164 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1181 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1189 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_12_1191 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1215 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_122 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1241 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1249 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1255 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1270 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1296 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_1308 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1313 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1317 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_1325 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_133 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1346 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1357 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_1369 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1392 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1404 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_141 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1423 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_1431 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_145 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1453 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1464 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1475 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1486 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1494 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_15 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1514 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1525 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1537 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_154 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1541 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_1553 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1560 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1572 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1591 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_160 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1602 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_1614 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1618 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1622 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1633 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1644 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1670 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1697 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_1709 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1730 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1738 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1740 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1744 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1755 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1766 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1792 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1801 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1809 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1829 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1840 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1848 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1853 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1880 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1888 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_19 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_190 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1907 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_1919 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1941 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_1953 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1975 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_198 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1984 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1995 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_2003 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_202 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_2024 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_2035 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_2043 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_2063 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_2089 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_2101 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_2124 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_2135 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_2143 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_215 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_223 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_227 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_23 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_238 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_246 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_250 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_261 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_273 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_276 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_298 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_3 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_306 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_312 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_32 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_323 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_335 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_355 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_381 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_393 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_40 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_401 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_413 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_425 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_437 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_445 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_450 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_12_459 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_483 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_509 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_517 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_523 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_534 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_546 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_553 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_564 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_576 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_581 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_587 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_598 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_60 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_610 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_622 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_633 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_660 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_677 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_694 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_706 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_71 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_718 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_731 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_742 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_753 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_761 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_773 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_781 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_792 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_800 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_812 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_82 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_828 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_845 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_857 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_869 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_881 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_895 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_90 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_907 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_920 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_937 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_945 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_956 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_96 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_968 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_972 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_982 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_999 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1009 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1026 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_13_1034 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_13_104 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1047 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_13_1059 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1083 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_13_1095 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_110 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1102 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_1110 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1129 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_1137 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_114 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1147 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1163 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1171 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1191 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1208 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1224 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1232 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1252 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_126 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1267 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1279 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1285 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1293 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1298 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1309 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1320 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_13_1328 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1334 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_1343 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_1347 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1366 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_13_1374 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_13_138 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1395 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1404 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1430 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1456 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_13_1465 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_1471 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1490 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_15 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1516 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_1524 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1529 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1540 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1551 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_1559 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1578 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_1587 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1606 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1617 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_162 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1628 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1639 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_1648 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1652 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1678 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1689 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1700 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1727 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_173 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_1739 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1761 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_13_1770 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1779 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_13_1787 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1808 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_181 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_13_1816 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1822 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_1831 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1835 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_184 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1861 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1872 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1883 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_1892 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1911 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1937 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_13_1949 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_13_1953 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_1959 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_196 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1978 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_1986 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_2005 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_2032 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_2058 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_2070 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_2078 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_208 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_2090 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_2110 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_2121 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_2133 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_2136 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_2144 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_228 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_23 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_240 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_245 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_257 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_27 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_277 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_288 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_3 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_300 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_304 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_324 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_13_332 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_353 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_365 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_370 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_382 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_386 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_405 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_416 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_13_424 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_428 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_432 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_436 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_462 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_473 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_13_485 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_492 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_504 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_523 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_53 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_534 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_13_546 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_550 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_562 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_570 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_574 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_600 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_608 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_611 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_623 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_627 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_653 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_13_665 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_675 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_686 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_697 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_705 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_724 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_733 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_737 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_741 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_13_753 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_768 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_785 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_13_794 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_80 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_806 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_818 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_829 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_841 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_845 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_853 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_855 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_863 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_883 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_895 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_899 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_911 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_92 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_925 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_942 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_959 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_971 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_975 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_977 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_981 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_989 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_1003 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1011 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_1023 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1042 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_105 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1059 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_1067 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1072 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1083 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_109 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_1095 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1100 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1111 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_14_1123 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_14_1130 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1139 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1150 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1167 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1182 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1200 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_1212 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1234 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_1246 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_1250 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1252 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_1260 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1264 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_128 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1290 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1301 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_14_1309 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1331 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_1339 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1358 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_14_1370 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1374 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_1382 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_140 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1402 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1413 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1424 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_1432 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1438 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_145 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1468 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1479 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_1491 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_15 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1514 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1525 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1536 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1547 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_1555 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_157 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1575 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1601 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_1613 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1621 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_1629 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1633 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1644 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1670 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1697 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1708 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_1716 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1720 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1731 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1740 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1751 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1777 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1788 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_14_1801 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_1807 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1826 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_183 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_1834 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1853 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_1862 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1869 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1895 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_19 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_14_1907 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1913 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_1921 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1926 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_1938 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1943 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_195 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1969 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_1981 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1987 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_1995 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_2015 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_14_2027 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_2036 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_14_2045 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_2066 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_14_207 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_2092 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_2104 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_2124 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_213 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_2135 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_14_2143 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_215 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_219 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_223 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_23 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_235 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_247 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_259 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_271 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_276 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_283 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_3 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_309 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_14_32 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_321 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_14_333 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_340 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_351 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_363 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_375 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_387 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_395 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_416 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_428 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_450 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_459 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_481 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_507 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_523 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_535 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_547 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_559 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_56 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_571 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_579 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_14_581 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_605 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_617 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_629 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_633 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_651 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_662 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_67 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_673 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_684 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_14_696 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_703 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_708 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_719 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_730 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_14_738 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_744 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_755 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_773 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_78 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_785 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_807 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_819 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_823 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_834 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_14_846 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_861 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_872 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_884 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_889 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_90 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_901 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_923 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_93 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_934 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_950 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_961 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_969 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_973 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_981 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_991 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1015 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1033 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1044 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_1052 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1058 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_106 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1069 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_1081 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1089 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1100 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_1112 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1120 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1131 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_1143 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1148 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1159 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1170 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_1179 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_118 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1201 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1228 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1244 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1255 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_1267 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_128 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1290 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1306 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_1318 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1325 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_15_1334 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1355 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_1363 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_1365 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1387 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_140 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1414 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1430 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1441 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_1453 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1461 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1472 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_1484 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1492 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_15 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1503 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_1515 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_15_152 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1523 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1534 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_1546 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1554 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1565 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_1577 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1585 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1596 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_1608 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1616 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_1628 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1635 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1662 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1693 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1706 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1717 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1728 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1737 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_174 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1748 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1759 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1786 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1817 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_1830 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1852 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_187 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1879 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_15_1892 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_19 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1913 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_1921 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1923 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1934 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1945 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_1954 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1976 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_1985 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_199 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_2007 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_15_2016 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_2037 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_2045 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_2065 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_2078 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_2100 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_211 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_2127 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_2140 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_218 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_23 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_230 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_242 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_249 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_261 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_273 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_280 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_286 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_290 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_3 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_302 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_311 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_32 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_323 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_335 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_342 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_354 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_366 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_373 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_385 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_397 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_404 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_416 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_428 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_435 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_447 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_451 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_455 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_463 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_484 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_500 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_511 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_523 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_528 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_54 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_540 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_552 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_559 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_571 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_583 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_590 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_602 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_614 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_621 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_633 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_637 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_641 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_649 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_661 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_672 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_680 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_683 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_694 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_705 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_714 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_725 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_736 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_745 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_750 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_758 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_762 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_774 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_776 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_785 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_793 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_797 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_805 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_81 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_810 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_821 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_833 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_841 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_853 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_857 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_15_865 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_878 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_889 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_897 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_903 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_914 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_926 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_934 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_94 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_945 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_957 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_965 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_15_977 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_983 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_991 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_993 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1003 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_1015 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1027 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_1035 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1047 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_1055 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1067 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_1075 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1079 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1090 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_110 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1108 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_1_1120 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_1124 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1134 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_114 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1151 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1169 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1190 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_1202 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1208 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1224 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_123 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_1236 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1242 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1253 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1266 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_1278 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_1_1285 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_129 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_1291 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1297 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1308 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_1316 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1322 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1333 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_1341 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_1_1348 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_1352 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_1_1358 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1369 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_1377 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1382 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1393 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_140 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_1401 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1407 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1418 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_1430 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1434 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1445 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1456 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1468 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_1480 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1484 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1495 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_15 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1506 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1517 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_152 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1526 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1538 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_1550 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1555 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1566 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_1574 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1578 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1590 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1601 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1613 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1625 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1637 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_1645 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_1_1648 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1655 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1667 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_167 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_1679 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1684 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_1696 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1700 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_1_1709 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1716 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1727 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1738 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1749 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1760 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_1768 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_1_1770 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_1776 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1780 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_1_179 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1791 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_1_1803 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_1807 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1811 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1822 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1834 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_1_1846 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_1850 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1869 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_187 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1880 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_1888 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1895 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_1_1907 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1916 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_1924 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1930 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1941 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_1949 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_1953 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1957 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1968 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_1_1980 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1987 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_199 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_1999 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_2005 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_2017 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_2029 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_2033 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_2045 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_2051 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_2062 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_207 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_2075 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_2083 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_2087 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_2107 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_2118 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_213 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_1_2130 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_2134 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_2136 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_2144 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_221 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_225 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_236 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_248 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_1_260 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_269 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_27 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_280 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_292 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_3 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_304 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_306 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_314 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_319 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_330 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_341 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_352 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_364 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_370 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_385 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_1_39 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_397 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_401 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_413 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_418 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_426 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_1_428 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_437 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_445 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_450 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_458 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_462 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_473 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_48 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_485 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_489 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_493 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_504 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_515 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_527 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_535 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_541 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_559 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_576 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_584 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_594 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_60 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_1_606 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_614 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_626 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_636 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_65 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_653 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_1_665 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_681 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_698 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_715 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_1_727 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_731 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_742 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_76 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_763 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_780 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_792 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_803 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_811 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_823 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_840 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_852 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_864 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_87 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_881 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_898 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_1_910 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_914 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_925 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_933 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_944 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_961 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_973 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_98 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_986 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_1005 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_1008 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_1014 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1024 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1035 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_105 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1052 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_1064 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1078 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1095 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1112 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_1124 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_1128 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_1130 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1134 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_2_1142 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1154 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_116 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_1166 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1181 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_1189 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1200 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1211 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_1223 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_1227 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1231 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1242 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_1250 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1252 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_1260 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1264 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1275 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_128 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_1286 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_1292 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1298 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_1310 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1316 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_1328 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_1335 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_1346 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1357 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_136 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_1369 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1377 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_1388 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1399 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_2_1407 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_141 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1413 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1424 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_1432 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1438 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1468 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_1480 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1487 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1499 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_15 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1510 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1522 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1534 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1546 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_1554 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_1557 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1562 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_157 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1574 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1586 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1598 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_1610 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_1616 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1618 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1630 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1642 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1654 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1666 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1679 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_169 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_1691 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1698 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1709 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1720 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_173 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1731 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1743 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_1755 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1764 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_177 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_1776 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1781 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1792 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1801 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_1809 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1813 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_1825 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1830 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_1842 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1851 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_1859 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1880 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_189 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1891 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1902 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_1910 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1914 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1923 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1949 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1975 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_2002 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_201 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_2028 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_2040 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_2048 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_2_2056 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_2062 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_2073 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_2084 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_2092 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_2097 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_2109 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_2120 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_213 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_2131 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_2_2143 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_218 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_229 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_241 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_250 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_258 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_263 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_27 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_279 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_291 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_3 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_303 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_315 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_32 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_327 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_335 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_337 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_352 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_364 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_376 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_380 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_392 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_396 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_398 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_402 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_414 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_426 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_438 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_2_44 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_446 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_450 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_462 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_2_470 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_476 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_487 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_498 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_50 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_509 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_517 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_520 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_2_532 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_538 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_553 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_564 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_576 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_581 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_585 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_596 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_608 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_61 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_618 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_630 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_2_638 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_642 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_655 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_2_667 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_679 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_691 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_2_699 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_703 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_709 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_719 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_72 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_736 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_744 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_755 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_764 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_770 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_780 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_2_788 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_800 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_811 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_823 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_825 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_83 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_835 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_852 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_869 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_881 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_886 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_893 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_91 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_910 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_922 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_93 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_933 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_945 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_950 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_958 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_969 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_986 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_997 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1007 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1024 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_1036 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1041 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_1053 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1064 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_1072 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1083 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_1095 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_1099 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1111 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_1123 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1128 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_1136 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_114 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1146 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_1158 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1169 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1186 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1197 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1208 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1226 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_1238 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1242 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_1250 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1256 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_126 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_1264 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1270 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_1278 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_3_1282 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_1286 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1290 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1301 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1312 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_3_1324 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1333 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_1341 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1343 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1354 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_137 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_3_1380 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1391 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1404 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_1412 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1417 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_1425 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1445 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1456 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1468 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_1476 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1484 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1495 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_15 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1506 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1517 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_152 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1529 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1541 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1553 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_1561 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1568 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_3_1580 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1587 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1599 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1611 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1623 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_1631 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1636 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_164 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_1644 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1648 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_3_1660 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_1664 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_3_176 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_182 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_184 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_196 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_207 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_215 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_219 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_231 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_243 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_245 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_256 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_267 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_27 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_279 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_284 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_296 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_3 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_304 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_309 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_321 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_3_333 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_337 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_341 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_35 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_352 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_364 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_367 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_379 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_391 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_40 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_403 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_415 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_3_428 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_434 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_438 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_450 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_455 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_466 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_477 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_485 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_492 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_504 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_51 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_512 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_518 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_530 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_541 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_550 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_561 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_572 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_583 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_59 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_595 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_607 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_3_611 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_615 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_619 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_631 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_65 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_652 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_3_664 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_670 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_681 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_689 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_701 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_718 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_730 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_742 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_76 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_763 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_780 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_792 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_797 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_818 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_835 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_846 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_864 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_87 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_875 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_3_887 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_902 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_914 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_925 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_933 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_938 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_955 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_966 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_974 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_986 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_99 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_4_1003 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1017 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1028 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1039 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_1047 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1057 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_4_1065 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1078 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_4_108 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1089 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1100 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1111 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_4_1123 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_1130 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1140 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1157 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1174 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_4_1186 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1194 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1205 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1216 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1227 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_1239 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1243 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1252 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1263 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1274 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_128 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_4_1282 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1287 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1298 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_4_1310 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_4_1313 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1318 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_4_1348 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_1354 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1360 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_1372 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1374 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_4_1382 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1387 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_140 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1417 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_4_1429 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_1433 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1438 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1449 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_4_1475 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1486 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_1494 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1499 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_15 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1510 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_152 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1521 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1536 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_154 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1548 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1562 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1574 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1586 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1598 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1609 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1618 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1630 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1642 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1654 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_166 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_4_1662 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_178 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_4_190 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_195 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_206 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_215 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_227 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_235 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_239 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_250 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_261 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_4_27 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_4_273 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_4_276 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_282 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_286 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_4_294 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_299 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_3 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_311 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_4_32 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_323 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_335 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_4_337 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_359 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_36 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_371 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_383 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_4_395 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_40 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_401 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_413 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_425 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_440 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_4_452 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_462 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_4_470 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_491 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_503 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_51 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_4_515 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_520 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_532 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_540 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_544 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_555 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_566 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_4_578 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_581 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_4_589 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_594 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_4_606 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_612 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_62 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_4_624 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_633 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_645 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_4_653 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_665 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_677 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_689 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_4_70 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_701 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_703 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_713 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_725 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_4_733 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_739 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_750 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_76 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_762 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_4_764 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_770 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_780 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_791 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_4_803 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_816 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_828 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_4_840 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_852 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_869 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_4_88 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_4_881 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_4_886 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_895 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_912 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_929 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_4_941 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_945 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_947 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_96 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_964 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_4_976 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_991 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1001 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1012 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1023 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1035 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_1038 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1050 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1062 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1073 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1090 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1102 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_111 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_1110 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1114 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1140 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1151 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1169 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1180 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_119 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1191 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1203 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1208 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1224 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_1232 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1251 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_126 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1262 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1273 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_5_1282 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1289 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1315 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_1327 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1333 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_1341 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_1343 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1349 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_137 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1375 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1386 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_5_1398 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_1402 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1404 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1424 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1450 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1462 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1468 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1479 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_1487 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_149 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_15 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1506 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1517 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1529 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1540 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1552 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1564 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1576 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1584 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1587 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1599 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_161 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1611 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1623 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1635 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1648 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_5_1660 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_1664 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_173 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_181 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_184 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_5_196 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_218 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_230 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_236 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_26 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_263 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_275 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_294 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_3 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_302 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_5_306 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_313 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_325 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_344 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_355 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_363 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_367 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_37 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_379 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_391 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_403 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_415 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_431 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_5_443 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_465 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_473 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_477 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_48 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_485 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_489 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_495 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_506 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_514 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_519 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_5_531 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_537 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_541 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_568 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_579 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_590 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_60 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_601 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_609 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_5_611 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_5_62 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_624 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_650 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_66 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_661 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_669 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_5_672 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_685 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_697 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_709 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_724 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_742 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_759 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_770 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_781 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_803 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_811 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_822 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_834 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_846 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_85 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_858 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_866 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_871 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_882 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_894 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_904 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_912 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_919 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_5_931 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_946 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_963 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_975 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_980 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_6_1001 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1017 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_104 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1047 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_6_1055 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1060 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1087 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_1099 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1120 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_1128 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1139 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_1147 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1151 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1177 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_1189 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1191 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1202 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1228 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1239 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_125 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1252 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_1260 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1279 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_1291 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1295 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_6_1307 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_1311 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1313 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1339 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_136 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1365 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1374 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_1382 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1401 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1412 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1423 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_1431 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1435 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1446 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_1454 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1473 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_6_148 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1484 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_1492 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1499 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_6_15 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_1507 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_152 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1528 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1539 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_6_1551 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_1555 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1557 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1569 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_157 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1581 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1593 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1605 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1618 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1630 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1642 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1654 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_1662 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_169 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_173 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_185 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_19 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_197 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_201 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_213 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_218 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_229 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_23 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_6_237 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_257 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_6_269 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_6_276 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_280 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_284 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_292 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_3 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_313 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_6_32 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_321 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_325 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_333 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_6_337 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_361 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_372 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_383 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_6_395 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_401 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_413 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_6_425 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_449 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_457 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_462 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_6_474 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_496 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_507 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_538 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_56 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_568 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_581 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_600 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_611 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_622 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_633 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_660 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_671 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_682 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_694 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_703 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_718 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_729 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_755 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_782 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_794 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_806 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_6_818 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_82 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_834 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_6_846 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_870 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_882 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_889 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_897 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_6_90 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_909 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_926 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_934 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_938 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_956 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_96 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_968 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_989 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1020 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_7_103 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_7_1032 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_1036 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_1047 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1058 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_1070 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_1089 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_109 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_1097 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_1099 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_11 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_1110 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_1136 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1147 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1169 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_7_1181 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_1185 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1195 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1207 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_121 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_1212 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_1239 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_1247 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1266 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_7_1278 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1282 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_1287 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1313 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_7_1325 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_1334 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_1361 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1369 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1389 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1401 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_1404 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_141 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_1412 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_1431 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_1442 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_1453 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_7_1461 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_1483 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1509 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_7_1521 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1529 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_7_1541 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1562 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1574 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1587 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1599 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_16 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1611 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1623 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1635 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_7_1648 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_1657 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_167 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_7_179 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_184 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_196 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_215 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_226 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_7_238 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_263 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_27 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_275 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_287 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_7_299 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_3 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_306 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_325 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_351 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_7_363 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_370 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_7_378 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_399 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_411 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_7_423 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_446 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_7_458 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_480 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_507 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_7_519 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_526 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_53 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_541 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_7_550 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_574 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_582 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_602 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_7_611 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_626 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_652 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_663 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_681 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_692 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_707 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_724 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_7_733 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_746 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_763 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_780 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_792 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_80 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_803 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_818 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_829 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_846 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_864 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_881 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_892 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_907 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_91 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_934 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_7_946 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_968 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_986 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_7_998 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_8_1001 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_8_1008 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1030 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_8_1038 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1059 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_1067 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1072 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1083 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1098 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_111 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_1110 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1121 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1133 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_1141 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1160 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1177 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_1189 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_12 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1209 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1235 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_8_1247 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1255 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1266 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1292 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_1300 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1304 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_1313 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1318 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1344 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_8_1356 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1365 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_137 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_1374 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1393 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_8_1405 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1426 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1453 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1479 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_8_149 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_8_1491 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1514 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1525 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1536 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_1544 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1548 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1560 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1571 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1583 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1595 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1607 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_1615 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1618 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1630 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_1638 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1657 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_172 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_8_184 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_206 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_8_215 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_23 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_237 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_263 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_279 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_287 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_291 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_8_3 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_317 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_32 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_328 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_8_337 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_343 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_369 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_8_377 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_383 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_395 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_40 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_416 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_427 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_8_439 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_443 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_447 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_8_455 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_8_459 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_465 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_469 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_495 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_506 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_518 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_523 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_535 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_555 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_566 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_578 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_59 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_599 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_8_611 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_633 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_642 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_662 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_679 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_690 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_70 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_8_703 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_709 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_713 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_739 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_754 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_762 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_782 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_799 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_81 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_816 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_8_825 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_849 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_875 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_883 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_8_89 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_895 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_906 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_917 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_929 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_934 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_965 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_8_977 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_989 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1007 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_1015 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_102 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1027 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1035 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_1038 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1050 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1067 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1078 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1089 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_1097 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_110 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1108 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_1116 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1135 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_114 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1146 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_1158 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1169 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1186 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1203 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_1215 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_1219 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_1221 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1228 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1254 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1266 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1271 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1279 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1300 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1326 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_1338 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1361 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_1369 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1388 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_1400 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1407 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_141 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_1415 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1434 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1445 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1456 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1465 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1485 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_15 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1511 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1523 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1529 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_153 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1540 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1570 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_1582 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1590 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1602 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1614 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_1622 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1628 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1639 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_9_1648 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1657 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_175 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_202 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_23 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_232 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_263 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_27 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_275 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_297 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_3 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_306 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_328 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_354 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_9_367 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_391 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_417 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_425 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_428 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_440 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_448 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_454 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_480 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_507 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_53 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_533 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_545 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_553 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_561 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_582 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_593 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_605 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_609 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_614 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_626 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_630 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_649 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_660 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_668 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_9_672 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_678 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_688 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_699 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_710 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_721 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_729 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_742 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_759 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_776 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_788 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_792 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_9_794 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_80 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_800 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_810 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_827 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_835 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_846 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_864 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_881 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_898 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_91 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_910 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_914 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_925 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_933 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_944 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_961 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_973 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_977 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_987 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_995 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_0 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_1 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_10 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_100 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_101 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_102 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_103 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_104 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_105 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_106 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_107 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_108 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_109 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_11 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_110 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_111 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_112 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_113 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_114 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_115 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_116 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_117 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_118 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_119 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_12 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_120 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_121 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_122 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_123 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_124 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_125 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_126 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_127 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_128 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_129 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_13 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_130 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_131 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_132 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_133 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_134 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_135 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_136 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_137 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_138 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_139 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_14 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_140 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_141 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_142 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_143 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_144 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_145 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_146 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_147 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_148 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_149 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_15 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_150 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_151 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_152 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_153 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_154 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_155 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_156 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_157 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_158 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_159 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_16 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_160 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_161 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_162 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_163 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_164 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_165 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_166 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_167 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_168 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_169 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_17 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_170 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_171 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_172 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_173 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_174 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_175 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_176 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_177 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_178 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_179 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_18 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_180 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_181 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_182 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_183 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_184 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_185 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_186 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_187 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_188 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_189 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_19 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_190 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_191 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_192 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_193 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_194 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_195 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_196 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_197 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_198 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_199 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_2 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_20 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_200 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_201 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_202 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_203 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_204 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_205 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_206 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_207 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_208 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_209 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_21 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_210 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_211 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_212 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_213 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_214 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_215 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_216 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_217 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_218 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_219 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_22 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_220 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_221 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_222 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_223 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_224 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_225 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_226 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_227 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_228 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_229 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_23 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_230 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_231 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_232 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_233 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_234 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_235 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_236 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_237 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_238 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_239 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_24 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_240 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_241 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_242 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_243 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_244 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_245 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_246 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_247 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_248 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_249 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_25 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_250 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_251 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_252 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_253 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_254 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_255 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_256 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_257 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_258 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_259 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_26 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_260 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_261 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_262 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_263 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_264 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_265 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_266 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_267 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_268 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_269 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_27 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_270 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_271 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_272 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_273 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_274 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_275 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_276 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_277 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_278 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_279 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_28 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_280 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_281 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_282 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_283 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_284 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_285 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_286 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_287 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_288 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_289 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_29 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_290 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_291 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_292 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_293 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_294 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_295 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_296 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_297 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_298 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_299 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_3 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_30 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_300 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_301 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_302 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_303 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_304 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_305 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_306 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_307 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_308 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_309 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_31 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_310 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_311 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_312 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_313 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_314 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_315 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_316 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_317 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_318 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_319 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_32 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_320 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_321 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_322 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_323 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_324 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_325 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_326 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_327 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_328 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_329 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_33 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_330 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_331 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_332 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_333 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_334 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_335 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_336 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_337 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_338 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_339 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_34 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_340 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_341 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_342 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_343 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_344 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_345 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_346 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_347 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_348 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_349 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_35 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_350 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_351 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_352 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_353 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_354 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_355 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_356 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_357 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_358 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_359 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_36 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_360 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_361 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_362 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_363 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_364 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_365 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_366 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_367 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_368 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_369 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_37 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_370 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_371 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_372 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_373 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_374 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_375 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_376 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_377 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_378 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_379 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_38 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_380 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_381 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_382 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_383 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_384 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_385 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_386 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_387 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_388 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_389 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_39 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_390 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_391 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_392 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_393 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_394 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_395 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_396 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_397 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_398 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_399 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_4 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_40 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_400 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_401 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_402 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_403 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_404 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_405 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_406 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_407 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_408 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_409 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_41 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_410 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_411 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_412 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_413 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_414 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_415 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_416 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_417 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_418 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_419 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_42 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_420 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_421 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_422 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_423 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_424 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_425 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_426 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_427 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_428 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_429 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_43 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_430 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_431 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_432 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_433 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_434 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_435 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_436 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_437 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_438 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_439 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_44 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_440 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_441 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_442 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_443 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_444 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_445 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_446 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_447 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_448 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_449 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_45 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_450 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_451 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_452 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_453 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_454 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_455 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_456 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_457 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_458 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_459 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_46 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_460 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_461 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_462 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_463 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_464 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_465 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_466 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_467 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_468 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_469 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_47 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_470 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_471 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_472 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_473 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_474 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_475 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_476 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_477 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_478 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_479 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_48 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_480 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_481 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_482 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_483 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_484 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_485 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_486 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_487 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_488 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_489 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_49 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_490 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_491 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_492 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_493 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_494 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_495 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_496 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_497 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_498 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_499 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_5 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_50 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_500 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_501 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_502 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_503 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_504 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_505 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_506 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_507 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_508 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_509 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_51 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_510 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_511 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_512 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_513 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_514 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_515 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_516 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_517 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_518 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_519 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_52 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_520 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_521 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_522 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_523 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_524 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_525 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_526 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_527 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_528 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_529 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_53 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_530 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_531 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_532 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_533 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_534 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_535 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_536 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_537 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_538 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_539 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_54 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_540 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_541 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_542 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_543 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_544 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_545 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_546 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_547 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_548 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_549 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_55 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_550 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_551 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_552 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_553 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_554 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_555 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_556 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_557 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_558 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_559 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_56 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_560 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_561 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_562 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_563 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_564 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_565 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_566 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_567 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_568 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_569 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_57 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_570 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_571 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_572 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_573 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_574 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_575 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_576 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_577 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_578 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_579 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_58 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_580 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_581 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_582 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_583 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_584 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_585 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_586 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_587 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_59 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_6 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_60 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_61 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_62 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_63 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_64 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_65 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_66 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_67 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_68 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_69 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_7 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_70 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_71 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_72 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_73 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_74 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_75 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_76 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_77 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_78 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_79 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_8 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_80 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_81 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_82 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_83 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_84 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_85 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_86 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_87 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_88 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_89 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__decap_3 PHY_9 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_90 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_91 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_92 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_93 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_94 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_95 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_96 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_97 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_98 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_99 (
    .VGND(vssa2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__inv_2 _330_ (
    .A(la_oen_mprj[62]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_288_)
  );
  sky130_fd_sc_hd__inv_2 _331_ (
    .A(la_oen_mprj[63]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_289_)
  );
  sky130_fd_sc_hd__inv_2 _332_ (
    .A(la_oen_mprj[64]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_290_)
  );
  sky130_fd_sc_hd__inv_2 _333_ (
    .A(la_oen_mprj[65]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_291_)
  );
  sky130_fd_sc_hd__inv_2 _334_ (
    .A(la_oen_mprj[66]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_292_)
  );
  sky130_fd_sc_hd__inv_2 _335_ (
    .A(la_oen_mprj[67]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_293_)
  );
  sky130_fd_sc_hd__inv_2 _336_ (
    .A(la_oen_mprj[68]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_294_)
  );
  sky130_fd_sc_hd__inv_2 _337_ (
    .A(la_oen_mprj[69]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_295_)
  );
  sky130_fd_sc_hd__inv_2 _338_ (
    .A(la_oen_mprj[70]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_297_)
  );
  sky130_fd_sc_hd__inv_2 _339_ (
    .A(la_oen_mprj[71]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_298_)
  );
  sky130_fd_sc_hd__inv_2 _340_ (
    .A(la_oen_mprj[72]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_299_)
  );
  sky130_fd_sc_hd__inv_2 _341_ (
    .A(la_oen_mprj[73]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_300_)
  );
  sky130_fd_sc_hd__inv_2 _342_ (
    .A(la_oen_mprj[74]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_301_)
  );
  sky130_fd_sc_hd__inv_2 _343_ (
    .A(la_oen_mprj[75]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_302_)
  );
  sky130_fd_sc_hd__inv_2 _344_ (
    .A(la_oen_mprj[76]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_303_)
  );
  sky130_fd_sc_hd__inv_2 _345_ (
    .A(la_oen_mprj[77]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_304_)
  );
  sky130_fd_sc_hd__inv_2 _346_ (
    .A(la_oen_mprj[78]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_305_)
  );
  sky130_fd_sc_hd__inv_2 _347_ (
    .A(la_oen_mprj[79]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_306_)
  );
  sky130_fd_sc_hd__inv_2 _348_ (
    .A(la_oen_mprj[80]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_308_)
  );
  sky130_fd_sc_hd__inv_2 _349_ (
    .A(la_oen_mprj[81]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_309_)
  );
  sky130_fd_sc_hd__inv_2 _350_ (
    .A(la_oen_mprj[82]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_310_)
  );
  sky130_fd_sc_hd__inv_2 _351_ (
    .A(la_oen_mprj[83]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_311_)
  );
  sky130_fd_sc_hd__inv_2 _352_ (
    .A(la_oen_mprj[84]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_312_)
  );
  sky130_fd_sc_hd__inv_2 _353_ (
    .A(la_oen_mprj[85]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_313_)
  );
  sky130_fd_sc_hd__inv_2 _354_ (
    .A(la_oen_mprj[86]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_314_)
  );
  sky130_fd_sc_hd__inv_2 _355_ (
    .A(la_oen_mprj[87]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_315_)
  );
  sky130_fd_sc_hd__inv_2 _356_ (
    .A(la_oen_mprj[88]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_316_)
  );
  sky130_fd_sc_hd__inv_2 _357_ (
    .A(la_oen_mprj[89]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_317_)
  );
  sky130_fd_sc_hd__inv_2 _358_ (
    .A(la_oen_mprj[90]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_319_)
  );
  sky130_fd_sc_hd__inv_2 _359_ (
    .A(la_oen_mprj[91]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_320_)
  );
  sky130_fd_sc_hd__inv_2 _360_ (
    .A(la_oen_mprj[92]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_321_)
  );
  sky130_fd_sc_hd__inv_2 _361_ (
    .A(la_oen_mprj[93]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_322_)
  );
  sky130_fd_sc_hd__inv_2 _362_ (
    .A(la_oen_mprj[94]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_323_)
  );
  sky130_fd_sc_hd__inv_2 _363_ (
    .A(la_oen_mprj[95]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_324_)
  );
  sky130_fd_sc_hd__inv_2 _364_ (
    .A(la_oen_mprj[96]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_325_)
  );
  sky130_fd_sc_hd__inv_2 _365_ (
    .A(la_oen_mprj[97]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_326_)
  );
  sky130_fd_sc_hd__inv_2 _366_ (
    .A(la_oen_mprj[98]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_327_)
  );
  sky130_fd_sc_hd__inv_2 _367_ (
    .A(la_oen_mprj[99]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_328_)
  );
  sky130_fd_sc_hd__inv_2 _368_ (
    .A(la_oen_mprj[100]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_203_)
  );
  sky130_fd_sc_hd__inv_2 _369_ (
    .A(la_oen_mprj[101]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_204_)
  );
  sky130_fd_sc_hd__inv_2 _370_ (
    .A(la_oen_mprj[102]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_205_)
  );
  sky130_fd_sc_hd__inv_2 _371_ (
    .A(la_oen_mprj[103]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_206_)
  );
  sky130_fd_sc_hd__inv_2 _372_ (
    .A(la_oen_mprj[104]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_207_)
  );
  sky130_fd_sc_hd__inv_2 _373_ (
    .A(la_oen_mprj[105]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_208_)
  );
  sky130_fd_sc_hd__inv_2 _374_ (
    .A(la_oen_mprj[106]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_209_)
  );
  sky130_fd_sc_hd__inv_2 _375_ (
    .A(la_oen_mprj[107]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_210_)
  );
  sky130_fd_sc_hd__inv_2 _376_ (
    .A(la_oen_mprj[108]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_211_)
  );
  sky130_fd_sc_hd__inv_2 _377_ (
    .A(la_oen_mprj[109]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_212_)
  );
  sky130_fd_sc_hd__inv_2 _378_ (
    .A(la_oen_mprj[110]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_214_)
  );
  sky130_fd_sc_hd__inv_2 _379_ (
    .A(la_oen_mprj[111]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_215_)
  );
  sky130_fd_sc_hd__inv_2 _380_ (
    .A(la_oen_mprj[112]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_216_)
  );
  sky130_fd_sc_hd__inv_2 _381_ (
    .A(la_oen_mprj[113]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_217_)
  );
  sky130_fd_sc_hd__inv_2 _382_ (
    .A(la_oen_mprj[114]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_218_)
  );
  sky130_fd_sc_hd__inv_2 _383_ (
    .A(la_oen_mprj[115]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_219_)
  );
  sky130_fd_sc_hd__inv_2 _384_ (
    .A(la_oen_mprj[116]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_220_)
  );
  sky130_fd_sc_hd__inv_2 _385_ (
    .A(la_oen_mprj[117]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_221_)
  );
  sky130_fd_sc_hd__inv_2 _386_ (
    .A(la_oen_mprj[118]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_222_)
  );
  sky130_fd_sc_hd__inv_2 _387_ (
    .A(la_oen_mprj[119]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_223_)
  );
  sky130_fd_sc_hd__inv_2 _388_ (
    .A(la_oen_mprj[120]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_225_)
  );
  sky130_fd_sc_hd__inv_2 _389_ (
    .A(la_oen_mprj[121]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_226_)
  );
  sky130_fd_sc_hd__inv_2 _390_ (
    .A(la_oen_mprj[122]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_227_)
  );
  sky130_fd_sc_hd__inv_2 _391_ (
    .A(la_oen_mprj[123]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_228_)
  );
  sky130_fd_sc_hd__inv_2 _392_ (
    .A(la_oen_mprj[124]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_229_)
  );
  sky130_fd_sc_hd__inv_2 _393_ (
    .A(la_oen_mprj[125]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_230_)
  );
  sky130_fd_sc_hd__inv_2 _394_ (
    .A(la_oen_mprj[126]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_231_)
  );
  sky130_fd_sc_hd__inv_2 _395_ (
    .A(la_oen_mprj[127]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_232_)
  );
  sky130_fd_sc_hd__inv_2 _396_ (
    .A(caravel_rstn),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_000_)
  );
  sky130_fd_sc_hd__inv_2 _397_ (
    .A(user_resetn),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(user_reset)
  );
  sky130_fd_sc_hd__inv_2 _398_ (
    .A(caravel_clk),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_001_)
  );
  sky130_fd_sc_hd__inv_2 _399_ (
    .A(caravel_clk2),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_002_)
  );
  sky130_fd_sc_hd__inv_2 _400_ (
    .A(mprj_cyc_o_core),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_003_)
  );
  sky130_fd_sc_hd__inv_2 _401_ (
    .A(mprj_stb_o_core),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_004_)
  );
  sky130_fd_sc_hd__inv_2 _402_ (
    .A(mprj_we_o_core),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_005_)
  );
  sky130_fd_sc_hd__inv_2 _403_ (
    .A(mprj_sel_o_core[0]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_006_)
  );
  sky130_fd_sc_hd__inv_2 _404_ (
    .A(mprj_sel_o_core[1]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_007_)
  );
  sky130_fd_sc_hd__inv_2 _405_ (
    .A(mprj_sel_o_core[2]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_008_)
  );
  sky130_fd_sc_hd__inv_2 _406_ (
    .A(mprj_sel_o_core[3]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_009_)
  );
  sky130_fd_sc_hd__inv_2 _407_ (
    .A(mprj_adr_o_core[0]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_010_)
  );
  sky130_fd_sc_hd__inv_2 _408_ (
    .A(mprj_adr_o_core[1]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_021_)
  );
  sky130_fd_sc_hd__inv_2 _409_ (
    .A(mprj_adr_o_core[2]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_032_)
  );
  sky130_fd_sc_hd__inv_2 _410_ (
    .A(mprj_adr_o_core[3]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_035_)
  );
  sky130_fd_sc_hd__inv_2 _411_ (
    .A(mprj_adr_o_core[4]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_036_)
  );
  sky130_fd_sc_hd__inv_2 _412_ (
    .A(mprj_adr_o_core[5]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_037_)
  );
  sky130_fd_sc_hd__inv_2 _413_ (
    .A(mprj_adr_o_core[6]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_038_)
  );
  sky130_fd_sc_hd__inv_2 _414_ (
    .A(mprj_adr_o_core[7]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_039_)
  );
  sky130_fd_sc_hd__inv_2 _415_ (
    .A(mprj_adr_o_core[8]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_040_)
  );
  sky130_fd_sc_hd__inv_2 _416_ (
    .A(mprj_adr_o_core[9]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_041_)
  );
  sky130_fd_sc_hd__inv_2 _417_ (
    .A(mprj_adr_o_core[10]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_011_)
  );
  sky130_fd_sc_hd__inv_2 _418_ (
    .A(mprj_adr_o_core[11]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_012_)
  );
  sky130_fd_sc_hd__inv_2 _419_ (
    .A(mprj_adr_o_core[12]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_013_)
  );
  sky130_fd_sc_hd__inv_2 _420_ (
    .A(mprj_adr_o_core[13]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_014_)
  );
  sky130_fd_sc_hd__inv_2 _421_ (
    .A(mprj_adr_o_core[14]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_015_)
  );
  sky130_fd_sc_hd__inv_2 _422_ (
    .A(mprj_adr_o_core[15]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_016_)
  );
  sky130_fd_sc_hd__inv_2 _423_ (
    .A(mprj_adr_o_core[16]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_017_)
  );
  sky130_fd_sc_hd__inv_2 _424_ (
    .A(mprj_adr_o_core[17]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_018_)
  );
  sky130_fd_sc_hd__inv_2 _425_ (
    .A(mprj_adr_o_core[18]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_019_)
  );
  sky130_fd_sc_hd__inv_2 _426_ (
    .A(mprj_adr_o_core[19]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_020_)
  );
  sky130_fd_sc_hd__inv_2 _427_ (
    .A(mprj_adr_o_core[20]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_022_)
  );
  sky130_fd_sc_hd__inv_2 _428_ (
    .A(mprj_adr_o_core[21]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_023_)
  );
  sky130_fd_sc_hd__inv_2 _429_ (
    .A(mprj_adr_o_core[22]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_024_)
  );
  sky130_fd_sc_hd__inv_2 _430_ (
    .A(mprj_adr_o_core[23]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_025_)
  );
  sky130_fd_sc_hd__inv_2 _431_ (
    .A(mprj_adr_o_core[24]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_026_)
  );
  sky130_fd_sc_hd__inv_2 _432_ (
    .A(mprj_adr_o_core[25]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_027_)
  );
  sky130_fd_sc_hd__inv_2 _433_ (
    .A(mprj_adr_o_core[26]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_028_)
  );
  sky130_fd_sc_hd__inv_2 _434_ (
    .A(mprj_adr_o_core[27]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_029_)
  );
  sky130_fd_sc_hd__inv_2 _435_ (
    .A(mprj_adr_o_core[28]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_030_)
  );
  sky130_fd_sc_hd__inv_2 _436_ (
    .A(mprj_adr_o_core[29]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_031_)
  );
  sky130_fd_sc_hd__inv_2 _437_ (
    .A(mprj_adr_o_core[30]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_033_)
  );
  sky130_fd_sc_hd__inv_2 _438_ (
    .A(mprj_adr_o_core[31]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_034_)
  );
  sky130_fd_sc_hd__inv_2 _439_ (
    .A(mprj_dat_o_core[0]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_042_)
  );
  sky130_fd_sc_hd__inv_2 _440_ (
    .A(mprj_dat_o_core[1]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_053_)
  );
  sky130_fd_sc_hd__inv_2 _441_ (
    .A(mprj_dat_o_core[2]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_064_)
  );
  sky130_fd_sc_hd__inv_2 _442_ (
    .A(mprj_dat_o_core[3]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_067_)
  );
  sky130_fd_sc_hd__inv_2 _443_ (
    .A(mprj_dat_o_core[4]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_068_)
  );
  sky130_fd_sc_hd__inv_2 _444_ (
    .A(mprj_dat_o_core[5]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_069_)
  );
  sky130_fd_sc_hd__inv_2 _445_ (
    .A(mprj_dat_o_core[6]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_070_)
  );
  sky130_fd_sc_hd__inv_2 _446_ (
    .A(mprj_dat_o_core[7]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_071_)
  );
  sky130_fd_sc_hd__inv_2 _447_ (
    .A(mprj_dat_o_core[8]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_072_)
  );
  sky130_fd_sc_hd__inv_2 _448_ (
    .A(mprj_dat_o_core[9]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_073_)
  );
  sky130_fd_sc_hd__inv_2 _449_ (
    .A(mprj_dat_o_core[10]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_043_)
  );
  sky130_fd_sc_hd__inv_2 _450_ (
    .A(mprj_dat_o_core[11]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_044_)
  );
  sky130_fd_sc_hd__inv_2 _451_ (
    .A(mprj_dat_o_core[12]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_045_)
  );
  sky130_fd_sc_hd__inv_2 _452_ (
    .A(mprj_dat_o_core[13]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_046_)
  );
  sky130_fd_sc_hd__inv_2 _453_ (
    .A(mprj_dat_o_core[14]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_047_)
  );
  sky130_fd_sc_hd__inv_2 _454_ (
    .A(mprj_dat_o_core[15]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_048_)
  );
  sky130_fd_sc_hd__inv_2 _455_ (
    .A(mprj_dat_o_core[16]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_049_)
  );
  sky130_fd_sc_hd__inv_2 _456_ (
    .A(mprj_dat_o_core[17]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_050_)
  );
  sky130_fd_sc_hd__inv_2 _457_ (
    .A(mprj_dat_o_core[18]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_051_)
  );
  sky130_fd_sc_hd__inv_2 _458_ (
    .A(mprj_dat_o_core[19]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_052_)
  );
  sky130_fd_sc_hd__inv_2 _459_ (
    .A(mprj_dat_o_core[20]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_054_)
  );
  sky130_fd_sc_hd__inv_2 _460_ (
    .A(mprj_dat_o_core[21]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_055_)
  );
  sky130_fd_sc_hd__inv_2 _461_ (
    .A(mprj_dat_o_core[22]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_056_)
  );
  sky130_fd_sc_hd__inv_2 _462_ (
    .A(mprj_dat_o_core[23]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_057_)
  );
  sky130_fd_sc_hd__inv_2 _463_ (
    .A(mprj_dat_o_core[24]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_058_)
  );
  sky130_fd_sc_hd__inv_2 _464_ (
    .A(mprj_dat_o_core[25]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_059_)
  );
  sky130_fd_sc_hd__inv_2 _465_ (
    .A(mprj_dat_o_core[26]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_060_)
  );
  sky130_fd_sc_hd__inv_2 _466_ (
    .A(mprj_dat_o_core[27]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_061_)
  );
  sky130_fd_sc_hd__inv_2 _467_ (
    .A(mprj_dat_o_core[28]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_062_)
  );
  sky130_fd_sc_hd__inv_2 _468_ (
    .A(mprj_dat_o_core[29]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_063_)
  );
  sky130_fd_sc_hd__inv_2 _469_ (
    .A(mprj_dat_o_core[30]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_065_)
  );
  sky130_fd_sc_hd__inv_2 _470_ (
    .A(mprj_dat_o_core[31]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_066_)
  );
  sky130_fd_sc_hd__inv_2 _471_ (
    .A(la_data_out_mprj[0]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_074_)
  );
  sky130_fd_sc_hd__inv_2 _472_ (
    .A(la_data_out_mprj[1]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_113_)
  );
  sky130_fd_sc_hd__inv_2 _473_ (
    .A(la_data_out_mprj[2]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_124_)
  );
  sky130_fd_sc_hd__inv_2 _474_ (
    .A(la_data_out_mprj[3]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_135_)
  );
  sky130_fd_sc_hd__inv_2 _475_ (
    .A(la_data_out_mprj[4]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_146_)
  );
  sky130_fd_sc_hd__inv_2 _476_ (
    .A(la_data_out_mprj[5]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_157_)
  );
  sky130_fd_sc_hd__inv_2 _477_ (
    .A(la_data_out_mprj[6]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_168_)
  );
  sky130_fd_sc_hd__inv_2 _478_ (
    .A(la_data_out_mprj[7]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_179_)
  );
  sky130_fd_sc_hd__inv_2 _479_ (
    .A(la_data_out_mprj[8]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_190_)
  );
  sky130_fd_sc_hd__inv_2 _480_ (
    .A(la_data_out_mprj[9]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_201_)
  );
  sky130_fd_sc_hd__inv_2 _481_ (
    .A(la_data_out_mprj[10]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_085_)
  );
  sky130_fd_sc_hd__inv_2 _482_ (
    .A(la_data_out_mprj[11]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_096_)
  );
  sky130_fd_sc_hd__inv_2 _483_ (
    .A(la_data_out_mprj[12]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_105_)
  );
  sky130_fd_sc_hd__inv_2 _484_ (
    .A(la_data_out_mprj[13]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_106_)
  );
  sky130_fd_sc_hd__inv_2 _485_ (
    .A(la_data_out_mprj[14]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_107_)
  );
  sky130_fd_sc_hd__inv_2 _486_ (
    .A(la_data_out_mprj[15]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_108_)
  );
  sky130_fd_sc_hd__inv_2 _487_ (
    .A(la_data_out_mprj[16]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_109_)
  );
  sky130_fd_sc_hd__inv_2 _488_ (
    .A(la_data_out_mprj[17]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_110_)
  );
  sky130_fd_sc_hd__inv_2 _489_ (
    .A(la_data_out_mprj[18]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_111_)
  );
  sky130_fd_sc_hd__inv_2 _490_ (
    .A(la_data_out_mprj[19]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_112_)
  );
  sky130_fd_sc_hd__inv_2 _491_ (
    .A(la_data_out_mprj[20]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_114_)
  );
  sky130_fd_sc_hd__inv_2 _492_ (
    .A(la_data_out_mprj[21]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_115_)
  );
  sky130_fd_sc_hd__inv_2 _493_ (
    .A(la_data_out_mprj[22]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_116_)
  );
  sky130_fd_sc_hd__inv_2 _494_ (
    .A(la_data_out_mprj[23]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_117_)
  );
  sky130_fd_sc_hd__inv_2 _495_ (
    .A(la_data_out_mprj[24]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_118_)
  );
  sky130_fd_sc_hd__inv_2 _496_ (
    .A(la_data_out_mprj[25]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_119_)
  );
  sky130_fd_sc_hd__inv_2 _497_ (
    .A(la_data_out_mprj[26]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_120_)
  );
  sky130_fd_sc_hd__inv_2 _498_ (
    .A(la_data_out_mprj[27]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_121_)
  );
  sky130_fd_sc_hd__inv_2 _499_ (
    .A(la_data_out_mprj[28]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_122_)
  );
  sky130_fd_sc_hd__inv_2 _500_ (
    .A(la_data_out_mprj[29]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_123_)
  );
  sky130_fd_sc_hd__inv_2 _501_ (
    .A(la_data_out_mprj[30]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_125_)
  );
  sky130_fd_sc_hd__inv_2 _502_ (
    .A(la_data_out_mprj[31]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_126_)
  );
  sky130_fd_sc_hd__inv_2 _503_ (
    .A(la_data_out_mprj[32]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_127_)
  );
  sky130_fd_sc_hd__inv_2 _504_ (
    .A(la_data_out_mprj[33]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_128_)
  );
  sky130_fd_sc_hd__inv_2 _505_ (
    .A(la_data_out_mprj[34]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_129_)
  );
  sky130_fd_sc_hd__inv_2 _506_ (
    .A(la_data_out_mprj[35]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_130_)
  );
  sky130_fd_sc_hd__inv_2 _507_ (
    .A(la_data_out_mprj[36]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_131_)
  );
  sky130_fd_sc_hd__inv_2 _508_ (
    .A(la_data_out_mprj[37]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_132_)
  );
  sky130_fd_sc_hd__inv_2 _509_ (
    .A(la_data_out_mprj[38]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_133_)
  );
  sky130_fd_sc_hd__inv_2 _510_ (
    .A(la_data_out_mprj[39]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_134_)
  );
  sky130_fd_sc_hd__inv_2 _511_ (
    .A(la_data_out_mprj[40]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_136_)
  );
  sky130_fd_sc_hd__inv_2 _512_ (
    .A(la_data_out_mprj[41]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_137_)
  );
  sky130_fd_sc_hd__inv_2 _513_ (
    .A(la_data_out_mprj[42]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_138_)
  );
  sky130_fd_sc_hd__inv_2 _514_ (
    .A(la_data_out_mprj[43]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_139_)
  );
  sky130_fd_sc_hd__inv_2 _515_ (
    .A(la_data_out_mprj[44]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_140_)
  );
  sky130_fd_sc_hd__inv_2 _516_ (
    .A(la_data_out_mprj[45]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_141_)
  );
  sky130_fd_sc_hd__inv_2 _517_ (
    .A(la_data_out_mprj[46]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_142_)
  );
  sky130_fd_sc_hd__inv_2 _518_ (
    .A(la_data_out_mprj[47]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_143_)
  );
  sky130_fd_sc_hd__inv_2 _519_ (
    .A(la_data_out_mprj[48]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_144_)
  );
  sky130_fd_sc_hd__inv_2 _520_ (
    .A(la_data_out_mprj[49]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_145_)
  );
  sky130_fd_sc_hd__inv_2 _521_ (
    .A(la_data_out_mprj[50]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_147_)
  );
  sky130_fd_sc_hd__inv_2 _522_ (
    .A(la_data_out_mprj[51]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_148_)
  );
  sky130_fd_sc_hd__inv_2 _523_ (
    .A(la_data_out_mprj[52]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_149_)
  );
  sky130_fd_sc_hd__inv_2 _524_ (
    .A(la_data_out_mprj[53]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_150_)
  );
  sky130_fd_sc_hd__inv_2 _525_ (
    .A(la_data_out_mprj[54]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_151_)
  );
  sky130_fd_sc_hd__inv_2 _526_ (
    .A(la_data_out_mprj[55]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_152_)
  );
  sky130_fd_sc_hd__inv_2 _527_ (
    .A(la_data_out_mprj[56]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_153_)
  );
  sky130_fd_sc_hd__inv_2 _528_ (
    .A(la_data_out_mprj[57]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_154_)
  );
  sky130_fd_sc_hd__inv_2 _529_ (
    .A(la_data_out_mprj[58]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_155_)
  );
  sky130_fd_sc_hd__inv_2 _530_ (
    .A(la_data_out_mprj[59]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_156_)
  );
  sky130_fd_sc_hd__inv_2 _531_ (
    .A(la_data_out_mprj[60]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_158_)
  );
  sky130_fd_sc_hd__inv_2 _532_ (
    .A(la_data_out_mprj[61]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_159_)
  );
  sky130_fd_sc_hd__inv_2 _533_ (
    .A(la_data_out_mprj[62]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_160_)
  );
  sky130_fd_sc_hd__inv_2 _534_ (
    .A(la_data_out_mprj[63]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_161_)
  );
  sky130_fd_sc_hd__inv_2 _535_ (
    .A(la_data_out_mprj[64]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_162_)
  );
  sky130_fd_sc_hd__inv_2 _536_ (
    .A(la_data_out_mprj[65]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_163_)
  );
  sky130_fd_sc_hd__inv_2 _537_ (
    .A(la_data_out_mprj[66]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_164_)
  );
  sky130_fd_sc_hd__inv_2 _538_ (
    .A(la_data_out_mprj[67]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_165_)
  );
  sky130_fd_sc_hd__inv_2 _539_ (
    .A(la_data_out_mprj[68]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_166_)
  );
  sky130_fd_sc_hd__inv_2 _540_ (
    .A(la_data_out_mprj[69]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_167_)
  );
  sky130_fd_sc_hd__inv_2 _541_ (
    .A(la_data_out_mprj[70]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_169_)
  );
  sky130_fd_sc_hd__inv_2 _542_ (
    .A(la_data_out_mprj[71]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_170_)
  );
  sky130_fd_sc_hd__inv_2 _543_ (
    .A(la_data_out_mprj[72]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_171_)
  );
  sky130_fd_sc_hd__inv_2 _544_ (
    .A(la_data_out_mprj[73]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_172_)
  );
  sky130_fd_sc_hd__inv_2 _545_ (
    .A(la_data_out_mprj[74]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_173_)
  );
  sky130_fd_sc_hd__inv_2 _546_ (
    .A(la_data_out_mprj[75]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_174_)
  );
  sky130_fd_sc_hd__inv_2 _547_ (
    .A(la_data_out_mprj[76]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_175_)
  );
  sky130_fd_sc_hd__inv_2 _548_ (
    .A(la_data_out_mprj[77]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_176_)
  );
  sky130_fd_sc_hd__inv_2 _549_ (
    .A(la_data_out_mprj[78]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_177_)
  );
  sky130_fd_sc_hd__inv_2 _550_ (
    .A(la_data_out_mprj[79]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_178_)
  );
  sky130_fd_sc_hd__inv_2 _551_ (
    .A(la_data_out_mprj[80]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_180_)
  );
  sky130_fd_sc_hd__inv_2 _552_ (
    .A(la_data_out_mprj[81]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_181_)
  );
  sky130_fd_sc_hd__inv_2 _553_ (
    .A(la_data_out_mprj[82]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_182_)
  );
  sky130_fd_sc_hd__inv_2 _554_ (
    .A(la_data_out_mprj[83]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_183_)
  );
  sky130_fd_sc_hd__inv_2 _555_ (
    .A(la_data_out_mprj[84]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_184_)
  );
  sky130_fd_sc_hd__inv_2 _556_ (
    .A(la_data_out_mprj[85]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_185_)
  );
  sky130_fd_sc_hd__inv_2 _557_ (
    .A(la_data_out_mprj[86]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_186_)
  );
  sky130_fd_sc_hd__inv_2 _558_ (
    .A(la_data_out_mprj[87]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_187_)
  );
  sky130_fd_sc_hd__inv_2 _559_ (
    .A(la_data_out_mprj[88]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_188_)
  );
  sky130_fd_sc_hd__inv_2 _560_ (
    .A(la_data_out_mprj[89]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_189_)
  );
  sky130_fd_sc_hd__inv_2 _561_ (
    .A(la_data_out_mprj[90]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_191_)
  );
  sky130_fd_sc_hd__inv_2 _562_ (
    .A(la_data_out_mprj[91]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_192_)
  );
  sky130_fd_sc_hd__inv_2 _563_ (
    .A(la_data_out_mprj[92]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_193_)
  );
  sky130_fd_sc_hd__inv_2 _564_ (
    .A(la_data_out_mprj[93]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_194_)
  );
  sky130_fd_sc_hd__inv_2 _565_ (
    .A(la_data_out_mprj[94]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_195_)
  );
  sky130_fd_sc_hd__inv_2 _566_ (
    .A(la_data_out_mprj[95]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_196_)
  );
  sky130_fd_sc_hd__inv_2 _567_ (
    .A(la_data_out_mprj[96]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_197_)
  );
  sky130_fd_sc_hd__inv_2 _568_ (
    .A(la_data_out_mprj[97]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_198_)
  );
  sky130_fd_sc_hd__inv_2 _569_ (
    .A(la_data_out_mprj[98]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_199_)
  );
  sky130_fd_sc_hd__inv_2 _570_ (
    .A(la_data_out_mprj[99]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_200_)
  );
  sky130_fd_sc_hd__inv_2 _571_ (
    .A(la_data_out_mprj[100]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_075_)
  );
  sky130_fd_sc_hd__inv_2 _572_ (
    .A(la_data_out_mprj[101]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_076_)
  );
  sky130_fd_sc_hd__inv_2 _573_ (
    .A(la_data_out_mprj[102]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_077_)
  );
  sky130_fd_sc_hd__inv_2 _574_ (
    .A(la_data_out_mprj[103]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_078_)
  );
  sky130_fd_sc_hd__inv_2 _575_ (
    .A(la_data_out_mprj[104]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_079_)
  );
  sky130_fd_sc_hd__inv_2 _576_ (
    .A(la_data_out_mprj[105]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_080_)
  );
  sky130_fd_sc_hd__inv_2 _577_ (
    .A(la_data_out_mprj[106]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_081_)
  );
  sky130_fd_sc_hd__inv_2 _578_ (
    .A(la_data_out_mprj[107]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_082_)
  );
  sky130_fd_sc_hd__inv_2 _579_ (
    .A(la_data_out_mprj[108]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_083_)
  );
  sky130_fd_sc_hd__inv_2 _580_ (
    .A(la_data_out_mprj[109]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_084_)
  );
  sky130_fd_sc_hd__inv_2 _581_ (
    .A(la_data_out_mprj[110]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_086_)
  );
  sky130_fd_sc_hd__inv_2 _582_ (
    .A(la_data_out_mprj[111]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_087_)
  );
  sky130_fd_sc_hd__inv_2 _583_ (
    .A(la_data_out_mprj[112]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_088_)
  );
  sky130_fd_sc_hd__inv_2 _584_ (
    .A(la_data_out_mprj[113]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_089_)
  );
  sky130_fd_sc_hd__inv_2 _585_ (
    .A(la_data_out_mprj[114]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_090_)
  );
  sky130_fd_sc_hd__inv_2 _586_ (
    .A(la_data_out_mprj[115]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_091_)
  );
  sky130_fd_sc_hd__inv_2 _587_ (
    .A(la_data_out_mprj[116]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_092_)
  );
  sky130_fd_sc_hd__inv_2 _588_ (
    .A(la_data_out_mprj[117]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_093_)
  );
  sky130_fd_sc_hd__inv_2 _589_ (
    .A(la_data_out_mprj[118]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_094_)
  );
  sky130_fd_sc_hd__inv_2 _590_ (
    .A(la_data_out_mprj[119]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_095_)
  );
  sky130_fd_sc_hd__inv_2 _591_ (
    .A(la_data_out_mprj[120]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_097_)
  );
  sky130_fd_sc_hd__inv_2 _592_ (
    .A(la_data_out_mprj[121]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_098_)
  );
  sky130_fd_sc_hd__inv_2 _593_ (
    .A(la_data_out_mprj[122]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_099_)
  );
  sky130_fd_sc_hd__inv_2 _594_ (
    .A(la_data_out_mprj[123]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_100_)
  );
  sky130_fd_sc_hd__inv_2 _595_ (
    .A(la_data_out_mprj[124]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_101_)
  );
  sky130_fd_sc_hd__inv_2 _596_ (
    .A(la_data_out_mprj[125]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_102_)
  );
  sky130_fd_sc_hd__inv_2 _597_ (
    .A(la_data_out_mprj[126]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_103_)
  );
  sky130_fd_sc_hd__inv_2 _598_ (
    .A(la_data_out_mprj[127]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_104_)
  );
  sky130_fd_sc_hd__inv_2 _599_ (
    .A(la_oen_mprj[0]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_202_)
  );
  sky130_fd_sc_hd__inv_2 _600_ (
    .A(la_oen_mprj[1]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_241_)
  );
  sky130_fd_sc_hd__inv_2 _601_ (
    .A(la_oen_mprj[2]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_252_)
  );
  sky130_fd_sc_hd__inv_2 _602_ (
    .A(la_oen_mprj[3]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_263_)
  );
  sky130_fd_sc_hd__inv_2 _603_ (
    .A(la_oen_mprj[4]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_274_)
  );
  sky130_fd_sc_hd__inv_2 _604_ (
    .A(la_oen_mprj[5]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_285_)
  );
  sky130_fd_sc_hd__inv_2 _605_ (
    .A(la_oen_mprj[6]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_296_)
  );
  sky130_fd_sc_hd__inv_2 _606_ (
    .A(la_oen_mprj[7]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_307_)
  );
  sky130_fd_sc_hd__inv_2 _607_ (
    .A(la_oen_mprj[8]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_318_)
  );
  sky130_fd_sc_hd__inv_2 _608_ (
    .A(la_oen_mprj[9]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_329_)
  );
  sky130_fd_sc_hd__inv_2 _609_ (
    .A(la_oen_mprj[10]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_213_)
  );
  sky130_fd_sc_hd__inv_2 _610_ (
    .A(la_oen_mprj[11]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_224_)
  );
  sky130_fd_sc_hd__inv_2 _611_ (
    .A(la_oen_mprj[12]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_233_)
  );
  sky130_fd_sc_hd__inv_2 _612_ (
    .A(la_oen_mprj[13]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_234_)
  );
  sky130_fd_sc_hd__inv_2 _613_ (
    .A(la_oen_mprj[14]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_235_)
  );
  sky130_fd_sc_hd__inv_2 _614_ (
    .A(la_oen_mprj[15]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_236_)
  );
  sky130_fd_sc_hd__inv_2 _615_ (
    .A(la_oen_mprj[16]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_237_)
  );
  sky130_fd_sc_hd__inv_2 _616_ (
    .A(la_oen_mprj[17]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_238_)
  );
  sky130_fd_sc_hd__inv_2 _617_ (
    .A(la_oen_mprj[18]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_239_)
  );
  sky130_fd_sc_hd__inv_2 _618_ (
    .A(la_oen_mprj[19]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_240_)
  );
  sky130_fd_sc_hd__inv_2 _619_ (
    .A(la_oen_mprj[20]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_242_)
  );
  sky130_fd_sc_hd__inv_2 _620_ (
    .A(la_oen_mprj[21]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_243_)
  );
  sky130_fd_sc_hd__inv_2 _621_ (
    .A(la_oen_mprj[22]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_244_)
  );
  sky130_fd_sc_hd__inv_2 _622_ (
    .A(la_oen_mprj[23]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_245_)
  );
  sky130_fd_sc_hd__inv_2 _623_ (
    .A(la_oen_mprj[24]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_246_)
  );
  sky130_fd_sc_hd__inv_2 _624_ (
    .A(la_oen_mprj[25]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_247_)
  );
  sky130_fd_sc_hd__inv_2 _625_ (
    .A(la_oen_mprj[26]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_248_)
  );
  sky130_fd_sc_hd__inv_2 _626_ (
    .A(la_oen_mprj[27]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_249_)
  );
  sky130_fd_sc_hd__inv_2 _627_ (
    .A(la_oen_mprj[28]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_250_)
  );
  sky130_fd_sc_hd__inv_2 _628_ (
    .A(la_oen_mprj[29]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_251_)
  );
  sky130_fd_sc_hd__inv_2 _629_ (
    .A(la_oen_mprj[30]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_253_)
  );
  sky130_fd_sc_hd__inv_2 _630_ (
    .A(la_oen_mprj[31]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_254_)
  );
  sky130_fd_sc_hd__inv_2 _631_ (
    .A(la_oen_mprj[32]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_255_)
  );
  sky130_fd_sc_hd__inv_2 _632_ (
    .A(la_oen_mprj[33]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_256_)
  );
  sky130_fd_sc_hd__inv_2 _633_ (
    .A(la_oen_mprj[34]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_257_)
  );
  sky130_fd_sc_hd__inv_2 _634_ (
    .A(la_oen_mprj[35]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_258_)
  );
  sky130_fd_sc_hd__inv_2 _635_ (
    .A(la_oen_mprj[36]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_259_)
  );
  sky130_fd_sc_hd__inv_2 _636_ (
    .A(la_oen_mprj[37]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_260_)
  );
  sky130_fd_sc_hd__inv_2 _637_ (
    .A(la_oen_mprj[38]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_261_)
  );
  sky130_fd_sc_hd__inv_2 _638_ (
    .A(la_oen_mprj[39]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_262_)
  );
  sky130_fd_sc_hd__inv_2 _639_ (
    .A(la_oen_mprj[40]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_264_)
  );
  sky130_fd_sc_hd__inv_2 _640_ (
    .A(la_oen_mprj[41]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_265_)
  );
  sky130_fd_sc_hd__inv_2 _641_ (
    .A(la_oen_mprj[42]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_266_)
  );
  sky130_fd_sc_hd__inv_2 _642_ (
    .A(la_oen_mprj[43]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_267_)
  );
  sky130_fd_sc_hd__inv_2 _643_ (
    .A(la_oen_mprj[44]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_268_)
  );
  sky130_fd_sc_hd__inv_2 _644_ (
    .A(la_oen_mprj[45]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_269_)
  );
  sky130_fd_sc_hd__inv_2 _645_ (
    .A(la_oen_mprj[46]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_270_)
  );
  sky130_fd_sc_hd__inv_2 _646_ (
    .A(la_oen_mprj[47]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_271_)
  );
  sky130_fd_sc_hd__inv_2 _647_ (
    .A(la_oen_mprj[48]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_272_)
  );
  sky130_fd_sc_hd__inv_2 _648_ (
    .A(la_oen_mprj[49]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_273_)
  );
  sky130_fd_sc_hd__inv_2 _649_ (
    .A(la_oen_mprj[50]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_275_)
  );
  sky130_fd_sc_hd__inv_2 _650_ (
    .A(la_oen_mprj[51]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_276_)
  );
  sky130_fd_sc_hd__inv_2 _651_ (
    .A(la_oen_mprj[52]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_277_)
  );
  sky130_fd_sc_hd__inv_2 _652_ (
    .A(la_oen_mprj[53]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_278_)
  );
  sky130_fd_sc_hd__inv_2 _653_ (
    .A(la_oen_mprj[54]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_279_)
  );
  sky130_fd_sc_hd__inv_2 _654_ (
    .A(la_oen_mprj[55]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_280_)
  );
  sky130_fd_sc_hd__inv_2 _655_ (
    .A(la_oen_mprj[56]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_281_)
  );
  sky130_fd_sc_hd__inv_2 _656_ (
    .A(la_oen_mprj[57]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_282_)
  );
  sky130_fd_sc_hd__inv_2 _657_ (
    .A(la_oen_mprj[58]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_283_)
  );
  sky130_fd_sc_hd__inv_2 _658_ (
    .A(la_oen_mprj[59]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_284_)
  );
  sky130_fd_sc_hd__inv_2 _659_ (
    .A(la_oen_mprj[60]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_286_)
  );
  sky130_fd_sc_hd__inv_2 _660_ (
    .A(la_oen_mprj[61]),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(_287_)
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[0]  (
    .A(_074_),
    .TE(\mprj_logic1[74] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[0])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[100]  (
    .A(_075_),
    .TE(\mprj_logic1[174] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[100])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[101]  (
    .A(_076_),
    .TE(\mprj_logic1[175] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[101])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[102]  (
    .A(_077_),
    .TE(\mprj_logic1[176] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[102])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[103]  (
    .A(_078_),
    .TE(\mprj_logic1[177] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[103])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[104]  (
    .A(_079_),
    .TE(\mprj_logic1[178] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[104])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[105]  (
    .A(_080_),
    .TE(\mprj_logic1[179] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[105])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[106]  (
    .A(_081_),
    .TE(\mprj_logic1[180] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[106])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[107]  (
    .A(_082_),
    .TE(\mprj_logic1[181] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[107])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[108]  (
    .A(_083_),
    .TE(\mprj_logic1[182] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[108])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[109]  (
    .A(_084_),
    .TE(\mprj_logic1[183] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[109])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[10]  (
    .A(_085_),
    .TE(\mprj_logic1[84] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[10])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[110]  (
    .A(_086_),
    .TE(\mprj_logic1[184] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[110])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[111]  (
    .A(_087_),
    .TE(\mprj_logic1[185] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[111])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[112]  (
    .A(_088_),
    .TE(\mprj_logic1[186] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[112])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[113]  (
    .A(_089_),
    .TE(\mprj_logic1[187] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[113])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[114]  (
    .A(_090_),
    .TE(\mprj_logic1[188] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[114])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[115]  (
    .A(_091_),
    .TE(\mprj_logic1[189] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[115])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[116]  (
    .A(_092_),
    .TE(\mprj_logic1[190] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[116])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[117]  (
    .A(_093_),
    .TE(\mprj_logic1[191] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[117])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[118]  (
    .A(_094_),
    .TE(\mprj_logic1[192] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[118])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[119]  (
    .A(_095_),
    .TE(\mprj_logic1[193] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[119])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[11]  (
    .A(_096_),
    .TE(\mprj_logic1[85] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[11])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[120]  (
    .A(_097_),
    .TE(\mprj_logic1[194] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[120])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[121]  (
    .A(_098_),
    .TE(\mprj_logic1[195] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[121])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[122]  (
    .A(_099_),
    .TE(\mprj_logic1[196] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[122])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[123]  (
    .A(_100_),
    .TE(\mprj_logic1[197] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[123])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[124]  (
    .A(_101_),
    .TE(\mprj_logic1[198] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[124])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[125]  (
    .A(_102_),
    .TE(\mprj_logic1[199] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[125])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[126]  (
    .A(_103_),
    .TE(\mprj_logic1[200] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[126])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[127]  (
    .A(_104_),
    .TE(\mprj_logic1[201] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[127])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[12]  (
    .A(_105_),
    .TE(\mprj_logic1[86] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[12])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[13]  (
    .A(_106_),
    .TE(\mprj_logic1[87] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[13])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[14]  (
    .A(_107_),
    .TE(\mprj_logic1[88] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[14])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[15]  (
    .A(_108_),
    .TE(\mprj_logic1[89] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[15])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[16]  (
    .A(_109_),
    .TE(\mprj_logic1[90] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[16])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[17]  (
    .A(_110_),
    .TE(\mprj_logic1[91] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[17])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[18]  (
    .A(_111_),
    .TE(\mprj_logic1[92] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[18])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[19]  (
    .A(_112_),
    .TE(\mprj_logic1[93] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[19])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[1]  (
    .A(_113_),
    .TE(\mprj_logic1[75] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[1])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[20]  (
    .A(_114_),
    .TE(\mprj_logic1[94] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[20])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[21]  (
    .A(_115_),
    .TE(\mprj_logic1[95] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[21])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[22]  (
    .A(_116_),
    .TE(\mprj_logic1[96] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[22])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[23]  (
    .A(_117_),
    .TE(\mprj_logic1[97] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[23])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[24]  (
    .A(_118_),
    .TE(\mprj_logic1[98] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[24])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[25]  (
    .A(_119_),
    .TE(\mprj_logic1[99] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[25])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[26]  (
    .A(_120_),
    .TE(\mprj_logic1[100] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[26])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[27]  (
    .A(_121_),
    .TE(\mprj_logic1[101] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[27])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[28]  (
    .A(_122_),
    .TE(\mprj_logic1[102] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[28])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[29]  (
    .A(_123_),
    .TE(\mprj_logic1[103] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[29])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[2]  (
    .A(_124_),
    .TE(\mprj_logic1[76] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[2])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[30]  (
    .A(_125_),
    .TE(\mprj_logic1[104] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[30])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[31]  (
    .A(_126_),
    .TE(\mprj_logic1[105] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[31])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[32]  (
    .A(_127_),
    .TE(\mprj_logic1[106] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[32])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[33]  (
    .A(_128_),
    .TE(\mprj_logic1[107] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[33])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[34]  (
    .A(_129_),
    .TE(\mprj_logic1[108] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[34])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[35]  (
    .A(_130_),
    .TE(\mprj_logic1[109] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[35])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[36]  (
    .A(_131_),
    .TE(\mprj_logic1[110] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[36])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[37]  (
    .A(_132_),
    .TE(\mprj_logic1[111] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[37])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[38]  (
    .A(_133_),
    .TE(\mprj_logic1[112] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[38])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[39]  (
    .A(_134_),
    .TE(\mprj_logic1[113] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[39])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[3]  (
    .A(_135_),
    .TE(\mprj_logic1[77] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[3])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[40]  (
    .A(_136_),
    .TE(\mprj_logic1[114] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[40])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[41]  (
    .A(_137_),
    .TE(\mprj_logic1[115] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[41])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[42]  (
    .A(_138_),
    .TE(\mprj_logic1[116] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[42])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[43]  (
    .A(_139_),
    .TE(\mprj_logic1[117] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[43])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[44]  (
    .A(_140_),
    .TE(\mprj_logic1[118] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[44])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[45]  (
    .A(_141_),
    .TE(\mprj_logic1[119] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[45])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[46]  (
    .A(_142_),
    .TE(\mprj_logic1[120] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[46])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[47]  (
    .A(_143_),
    .TE(\mprj_logic1[121] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[47])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[48]  (
    .A(_144_),
    .TE(\mprj_logic1[122] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[48])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[49]  (
    .A(_145_),
    .TE(\mprj_logic1[123] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[49])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[4]  (
    .A(_146_),
    .TE(\mprj_logic1[78] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[4])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[50]  (
    .A(_147_),
    .TE(\mprj_logic1[124] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[50])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[51]  (
    .A(_148_),
    .TE(\mprj_logic1[125] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[51])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[52]  (
    .A(_149_),
    .TE(\mprj_logic1[126] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[52])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[53]  (
    .A(_150_),
    .TE(\mprj_logic1[127] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[53])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[54]  (
    .A(_151_),
    .TE(\mprj_logic1[128] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[54])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[55]  (
    .A(_152_),
    .TE(\mprj_logic1[129] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[55])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[56]  (
    .A(_153_),
    .TE(\mprj_logic1[130] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[56])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[57]  (
    .A(_154_),
    .TE(\mprj_logic1[131] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[57])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[58]  (
    .A(_155_),
    .TE(\mprj_logic1[132] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[58])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[59]  (
    .A(_156_),
    .TE(\mprj_logic1[133] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[59])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[5]  (
    .A(_157_),
    .TE(\mprj_logic1[79] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[5])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[60]  (
    .A(_158_),
    .TE(\mprj_logic1[134] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[60])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[61]  (
    .A(_159_),
    .TE(\mprj_logic1[135] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[61])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[62]  (
    .A(_160_),
    .TE(\mprj_logic1[136] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[62])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[63]  (
    .A(_161_),
    .TE(\mprj_logic1[137] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[63])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[64]  (
    .A(_162_),
    .TE(\mprj_logic1[138] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[64])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[65]  (
    .A(_163_),
    .TE(\mprj_logic1[139] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[65])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[66]  (
    .A(_164_),
    .TE(\mprj_logic1[140] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[66])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[67]  (
    .A(_165_),
    .TE(\mprj_logic1[141] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[67])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[68]  (
    .A(_166_),
    .TE(\mprj_logic1[142] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[68])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[69]  (
    .A(_167_),
    .TE(\mprj_logic1[143] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[69])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[6]  (
    .A(_168_),
    .TE(\mprj_logic1[80] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[6])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[70]  (
    .A(_169_),
    .TE(\mprj_logic1[144] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[70])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[71]  (
    .A(_170_),
    .TE(\mprj_logic1[145] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[71])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[72]  (
    .A(_171_),
    .TE(\mprj_logic1[146] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[72])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[73]  (
    .A(_172_),
    .TE(\mprj_logic1[147] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[73])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[74]  (
    .A(_173_),
    .TE(\mprj_logic1[148] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[74])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[75]  (
    .A(_174_),
    .TE(\mprj_logic1[149] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[75])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[76]  (
    .A(_175_),
    .TE(\mprj_logic1[150] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[76])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[77]  (
    .A(_176_),
    .TE(\mprj_logic1[151] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[77])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[78]  (
    .A(_177_),
    .TE(\mprj_logic1[152] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[78])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[79]  (
    .A(_178_),
    .TE(\mprj_logic1[153] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[79])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[7]  (
    .A(_179_),
    .TE(\mprj_logic1[81] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[7])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[80]  (
    .A(_180_),
    .TE(\mprj_logic1[154] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[80])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[81]  (
    .A(_181_),
    .TE(\mprj_logic1[155] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[81])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[82]  (
    .A(_182_),
    .TE(\mprj_logic1[156] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[82])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[83]  (
    .A(_183_),
    .TE(\mprj_logic1[157] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[83])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[84]  (
    .A(_184_),
    .TE(\mprj_logic1[158] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[84])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[85]  (
    .A(_185_),
    .TE(\mprj_logic1[159] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[85])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[86]  (
    .A(_186_),
    .TE(\mprj_logic1[160] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[86])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[87]  (
    .A(_187_),
    .TE(\mprj_logic1[161] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[87])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[88]  (
    .A(_188_),
    .TE(\mprj_logic1[162] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[88])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[89]  (
    .A(_189_),
    .TE(\mprj_logic1[163] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[89])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[8]  (
    .A(_190_),
    .TE(\mprj_logic1[82] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[8])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[90]  (
    .A(_191_),
    .TE(\mprj_logic1[164] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[90])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[91]  (
    .A(_192_),
    .TE(\mprj_logic1[165] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[91])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[92]  (
    .A(_193_),
    .TE(\mprj_logic1[166] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[92])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[93]  (
    .A(_194_),
    .TE(\mprj_logic1[167] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[93])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[94]  (
    .A(_195_),
    .TE(\mprj_logic1[168] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[94])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[95]  (
    .A(_196_),
    .TE(\mprj_logic1[169] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[95])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[96]  (
    .A(_197_),
    .TE(\mprj_logic1[170] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[96])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[97]  (
    .A(_198_),
    .TE(\mprj_logic1[171] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[97])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[98]  (
    .A(_199_),
    .TE(\mprj_logic1[172] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[98])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[99]  (
    .A(_200_),
    .TE(\mprj_logic1[173] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[99])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[9]  (
    .A(_201_),
    .TE(\mprj_logic1[83] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_data_in_core[9])
  );
  sky130_fd_sc_hd__buf_8 mprj2_pwrgood (
    .A(mprj2_vdd_logic1),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .X(user2_vcc_powergood)
  );
  sky130_fd_sc_hd__buf_8 mprj2_vdd_pwrgood (
    .A(mprj2_vdd_logic1),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .X(user2_vdd_powergood)
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[0]  (
    .A(_010_),
    .TE(\mprj_logic1[10] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[0])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[10]  (
    .A(_011_),
    .TE(\mprj_logic1[20] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[10])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[11]  (
    .A(_012_),
    .TE(\mprj_logic1[21] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[11])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[12]  (
    .A(_013_),
    .TE(\mprj_logic1[22] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[12])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[13]  (
    .A(_014_),
    .TE(\mprj_logic1[23] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[13])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[14]  (
    .A(_015_),
    .TE(\mprj_logic1[24] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[14])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[15]  (
    .A(_016_),
    .TE(\mprj_logic1[25] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[15])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[16]  (
    .A(_017_),
    .TE(\mprj_logic1[26] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[16])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[17]  (
    .A(_018_),
    .TE(\mprj_logic1[27] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[17])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[18]  (
    .A(_019_),
    .TE(\mprj_logic1[28] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[18])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[19]  (
    .A(_020_),
    .TE(\mprj_logic1[29] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[19])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[1]  (
    .A(_021_),
    .TE(\mprj_logic1[11] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[1])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[20]  (
    .A(_022_),
    .TE(\mprj_logic1[30] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[20])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[21]  (
    .A(_023_),
    .TE(\mprj_logic1[31] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[21])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[22]  (
    .A(_024_),
    .TE(\mprj_logic1[32] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[22])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[23]  (
    .A(_025_),
    .TE(\mprj_logic1[33] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[23])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[24]  (
    .A(_026_),
    .TE(\mprj_logic1[34] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[24])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[25]  (
    .A(_027_),
    .TE(\mprj_logic1[35] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[25])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[26]  (
    .A(_028_),
    .TE(\mprj_logic1[36] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[26])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[27]  (
    .A(_029_),
    .TE(\mprj_logic1[37] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[27])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[28]  (
    .A(_030_),
    .TE(\mprj_logic1[38] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[28])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[29]  (
    .A(_031_),
    .TE(\mprj_logic1[39] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[29])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[2]  (
    .A(_032_),
    .TE(\mprj_logic1[12] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[2])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[30]  (
    .A(_033_),
    .TE(\mprj_logic1[40] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[30])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[31]  (
    .A(_034_),
    .TE(\mprj_logic1[41] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[31])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[3]  (
    .A(_035_),
    .TE(\mprj_logic1[13] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[3])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[4]  (
    .A(_036_),
    .TE(\mprj_logic1[14] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[4])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[5]  (
    .A(_037_),
    .TE(\mprj_logic1[15] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[5])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[6]  (
    .A(_038_),
    .TE(\mprj_logic1[16] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[6])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[7]  (
    .A(_039_),
    .TE(\mprj_logic1[17] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[7])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[8]  (
    .A(_040_),
    .TE(\mprj_logic1[18] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[8])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[9]  (
    .A(_041_),
    .TE(\mprj_logic1[19] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_adr_o_user[9])
  );
  sky130_fd_sc_hd__einvp_8 mprj_clk2_buf (
    .A(_002_),
    .TE(\mprj_logic1[2] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(user_clock2)
  );
  sky130_fd_sc_hd__einvp_8 mprj_clk_buf (
    .A(_001_),
    .TE(\mprj_logic1[1] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(user_clock)
  );
  sky130_fd_sc_hd__einvp_8 mprj_cyc_buf (
    .A(_003_),
    .TE(\mprj_logic1[3] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_cyc_o_user)
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[0]  (
    .A(_042_),
    .TE(\mprj_logic1[42] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[0])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[10]  (
    .A(_043_),
    .TE(\mprj_logic1[52] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[10])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[11]  (
    .A(_044_),
    .TE(\mprj_logic1[53] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[11])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[12]  (
    .A(_045_),
    .TE(\mprj_logic1[54] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[12])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[13]  (
    .A(_046_),
    .TE(\mprj_logic1[55] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[13])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[14]  (
    .A(_047_),
    .TE(\mprj_logic1[56] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[14])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[15]  (
    .A(_048_),
    .TE(\mprj_logic1[57] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[15])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[16]  (
    .A(_049_),
    .TE(\mprj_logic1[58] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[16])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[17]  (
    .A(_050_),
    .TE(\mprj_logic1[59] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[17])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[18]  (
    .A(_051_),
    .TE(\mprj_logic1[60] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[18])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[19]  (
    .A(_052_),
    .TE(\mprj_logic1[61] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[19])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[1]  (
    .A(_053_),
    .TE(\mprj_logic1[43] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[1])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[20]  (
    .A(_054_),
    .TE(\mprj_logic1[62] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[20])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[21]  (
    .A(_055_),
    .TE(\mprj_logic1[63] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[21])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[22]  (
    .A(_056_),
    .TE(\mprj_logic1[64] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[22])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[23]  (
    .A(_057_),
    .TE(\mprj_logic1[65] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[23])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[24]  (
    .A(_058_),
    .TE(\mprj_logic1[66] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[24])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[25]  (
    .A(_059_),
    .TE(\mprj_logic1[67] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[25])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[26]  (
    .A(_060_),
    .TE(\mprj_logic1[68] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[26])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[27]  (
    .A(_061_),
    .TE(\mprj_logic1[69] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[27])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[28]  (
    .A(_062_),
    .TE(\mprj_logic1[70] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[28])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[29]  (
    .A(_063_),
    .TE(\mprj_logic1[71] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[29])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[2]  (
    .A(_064_),
    .TE(\mprj_logic1[44] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[2])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[30]  (
    .A(_065_),
    .TE(\mprj_logic1[72] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[30])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[31]  (
    .A(_066_),
    .TE(\mprj_logic1[73] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[31])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[3]  (
    .A(_067_),
    .TE(\mprj_logic1[45] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[3])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[4]  (
    .A(_068_),
    .TE(\mprj_logic1[46] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[4])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[5]  (
    .A(_069_),
    .TE(\mprj_logic1[47] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[5])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[6]  (
    .A(_070_),
    .TE(\mprj_logic1[48] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[6])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[7]  (
    .A(_071_),
    .TE(\mprj_logic1[49] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[7])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[8]  (
    .A(_072_),
    .TE(\mprj_logic1[50] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[8])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[9]  (
    .A(_073_),
    .TE(\mprj_logic1[51] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_dat_o_user[9])
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[0]  (
    .HI(\mprj_logic1[0] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[100]  (
    .HI(\mprj_logic1[100] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[101]  (
    .HI(\mprj_logic1[101] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[102]  (
    .HI(\mprj_logic1[102] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[103]  (
    .HI(\mprj_logic1[103] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[104]  (
    .HI(\mprj_logic1[104] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[105]  (
    .HI(\mprj_logic1[105] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[106]  (
    .HI(\mprj_logic1[106] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[107]  (
    .HI(\mprj_logic1[107] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[108]  (
    .HI(\mprj_logic1[108] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[109]  (
    .HI(\mprj_logic1[109] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[10]  (
    .HI(\mprj_logic1[10] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[110]  (
    .HI(\mprj_logic1[110] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[111]  (
    .HI(\mprj_logic1[111] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[112]  (
    .HI(\mprj_logic1[112] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[113]  (
    .HI(\mprj_logic1[113] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[114]  (
    .HI(\mprj_logic1[114] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[115]  (
    .HI(\mprj_logic1[115] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[116]  (
    .HI(\mprj_logic1[116] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[117]  (
    .HI(\mprj_logic1[117] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[118]  (
    .HI(\mprj_logic1[118] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[119]  (
    .HI(\mprj_logic1[119] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[11]  (
    .HI(\mprj_logic1[11] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[120]  (
    .HI(\mprj_logic1[120] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[121]  (
    .HI(\mprj_logic1[121] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[122]  (
    .HI(\mprj_logic1[122] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[123]  (
    .HI(\mprj_logic1[123] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[124]  (
    .HI(\mprj_logic1[124] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[125]  (
    .HI(\mprj_logic1[125] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[126]  (
    .HI(\mprj_logic1[126] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[127]  (
    .HI(\mprj_logic1[127] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[128]  (
    .HI(\mprj_logic1[128] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[129]  (
    .HI(\mprj_logic1[129] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[12]  (
    .HI(\mprj_logic1[12] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[130]  (
    .HI(\mprj_logic1[130] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[131]  (
    .HI(\mprj_logic1[131] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[132]  (
    .HI(\mprj_logic1[132] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[133]  (
    .HI(\mprj_logic1[133] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[134]  (
    .HI(\mprj_logic1[134] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[135]  (
    .HI(\mprj_logic1[135] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[136]  (
    .HI(\mprj_logic1[136] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[137]  (
    .HI(\mprj_logic1[137] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[138]  (
    .HI(\mprj_logic1[138] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[139]  (
    .HI(\mprj_logic1[139] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[13]  (
    .HI(\mprj_logic1[13] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[140]  (
    .HI(\mprj_logic1[140] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[141]  (
    .HI(\mprj_logic1[141] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[142]  (
    .HI(\mprj_logic1[142] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[143]  (
    .HI(\mprj_logic1[143] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[144]  (
    .HI(\mprj_logic1[144] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[145]  (
    .HI(\mprj_logic1[145] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[146]  (
    .HI(\mprj_logic1[146] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[147]  (
    .HI(\mprj_logic1[147] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[148]  (
    .HI(\mprj_logic1[148] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[149]  (
    .HI(\mprj_logic1[149] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[14]  (
    .HI(\mprj_logic1[14] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[150]  (
    .HI(\mprj_logic1[150] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[151]  (
    .HI(\mprj_logic1[151] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[152]  (
    .HI(\mprj_logic1[152] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[153]  (
    .HI(\mprj_logic1[153] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[154]  (
    .HI(\mprj_logic1[154] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[155]  (
    .HI(\mprj_logic1[155] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[156]  (
    .HI(\mprj_logic1[156] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[157]  (
    .HI(\mprj_logic1[157] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[158]  (
    .HI(\mprj_logic1[158] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[159]  (
    .HI(\mprj_logic1[159] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[15]  (
    .HI(\mprj_logic1[15] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[160]  (
    .HI(\mprj_logic1[160] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[161]  (
    .HI(\mprj_logic1[161] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[162]  (
    .HI(\mprj_logic1[162] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[163]  (
    .HI(\mprj_logic1[163] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[164]  (
    .HI(\mprj_logic1[164] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[165]  (
    .HI(\mprj_logic1[165] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[166]  (
    .HI(\mprj_logic1[166] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[167]  (
    .HI(\mprj_logic1[167] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[168]  (
    .HI(\mprj_logic1[168] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[169]  (
    .HI(\mprj_logic1[169] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[16]  (
    .HI(\mprj_logic1[16] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[170]  (
    .HI(\mprj_logic1[170] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[171]  (
    .HI(\mprj_logic1[171] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[172]  (
    .HI(\mprj_logic1[172] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[173]  (
    .HI(\mprj_logic1[173] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[174]  (
    .HI(\mprj_logic1[174] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[175]  (
    .HI(\mprj_logic1[175] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[176]  (
    .HI(\mprj_logic1[176] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[177]  (
    .HI(\mprj_logic1[177] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[178]  (
    .HI(\mprj_logic1[178] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[179]  (
    .HI(\mprj_logic1[179] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[17]  (
    .HI(\mprj_logic1[17] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[180]  (
    .HI(\mprj_logic1[180] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[181]  (
    .HI(\mprj_logic1[181] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[182]  (
    .HI(\mprj_logic1[182] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[183]  (
    .HI(\mprj_logic1[183] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[184]  (
    .HI(\mprj_logic1[184] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[185]  (
    .HI(\mprj_logic1[185] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[186]  (
    .HI(\mprj_logic1[186] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[187]  (
    .HI(\mprj_logic1[187] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[188]  (
    .HI(\mprj_logic1[188] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[189]  (
    .HI(\mprj_logic1[189] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[18]  (
    .HI(\mprj_logic1[18] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[190]  (
    .HI(\mprj_logic1[190] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[191]  (
    .HI(\mprj_logic1[191] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[192]  (
    .HI(\mprj_logic1[192] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[193]  (
    .HI(\mprj_logic1[193] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[194]  (
    .HI(\mprj_logic1[194] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[195]  (
    .HI(\mprj_logic1[195] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[196]  (
    .HI(\mprj_logic1[196] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[197]  (
    .HI(\mprj_logic1[197] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[198]  (
    .HI(\mprj_logic1[198] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[199]  (
    .HI(\mprj_logic1[199] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[19]  (
    .HI(\mprj_logic1[19] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[1]  (
    .HI(\mprj_logic1[1] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[200]  (
    .HI(\mprj_logic1[200] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[201]  (
    .HI(\mprj_logic1[201] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[202]  (
    .HI(\mprj_logic1[202] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[203]  (
    .HI(\mprj_logic1[203] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[204]  (
    .HI(\mprj_logic1[204] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[205]  (
    .HI(\mprj_logic1[205] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[206]  (
    .HI(\mprj_logic1[206] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[207]  (
    .HI(\mprj_logic1[207] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[208]  (
    .HI(\mprj_logic1[208] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[209]  (
    .HI(\mprj_logic1[209] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[20]  (
    .HI(\mprj_logic1[20] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[210]  (
    .HI(\mprj_logic1[210] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[211]  (
    .HI(\mprj_logic1[211] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[212]  (
    .HI(\mprj_logic1[212] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[213]  (
    .HI(\mprj_logic1[213] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[214]  (
    .HI(\mprj_logic1[214] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[215]  (
    .HI(\mprj_logic1[215] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[216]  (
    .HI(\mprj_logic1[216] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[217]  (
    .HI(\mprj_logic1[217] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[218]  (
    .HI(\mprj_logic1[218] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[219]  (
    .HI(\mprj_logic1[219] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[21]  (
    .HI(\mprj_logic1[21] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[220]  (
    .HI(\mprj_logic1[220] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[221]  (
    .HI(\mprj_logic1[221] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[222]  (
    .HI(\mprj_logic1[222] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[223]  (
    .HI(\mprj_logic1[223] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[224]  (
    .HI(\mprj_logic1[224] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[225]  (
    .HI(\mprj_logic1[225] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[226]  (
    .HI(\mprj_logic1[226] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[227]  (
    .HI(\mprj_logic1[227] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[228]  (
    .HI(\mprj_logic1[228] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[229]  (
    .HI(\mprj_logic1[229] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[22]  (
    .HI(\mprj_logic1[22] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[230]  (
    .HI(\mprj_logic1[230] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[231]  (
    .HI(\mprj_logic1[231] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[232]  (
    .HI(\mprj_logic1[232] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[233]  (
    .HI(\mprj_logic1[233] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[234]  (
    .HI(\mprj_logic1[234] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[235]  (
    .HI(\mprj_logic1[235] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[236]  (
    .HI(\mprj_logic1[236] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[237]  (
    .HI(\mprj_logic1[237] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[238]  (
    .HI(\mprj_logic1[238] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[239]  (
    .HI(\mprj_logic1[239] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[23]  (
    .HI(\mprj_logic1[23] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[240]  (
    .HI(\mprj_logic1[240] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[241]  (
    .HI(\mprj_logic1[241] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[242]  (
    .HI(\mprj_logic1[242] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[243]  (
    .HI(\mprj_logic1[243] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[244]  (
    .HI(\mprj_logic1[244] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[245]  (
    .HI(\mprj_logic1[245] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[246]  (
    .HI(\mprj_logic1[246] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[247]  (
    .HI(\mprj_logic1[247] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[248]  (
    .HI(\mprj_logic1[248] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[249]  (
    .HI(\mprj_logic1[249] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[24]  (
    .HI(\mprj_logic1[24] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[250]  (
    .HI(\mprj_logic1[250] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[251]  (
    .HI(\mprj_logic1[251] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[252]  (
    .HI(\mprj_logic1[252] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[253]  (
    .HI(\mprj_logic1[253] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[254]  (
    .HI(\mprj_logic1[254] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[255]  (
    .HI(\mprj_logic1[255] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[256]  (
    .HI(\mprj_logic1[256] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[257]  (
    .HI(\mprj_logic1[257] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[258]  (
    .HI(\mprj_logic1[258] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[259]  (
    .HI(\mprj_logic1[259] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[25]  (
    .HI(\mprj_logic1[25] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[260]  (
    .HI(\mprj_logic1[260] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[261]  (
    .HI(\mprj_logic1[261] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[262]  (
    .HI(\mprj_logic1[262] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[263]  (
    .HI(\mprj_logic1[263] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[264]  (
    .HI(\mprj_logic1[264] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[265]  (
    .HI(\mprj_logic1[265] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[266]  (
    .HI(\mprj_logic1[266] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[267]  (
    .HI(\mprj_logic1[267] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[268]  (
    .HI(\mprj_logic1[268] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[269]  (
    .HI(\mprj_logic1[269] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[26]  (
    .HI(\mprj_logic1[26] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[270]  (
    .HI(\mprj_logic1[270] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[271]  (
    .HI(\mprj_logic1[271] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[272]  (
    .HI(\mprj_logic1[272] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[273]  (
    .HI(\mprj_logic1[273] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[274]  (
    .HI(\mprj_logic1[274] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[275]  (
    .HI(\mprj_logic1[275] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[276]  (
    .HI(\mprj_logic1[276] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[277]  (
    .HI(\mprj_logic1[277] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[278]  (
    .HI(\mprj_logic1[278] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[279]  (
    .HI(\mprj_logic1[279] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[27]  (
    .HI(\mprj_logic1[27] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[280]  (
    .HI(\mprj_logic1[280] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[281]  (
    .HI(\mprj_logic1[281] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[282]  (
    .HI(\mprj_logic1[282] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[283]  (
    .HI(\mprj_logic1[283] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[284]  (
    .HI(\mprj_logic1[284] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[285]  (
    .HI(\mprj_logic1[285] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[286]  (
    .HI(\mprj_logic1[286] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[287]  (
    .HI(\mprj_logic1[287] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[288]  (
    .HI(\mprj_logic1[288] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[289]  (
    .HI(\mprj_logic1[289] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[28]  (
    .HI(\mprj_logic1[28] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[290]  (
    .HI(\mprj_logic1[290] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[291]  (
    .HI(\mprj_logic1[291] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[292]  (
    .HI(\mprj_logic1[292] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[293]  (
    .HI(\mprj_logic1[293] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[294]  (
    .HI(\mprj_logic1[294] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[295]  (
    .HI(\mprj_logic1[295] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[296]  (
    .HI(\mprj_logic1[296] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[297]  (
    .HI(\mprj_logic1[297] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[298]  (
    .HI(\mprj_logic1[298] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[299]  (
    .HI(\mprj_logic1[299] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[29]  (
    .HI(\mprj_logic1[29] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[2]  (
    .HI(\mprj_logic1[2] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[300]  (
    .HI(\mprj_logic1[300] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[301]  (
    .HI(\mprj_logic1[301] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[302]  (
    .HI(\mprj_logic1[302] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[303]  (
    .HI(\mprj_logic1[303] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[304]  (
    .HI(\mprj_logic1[304] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[305]  (
    .HI(\mprj_logic1[305] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[306]  (
    .HI(\mprj_logic1[306] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[307]  (
    .HI(\mprj_logic1[307] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[308]  (
    .HI(\mprj_logic1[308] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[309]  (
    .HI(\mprj_logic1[309] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[30]  (
    .HI(\mprj_logic1[30] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[310]  (
    .HI(\mprj_logic1[310] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[311]  (
    .HI(\mprj_logic1[311] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[312]  (
    .HI(\mprj_logic1[312] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[313]  (
    .HI(\mprj_logic1[313] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[314]  (
    .HI(\mprj_logic1[314] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[315]  (
    .HI(\mprj_logic1[315] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[316]  (
    .HI(\mprj_logic1[316] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[317]  (
    .HI(\mprj_logic1[317] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[318]  (
    .HI(\mprj_logic1[318] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[319]  (
    .HI(\mprj_logic1[319] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[31]  (
    .HI(\mprj_logic1[31] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[320]  (
    .HI(\mprj_logic1[320] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[321]  (
    .HI(\mprj_logic1[321] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[322]  (
    .HI(\mprj_logic1[322] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[323]  (
    .HI(\mprj_logic1[323] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[324]  (
    .HI(\mprj_logic1[324] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[325]  (
    .HI(\mprj_logic1[325] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[326]  (
    .HI(\mprj_logic1[326] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[327]  (
    .HI(\mprj_logic1[327] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[328]  (
    .HI(\mprj_logic1[328] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[329]  (
    .HI(\mprj_logic1[329] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[32]  (
    .HI(\mprj_logic1[32] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[330]  (
    .HI(\mprj_logic1[330] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[331]  (
    .HI(\mprj_logic1[331] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[332]  (
    .HI(\mprj_logic1[332] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[333]  (
    .HI(\mprj_logic1[333] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[334]  (
    .HI(\mprj_logic1[334] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[335]  (
    .HI(\mprj_logic1[335] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[336]  (
    .HI(\mprj_logic1[336] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[337]  (
    .HI(\mprj_logic1[337] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[338]  (
    .HI(\mprj_logic1[338] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[339]  (
    .HI(\mprj_logic1[339] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[33]  (
    .HI(\mprj_logic1[33] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[340]  (
    .HI(\mprj_logic1[340] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[341]  (
    .HI(\mprj_logic1[341] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[342]  (
    .HI(\mprj_logic1[342] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[343]  (
    .HI(\mprj_logic1[343] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[344]  (
    .HI(\mprj_logic1[344] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[345]  (
    .HI(\mprj_logic1[345] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[346]  (
    .HI(\mprj_logic1[346] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[347]  (
    .HI(\mprj_logic1[347] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[348]  (
    .HI(\mprj_logic1[348] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[349]  (
    .HI(\mprj_logic1[349] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[34]  (
    .HI(\mprj_logic1[34] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[350]  (
    .HI(\mprj_logic1[350] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[351]  (
    .HI(\mprj_logic1[351] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[352]  (
    .HI(\mprj_logic1[352] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[353]  (
    .HI(\mprj_logic1[353] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[354]  (
    .HI(\mprj_logic1[354] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[355]  (
    .HI(\mprj_logic1[355] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[356]  (
    .HI(\mprj_logic1[356] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[357]  (
    .HI(\mprj_logic1[357] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[358]  (
    .HI(\mprj_logic1[358] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[359]  (
    .HI(\mprj_logic1[359] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[35]  (
    .HI(\mprj_logic1[35] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[360]  (
    .HI(\mprj_logic1[360] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[361]  (
    .HI(\mprj_logic1[361] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[362]  (
    .HI(\mprj_logic1[362] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[363]  (
    .HI(\mprj_logic1[363] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[364]  (
    .HI(\mprj_logic1[364] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[365]  (
    .HI(\mprj_logic1[365] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[366]  (
    .HI(\mprj_logic1[366] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[367]  (
    .HI(\mprj_logic1[367] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[368]  (
    .HI(\mprj_logic1[368] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[369]  (
    .HI(\mprj_logic1[369] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[36]  (
    .HI(\mprj_logic1[36] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[370]  (
    .HI(\mprj_logic1[370] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[371]  (
    .HI(\mprj_logic1[371] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[372]  (
    .HI(\mprj_logic1[372] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[373]  (
    .HI(\mprj_logic1[373] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[374]  (
    .HI(\mprj_logic1[374] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[375]  (
    .HI(\mprj_logic1[375] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[376]  (
    .HI(\mprj_logic1[376] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[377]  (
    .HI(\mprj_logic1[377] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[378]  (
    .HI(\mprj_logic1[378] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[379]  (
    .HI(\mprj_logic1[379] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[37]  (
    .HI(\mprj_logic1[37] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[380]  (
    .HI(\mprj_logic1[380] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[381]  (
    .HI(\mprj_logic1[381] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[382]  (
    .HI(\mprj_logic1[382] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[383]  (
    .HI(\mprj_logic1[383] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[384]  (
    .HI(\mprj_logic1[384] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[385]  (
    .HI(\mprj_logic1[385] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[386]  (
    .HI(\mprj_logic1[386] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[387]  (
    .HI(\mprj_logic1[387] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[388]  (
    .HI(\mprj_logic1[388] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[389]  (
    .HI(\mprj_logic1[389] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[38]  (
    .HI(\mprj_logic1[38] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[390]  (
    .HI(\mprj_logic1[390] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[391]  (
    .HI(\mprj_logic1[391] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[392]  (
    .HI(\mprj_logic1[392] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[393]  (
    .HI(\mprj_logic1[393] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[394]  (
    .HI(\mprj_logic1[394] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[395]  (
    .HI(\mprj_logic1[395] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[396]  (
    .HI(\mprj_logic1[396] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[397]  (
    .HI(\mprj_logic1[397] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[398]  (
    .HI(\mprj_logic1[398] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[399]  (
    .HI(\mprj_logic1[399] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[39]  (
    .HI(\mprj_logic1[39] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[3]  (
    .HI(\mprj_logic1[3] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[400]  (
    .HI(\mprj_logic1[400] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[401]  (
    .HI(\mprj_logic1[401] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[402]  (
    .HI(\mprj_logic1[402] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[403]  (
    .HI(\mprj_logic1[403] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[404]  (
    .HI(\mprj_logic1[404] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[405]  (
    .HI(\mprj_logic1[405] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[406]  (
    .HI(\mprj_logic1[406] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[407]  (
    .HI(\mprj_logic1[407] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[408]  (
    .HI(\mprj_logic1[408] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[409]  (
    .HI(\mprj_logic1[409] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[40]  (
    .HI(\mprj_logic1[40] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[410]  (
    .HI(\mprj_logic1[410] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[411]  (
    .HI(\mprj_logic1[411] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[412]  (
    .HI(\mprj_logic1[412] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[413]  (
    .HI(\mprj_logic1[413] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[414]  (
    .HI(\mprj_logic1[414] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[415]  (
    .HI(\mprj_logic1[415] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[416]  (
    .HI(\mprj_logic1[416] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[417]  (
    .HI(\mprj_logic1[417] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[418]  (
    .HI(\mprj_logic1[418] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[419]  (
    .HI(\mprj_logic1[419] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[41]  (
    .HI(\mprj_logic1[41] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[420]  (
    .HI(\mprj_logic1[420] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[421]  (
    .HI(\mprj_logic1[421] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[422]  (
    .HI(\mprj_logic1[422] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[423]  (
    .HI(\mprj_logic1[423] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[424]  (
    .HI(\mprj_logic1[424] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[425]  (
    .HI(\mprj_logic1[425] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[426]  (
    .HI(\mprj_logic1[426] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[427]  (
    .HI(\mprj_logic1[427] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[428]  (
    .HI(\mprj_logic1[428] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[429]  (
    .HI(\mprj_logic1[429] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[42]  (
    .HI(\mprj_logic1[42] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[430]  (
    .HI(\mprj_logic1[430] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[431]  (
    .HI(\mprj_logic1[431] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[432]  (
    .HI(\mprj_logic1[432] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[433]  (
    .HI(\mprj_logic1[433] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[434]  (
    .HI(\mprj_logic1[434] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[435]  (
    .HI(\mprj_logic1[435] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[436]  (
    .HI(\mprj_logic1[436] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[437]  (
    .HI(\mprj_logic1[437] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[438]  (
    .HI(\mprj_logic1[438] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[439]  (
    .HI(\mprj_logic1[439] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[43]  (
    .HI(\mprj_logic1[43] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[440]  (
    .HI(\mprj_logic1[440] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[441]  (
    .HI(\mprj_logic1[441] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[442]  (
    .HI(\mprj_logic1[442] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[443]  (
    .HI(\mprj_logic1[443] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[444]  (
    .HI(\mprj_logic1[444] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[445]  (
    .HI(\mprj_logic1[445] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[446]  (
    .HI(\mprj_logic1[446] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[447]  (
    .HI(\mprj_logic1[447] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[448]  (
    .HI(\mprj_logic1[448] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[449]  (
    .HI(\mprj_logic1[449] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[44]  (
    .HI(\mprj_logic1[44] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[450]  (
    .HI(\mprj_logic1[450] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[451]  (
    .HI(\mprj_logic1[451] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[452]  (
    .HI(\mprj_logic1[452] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[453]  (
    .HI(\mprj_logic1[453] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[454]  (
    .HI(\mprj_logic1[454] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[455]  (
    .HI(\mprj_logic1[455] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[456]  (
    .HI(\mprj_logic1[456] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[457]  (
    .HI(\mprj_logic1[457] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[458]  (
    .HI(\mprj_logic1[458] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[45]  (
    .HI(\mprj_logic1[45] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[46]  (
    .HI(\mprj_logic1[46] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[47]  (
    .HI(\mprj_logic1[47] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[48]  (
    .HI(\mprj_logic1[48] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[49]  (
    .HI(\mprj_logic1[49] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[4]  (
    .HI(\mprj_logic1[4] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[50]  (
    .HI(\mprj_logic1[50] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[51]  (
    .HI(\mprj_logic1[51] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[52]  (
    .HI(\mprj_logic1[52] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[53]  (
    .HI(\mprj_logic1[53] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[54]  (
    .HI(\mprj_logic1[54] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[55]  (
    .HI(\mprj_logic1[55] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[56]  (
    .HI(\mprj_logic1[56] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[57]  (
    .HI(\mprj_logic1[57] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[58]  (
    .HI(\mprj_logic1[58] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[59]  (
    .HI(\mprj_logic1[59] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[5]  (
    .HI(\mprj_logic1[5] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[60]  (
    .HI(\mprj_logic1[60] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[61]  (
    .HI(\mprj_logic1[61] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[62]  (
    .HI(\mprj_logic1[62] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[63]  (
    .HI(\mprj_logic1[63] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[64]  (
    .HI(\mprj_logic1[64] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[65]  (
    .HI(\mprj_logic1[65] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[66]  (
    .HI(\mprj_logic1[66] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[67]  (
    .HI(\mprj_logic1[67] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[68]  (
    .HI(\mprj_logic1[68] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[69]  (
    .HI(\mprj_logic1[69] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[6]  (
    .HI(\mprj_logic1[6] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[70]  (
    .HI(\mprj_logic1[70] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[71]  (
    .HI(\mprj_logic1[71] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[72]  (
    .HI(\mprj_logic1[72] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[73]  (
    .HI(\mprj_logic1[73] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[74]  (
    .HI(\mprj_logic1[74] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[75]  (
    .HI(\mprj_logic1[75] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[76]  (
    .HI(\mprj_logic1[76] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[77]  (
    .HI(\mprj_logic1[77] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[78]  (
    .HI(\mprj_logic1[78] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[79]  (
    .HI(\mprj_logic1[79] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[7]  (
    .HI(\mprj_logic1[7] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[80]  (
    .HI(\mprj_logic1[80] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[81]  (
    .HI(\mprj_logic1[81] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[82]  (
    .HI(\mprj_logic1[82] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[83]  (
    .HI(\mprj_logic1[83] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[84]  (
    .HI(\mprj_logic1[84] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[85]  (
    .HI(\mprj_logic1[85] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[86]  (
    .HI(\mprj_logic1[86] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[87]  (
    .HI(\mprj_logic1[87] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[88]  (
    .HI(\mprj_logic1[88] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[89]  (
    .HI(\mprj_logic1[89] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[8]  (
    .HI(\mprj_logic1[8] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[90]  (
    .HI(\mprj_logic1[90] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[91]  (
    .HI(\mprj_logic1[91] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[92]  (
    .HI(\mprj_logic1[92] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[93]  (
    .HI(\mprj_logic1[93] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[94]  (
    .HI(\mprj_logic1[94] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[95]  (
    .HI(\mprj_logic1[95] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[96]  (
    .HI(\mprj_logic1[96] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[97]  (
    .HI(\mprj_logic1[97] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[98]  (
    .HI(\mprj_logic1[98] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[99]  (
    .HI(\mprj_logic1[99] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__conb_1 \mprj_logic_high[9]  (
    .HI(\mprj_logic1[9] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hd__buf_8 mprj_pwrgood (
    .A(\mprj_logic1[458] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .X(user1_vcc_powergood)
  );
  sky130_fd_sc_hd__einvp_8 mprj_rstn_buf (
    .A(_000_),
    .TE(\mprj_logic1[0] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(user_resetn)
  );
  sky130_fd_sc_hd__einvp_8 \mprj_sel_buf[0]  (
    .A(_006_),
    .TE(\mprj_logic1[6] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_sel_o_user[0])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_sel_buf[1]  (
    .A(_007_),
    .TE(\mprj_logic1[7] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_sel_o_user[1])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_sel_buf[2]  (
    .A(_008_),
    .TE(\mprj_logic1[8] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_sel_o_user[2])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_sel_buf[3]  (
    .A(_009_),
    .TE(\mprj_logic1[9] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_sel_o_user[3])
  );
  sky130_fd_sc_hd__einvp_8 mprj_stb_buf (
    .A(_004_),
    .TE(\mprj_logic1[4] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_stb_o_user)
  );
  sky130_fd_sc_hd__buf_8 mprj_vdd_pwrgood (
    .A(mprj_vdd_logic1),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .X(user1_vdd_powergood)
  );
  sky130_fd_sc_hd__einvp_8 mprj_we_buf (
    .A(_005_),
    .TE(\mprj_logic1[5] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(mprj_we_o_user)
  );
  mgmt_protect_hv powergood_check (
    .mprj2_vdd_logic1(mprj2_vdd_logic1),
    .mprj_vdd_logic1(mprj_vdd_logic1),
    .vccd(vdda2),
    .vdda1(vdda2),
    .vdda2(vdda2),
    .vssa1(vssa2),
    .vssa2(vssa2),
    .vssd(vssa2)
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[0]  (
    .A(\la_data_in_mprj_bar[0] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[0])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[100]  (
    .A(\la_data_in_mprj_bar[100] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[100])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[101]  (
    .A(\la_data_in_mprj_bar[101] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[101])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[102]  (
    .A(\la_data_in_mprj_bar[102] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[102])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[103]  (
    .A(\la_data_in_mprj_bar[103] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[103])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[104]  (
    .A(\la_data_in_mprj_bar[104] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[104])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[105]  (
    .A(\la_data_in_mprj_bar[105] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[105])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[106]  (
    .A(\la_data_in_mprj_bar[106] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[106])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[107]  (
    .A(\la_data_in_mprj_bar[107] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[107])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[108]  (
    .A(\la_data_in_mprj_bar[108] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[108])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[109]  (
    .A(\la_data_in_mprj_bar[109] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[109])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[10]  (
    .A(\la_data_in_mprj_bar[10] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[10])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[110]  (
    .A(\la_data_in_mprj_bar[110] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[110])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[111]  (
    .A(\la_data_in_mprj_bar[111] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[111])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[112]  (
    .A(\la_data_in_mprj_bar[112] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[112])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[113]  (
    .A(\la_data_in_mprj_bar[113] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[113])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[114]  (
    .A(\la_data_in_mprj_bar[114] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[114])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[115]  (
    .A(\la_data_in_mprj_bar[115] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[115])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[116]  (
    .A(\la_data_in_mprj_bar[116] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[116])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[117]  (
    .A(\la_data_in_mprj_bar[117] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[117])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[118]  (
    .A(\la_data_in_mprj_bar[118] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[118])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[119]  (
    .A(\la_data_in_mprj_bar[119] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[119])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[11]  (
    .A(\la_data_in_mprj_bar[11] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[11])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[120]  (
    .A(\la_data_in_mprj_bar[120] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[120])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[121]  (
    .A(\la_data_in_mprj_bar[121] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[121])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[122]  (
    .A(\la_data_in_mprj_bar[122] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[122])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[123]  (
    .A(\la_data_in_mprj_bar[123] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[123])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[124]  (
    .A(\la_data_in_mprj_bar[124] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[124])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[125]  (
    .A(\la_data_in_mprj_bar[125] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[125])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[126]  (
    .A(\la_data_in_mprj_bar[126] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[126])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[127]  (
    .A(\la_data_in_mprj_bar[127] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[127])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[12]  (
    .A(\la_data_in_mprj_bar[12] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[12])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[13]  (
    .A(\la_data_in_mprj_bar[13] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[13])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[14]  (
    .A(\la_data_in_mprj_bar[14] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[14])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[15]  (
    .A(\la_data_in_mprj_bar[15] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[15])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[16]  (
    .A(\la_data_in_mprj_bar[16] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[16])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[17]  (
    .A(\la_data_in_mprj_bar[17] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[17])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[18]  (
    .A(\la_data_in_mprj_bar[18] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[18])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[19]  (
    .A(\la_data_in_mprj_bar[19] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[19])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[1]  (
    .A(\la_data_in_mprj_bar[1] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[1])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[20]  (
    .A(\la_data_in_mprj_bar[20] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[20])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[21]  (
    .A(\la_data_in_mprj_bar[21] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[21])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[22]  (
    .A(\la_data_in_mprj_bar[22] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[22])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[23]  (
    .A(\la_data_in_mprj_bar[23] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[23])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[24]  (
    .A(\la_data_in_mprj_bar[24] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[24])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[25]  (
    .A(\la_data_in_mprj_bar[25] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[25])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[26]  (
    .A(\la_data_in_mprj_bar[26] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[26])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[27]  (
    .A(\la_data_in_mprj_bar[27] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[27])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[28]  (
    .A(\la_data_in_mprj_bar[28] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[28])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[29]  (
    .A(\la_data_in_mprj_bar[29] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[29])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[2]  (
    .A(\la_data_in_mprj_bar[2] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[2])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[30]  (
    .A(\la_data_in_mprj_bar[30] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[30])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[31]  (
    .A(\la_data_in_mprj_bar[31] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[31])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[32]  (
    .A(\la_data_in_mprj_bar[32] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[32])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[33]  (
    .A(\la_data_in_mprj_bar[33] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[33])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[34]  (
    .A(\la_data_in_mprj_bar[34] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[34])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[35]  (
    .A(\la_data_in_mprj_bar[35] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[35])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[36]  (
    .A(\la_data_in_mprj_bar[36] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[36])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[37]  (
    .A(\la_data_in_mprj_bar[37] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[37])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[38]  (
    .A(\la_data_in_mprj_bar[38] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[38])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[39]  (
    .A(\la_data_in_mprj_bar[39] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[39])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[3]  (
    .A(\la_data_in_mprj_bar[3] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[3])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[40]  (
    .A(\la_data_in_mprj_bar[40] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[40])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[41]  (
    .A(\la_data_in_mprj_bar[41] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[41])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[42]  (
    .A(\la_data_in_mprj_bar[42] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[42])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[43]  (
    .A(\la_data_in_mprj_bar[43] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[43])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[44]  (
    .A(\la_data_in_mprj_bar[44] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[44])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[45]  (
    .A(\la_data_in_mprj_bar[45] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[45])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[46]  (
    .A(\la_data_in_mprj_bar[46] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[46])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[47]  (
    .A(\la_data_in_mprj_bar[47] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[47])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[48]  (
    .A(\la_data_in_mprj_bar[48] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[48])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[49]  (
    .A(\la_data_in_mprj_bar[49] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[49])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[4]  (
    .A(\la_data_in_mprj_bar[4] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[4])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[50]  (
    .A(\la_data_in_mprj_bar[50] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[50])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[51]  (
    .A(\la_data_in_mprj_bar[51] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[51])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[52]  (
    .A(\la_data_in_mprj_bar[52] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[52])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[53]  (
    .A(\la_data_in_mprj_bar[53] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[53])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[54]  (
    .A(\la_data_in_mprj_bar[54] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[54])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[55]  (
    .A(\la_data_in_mprj_bar[55] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[55])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[56]  (
    .A(\la_data_in_mprj_bar[56] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[56])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[57]  (
    .A(\la_data_in_mprj_bar[57] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[57])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[58]  (
    .A(\la_data_in_mprj_bar[58] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[58])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[59]  (
    .A(\la_data_in_mprj_bar[59] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[59])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[5]  (
    .A(\la_data_in_mprj_bar[5] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[5])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[60]  (
    .A(\la_data_in_mprj_bar[60] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[60])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[61]  (
    .A(\la_data_in_mprj_bar[61] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[61])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[62]  (
    .A(\la_data_in_mprj_bar[62] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[62])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[63]  (
    .A(\la_data_in_mprj_bar[63] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[63])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[64]  (
    .A(\la_data_in_mprj_bar[64] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[64])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[65]  (
    .A(\la_data_in_mprj_bar[65] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[65])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[66]  (
    .A(\la_data_in_mprj_bar[66] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[66])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[67]  (
    .A(\la_data_in_mprj_bar[67] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[67])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[68]  (
    .A(\la_data_in_mprj_bar[68] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[68])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[69]  (
    .A(\la_data_in_mprj_bar[69] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[69])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[6]  (
    .A(\la_data_in_mprj_bar[6] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[6])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[70]  (
    .A(\la_data_in_mprj_bar[70] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[70])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[71]  (
    .A(\la_data_in_mprj_bar[71] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[71])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[72]  (
    .A(\la_data_in_mprj_bar[72] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[72])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[73]  (
    .A(\la_data_in_mprj_bar[73] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[73])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[74]  (
    .A(\la_data_in_mprj_bar[74] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[74])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[75]  (
    .A(\la_data_in_mprj_bar[75] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[75])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[76]  (
    .A(\la_data_in_mprj_bar[76] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[76])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[77]  (
    .A(\la_data_in_mprj_bar[77] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[77])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[78]  (
    .A(\la_data_in_mprj_bar[78] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[78])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[79]  (
    .A(\la_data_in_mprj_bar[79] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[79])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[7]  (
    .A(\la_data_in_mprj_bar[7] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[7])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[80]  (
    .A(\la_data_in_mprj_bar[80] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[80])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[81]  (
    .A(\la_data_in_mprj_bar[81] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[81])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[82]  (
    .A(\la_data_in_mprj_bar[82] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[82])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[83]  (
    .A(\la_data_in_mprj_bar[83] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[83])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[84]  (
    .A(\la_data_in_mprj_bar[84] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[84])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[85]  (
    .A(\la_data_in_mprj_bar[85] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[85])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[86]  (
    .A(\la_data_in_mprj_bar[86] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[86])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[87]  (
    .A(\la_data_in_mprj_bar[87] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[87])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[88]  (
    .A(\la_data_in_mprj_bar[88] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[88])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[89]  (
    .A(\la_data_in_mprj_bar[89] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[89])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[8]  (
    .A(\la_data_in_mprj_bar[8] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[8])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[90]  (
    .A(\la_data_in_mprj_bar[90] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[90])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[91]  (
    .A(\la_data_in_mprj_bar[91] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[91])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[92]  (
    .A(\la_data_in_mprj_bar[92] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[92])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[93]  (
    .A(\la_data_in_mprj_bar[93] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[93])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[94]  (
    .A(\la_data_in_mprj_bar[94] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[94])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[95]  (
    .A(\la_data_in_mprj_bar[95] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[95])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[96]  (
    .A(\la_data_in_mprj_bar[96] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[96])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[97]  (
    .A(\la_data_in_mprj_bar[97] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[97])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[98]  (
    .A(\la_data_in_mprj_bar[98] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[98])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[99]  (
    .A(\la_data_in_mprj_bar[99] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[99])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[9]  (
    .A(\la_data_in_mprj_bar[9] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(la_data_in_mprj[9])
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[0]  (
    .A(la_data_out_core[0]),
    .B(\mprj_logic1[330] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[0] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[100]  (
    .A(la_data_out_core[100]),
    .B(\mprj_logic1[430] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[100] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[101]  (
    .A(la_data_out_core[101]),
    .B(\mprj_logic1[431] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[101] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[102]  (
    .A(la_data_out_core[102]),
    .B(\mprj_logic1[432] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[102] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[103]  (
    .A(la_data_out_core[103]),
    .B(\mprj_logic1[433] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[103] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[104]  (
    .A(la_data_out_core[104]),
    .B(\mprj_logic1[434] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[104] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[105]  (
    .A(la_data_out_core[105]),
    .B(\mprj_logic1[435] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[105] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[106]  (
    .A(la_data_out_core[106]),
    .B(\mprj_logic1[436] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[106] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[107]  (
    .A(la_data_out_core[107]),
    .B(\mprj_logic1[437] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[107] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[108]  (
    .A(la_data_out_core[108]),
    .B(\mprj_logic1[438] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[108] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[109]  (
    .A(la_data_out_core[109]),
    .B(\mprj_logic1[439] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[109] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[10]  (
    .A(la_data_out_core[10]),
    .B(\mprj_logic1[340] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[10] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[110]  (
    .A(la_data_out_core[110]),
    .B(\mprj_logic1[440] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[110] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[111]  (
    .A(la_data_out_core[111]),
    .B(\mprj_logic1[441] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[111] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[112]  (
    .A(la_data_out_core[112]),
    .B(\mprj_logic1[442] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[112] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[113]  (
    .A(la_data_out_core[113]),
    .B(\mprj_logic1[443] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[113] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[114]  (
    .A(la_data_out_core[114]),
    .B(\mprj_logic1[444] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[114] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[115]  (
    .A(la_data_out_core[115]),
    .B(\mprj_logic1[445] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[115] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[116]  (
    .A(la_data_out_core[116]),
    .B(\mprj_logic1[446] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[116] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[117]  (
    .A(la_data_out_core[117]),
    .B(\mprj_logic1[447] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[117] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[118]  (
    .A(la_data_out_core[118]),
    .B(\mprj_logic1[448] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[118] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[119]  (
    .A(la_data_out_core[119]),
    .B(\mprj_logic1[449] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[119] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[11]  (
    .A(la_data_out_core[11]),
    .B(\mprj_logic1[341] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[11] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[120]  (
    .A(la_data_out_core[120]),
    .B(\mprj_logic1[450] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[120] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[121]  (
    .A(la_data_out_core[121]),
    .B(\mprj_logic1[451] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[121] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[122]  (
    .A(la_data_out_core[122]),
    .B(\mprj_logic1[452] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[122] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[123]  (
    .A(la_data_out_core[123]),
    .B(\mprj_logic1[453] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[123] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[124]  (
    .A(la_data_out_core[124]),
    .B(\mprj_logic1[454] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[124] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[125]  (
    .A(la_data_out_core[125]),
    .B(\mprj_logic1[455] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[125] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[126]  (
    .A(la_data_out_core[126]),
    .B(\mprj_logic1[456] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[126] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[127]  (
    .A(la_data_out_core[127]),
    .B(\mprj_logic1[457] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[127] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[12]  (
    .A(la_data_out_core[12]),
    .B(\mprj_logic1[342] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[12] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[13]  (
    .A(la_data_out_core[13]),
    .B(\mprj_logic1[343] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[13] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[14]  (
    .A(la_data_out_core[14]),
    .B(\mprj_logic1[344] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[14] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[15]  (
    .A(la_data_out_core[15]),
    .B(\mprj_logic1[345] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[15] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[16]  (
    .A(la_data_out_core[16]),
    .B(\mprj_logic1[346] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[16] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[17]  (
    .A(la_data_out_core[17]),
    .B(\mprj_logic1[347] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[17] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[18]  (
    .A(la_data_out_core[18]),
    .B(\mprj_logic1[348] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[18] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[19]  (
    .A(la_data_out_core[19]),
    .B(\mprj_logic1[349] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[19] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[1]  (
    .A(la_data_out_core[1]),
    .B(\mprj_logic1[331] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[1] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[20]  (
    .A(la_data_out_core[20]),
    .B(\mprj_logic1[350] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[20] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[21]  (
    .A(la_data_out_core[21]),
    .B(\mprj_logic1[351] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[21] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[22]  (
    .A(la_data_out_core[22]),
    .B(\mprj_logic1[352] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[22] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[23]  (
    .A(la_data_out_core[23]),
    .B(\mprj_logic1[353] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[23] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[24]  (
    .A(la_data_out_core[24]),
    .B(\mprj_logic1[354] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[24] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[25]  (
    .A(la_data_out_core[25]),
    .B(\mprj_logic1[355] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[25] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[26]  (
    .A(la_data_out_core[26]),
    .B(\mprj_logic1[356] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[26] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[27]  (
    .A(la_data_out_core[27]),
    .B(\mprj_logic1[357] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[27] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[28]  (
    .A(la_data_out_core[28]),
    .B(\mprj_logic1[358] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[28] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[29]  (
    .A(la_data_out_core[29]),
    .B(\mprj_logic1[359] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[29] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[2]  (
    .A(la_data_out_core[2]),
    .B(\mprj_logic1[332] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[2] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[30]  (
    .A(la_data_out_core[30]),
    .B(\mprj_logic1[360] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[30] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[31]  (
    .A(la_data_out_core[31]),
    .B(\mprj_logic1[361] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[31] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[32]  (
    .A(la_data_out_core[32]),
    .B(\mprj_logic1[362] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[32] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[33]  (
    .A(la_data_out_core[33]),
    .B(\mprj_logic1[363] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[33] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[34]  (
    .A(la_data_out_core[34]),
    .B(\mprj_logic1[364] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[34] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[35]  (
    .A(la_data_out_core[35]),
    .B(\mprj_logic1[365] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[35] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[36]  (
    .A(la_data_out_core[36]),
    .B(\mprj_logic1[366] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[36] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[37]  (
    .A(la_data_out_core[37]),
    .B(\mprj_logic1[367] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[37] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[38]  (
    .A(la_data_out_core[38]),
    .B(\mprj_logic1[368] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[38] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[39]  (
    .A(la_data_out_core[39]),
    .B(\mprj_logic1[369] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[39] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[3]  (
    .A(la_data_out_core[3]),
    .B(\mprj_logic1[333] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[3] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[40]  (
    .A(la_data_out_core[40]),
    .B(\mprj_logic1[370] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[40] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[41]  (
    .A(la_data_out_core[41]),
    .B(\mprj_logic1[371] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[41] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[42]  (
    .A(la_data_out_core[42]),
    .B(\mprj_logic1[372] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[42] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[43]  (
    .A(la_data_out_core[43]),
    .B(\mprj_logic1[373] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[43] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[44]  (
    .A(la_data_out_core[44]),
    .B(\mprj_logic1[374] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[44] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[45]  (
    .A(la_data_out_core[45]),
    .B(\mprj_logic1[375] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[45] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[46]  (
    .A(la_data_out_core[46]),
    .B(\mprj_logic1[376] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[46] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[47]  (
    .A(la_data_out_core[47]),
    .B(\mprj_logic1[377] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[47] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[48]  (
    .A(la_data_out_core[48]),
    .B(\mprj_logic1[378] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[48] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[49]  (
    .A(la_data_out_core[49]),
    .B(\mprj_logic1[379] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[49] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[4]  (
    .A(la_data_out_core[4]),
    .B(\mprj_logic1[334] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[4] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[50]  (
    .A(la_data_out_core[50]),
    .B(\mprj_logic1[380] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[50] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[51]  (
    .A(la_data_out_core[51]),
    .B(\mprj_logic1[381] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[51] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[52]  (
    .A(la_data_out_core[52]),
    .B(\mprj_logic1[382] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[52] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[53]  (
    .A(la_data_out_core[53]),
    .B(\mprj_logic1[383] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[53] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[54]  (
    .A(la_data_out_core[54]),
    .B(\mprj_logic1[384] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[54] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[55]  (
    .A(la_data_out_core[55]),
    .B(\mprj_logic1[385] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[55] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[56]  (
    .A(la_data_out_core[56]),
    .B(\mprj_logic1[386] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[56] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[57]  (
    .A(la_data_out_core[57]),
    .B(\mprj_logic1[387] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[57] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[58]  (
    .A(la_data_out_core[58]),
    .B(\mprj_logic1[388] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[58] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[59]  (
    .A(la_data_out_core[59]),
    .B(\mprj_logic1[389] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[59] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[5]  (
    .A(la_data_out_core[5]),
    .B(\mprj_logic1[335] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[5] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[60]  (
    .A(la_data_out_core[60]),
    .B(\mprj_logic1[390] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[60] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[61]  (
    .A(la_data_out_core[61]),
    .B(\mprj_logic1[391] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[61] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[62]  (
    .A(la_data_out_core[62]),
    .B(\mprj_logic1[392] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[62] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[63]  (
    .A(la_data_out_core[63]),
    .B(\mprj_logic1[393] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[63] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[64]  (
    .A(la_data_out_core[64]),
    .B(\mprj_logic1[394] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[64] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[65]  (
    .A(la_data_out_core[65]),
    .B(\mprj_logic1[395] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[65] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[66]  (
    .A(la_data_out_core[66]),
    .B(\mprj_logic1[396] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[66] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[67]  (
    .A(la_data_out_core[67]),
    .B(\mprj_logic1[397] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[67] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[68]  (
    .A(la_data_out_core[68]),
    .B(\mprj_logic1[398] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[68] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[69]  (
    .A(la_data_out_core[69]),
    .B(\mprj_logic1[399] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[69] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[6]  (
    .A(la_data_out_core[6]),
    .B(\mprj_logic1[336] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[6] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[70]  (
    .A(la_data_out_core[70]),
    .B(\mprj_logic1[400] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[70] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[71]  (
    .A(la_data_out_core[71]),
    .B(\mprj_logic1[401] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[71] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[72]  (
    .A(la_data_out_core[72]),
    .B(\mprj_logic1[402] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[72] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[73]  (
    .A(la_data_out_core[73]),
    .B(\mprj_logic1[403] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[73] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[74]  (
    .A(la_data_out_core[74]),
    .B(\mprj_logic1[404] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[74] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[75]  (
    .A(la_data_out_core[75]),
    .B(\mprj_logic1[405] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[75] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[76]  (
    .A(la_data_out_core[76]),
    .B(\mprj_logic1[406] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[76] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[77]  (
    .A(la_data_out_core[77]),
    .B(\mprj_logic1[407] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[77] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[78]  (
    .A(la_data_out_core[78]),
    .B(\mprj_logic1[408] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[78] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[79]  (
    .A(la_data_out_core[79]),
    .B(\mprj_logic1[409] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[79] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[7]  (
    .A(la_data_out_core[7]),
    .B(\mprj_logic1[337] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[7] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[80]  (
    .A(la_data_out_core[80]),
    .B(\mprj_logic1[410] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[80] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[81]  (
    .A(la_data_out_core[81]),
    .B(\mprj_logic1[411] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[81] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[82]  (
    .A(la_data_out_core[82]),
    .B(\mprj_logic1[412] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[82] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[83]  (
    .A(la_data_out_core[83]),
    .B(\mprj_logic1[413] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[83] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[84]  (
    .A(la_data_out_core[84]),
    .B(\mprj_logic1[414] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[84] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[85]  (
    .A(la_data_out_core[85]),
    .B(\mprj_logic1[415] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[85] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[86]  (
    .A(la_data_out_core[86]),
    .B(\mprj_logic1[416] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[86] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[87]  (
    .A(la_data_out_core[87]),
    .B(\mprj_logic1[417] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[87] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[88]  (
    .A(la_data_out_core[88]),
    .B(\mprj_logic1[418] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[88] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[89]  (
    .A(la_data_out_core[89]),
    .B(\mprj_logic1[419] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[89] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[8]  (
    .A(la_data_out_core[8]),
    .B(\mprj_logic1[338] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[8] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[90]  (
    .A(la_data_out_core[90]),
    .B(\mprj_logic1[420] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[90] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[91]  (
    .A(la_data_out_core[91]),
    .B(\mprj_logic1[421] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[91] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[92]  (
    .A(la_data_out_core[92]),
    .B(\mprj_logic1[422] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[92] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[93]  (
    .A(la_data_out_core[93]),
    .B(\mprj_logic1[423] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[93] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[94]  (
    .A(la_data_out_core[94]),
    .B(\mprj_logic1[424] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[94] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[95]  (
    .A(la_data_out_core[95]),
    .B(\mprj_logic1[425] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[95] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[96]  (
    .A(la_data_out_core[96]),
    .B(\mprj_logic1[426] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[96] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[97]  (
    .A(la_data_out_core[97]),
    .B(\mprj_logic1[427] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[97] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[98]  (
    .A(la_data_out_core[98]),
    .B(\mprj_logic1[428] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[98] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[99]  (
    .A(la_data_out_core[99]),
    .B(\mprj_logic1[429] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[99] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[9]  (
    .A(la_data_out_core[9]),
    .B(\mprj_logic1[339] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Y(\la_data_in_mprj_bar[9] )
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[0]  (
    .A(_202_),
    .TE(\mprj_logic1[202] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[0])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[100]  (
    .A(_203_),
    .TE(\mprj_logic1[302] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[100])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[101]  (
    .A(_204_),
    .TE(\mprj_logic1[303] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[101])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[102]  (
    .A(_205_),
    .TE(\mprj_logic1[304] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[102])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[103]  (
    .A(_206_),
    .TE(\mprj_logic1[305] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[103])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[104]  (
    .A(_207_),
    .TE(\mprj_logic1[306] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[104])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[105]  (
    .A(_208_),
    .TE(\mprj_logic1[307] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[105])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[106]  (
    .A(_209_),
    .TE(\mprj_logic1[308] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[106])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[107]  (
    .A(_210_),
    .TE(\mprj_logic1[309] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[107])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[108]  (
    .A(_211_),
    .TE(\mprj_logic1[310] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[108])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[109]  (
    .A(_212_),
    .TE(\mprj_logic1[311] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[109])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[10]  (
    .A(_213_),
    .TE(\mprj_logic1[212] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[10])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[110]  (
    .A(_214_),
    .TE(\mprj_logic1[312] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[110])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[111]  (
    .A(_215_),
    .TE(\mprj_logic1[313] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[111])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[112]  (
    .A(_216_),
    .TE(\mprj_logic1[314] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[112])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[113]  (
    .A(_217_),
    .TE(\mprj_logic1[315] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[113])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[114]  (
    .A(_218_),
    .TE(\mprj_logic1[316] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[114])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[115]  (
    .A(_219_),
    .TE(\mprj_logic1[317] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[115])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[116]  (
    .A(_220_),
    .TE(\mprj_logic1[318] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[116])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[117]  (
    .A(_221_),
    .TE(\mprj_logic1[319] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[117])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[118]  (
    .A(_222_),
    .TE(\mprj_logic1[320] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[118])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[119]  (
    .A(_223_),
    .TE(\mprj_logic1[321] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[119])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[11]  (
    .A(_224_),
    .TE(\mprj_logic1[213] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[11])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[120]  (
    .A(_225_),
    .TE(\mprj_logic1[322] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[120])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[121]  (
    .A(_226_),
    .TE(\mprj_logic1[323] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[121])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[122]  (
    .A(_227_),
    .TE(\mprj_logic1[324] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[122])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[123]  (
    .A(_228_),
    .TE(\mprj_logic1[325] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[123])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[124]  (
    .A(_229_),
    .TE(\mprj_logic1[326] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[124])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[125]  (
    .A(_230_),
    .TE(\mprj_logic1[327] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[125])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[126]  (
    .A(_231_),
    .TE(\mprj_logic1[328] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[126])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[127]  (
    .A(_232_),
    .TE(\mprj_logic1[329] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[127])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[12]  (
    .A(_233_),
    .TE(\mprj_logic1[214] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[12])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[13]  (
    .A(_234_),
    .TE(\mprj_logic1[215] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[13])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[14]  (
    .A(_235_),
    .TE(\mprj_logic1[216] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[14])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[15]  (
    .A(_236_),
    .TE(\mprj_logic1[217] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[15])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[16]  (
    .A(_237_),
    .TE(\mprj_logic1[218] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[16])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[17]  (
    .A(_238_),
    .TE(\mprj_logic1[219] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[17])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[18]  (
    .A(_239_),
    .TE(\mprj_logic1[220] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[18])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[19]  (
    .A(_240_),
    .TE(\mprj_logic1[221] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[19])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[1]  (
    .A(_241_),
    .TE(\mprj_logic1[203] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[1])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[20]  (
    .A(_242_),
    .TE(\mprj_logic1[222] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[20])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[21]  (
    .A(_243_),
    .TE(\mprj_logic1[223] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[21])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[22]  (
    .A(_244_),
    .TE(\mprj_logic1[224] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[22])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[23]  (
    .A(_245_),
    .TE(\mprj_logic1[225] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[23])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[24]  (
    .A(_246_),
    .TE(\mprj_logic1[226] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[24])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[25]  (
    .A(_247_),
    .TE(\mprj_logic1[227] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[25])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[26]  (
    .A(_248_),
    .TE(\mprj_logic1[228] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[26])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[27]  (
    .A(_249_),
    .TE(\mprj_logic1[229] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[27])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[28]  (
    .A(_250_),
    .TE(\mprj_logic1[230] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[28])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[29]  (
    .A(_251_),
    .TE(\mprj_logic1[231] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[29])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[2]  (
    .A(_252_),
    .TE(\mprj_logic1[204] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[2])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[30]  (
    .A(_253_),
    .TE(\mprj_logic1[232] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[30])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[31]  (
    .A(_254_),
    .TE(\mprj_logic1[233] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[31])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[32]  (
    .A(_255_),
    .TE(\mprj_logic1[234] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[32])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[33]  (
    .A(_256_),
    .TE(\mprj_logic1[235] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[33])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[34]  (
    .A(_257_),
    .TE(\mprj_logic1[236] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[34])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[35]  (
    .A(_258_),
    .TE(\mprj_logic1[237] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[35])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[36]  (
    .A(_259_),
    .TE(\mprj_logic1[238] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[36])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[37]  (
    .A(_260_),
    .TE(\mprj_logic1[239] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[37])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[38]  (
    .A(_261_),
    .TE(\mprj_logic1[240] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[38])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[39]  (
    .A(_262_),
    .TE(\mprj_logic1[241] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[39])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[3]  (
    .A(_263_),
    .TE(\mprj_logic1[205] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[3])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[40]  (
    .A(_264_),
    .TE(\mprj_logic1[242] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[40])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[41]  (
    .A(_265_),
    .TE(\mprj_logic1[243] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[41])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[42]  (
    .A(_266_),
    .TE(\mprj_logic1[244] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[42])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[43]  (
    .A(_267_),
    .TE(\mprj_logic1[245] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[43])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[44]  (
    .A(_268_),
    .TE(\mprj_logic1[246] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[44])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[45]  (
    .A(_269_),
    .TE(\mprj_logic1[247] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[45])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[46]  (
    .A(_270_),
    .TE(\mprj_logic1[248] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[46])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[47]  (
    .A(_271_),
    .TE(\mprj_logic1[249] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[47])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[48]  (
    .A(_272_),
    .TE(\mprj_logic1[250] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[48])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[49]  (
    .A(_273_),
    .TE(\mprj_logic1[251] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[49])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[4]  (
    .A(_274_),
    .TE(\mprj_logic1[206] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[4])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[50]  (
    .A(_275_),
    .TE(\mprj_logic1[252] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[50])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[51]  (
    .A(_276_),
    .TE(\mprj_logic1[253] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[51])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[52]  (
    .A(_277_),
    .TE(\mprj_logic1[254] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[52])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[53]  (
    .A(_278_),
    .TE(\mprj_logic1[255] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[53])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[54]  (
    .A(_279_),
    .TE(\mprj_logic1[256] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[54])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[55]  (
    .A(_280_),
    .TE(\mprj_logic1[257] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[55])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[56]  (
    .A(_281_),
    .TE(\mprj_logic1[258] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[56])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[57]  (
    .A(_282_),
    .TE(\mprj_logic1[259] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[57])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[58]  (
    .A(_283_),
    .TE(\mprj_logic1[260] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[58])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[59]  (
    .A(_284_),
    .TE(\mprj_logic1[261] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[59])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[5]  (
    .A(_285_),
    .TE(\mprj_logic1[207] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[5])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[60]  (
    .A(_286_),
    .TE(\mprj_logic1[262] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[60])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[61]  (
    .A(_287_),
    .TE(\mprj_logic1[263] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[61])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[62]  (
    .A(_288_),
    .TE(\mprj_logic1[264] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[62])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[63]  (
    .A(_289_),
    .TE(\mprj_logic1[265] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[63])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[64]  (
    .A(_290_),
    .TE(\mprj_logic1[266] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[64])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[65]  (
    .A(_291_),
    .TE(\mprj_logic1[267] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[65])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[66]  (
    .A(_292_),
    .TE(\mprj_logic1[268] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[66])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[67]  (
    .A(_293_),
    .TE(\mprj_logic1[269] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[67])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[68]  (
    .A(_294_),
    .TE(\mprj_logic1[270] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[68])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[69]  (
    .A(_295_),
    .TE(\mprj_logic1[271] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[69])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[6]  (
    .A(_296_),
    .TE(\mprj_logic1[208] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[6])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[70]  (
    .A(_297_),
    .TE(\mprj_logic1[272] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[70])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[71]  (
    .A(_298_),
    .TE(\mprj_logic1[273] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[71])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[72]  (
    .A(_299_),
    .TE(\mprj_logic1[274] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[72])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[73]  (
    .A(_300_),
    .TE(\mprj_logic1[275] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[73])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[74]  (
    .A(_301_),
    .TE(\mprj_logic1[276] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[74])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[75]  (
    .A(_302_),
    .TE(\mprj_logic1[277] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[75])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[76]  (
    .A(_303_),
    .TE(\mprj_logic1[278] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[76])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[77]  (
    .A(_304_),
    .TE(\mprj_logic1[279] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[77])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[78]  (
    .A(_305_),
    .TE(\mprj_logic1[280] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[78])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[79]  (
    .A(_306_),
    .TE(\mprj_logic1[281] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[79])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[7]  (
    .A(_307_),
    .TE(\mprj_logic1[209] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[7])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[80]  (
    .A(_308_),
    .TE(\mprj_logic1[282] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[80])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[81]  (
    .A(_309_),
    .TE(\mprj_logic1[283] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[81])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[82]  (
    .A(_310_),
    .TE(\mprj_logic1[284] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[82])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[83]  (
    .A(_311_),
    .TE(\mprj_logic1[285] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[83])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[84]  (
    .A(_312_),
    .TE(\mprj_logic1[286] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[84])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[85]  (
    .A(_313_),
    .TE(\mprj_logic1[287] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[85])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[86]  (
    .A(_314_),
    .TE(\mprj_logic1[288] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[86])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[87]  (
    .A(_315_),
    .TE(\mprj_logic1[289] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[87])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[88]  (
    .A(_316_),
    .TE(\mprj_logic1[290] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[88])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[89]  (
    .A(_317_),
    .TE(\mprj_logic1[291] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[89])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[8]  (
    .A(_318_),
    .TE(\mprj_logic1[210] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[8])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[90]  (
    .A(_319_),
    .TE(\mprj_logic1[292] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[90])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[91]  (
    .A(_320_),
    .TE(\mprj_logic1[293] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[91])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[92]  (
    .A(_321_),
    .TE(\mprj_logic1[294] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[92])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[93]  (
    .A(_322_),
    .TE(\mprj_logic1[295] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[93])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[94]  (
    .A(_323_),
    .TE(\mprj_logic1[296] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[94])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[95]  (
    .A(_324_),
    .TE(\mprj_logic1[297] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[95])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[96]  (
    .A(_325_),
    .TE(\mprj_logic1[298] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[96])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[97]  (
    .A(_326_),
    .TE(\mprj_logic1[299] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[97])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[98]  (
    .A(_327_),
    .TE(\mprj_logic1[300] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[98])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[99]  (
    .A(_328_),
    .TE(\mprj_logic1[301] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[99])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[9]  (
    .A(_329_),
    .TE(\mprj_logic1[211] ),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .Z(la_oen_core[9])
  );
endmodule
