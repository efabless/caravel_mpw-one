magic
tech sky130A
timestamp 1623348513
<< obsli1 >>
rect 0 2272 5573 2305
rect 0 33 14 2258
rect 28 47 42 2272
rect 56 33 70 2258
rect 84 47 98 2272
rect 112 33 126 2258
rect 140 47 154 2272
rect 168 33 182 2258
rect 196 47 210 2272
rect 224 33 238 2258
rect 252 47 266 2272
rect 280 33 294 2258
rect 308 47 322 2272
rect 336 33 350 2258
rect 364 47 378 2272
rect 392 33 406 2258
rect 420 47 434 2272
rect 448 33 462 2258
rect 476 47 490 2272
rect 504 33 518 2258
rect 532 47 546 2272
rect 560 33 574 2258
rect 588 47 602 2272
rect 616 33 630 2258
rect 644 47 658 2272
rect 672 33 686 2258
rect 700 47 714 2272
rect 728 33 742 2258
rect 756 47 770 2272
rect 784 33 798 2258
rect 812 47 826 2272
rect 840 33 854 2258
rect 868 47 882 2272
rect 896 33 910 2258
rect 924 47 938 2272
rect 952 33 966 2258
rect 980 47 994 2272
rect 1008 33 1022 2258
rect 1036 47 1050 2272
rect 1064 33 1078 2258
rect 1092 47 1106 2272
rect 1120 33 1134 2258
rect 1148 47 1162 2272
rect 1176 33 1190 2258
rect 1204 47 1218 2272
rect 1232 33 1246 2258
rect 1260 47 1274 2272
rect 1288 33 1302 2258
rect 1316 47 1330 2272
rect 1344 33 1358 2258
rect 1372 47 1386 2272
rect 1400 33 1414 2258
rect 1428 47 1442 2272
rect 1456 33 1470 2258
rect 1484 47 1498 2272
rect 1512 33 1526 2258
rect 1540 47 1554 2272
rect 1568 33 1582 2258
rect 1596 47 1610 2272
rect 1624 33 1638 2258
rect 1652 47 1666 2272
rect 1680 33 1694 2258
rect 1708 47 1722 2272
rect 1736 33 1750 2258
rect 1764 47 1778 2272
rect 1792 33 1806 2258
rect 1820 47 1834 2272
rect 1848 33 1862 2258
rect 1876 47 1890 2272
rect 1904 33 1918 2258
rect 1932 47 1946 2272
rect 1960 33 1974 2258
rect 1988 47 2002 2272
rect 2016 33 2030 2258
rect 2044 47 2058 2272
rect 2072 33 2086 2258
rect 2100 47 2114 2272
rect 2128 33 2142 2258
rect 2156 47 2170 2272
rect 2184 33 2198 2258
rect 2212 47 2226 2272
rect 2240 33 2254 2258
rect 2268 47 2282 2272
rect 2296 33 2310 2258
rect 2324 47 2338 2272
rect 2352 33 2366 2258
rect 2380 47 2394 2272
rect 2408 33 2422 2258
rect 2436 47 2450 2272
rect 2464 33 2478 2258
rect 2492 47 2506 2272
rect 2520 33 2534 2258
rect 2548 47 2562 2272
rect 2576 33 2590 2258
rect 2604 47 2618 2272
rect 2632 33 2646 2258
rect 2660 47 2674 2272
rect 2688 33 2702 2258
rect 2716 47 2730 2272
rect 2744 33 2758 2258
rect 2772 47 2786 2272
rect 2800 33 2814 2258
rect 2828 47 2842 2272
rect 2856 33 2870 2258
rect 2884 47 2898 2272
rect 2912 33 2926 2258
rect 2940 47 2954 2272
rect 2968 33 2982 2258
rect 2996 47 3010 2272
rect 3024 33 3038 2258
rect 3052 47 3066 2272
rect 3080 33 3094 2258
rect 3108 47 3122 2272
rect 3136 33 3150 2258
rect 3164 47 3178 2272
rect 3192 33 3206 2258
rect 3220 47 3234 2272
rect 3248 33 3262 2258
rect 3276 47 3290 2272
rect 3304 33 3318 2258
rect 3332 47 3346 2272
rect 3360 33 3374 2258
rect 3388 47 3402 2272
rect 3416 33 3430 2258
rect 3444 47 3458 2272
rect 3472 33 3486 2258
rect 3500 47 3514 2272
rect 3528 33 3542 2258
rect 3556 47 3570 2272
rect 3584 33 3598 2258
rect 3612 47 3626 2272
rect 3640 33 3654 2258
rect 3668 47 3682 2272
rect 3696 33 3710 2258
rect 3724 47 3738 2272
rect 3752 33 3766 2258
rect 3780 47 3794 2272
rect 3808 33 3822 2258
rect 3836 47 3850 2272
rect 3864 33 3878 2258
rect 3892 47 3906 2272
rect 3920 33 3934 2258
rect 3948 47 3962 2272
rect 3976 33 3990 2258
rect 4004 47 4018 2272
rect 4032 33 4046 2258
rect 4060 47 4074 2272
rect 4088 33 4102 2258
rect 4116 47 4130 2272
rect 4144 33 4158 2258
rect 4172 47 4186 2272
rect 4200 33 4214 2258
rect 4228 47 4242 2272
rect 4256 33 4270 2258
rect 4284 47 4298 2272
rect 4312 33 4326 2258
rect 4340 47 4354 2272
rect 4368 33 4382 2258
rect 4396 47 4410 2272
rect 4424 33 4438 2258
rect 4452 47 4466 2272
rect 4480 33 4494 2258
rect 4508 47 4522 2272
rect 4536 33 4550 2258
rect 4564 47 4578 2272
rect 4592 33 4606 2258
rect 4620 47 4634 2272
rect 4648 33 4662 2258
rect 4676 47 4690 2272
rect 4704 33 4718 2258
rect 4732 47 4746 2272
rect 4760 33 4774 2258
rect 4788 47 4802 2272
rect 4816 33 4830 2258
rect 4844 47 4858 2272
rect 4872 33 4886 2258
rect 4900 47 4914 2272
rect 4928 33 4942 2258
rect 4956 47 4970 2272
rect 4984 33 4998 2258
rect 5012 47 5026 2272
rect 5040 33 5054 2258
rect 5068 47 5082 2272
rect 5096 33 5110 2258
rect 5124 47 5138 2272
rect 5152 33 5166 2258
rect 5180 47 5194 2272
rect 5208 33 5222 2258
rect 5236 47 5250 2272
rect 5264 33 5278 2258
rect 5292 47 5306 2272
rect 5320 33 5334 2258
rect 5348 47 5362 2272
rect 5376 33 5390 2258
rect 5404 47 5418 2272
rect 5432 33 5446 2258
rect 5460 47 5474 2272
rect 5488 33 5502 2258
rect 5516 47 5530 2272
rect 5544 33 5573 2258
rect 0 0 5573 33
<< obsm1 >>
rect 0 2272 5573 2305
rect 0 47 14 2272
rect 28 33 42 2258
rect 56 47 70 2272
rect 84 33 98 2258
rect 112 47 126 2272
rect 140 33 154 2258
rect 168 47 182 2272
rect 196 33 210 2258
rect 224 47 238 2272
rect 252 33 266 2258
rect 280 47 294 2272
rect 308 33 322 2258
rect 336 47 350 2272
rect 364 33 378 2258
rect 392 47 406 2272
rect 420 33 434 2258
rect 448 47 462 2272
rect 476 33 490 2258
rect 504 47 518 2272
rect 532 33 546 2258
rect 560 47 574 2272
rect 588 33 602 2258
rect 616 47 630 2272
rect 644 33 658 2258
rect 672 47 686 2272
rect 700 33 714 2258
rect 728 47 742 2272
rect 756 33 770 2258
rect 784 47 798 2272
rect 812 33 826 2258
rect 840 47 854 2272
rect 868 33 882 2258
rect 896 47 910 2272
rect 924 33 938 2258
rect 952 47 966 2272
rect 980 33 994 2258
rect 1008 47 1022 2272
rect 1036 33 1050 2258
rect 1064 47 1078 2272
rect 1092 33 1106 2258
rect 1120 47 1134 2272
rect 1148 33 1162 2258
rect 1176 47 1190 2272
rect 1204 33 1218 2258
rect 1232 47 1246 2272
rect 1260 33 1274 2258
rect 1288 47 1302 2272
rect 1316 33 1330 2258
rect 1344 47 1358 2272
rect 1372 33 1386 2258
rect 1400 47 1414 2272
rect 1428 33 1442 2258
rect 1456 47 1470 2272
rect 1484 33 1498 2258
rect 1512 47 1526 2272
rect 1540 33 1554 2258
rect 1568 47 1582 2272
rect 1596 33 1610 2258
rect 1624 47 1638 2272
rect 1652 33 1666 2258
rect 1680 47 1694 2272
rect 1708 33 1722 2258
rect 1736 47 1750 2272
rect 1764 33 1778 2258
rect 1792 47 1806 2272
rect 1820 33 1834 2258
rect 1848 47 1862 2272
rect 1876 33 1890 2258
rect 1904 47 1918 2272
rect 1932 33 1946 2258
rect 1960 47 1974 2272
rect 1988 33 2002 2258
rect 2016 47 2030 2272
rect 2044 33 2058 2258
rect 2072 47 2086 2272
rect 2100 33 2114 2258
rect 2128 47 2142 2272
rect 2156 33 2170 2258
rect 2184 47 2198 2272
rect 2212 33 2226 2258
rect 2240 47 2254 2272
rect 2268 33 2282 2258
rect 2296 47 2310 2272
rect 2324 33 2338 2258
rect 2352 47 2366 2272
rect 2380 33 2394 2258
rect 2408 47 2422 2272
rect 2436 33 2450 2258
rect 2464 47 2478 2272
rect 2492 33 2506 2258
rect 2520 47 2534 2272
rect 2548 33 2562 2258
rect 2576 47 2590 2272
rect 2604 33 2618 2258
rect 2632 47 2646 2272
rect 2660 33 2674 2258
rect 2688 47 2702 2272
rect 2716 33 2730 2258
rect 2744 47 2758 2272
rect 2772 33 2786 2258
rect 2800 47 2814 2272
rect 2828 33 2842 2258
rect 2856 47 2870 2272
rect 2884 33 2898 2258
rect 2912 47 2926 2272
rect 2940 33 2954 2258
rect 2968 47 2982 2272
rect 2996 33 3010 2258
rect 3024 47 3038 2272
rect 3052 33 3066 2258
rect 3080 47 3094 2272
rect 3108 33 3122 2258
rect 3136 47 3150 2272
rect 3164 33 3178 2258
rect 3192 47 3206 2272
rect 3220 33 3234 2258
rect 3248 47 3262 2272
rect 3276 33 3290 2258
rect 3304 47 3318 2272
rect 3332 33 3346 2258
rect 3360 47 3374 2272
rect 3388 33 3402 2258
rect 3416 47 3430 2272
rect 3444 33 3458 2258
rect 3472 47 3486 2272
rect 3500 33 3514 2258
rect 3528 47 3542 2272
rect 3556 33 3570 2258
rect 3584 47 3598 2272
rect 3612 33 3626 2258
rect 3640 47 3654 2272
rect 3668 33 3682 2258
rect 3696 47 3710 2272
rect 3724 33 3738 2258
rect 3752 47 3766 2272
rect 3780 33 3794 2258
rect 3808 47 3822 2272
rect 3836 33 3850 2258
rect 3864 47 3878 2272
rect 3892 33 3906 2258
rect 3920 47 3934 2272
rect 3948 33 3962 2258
rect 3976 47 3990 2272
rect 4004 33 4018 2258
rect 4032 47 4046 2272
rect 4060 33 4074 2258
rect 4088 47 4102 2272
rect 4116 33 4130 2258
rect 4144 47 4158 2272
rect 4172 33 4186 2258
rect 4200 47 4214 2272
rect 4228 33 4242 2258
rect 4256 47 4270 2272
rect 4284 33 4298 2258
rect 4312 47 4326 2272
rect 4340 33 4354 2258
rect 4368 47 4382 2272
rect 4396 33 4410 2258
rect 4424 47 4438 2272
rect 4452 33 4466 2258
rect 4480 47 4494 2272
rect 4508 33 4522 2258
rect 4536 47 4550 2272
rect 4564 33 4578 2258
rect 4592 47 4606 2272
rect 4620 33 4634 2258
rect 4648 47 4662 2272
rect 4676 33 4690 2258
rect 4704 47 4718 2272
rect 4732 33 4746 2258
rect 4760 47 4774 2272
rect 4788 33 4802 2258
rect 4816 47 4830 2272
rect 4844 33 4858 2258
rect 4872 47 4886 2272
rect 4900 33 4914 2258
rect 4928 47 4942 2272
rect 4956 33 4970 2258
rect 4984 47 4998 2272
rect 5012 33 5026 2258
rect 5040 47 5054 2272
rect 5068 33 5082 2258
rect 5096 47 5110 2272
rect 5124 33 5138 2258
rect 5152 47 5166 2272
rect 5180 33 5194 2258
rect 5208 47 5222 2272
rect 5236 33 5250 2258
rect 5264 47 5278 2272
rect 5292 33 5306 2258
rect 5320 47 5334 2272
rect 5348 33 5362 2258
rect 5376 47 5390 2272
rect 5404 33 5418 2258
rect 5432 47 5446 2272
rect 5460 33 5474 2258
rect 5488 47 5502 2272
rect 5516 33 5530 2258
rect 5544 47 5573 2272
rect 0 0 5573 33
<< obsm2 >>
rect 0 33 14 2305
rect 28 2272 98 2305
rect 28 47 42 2272
rect 56 33 70 2258
rect 0 0 70 33
rect 84 0 98 2272
rect 112 33 126 2305
rect 140 2272 210 2305
rect 140 47 154 2272
rect 168 33 182 2258
rect 112 0 182 33
rect 196 0 210 2272
rect 224 33 238 2305
rect 252 2272 322 2305
rect 252 47 266 2272
rect 280 33 294 2258
rect 224 0 294 33
rect 308 0 322 2272
rect 336 33 350 2305
rect 364 2272 434 2305
rect 364 47 378 2272
rect 392 33 406 2258
rect 336 0 406 33
rect 420 0 434 2272
rect 448 33 462 2305
rect 476 2272 546 2305
rect 476 47 490 2272
rect 504 33 518 2258
rect 448 0 518 33
rect 532 0 546 2272
rect 560 33 574 2305
rect 588 2272 658 2305
rect 588 47 602 2272
rect 616 33 630 2258
rect 560 0 630 33
rect 644 0 658 2272
rect 672 33 686 2305
rect 700 2272 770 2305
rect 700 47 714 2272
rect 728 33 742 2258
rect 672 0 742 33
rect 756 0 770 2272
rect 784 33 798 2305
rect 812 2272 882 2305
rect 812 47 826 2272
rect 840 33 854 2258
rect 784 0 854 33
rect 868 0 882 2272
rect 896 33 910 2305
rect 924 2272 994 2305
rect 924 47 938 2272
rect 952 33 966 2258
rect 896 0 966 33
rect 980 0 994 2272
rect 1008 33 1022 2305
rect 1036 2272 1106 2305
rect 1036 47 1050 2272
rect 1064 33 1078 2258
rect 1008 0 1078 33
rect 1092 0 1106 2272
rect 1120 33 1134 2305
rect 1148 2272 1218 2305
rect 1148 47 1162 2272
rect 1176 33 1190 2258
rect 1120 0 1190 33
rect 1204 0 1218 2272
rect 1232 33 1246 2305
rect 1260 2272 1330 2305
rect 1260 47 1274 2272
rect 1288 33 1302 2258
rect 1232 0 1302 33
rect 1316 0 1330 2272
rect 1344 33 1358 2305
rect 1372 2272 1442 2305
rect 1372 47 1386 2272
rect 1400 33 1414 2258
rect 1344 0 1414 33
rect 1428 0 1442 2272
rect 1456 33 1470 2305
rect 1484 2272 1554 2305
rect 1484 47 1498 2272
rect 1512 33 1526 2258
rect 1456 0 1526 33
rect 1540 0 1554 2272
rect 1568 33 1582 2305
rect 1596 2272 1666 2305
rect 1596 47 1610 2272
rect 1624 33 1638 2258
rect 1568 0 1638 33
rect 1652 0 1666 2272
rect 1680 33 1694 2305
rect 1708 2272 1778 2305
rect 1708 47 1722 2272
rect 1736 33 1750 2258
rect 1680 0 1750 33
rect 1764 0 1778 2272
rect 1792 33 1806 2305
rect 1820 2272 1890 2305
rect 1820 47 1834 2272
rect 1848 33 1862 2258
rect 1792 0 1862 33
rect 1876 0 1890 2272
rect 1904 33 1918 2305
rect 1932 2272 2002 2305
rect 1932 47 1946 2272
rect 1960 33 1974 2258
rect 1904 0 1974 33
rect 1988 0 2002 2272
rect 2016 33 2030 2305
rect 2044 2272 2114 2305
rect 2044 47 2058 2272
rect 2072 33 2086 2258
rect 2016 0 2086 33
rect 2100 0 2114 2272
rect 2128 33 2142 2305
rect 2156 2272 2226 2305
rect 2156 47 2170 2272
rect 2184 33 2198 2258
rect 2128 0 2198 33
rect 2212 0 2226 2272
rect 2240 33 2254 2305
rect 2268 2272 2338 2305
rect 2268 47 2282 2272
rect 2296 33 2310 2258
rect 2240 0 2310 33
rect 2324 0 2338 2272
rect 2352 33 2366 2305
rect 2380 2272 2450 2305
rect 2380 47 2394 2272
rect 2408 33 2422 2258
rect 2352 0 2422 33
rect 2436 0 2450 2272
rect 2464 33 2478 2305
rect 2492 2272 2562 2305
rect 2492 47 2506 2272
rect 2520 33 2534 2258
rect 2464 0 2534 33
rect 2548 0 2562 2272
rect 2576 33 2590 2305
rect 2604 2272 2674 2305
rect 2604 47 2618 2272
rect 2632 33 2646 2258
rect 2576 0 2646 33
rect 2660 0 2674 2272
rect 2688 33 2702 2305
rect 2716 2272 2786 2305
rect 2716 47 2730 2272
rect 2744 33 2758 2258
rect 2688 0 2758 33
rect 2772 0 2786 2272
rect 2800 33 2814 2305
rect 2828 2272 2898 2305
rect 2828 47 2842 2272
rect 2856 33 2870 2258
rect 2800 0 2870 33
rect 2884 0 2898 2272
rect 2912 33 2926 2305
rect 2940 2272 3010 2305
rect 2940 47 2954 2272
rect 2968 33 2982 2258
rect 2912 0 2982 33
rect 2996 0 3010 2272
rect 3024 33 3038 2305
rect 3052 2272 3122 2305
rect 3052 47 3066 2272
rect 3080 33 3094 2258
rect 3024 0 3094 33
rect 3108 0 3122 2272
rect 3136 33 3150 2305
rect 3164 2272 3234 2305
rect 3164 47 3178 2272
rect 3192 33 3206 2258
rect 3136 0 3206 33
rect 3220 0 3234 2272
rect 3248 33 3262 2305
rect 3276 2272 3346 2305
rect 3276 47 3290 2272
rect 3304 33 3318 2258
rect 3248 0 3318 33
rect 3332 0 3346 2272
rect 3360 33 3374 2305
rect 3388 2272 3458 2305
rect 3388 47 3402 2272
rect 3416 33 3430 2258
rect 3360 0 3430 33
rect 3444 0 3458 2272
rect 3472 33 3486 2305
rect 3500 2272 3570 2305
rect 3500 47 3514 2272
rect 3528 33 3542 2258
rect 3472 0 3542 33
rect 3556 0 3570 2272
rect 3584 33 3598 2305
rect 3612 2272 3682 2305
rect 3612 47 3626 2272
rect 3640 33 3654 2258
rect 3584 0 3654 33
rect 3668 0 3682 2272
rect 3696 33 3710 2305
rect 3724 2272 3794 2305
rect 3724 47 3738 2272
rect 3752 33 3766 2258
rect 3696 0 3766 33
rect 3780 0 3794 2272
rect 3808 33 3822 2305
rect 3836 2272 3906 2305
rect 3836 47 3850 2272
rect 3864 33 3878 2258
rect 3808 0 3878 33
rect 3892 0 3906 2272
rect 3920 33 3934 2305
rect 3948 2272 4018 2305
rect 3948 47 3962 2272
rect 3976 33 3990 2258
rect 3920 0 3990 33
rect 4004 0 4018 2272
rect 4032 33 4046 2305
rect 4060 2272 4130 2305
rect 4060 47 4074 2272
rect 4088 33 4102 2258
rect 4032 0 4102 33
rect 4116 0 4130 2272
rect 4144 33 4158 2305
rect 4172 2272 4242 2305
rect 4172 47 4186 2272
rect 4200 33 4214 2258
rect 4144 0 4214 33
rect 4228 0 4242 2272
rect 4256 33 4270 2305
rect 4284 2272 4354 2305
rect 4284 47 4298 2272
rect 4312 33 4326 2258
rect 4256 0 4326 33
rect 4340 0 4354 2272
rect 4368 33 4382 2305
rect 4396 2272 4466 2305
rect 4396 47 4410 2272
rect 4424 33 4438 2258
rect 4368 0 4438 33
rect 4452 0 4466 2272
rect 4480 33 4494 2305
rect 4508 2272 4578 2305
rect 4508 47 4522 2272
rect 4536 33 4550 2258
rect 4480 0 4550 33
rect 4564 0 4578 2272
rect 4592 33 4606 2305
rect 4620 2272 4690 2305
rect 4620 47 4634 2272
rect 4648 33 4662 2258
rect 4592 0 4662 33
rect 4676 0 4690 2272
rect 4704 33 4718 2305
rect 4732 2272 4802 2305
rect 4732 47 4746 2272
rect 4760 33 4774 2258
rect 4704 0 4774 33
rect 4788 0 4802 2272
rect 4816 33 4830 2305
rect 4844 2272 4914 2305
rect 4844 47 4858 2272
rect 4872 33 4886 2258
rect 4816 0 4886 33
rect 4900 0 4914 2272
rect 4928 33 4942 2305
rect 4956 2272 5026 2305
rect 4956 47 4970 2272
rect 4984 33 4998 2258
rect 4928 0 4998 33
rect 5012 0 5026 2272
rect 5040 33 5054 2305
rect 5068 2272 5138 2305
rect 5068 47 5082 2272
rect 5096 33 5110 2258
rect 5040 0 5110 33
rect 5124 0 5138 2272
rect 5152 33 5166 2305
rect 5180 2272 5250 2305
rect 5180 47 5194 2272
rect 5208 33 5222 2258
rect 5152 0 5222 33
rect 5236 0 5250 2272
rect 5264 33 5278 2305
rect 5292 2272 5362 2305
rect 5292 47 5306 2272
rect 5320 33 5334 2258
rect 5264 0 5334 33
rect 5348 0 5362 2272
rect 5376 33 5390 2305
rect 5404 2272 5573 2305
rect 5404 47 5418 2272
rect 5432 33 5446 2258
rect 5376 0 5446 33
rect 5460 0 5474 2272
rect 5488 33 5502 2258
rect 5516 47 5530 2272
rect 5544 33 5573 2258
rect 5488 0 5573 33
<< obsm3 >>
rect 0 2272 5573 2305
rect 0 63 30 2272
rect 60 33 90 2242
rect 120 63 150 2272
rect 180 33 210 2242
rect 240 63 270 2272
rect 300 33 330 2242
rect 360 63 390 2272
rect 420 33 450 2242
rect 480 63 510 2272
rect 540 33 570 2242
rect 600 63 630 2272
rect 660 33 690 2242
rect 720 63 750 2272
rect 780 33 810 2242
rect 840 63 870 2272
rect 900 33 930 2242
rect 960 63 990 2272
rect 1020 33 1050 2242
rect 1080 63 1110 2272
rect 1140 33 1170 2242
rect 1200 63 1230 2272
rect 1260 33 1290 2242
rect 1320 63 1350 2272
rect 1380 33 1410 2242
rect 1440 63 1470 2272
rect 1500 33 1530 2242
rect 1560 63 1590 2272
rect 1620 33 1650 2242
rect 1680 63 1710 2272
rect 1740 33 1770 2242
rect 1800 63 1830 2272
rect 1860 33 1890 2242
rect 1920 63 1950 2272
rect 1980 33 2010 2242
rect 2040 63 2070 2272
rect 2100 33 2130 2242
rect 2160 63 2190 2272
rect 2220 33 2250 2242
rect 2280 63 2310 2272
rect 2340 33 2370 2242
rect 2400 63 2430 2272
rect 2460 33 2490 2242
rect 2520 63 2550 2272
rect 2580 33 2610 2242
rect 2640 63 2670 2272
rect 2700 33 2730 2242
rect 2760 63 2790 2272
rect 2820 33 2850 2242
rect 2880 63 2910 2272
rect 2940 33 2970 2242
rect 3000 63 3030 2272
rect 3060 33 3090 2242
rect 3120 63 3150 2272
rect 3180 33 3210 2242
rect 3240 63 3270 2272
rect 3300 33 3330 2242
rect 3360 63 3390 2272
rect 3420 33 3450 2242
rect 3480 63 3510 2272
rect 3540 33 3570 2242
rect 3600 63 3630 2272
rect 3660 33 3690 2242
rect 3720 63 3750 2272
rect 3780 33 3810 2242
rect 3840 63 3870 2272
rect 3900 33 3930 2242
rect 3960 63 3990 2272
rect 4020 33 4050 2242
rect 4080 63 4110 2272
rect 4140 33 4170 2242
rect 4200 63 4230 2272
rect 4260 33 4290 2242
rect 4320 63 4350 2272
rect 4380 33 4410 2242
rect 4440 63 4470 2272
rect 4500 33 4530 2242
rect 4560 63 4590 2272
rect 4620 33 4650 2242
rect 4680 63 4710 2272
rect 4740 33 4770 2242
rect 4800 63 4830 2272
rect 4860 33 4890 2242
rect 4920 63 4950 2272
rect 4980 33 5010 2242
rect 5040 63 5070 2272
rect 5100 33 5130 2242
rect 5160 63 5190 2272
rect 5220 33 5250 2242
rect 5280 63 5310 2272
rect 5340 33 5370 2242
rect 5400 63 5430 2272
rect 5460 33 5490 2242
rect 5520 63 5573 2272
rect 0 0 5573 33
<< obsm4 >>
rect 0 2272 5573 2305
rect 0 33 30 2242
rect 60 2135 210 2272
rect 60 63 90 2135
rect 120 170 150 2105
rect 180 200 210 2135
rect 240 170 270 2242
rect 120 33 270 170
rect 300 63 330 2272
rect 360 33 390 2242
rect 420 63 450 2272
rect 480 33 510 2242
rect 540 63 570 2272
rect 600 33 630 2242
rect 660 63 690 2272
rect 720 33 750 2242
rect 780 2135 930 2272
rect 780 63 810 2135
rect 840 170 870 2105
rect 900 200 930 2135
rect 960 170 990 2242
rect 840 33 990 170
rect 1020 63 1050 2272
rect 1080 33 1110 2242
rect 1140 63 1170 2272
rect 1200 33 1230 2242
rect 1260 63 1290 2272
rect 1320 33 1350 2242
rect 1380 63 1410 2272
rect 1440 33 1470 2242
rect 1500 2135 1650 2272
rect 1500 63 1530 2135
rect 1560 170 1590 2105
rect 1620 200 1650 2135
rect 1680 170 1710 2242
rect 1560 33 1710 170
rect 1740 63 1770 2272
rect 1800 33 1830 2242
rect 1860 63 1890 2272
rect 1920 33 1950 2242
rect 1980 63 2010 2272
rect 2040 33 2070 2242
rect 2100 63 2130 2272
rect 2160 33 2190 2242
rect 2220 2135 2370 2272
rect 2220 63 2250 2135
rect 2280 170 2310 2105
rect 2340 200 2370 2135
rect 2400 170 2430 2242
rect 2280 33 2430 170
rect 2460 63 2490 2272
rect 2520 33 2550 2242
rect 2580 63 2610 2272
rect 2640 33 2670 2242
rect 2700 63 2730 2272
rect 2760 33 2790 2242
rect 2820 63 2850 2272
rect 2880 33 2910 2242
rect 2940 2135 3090 2272
rect 2940 63 2970 2135
rect 3000 170 3030 2105
rect 3060 200 3090 2135
rect 3120 170 3150 2242
rect 3000 33 3150 170
rect 3180 63 3210 2272
rect 3240 33 3270 2242
rect 3300 63 3330 2272
rect 3360 33 3390 2242
rect 3420 63 3450 2272
rect 3480 33 3510 2242
rect 3540 63 3570 2272
rect 3600 33 3630 2242
rect 3660 2135 3810 2272
rect 3660 63 3690 2135
rect 3720 170 3750 2105
rect 3780 200 3810 2135
rect 3840 170 3870 2242
rect 3720 33 3870 170
rect 3900 63 3930 2272
rect 3960 33 3990 2242
rect 4020 63 4050 2272
rect 4080 33 4110 2242
rect 4140 63 4170 2272
rect 4200 33 4230 2242
rect 4260 63 4290 2272
rect 4320 33 4350 2242
rect 4380 2135 4530 2272
rect 4380 63 4410 2135
rect 4440 170 4470 2105
rect 4500 200 4530 2135
rect 4560 170 4590 2242
rect 4440 33 4590 170
rect 4620 63 4650 2272
rect 4680 33 4710 2242
rect 4740 63 4770 2272
rect 4800 33 4830 2242
rect 4860 63 4890 2272
rect 4920 33 4950 2242
rect 4980 63 5010 2272
rect 5040 33 5070 2242
rect 5100 2135 5250 2272
rect 5100 63 5130 2135
rect 5160 170 5190 2105
rect 5220 200 5250 2135
rect 5280 170 5310 2242
rect 5160 33 5310 170
rect 5340 63 5370 2272
rect 5400 33 5430 2242
rect 5460 63 5490 2272
rect 5520 33 5573 2242
rect 0 0 5573 33
<< obsm5 >>
rect 0 2105 5493 2265
rect 0 360 160 2105
rect 320 200 480 1945
rect 640 360 800 2105
rect 960 200 1120 1945
rect 1280 360 1440 2105
rect 1600 200 1760 1945
rect 1920 360 2080 2105
rect 2240 200 2400 1945
rect 2560 360 2720 2105
rect 2880 200 3040 1945
rect 3200 360 3360 2105
rect 3520 200 3680 1945
rect 3840 360 4000 2105
rect 4160 200 4320 1945
rect 4480 360 4640 2105
rect 4800 200 4960 1945
rect 5120 360 5493 2105
rect 0 40 5493 200
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 5573 2305
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 4338416
string GDS_START 4182380
<< end >>
