magic
tech sky130A
magscale 1 2
timestamp 1624446551
<< locali >>
rect 5273 96815 5307 97597
rect 6561 96951 6595 97189
rect 6837 96747 6871 97801
rect 15577 97325 15945 97359
rect 6929 97257 7021 97291
rect 6745 96679 6779 96713
rect 6929 96679 6963 97257
rect 15577 97019 15611 97325
rect 22879 97257 23063 97291
rect 15669 97019 15703 97189
rect 22017 97019 22051 97189
rect 6745 96645 6963 96679
rect 23029 96679 23063 97257
rect 5365 95863 5399 96441
rect 5273 95523 5307 95829
rect 8493 95659 8527 96373
rect 39681 96271 39715 96509
rect 76757 96475 76791 96645
rect 80161 96475 80195 96713
rect 82461 96617 82495 97393
rect 82093 96583 82495 96617
rect 82093 96475 82127 96583
rect 8585 95727 8619 95829
rect 74549 95251 74583 96101
rect 74641 95115 74675 96441
rect 74549 95081 74675 95115
rect 74549 94775 74583 95081
rect 74641 94299 74675 94877
rect 74825 94639 74859 94741
rect 75009 94707 75043 96237
rect 76573 94979 76607 96237
rect 76665 95727 76699 96237
rect 80253 96067 80287 96101
rect 76757 95727 76791 95965
rect 79241 95795 79275 96033
rect 79149 95251 79183 95761
rect 79333 95591 79367 96033
rect 79977 96033 80287 96067
rect 79977 95795 80011 96033
rect 80345 95999 80379 96441
rect 80287 95965 80379 95999
rect 79919 95693 80069 95727
rect 79425 95183 79459 95557
rect 80161 95455 80195 95761
rect 80103 95421 80195 95455
rect 79977 95353 80345 95387
rect 79977 95319 80011 95353
rect 80069 95285 80437 95319
rect 74583 94265 74675 94299
rect 76205 94231 76239 94741
rect 76481 94639 76515 94945
rect 78321 94843 78355 95149
rect 76389 94163 76423 94605
rect 79241 94231 79275 94401
rect 79333 94299 79367 94401
rect 79425 94231 79459 94265
rect 79241 94197 79459 94231
rect 79517 94163 79551 95149
rect 80069 94979 80103 95285
rect 80069 94503 80103 94741
rect 80345 94707 80379 95217
rect 82277 94911 82311 96101
rect 82553 94979 82587 99161
rect 82645 96271 82679 97529
rect 82495 94945 82587 94979
rect 82277 94877 82679 94911
rect 80195 94673 80379 94707
rect 80437 94571 80471 94673
rect 82461 94571 82495 94741
rect 80437 94537 80529 94571
rect 82553 94503 82587 94537
rect 80069 94469 82587 94503
rect 79183 94129 79551 94163
rect 76239 94061 76423 94095
rect 76389 94027 76423 94061
rect 5273 90423 5307 93857
rect 78229 93517 78597 93551
rect 78229 93415 78263 93517
rect 77401 93279 77435 93381
rect 78413 93347 78447 93449
rect 79333 93415 79367 93653
rect 79241 93279 79275 93381
rect 78229 93245 78631 93279
rect 79241 93245 79609 93279
rect 78229 93211 78263 93245
rect 78321 93075 78355 93177
rect 78413 92939 78447 93041
rect 78597 93007 78631 93245
rect 82369 92871 82403 93041
rect 82277 92803 82311 92837
rect 82277 92769 82495 92803
rect 82461 92667 82495 92769
rect 82645 91783 82679 94877
rect 82737 94843 82771 98277
rect 82829 96135 82863 97597
rect 82921 96747 82955 104261
rect 83013 97291 83047 98889
rect 83473 97359 83507 104329
rect 83473 97325 83565 97359
rect 82829 92123 82863 93313
rect 82921 92327 82955 95693
rect 83013 92395 83047 95489
rect 83473 93619 83507 97325
rect 83657 96883 83691 98005
rect 84025 97087 84059 105689
rect 84853 97495 84887 97801
rect 84025 96815 84059 97053
rect 83657 3723 83691 4301
rect 6745 3111 6779 3417
rect 6837 3179 6871 3553
rect 15151 3213 15393 3247
rect 6837 3145 6929 3179
rect 15059 3145 15485 3179
rect 15151 3077 15393 3111
rect 82461 2839 82495 3553
rect 82403 2805 82495 2839
rect 82553 2703 82587 3621
rect 83105 3043 83139 3485
rect 83565 2771 83599 3213
rect 83105 1751 83139 2533
rect 83197 2431 83231 2533
rect 83013 1615 83047 1717
rect 83013 1581 83289 1615
<< viali >>
rect 85037 187357 85071 187391
rect 84669 187221 84703 187255
rect 84669 186337 84703 186371
rect 4813 182937 4847 182971
rect 4813 181849 4847 181883
rect 4721 180149 4755 180183
rect 84485 179605 84519 179639
rect 4721 179061 4755 179095
rect 4721 176885 4755 176919
rect 4813 176137 4847 176171
rect 4813 174505 4847 174539
rect 84485 167433 84519 167467
rect 84669 162401 84703 162435
rect 85129 162333 85163 162367
rect 84669 161993 84703 162027
rect 84485 160089 84519 160123
rect 84669 153833 84703 153867
rect 84945 141117 84979 141151
rect 84669 141049 84703 141083
rect 85221 140981 85255 141015
rect 84669 125749 84703 125783
rect 84669 124457 84703 124491
rect 84669 123369 84703 123403
rect 84669 120853 84703 120887
rect 84669 120037 84703 120071
rect 84669 118133 84703 118167
rect 84669 117045 84703 117079
rect 4813 116569 4847 116603
rect 4813 114937 4847 114971
rect 4445 105825 4479 105859
rect 84025 105689 84059 105723
rect 83473 104329 83507 104363
rect 82921 104261 82955 104295
rect 82553 99161 82587 99195
rect 4353 98549 4387 98583
rect 4813 98549 4847 98583
rect 3709 98073 3743 98107
rect 4445 98005 4479 98039
rect 4721 98005 4755 98039
rect 6837 97801 6871 97835
rect 3709 97733 3743 97767
rect 4077 97665 4111 97699
rect 4445 97597 4479 97631
rect 5273 97597 5307 97631
rect 2973 97529 3007 97563
rect 3341 97461 3375 97495
rect 4813 97461 4847 97495
rect 2605 97257 2639 97291
rect 3341 97257 3375 97291
rect 3709 97189 3743 97223
rect 4445 97053 4479 97087
rect 2237 96985 2271 97019
rect 2973 96917 3007 96951
rect 4813 96917 4847 96951
rect 6561 97189 6595 97223
rect 6561 96917 6595 96951
rect 5273 96781 5307 96815
rect 82461 97393 82495 97427
rect 15945 97325 15979 97359
rect 6745 96713 6779 96747
rect 6837 96713 6871 96747
rect 7021 97257 7055 97291
rect 22845 97257 22879 97291
rect 15577 96985 15611 97019
rect 15669 97189 15703 97223
rect 15669 96985 15703 97019
rect 22017 97189 22051 97223
rect 22017 96985 22051 97019
rect 80161 96713 80195 96747
rect 23029 96645 23063 96679
rect 76757 96645 76791 96679
rect 4077 96509 4111 96543
rect 39681 96509 39715 96543
rect 4445 96441 4479 96475
rect 5365 96441 5399 96475
rect 3341 96373 3375 96407
rect 3709 96373 3743 96407
rect 4813 96373 4847 96407
rect 3709 96169 3743 96203
rect 4445 95965 4479 95999
rect 4813 95829 4847 95863
rect 5273 95829 5307 95863
rect 5365 95829 5399 95863
rect 8493 96373 8527 96407
rect 4445 95625 4479 95659
rect 39681 96237 39715 96271
rect 74641 96441 74675 96475
rect 76757 96441 76791 96475
rect 80161 96441 80195 96475
rect 80345 96441 80379 96475
rect 82093 96441 82127 96475
rect 74549 96101 74583 96135
rect 8585 95829 8619 95863
rect 8585 95693 8619 95727
rect 8493 95625 8527 95659
rect 5273 95489 5307 95523
rect 4813 95285 4847 95319
rect 74549 95217 74583 95251
rect 75009 96237 75043 96271
rect 74549 94741 74583 94775
rect 74641 94877 74675 94911
rect 74825 94741 74859 94775
rect 76573 96237 76607 96271
rect 76665 96237 76699 96271
rect 80253 96101 80287 96135
rect 79241 96033 79275 96067
rect 76665 95693 76699 95727
rect 76757 95965 76791 95999
rect 76757 95693 76791 95727
rect 79149 95761 79183 95795
rect 79241 95761 79275 95795
rect 79333 96033 79367 96067
rect 80253 95965 80287 95999
rect 82277 96101 82311 96135
rect 79977 95761 80011 95795
rect 80161 95761 80195 95795
rect 79885 95693 79919 95727
rect 80069 95693 80103 95727
rect 79333 95557 79367 95591
rect 79425 95557 79459 95591
rect 79149 95217 79183 95251
rect 80069 95421 80103 95455
rect 80345 95353 80379 95387
rect 79977 95285 80011 95319
rect 80437 95285 80471 95319
rect 76481 94945 76515 94979
rect 76573 94945 76607 94979
rect 78321 95149 78355 95183
rect 79425 95149 79459 95183
rect 79517 95149 79551 95183
rect 75009 94673 75043 94707
rect 76205 94741 76239 94775
rect 74825 94605 74859 94639
rect 74549 94265 74583 94299
rect 78321 94809 78355 94843
rect 76205 94197 76239 94231
rect 76389 94605 76423 94639
rect 76481 94605 76515 94639
rect 79241 94401 79275 94435
rect 79333 94401 79367 94435
rect 79333 94265 79367 94299
rect 79425 94265 79459 94299
rect 80069 94945 80103 94979
rect 80345 95217 80379 95251
rect 80069 94741 80103 94775
rect 82737 98277 82771 98311
rect 82645 97529 82679 97563
rect 82645 96237 82679 96271
rect 82461 94945 82495 94979
rect 82461 94741 82495 94775
rect 80161 94673 80195 94707
rect 80437 94673 80471 94707
rect 80529 94537 80563 94571
rect 82461 94537 82495 94571
rect 82553 94537 82587 94571
rect 76389 94129 76423 94163
rect 79149 94129 79183 94163
rect 76205 94061 76239 94095
rect 76389 93993 76423 94027
rect 5273 93857 5307 93891
rect 79333 93653 79367 93687
rect 78597 93517 78631 93551
rect 77401 93381 77435 93415
rect 78229 93381 78263 93415
rect 78413 93449 78447 93483
rect 78413 93313 78447 93347
rect 79241 93381 79275 93415
rect 79333 93381 79367 93415
rect 77401 93245 77435 93279
rect 79609 93245 79643 93279
rect 78229 93177 78263 93211
rect 78321 93177 78355 93211
rect 78321 93041 78355 93075
rect 78413 93041 78447 93075
rect 78597 92973 78631 93007
rect 82369 93041 82403 93075
rect 78413 92905 78447 92939
rect 82277 92837 82311 92871
rect 82369 92837 82403 92871
rect 82461 92633 82495 92667
rect 82829 97597 82863 97631
rect 83013 98889 83047 98923
rect 83013 97257 83047 97291
rect 83657 98005 83691 98039
rect 83565 97325 83599 97359
rect 82921 96713 82955 96747
rect 82829 96101 82863 96135
rect 82737 94809 82771 94843
rect 82921 95693 82955 95727
rect 82829 93313 82863 93347
rect 83013 95489 83047 95523
rect 83657 96849 83691 96883
rect 84669 98005 84703 98039
rect 84853 97801 84887 97835
rect 85129 97801 85163 97835
rect 84669 97461 84703 97495
rect 84853 97461 84887 97495
rect 84669 97257 84703 97291
rect 84025 97053 84059 97087
rect 85037 97053 85071 97087
rect 85865 97053 85899 97087
rect 85405 96917 85439 96951
rect 84025 96781 84059 96815
rect 84761 96373 84795 96407
rect 85129 96373 85163 96407
rect 84761 95829 84795 95863
rect 83473 93585 83507 93619
rect 84761 93381 84795 93415
rect 85129 93381 85163 93415
rect 83013 92361 83047 92395
rect 82921 92293 82955 92327
rect 82829 92089 82863 92123
rect 84761 92021 84795 92055
rect 82645 91749 82679 91783
rect 5273 90389 5307 90423
rect 4813 89029 4847 89063
rect 4813 88009 4847 88043
rect 4813 86377 4847 86411
rect 4721 85289 4755 85323
rect 4813 83317 4847 83351
rect 4813 82229 4847 82263
rect 4813 80393 4847 80427
rect 4445 57885 4479 57919
rect 4445 49929 4479 49963
rect 84485 39049 84519 39083
rect 84761 31977 84795 32011
rect 84761 30277 84795 30311
rect 84761 29257 84795 29291
rect 84761 27557 84795 27591
rect 84761 26537 84795 26571
rect 84761 24361 84795 24395
rect 84761 23273 84795 23307
rect 4721 22389 4755 22423
rect 4813 20825 4847 20859
rect 84485 17697 84519 17731
rect 84669 14569 84703 14603
rect 85313 13889 85347 13923
rect 84669 13821 84703 13855
rect 4445 10081 4479 10115
rect 4813 4981 4847 5015
rect 4813 4777 4847 4811
rect 4445 4709 4479 4743
rect 83657 4301 83691 4335
rect 3985 4097 4019 4131
rect 4445 4029 4479 4063
rect 3341 3961 3375 3995
rect 3709 3893 3743 3927
rect 4813 3893 4847 3927
rect 84669 4097 84703 4131
rect 3341 3689 3375 3723
rect 4813 3689 4847 3723
rect 83657 3689 83691 3723
rect 84669 3689 84703 3723
rect 85037 3689 85071 3723
rect 85405 3689 85439 3723
rect 4445 3621 4479 3655
rect 82553 3621 82587 3655
rect 6837 3553 6871 3587
rect 3709 3485 3743 3519
rect 2605 3417 2639 3451
rect 6745 3417 6779 3451
rect 2973 3349 3007 3383
rect 2237 3145 2271 3179
rect 3709 3145 3743 3179
rect 4445 3145 4479 3179
rect 82461 3553 82495 3587
rect 15117 3213 15151 3247
rect 15393 3213 15427 3247
rect 6929 3145 6963 3179
rect 15025 3145 15059 3179
rect 15485 3145 15519 3179
rect 2513 3077 2547 3111
rect 4077 3077 4111 3111
rect 6745 3077 6779 3111
rect 15117 3077 15151 3111
rect 15393 3077 15427 3111
rect 2973 2941 3007 2975
rect 3341 2805 3375 2839
rect 4721 2805 4755 2839
rect 82369 2805 82403 2839
rect 83105 3485 83139 3519
rect 83105 3009 83139 3043
rect 83565 3213 83599 3247
rect 85773 3145 85807 3179
rect 84669 3009 84703 3043
rect 85037 2873 85071 2907
rect 85405 2805 85439 2839
rect 83565 2737 83599 2771
rect 82553 2669 82587 2703
rect 3709 2601 3743 2635
rect 3341 2533 3375 2567
rect 83105 2533 83139 2567
rect 4445 2465 4479 2499
rect 2973 2397 3007 2431
rect 2605 2329 2639 2363
rect 4813 2261 4847 2295
rect 83197 2533 83231 2567
rect 83197 2397 83231 2431
rect 85037 2329 85071 2363
rect 84669 2261 84703 2295
rect 83013 1717 83047 1751
rect 83105 1717 83139 1751
rect 83289 1581 83323 1615
<< metal1 >>
rect 1104 189338 5152 189360
rect 1104 189286 1982 189338
rect 2034 189286 2046 189338
rect 2098 189286 2110 189338
rect 2162 189286 2174 189338
rect 2226 189286 5152 189338
rect 1104 189264 5152 189286
rect 84180 189338 90896 189360
rect 84180 189286 85982 189338
rect 86034 189286 86046 189338
rect 86098 189286 86110 189338
rect 86162 189286 86174 189338
rect 86226 189286 89982 189338
rect 90034 189286 90046 189338
rect 90098 189286 90110 189338
rect 90162 189286 90174 189338
rect 90226 189286 90896 189338
rect 84180 189264 90896 189286
rect 75822 189048 75828 189100
rect 75880 189088 75886 189100
rect 84470 189088 84476 189100
rect 75880 189060 84476 189088
rect 75880 189048 75886 189060
rect 84470 189048 84476 189060
rect 84528 189048 84534 189100
rect 1104 188794 5152 188816
rect 1104 188742 3982 188794
rect 4034 188742 4046 188794
rect 4098 188742 4110 188794
rect 4162 188742 4174 188794
rect 4226 188742 5152 188794
rect 1104 188720 5152 188742
rect 84180 188794 90896 188816
rect 84180 188742 87982 188794
rect 88034 188742 88046 188794
rect 88098 188742 88110 188794
rect 88162 188742 88174 188794
rect 88226 188742 90896 188794
rect 84180 188720 90896 188742
rect 1104 188250 5152 188272
rect 1104 188198 1982 188250
rect 2034 188198 2046 188250
rect 2098 188198 2110 188250
rect 2162 188198 2174 188250
rect 2226 188198 5152 188250
rect 1104 188176 5152 188198
rect 84180 188250 90896 188272
rect 84180 188198 85982 188250
rect 86034 188198 86046 188250
rect 86098 188198 86110 188250
rect 86162 188198 86174 188250
rect 86226 188198 89982 188250
rect 90034 188198 90046 188250
rect 90098 188198 90110 188250
rect 90162 188198 90174 188250
rect 90226 188198 90896 188250
rect 84180 188176 90896 188198
rect 1104 187706 5152 187728
rect 1104 187654 3982 187706
rect 4034 187654 4046 187706
rect 4098 187654 4110 187706
rect 4162 187654 4174 187706
rect 4226 187654 5152 187706
rect 1104 187632 5152 187654
rect 84180 187706 90896 187728
rect 84180 187654 87982 187706
rect 88034 187654 88046 187706
rect 88098 187654 88110 187706
rect 88162 187654 88174 187706
rect 88226 187654 90896 187706
rect 84180 187632 90896 187654
rect 79318 187348 79324 187400
rect 79376 187388 79382 187400
rect 85025 187391 85083 187397
rect 85025 187388 85037 187391
rect 79376 187360 85037 187388
rect 79376 187348 79382 187360
rect 85025 187357 85037 187360
rect 85071 187357 85083 187391
rect 85025 187351 85083 187357
rect 84470 187212 84476 187264
rect 84528 187252 84534 187264
rect 84657 187255 84715 187261
rect 84657 187252 84669 187255
rect 84528 187224 84669 187252
rect 84528 187212 84534 187224
rect 84657 187221 84669 187224
rect 84703 187221 84715 187255
rect 84657 187215 84715 187221
rect 1104 187162 5152 187184
rect 1104 187110 1982 187162
rect 2034 187110 2046 187162
rect 2098 187110 2110 187162
rect 2162 187110 2174 187162
rect 2226 187110 5152 187162
rect 1104 187088 5152 187110
rect 84180 187162 90896 187184
rect 84180 187110 85982 187162
rect 86034 187110 86046 187162
rect 86098 187110 86110 187162
rect 86162 187110 86174 187162
rect 86226 187110 89982 187162
rect 90034 187110 90046 187162
rect 90098 187110 90110 187162
rect 90162 187110 90174 187162
rect 90226 187110 90896 187162
rect 84180 187088 90896 187110
rect 79318 186844 79324 186856
rect 64846 186816 79324 186844
rect 4430 186736 4436 186788
rect 4488 186776 4494 186788
rect 64846 186776 64874 186816
rect 79318 186804 79324 186816
rect 79376 186804 79382 186856
rect 4488 186748 64874 186776
rect 4488 186736 4494 186748
rect 1104 186618 5152 186640
rect 1104 186566 3982 186618
rect 4034 186566 4046 186618
rect 4098 186566 4110 186618
rect 4162 186566 4174 186618
rect 4226 186566 5152 186618
rect 1104 186544 5152 186566
rect 84180 186618 90896 186640
rect 84180 186566 87982 186618
rect 88034 186566 88046 186618
rect 88098 186566 88110 186618
rect 88162 186566 88174 186618
rect 88226 186566 90896 186618
rect 84180 186544 90896 186566
rect 84378 186328 84384 186380
rect 84436 186368 84442 186380
rect 84657 186371 84715 186377
rect 84657 186368 84669 186371
rect 84436 186340 84669 186368
rect 84436 186328 84442 186340
rect 84657 186337 84669 186340
rect 84703 186337 84715 186371
rect 84657 186331 84715 186337
rect 1104 186074 5152 186096
rect 1104 186022 1982 186074
rect 2034 186022 2046 186074
rect 2098 186022 2110 186074
rect 2162 186022 2174 186074
rect 2226 186022 5152 186074
rect 1104 186000 5152 186022
rect 84180 186074 90896 186096
rect 84180 186022 85982 186074
rect 86034 186022 86046 186074
rect 86098 186022 86110 186074
rect 86162 186022 86174 186074
rect 86226 186022 89982 186074
rect 90034 186022 90046 186074
rect 90098 186022 90110 186074
rect 90162 186022 90174 186074
rect 90226 186022 90896 186074
rect 84180 186000 90896 186022
rect 1104 185530 5152 185552
rect 1104 185478 3982 185530
rect 4034 185478 4046 185530
rect 4098 185478 4110 185530
rect 4162 185478 4174 185530
rect 4226 185478 5152 185530
rect 1104 185456 5152 185478
rect 84180 185530 90896 185552
rect 84180 185478 87982 185530
rect 88034 185478 88046 185530
rect 88098 185478 88110 185530
rect 88162 185478 88174 185530
rect 88226 185478 90896 185530
rect 84180 185456 90896 185478
rect 1104 184986 5152 185008
rect 1104 184934 1982 184986
rect 2034 184934 2046 184986
rect 2098 184934 2110 184986
rect 2162 184934 2174 184986
rect 2226 184934 5152 184986
rect 1104 184912 5152 184934
rect 84180 184986 90896 185008
rect 84180 184934 85982 184986
rect 86034 184934 86046 184986
rect 86098 184934 86110 184986
rect 86162 184934 86174 184986
rect 86226 184934 89982 184986
rect 90034 184934 90046 184986
rect 90098 184934 90110 184986
rect 90162 184934 90174 184986
rect 90226 184934 90896 184986
rect 84180 184912 90896 184934
rect 1104 184442 5152 184464
rect 1104 184390 3982 184442
rect 4034 184390 4046 184442
rect 4098 184390 4110 184442
rect 4162 184390 4174 184442
rect 4226 184390 5152 184442
rect 1104 184368 5152 184390
rect 84180 184442 90896 184464
rect 84180 184390 87982 184442
rect 88034 184390 88046 184442
rect 88098 184390 88110 184442
rect 88162 184390 88174 184442
rect 88226 184390 90896 184442
rect 84180 184368 90896 184390
rect 1104 183898 5152 183920
rect 1104 183846 1982 183898
rect 2034 183846 2046 183898
rect 2098 183846 2110 183898
rect 2162 183846 2174 183898
rect 2226 183846 5152 183898
rect 1104 183824 5152 183846
rect 84180 183898 90896 183920
rect 84180 183846 85982 183898
rect 86034 183846 86046 183898
rect 86098 183846 86110 183898
rect 86162 183846 86174 183898
rect 86226 183846 89982 183898
rect 90034 183846 90046 183898
rect 90098 183846 90110 183898
rect 90162 183846 90174 183898
rect 90226 183846 90896 183898
rect 84180 183824 90896 183846
rect 1104 183354 5152 183376
rect 1104 183302 3982 183354
rect 4034 183302 4046 183354
rect 4098 183302 4110 183354
rect 4162 183302 4174 183354
rect 4226 183302 5152 183354
rect 1104 183280 5152 183302
rect 84180 183354 90896 183376
rect 84180 183302 87982 183354
rect 88034 183302 88046 183354
rect 88098 183302 88110 183354
rect 88162 183302 88174 183354
rect 88226 183302 90896 183354
rect 84180 183280 90896 183302
rect 4798 182968 4804 182980
rect 4759 182940 4804 182968
rect 4798 182928 4804 182940
rect 4856 182928 4862 182980
rect 1104 182810 5152 182832
rect 1104 182758 1982 182810
rect 2034 182758 2046 182810
rect 2098 182758 2110 182810
rect 2162 182758 2174 182810
rect 2226 182758 5152 182810
rect 1104 182736 5152 182758
rect 84180 182810 90896 182832
rect 84180 182758 85982 182810
rect 86034 182758 86046 182810
rect 86098 182758 86110 182810
rect 86162 182758 86174 182810
rect 86226 182758 89982 182810
rect 90034 182758 90046 182810
rect 90098 182758 90110 182810
rect 90162 182758 90174 182810
rect 90226 182758 90896 182810
rect 84180 182736 90896 182758
rect 1104 182266 5152 182288
rect 1104 182214 3982 182266
rect 4034 182214 4046 182266
rect 4098 182214 4110 182266
rect 4162 182214 4174 182266
rect 4226 182214 5152 182266
rect 1104 182192 5152 182214
rect 84180 182266 90896 182288
rect 84180 182214 87982 182266
rect 88034 182214 88046 182266
rect 88098 182214 88110 182266
rect 88162 182214 88174 182266
rect 88226 182214 90896 182266
rect 84180 182192 90896 182214
rect 4798 181880 4804 181892
rect 4759 181852 4804 181880
rect 4798 181840 4804 181852
rect 4856 181840 4862 181892
rect 1104 181722 5152 181744
rect 1104 181670 1982 181722
rect 2034 181670 2046 181722
rect 2098 181670 2110 181722
rect 2162 181670 2174 181722
rect 2226 181670 5152 181722
rect 1104 181648 5152 181670
rect 84180 181722 90896 181744
rect 84180 181670 85982 181722
rect 86034 181670 86046 181722
rect 86098 181670 86110 181722
rect 86162 181670 86174 181722
rect 86226 181670 89982 181722
rect 90034 181670 90046 181722
rect 90098 181670 90110 181722
rect 90162 181670 90174 181722
rect 90226 181670 90896 181722
rect 84180 181648 90896 181670
rect 1104 181178 5152 181200
rect 1104 181126 3982 181178
rect 4034 181126 4046 181178
rect 4098 181126 4110 181178
rect 4162 181126 4174 181178
rect 4226 181126 5152 181178
rect 1104 181104 5152 181126
rect 84180 181178 90896 181200
rect 84180 181126 87982 181178
rect 88034 181126 88046 181178
rect 88098 181126 88110 181178
rect 88162 181126 88174 181178
rect 88226 181126 90896 181178
rect 84180 181104 90896 181126
rect 83734 180820 83740 180872
rect 83792 180860 83798 180872
rect 87690 180860 87696 180872
rect 83792 180832 87696 180860
rect 83792 180820 83798 180832
rect 87690 180820 87696 180832
rect 87748 180820 87754 180872
rect 1104 180634 5152 180656
rect 1104 180582 1982 180634
rect 2034 180582 2046 180634
rect 2098 180582 2110 180634
rect 2162 180582 2174 180634
rect 2226 180582 5152 180634
rect 1104 180560 5152 180582
rect 84180 180634 90896 180656
rect 84180 180582 85982 180634
rect 86034 180582 86046 180634
rect 86098 180582 86110 180634
rect 86162 180582 86174 180634
rect 86226 180582 89982 180634
rect 90034 180582 90046 180634
rect 90098 180582 90110 180634
rect 90162 180582 90174 180634
rect 90226 180582 90896 180634
rect 84180 180560 90896 180582
rect 4614 180140 4620 180192
rect 4672 180180 4678 180192
rect 4709 180183 4767 180189
rect 4709 180180 4721 180183
rect 4672 180152 4721 180180
rect 4672 180140 4678 180152
rect 4709 180149 4721 180152
rect 4755 180149 4767 180183
rect 4709 180143 4767 180149
rect 1104 180090 5152 180112
rect 1104 180038 3982 180090
rect 4034 180038 4046 180090
rect 4098 180038 4110 180090
rect 4162 180038 4174 180090
rect 4226 180038 5152 180090
rect 1104 180016 5152 180038
rect 84180 180090 90896 180112
rect 84180 180038 87982 180090
rect 88034 180038 88046 180090
rect 88098 180038 88110 180090
rect 88162 180038 88174 180090
rect 88226 180038 90896 180090
rect 84180 180016 90896 180038
rect 84473 179639 84531 179645
rect 84473 179605 84485 179639
rect 84519 179636 84531 179639
rect 84562 179636 84568 179648
rect 84519 179608 84568 179636
rect 84519 179605 84531 179608
rect 84473 179599 84531 179605
rect 84562 179596 84568 179608
rect 84620 179596 84626 179648
rect 1104 179546 5152 179568
rect 1104 179494 1982 179546
rect 2034 179494 2046 179546
rect 2098 179494 2110 179546
rect 2162 179494 2174 179546
rect 2226 179494 5152 179546
rect 1104 179472 5152 179494
rect 84180 179546 90896 179568
rect 84180 179494 85982 179546
rect 86034 179494 86046 179546
rect 86098 179494 86110 179546
rect 86162 179494 86174 179546
rect 86226 179494 89982 179546
rect 90034 179494 90046 179546
rect 90098 179494 90110 179546
rect 90162 179494 90174 179546
rect 90226 179494 90896 179546
rect 84180 179472 90896 179494
rect 4522 179052 4528 179104
rect 4580 179092 4586 179104
rect 4709 179095 4767 179101
rect 4709 179092 4721 179095
rect 4580 179064 4721 179092
rect 4580 179052 4586 179064
rect 4709 179061 4721 179064
rect 4755 179061 4767 179095
rect 4709 179055 4767 179061
rect 1104 179002 5152 179024
rect 1104 178950 3982 179002
rect 4034 178950 4046 179002
rect 4098 178950 4110 179002
rect 4162 178950 4174 179002
rect 4226 178950 5152 179002
rect 1104 178928 5152 178950
rect 84180 179002 90896 179024
rect 84180 178950 87982 179002
rect 88034 178950 88046 179002
rect 88098 178950 88110 179002
rect 88162 178950 88174 179002
rect 88226 178950 90896 179002
rect 84180 178928 90896 178950
rect 1104 178458 5152 178480
rect 1104 178406 1982 178458
rect 2034 178406 2046 178458
rect 2098 178406 2110 178458
rect 2162 178406 2174 178458
rect 2226 178406 5152 178458
rect 1104 178384 5152 178406
rect 84180 178458 90896 178480
rect 84180 178406 85982 178458
rect 86034 178406 86046 178458
rect 86098 178406 86110 178458
rect 86162 178406 86174 178458
rect 86226 178406 89982 178458
rect 90034 178406 90046 178458
rect 90098 178406 90110 178458
rect 90162 178406 90174 178458
rect 90226 178406 90896 178458
rect 84180 178384 90896 178406
rect 1104 177914 5152 177936
rect 1104 177862 3982 177914
rect 4034 177862 4046 177914
rect 4098 177862 4110 177914
rect 4162 177862 4174 177914
rect 4226 177862 5152 177914
rect 1104 177840 5152 177862
rect 84180 177914 90896 177936
rect 84180 177862 87982 177914
rect 88034 177862 88046 177914
rect 88098 177862 88110 177914
rect 88162 177862 88174 177914
rect 88226 177862 90896 177914
rect 84180 177840 90896 177862
rect 1104 177370 5152 177392
rect 1104 177318 1982 177370
rect 2034 177318 2046 177370
rect 2098 177318 2110 177370
rect 2162 177318 2174 177370
rect 2226 177318 5152 177370
rect 1104 177296 5152 177318
rect 84180 177370 90896 177392
rect 84180 177318 85982 177370
rect 86034 177318 86046 177370
rect 86098 177318 86110 177370
rect 86162 177318 86174 177370
rect 86226 177318 89982 177370
rect 90034 177318 90046 177370
rect 90098 177318 90110 177370
rect 90162 177318 90174 177370
rect 90226 177318 90896 177370
rect 84180 177296 90896 177318
rect 4706 176916 4712 176928
rect 4667 176888 4712 176916
rect 4706 176876 4712 176888
rect 4764 176876 4770 176928
rect 1104 176826 5152 176848
rect 1104 176774 3982 176826
rect 4034 176774 4046 176826
rect 4098 176774 4110 176826
rect 4162 176774 4174 176826
rect 4226 176774 5152 176826
rect 1104 176752 5152 176774
rect 84180 176826 90896 176848
rect 84180 176774 87982 176826
rect 88034 176774 88046 176826
rect 88098 176774 88110 176826
rect 88162 176774 88174 176826
rect 88226 176774 90896 176826
rect 84180 176752 90896 176774
rect 1104 176282 5152 176304
rect 1104 176230 1982 176282
rect 2034 176230 2046 176282
rect 2098 176230 2110 176282
rect 2162 176230 2174 176282
rect 2226 176230 5152 176282
rect 1104 176208 5152 176230
rect 84180 176282 90896 176304
rect 84180 176230 85982 176282
rect 86034 176230 86046 176282
rect 86098 176230 86110 176282
rect 86162 176230 86174 176282
rect 86226 176230 89982 176282
rect 90034 176230 90046 176282
rect 90098 176230 90110 176282
rect 90162 176230 90174 176282
rect 90226 176230 90896 176282
rect 84180 176208 90896 176230
rect 4798 176168 4804 176180
rect 4759 176140 4804 176168
rect 4798 176128 4804 176140
rect 4856 176128 4862 176180
rect 1104 175738 5152 175760
rect 1104 175686 3982 175738
rect 4034 175686 4046 175738
rect 4098 175686 4110 175738
rect 4162 175686 4174 175738
rect 4226 175686 5152 175738
rect 1104 175664 5152 175686
rect 84180 175738 90896 175760
rect 84180 175686 87982 175738
rect 88034 175686 88046 175738
rect 88098 175686 88110 175738
rect 88162 175686 88174 175738
rect 88226 175686 90896 175738
rect 84180 175664 90896 175686
rect 1104 175194 5152 175216
rect 1104 175142 1982 175194
rect 2034 175142 2046 175194
rect 2098 175142 2110 175194
rect 2162 175142 2174 175194
rect 2226 175142 5152 175194
rect 1104 175120 5152 175142
rect 84180 175194 90896 175216
rect 84180 175142 85982 175194
rect 86034 175142 86046 175194
rect 86098 175142 86110 175194
rect 86162 175142 86174 175194
rect 86226 175142 89982 175194
rect 90034 175142 90046 175194
rect 90098 175142 90110 175194
rect 90162 175142 90174 175194
rect 90226 175142 90896 175194
rect 84180 175120 90896 175142
rect 1104 174650 5152 174672
rect 1104 174598 3982 174650
rect 4034 174598 4046 174650
rect 4098 174598 4110 174650
rect 4162 174598 4174 174650
rect 4226 174598 5152 174650
rect 1104 174576 5152 174598
rect 84180 174650 90896 174672
rect 84180 174598 87982 174650
rect 88034 174598 88046 174650
rect 88098 174598 88110 174650
rect 88162 174598 88174 174650
rect 88226 174598 90896 174650
rect 84180 174576 90896 174598
rect 4798 174536 4804 174548
rect 4759 174508 4804 174536
rect 4798 174496 4804 174508
rect 4856 174496 4862 174548
rect 4522 174360 4528 174412
rect 4580 174400 4586 174412
rect 4798 174400 4804 174412
rect 4580 174372 4804 174400
rect 4580 174360 4586 174372
rect 4798 174360 4804 174372
rect 4856 174360 4862 174412
rect 4614 174292 4620 174344
rect 4672 174332 4678 174344
rect 4982 174332 4988 174344
rect 4672 174304 4988 174332
rect 4672 174292 4678 174304
rect 4982 174292 4988 174304
rect 5040 174292 5046 174344
rect 1104 174106 5152 174128
rect 1104 174054 1982 174106
rect 2034 174054 2046 174106
rect 2098 174054 2110 174106
rect 2162 174054 2174 174106
rect 2226 174054 5152 174106
rect 1104 174032 5152 174054
rect 84180 174106 90896 174128
rect 84180 174054 85982 174106
rect 86034 174054 86046 174106
rect 86098 174054 86110 174106
rect 86162 174054 86174 174106
rect 86226 174054 89982 174106
rect 90034 174054 90046 174106
rect 90098 174054 90110 174106
rect 90162 174054 90174 174106
rect 90226 174054 90896 174106
rect 84180 174032 90896 174054
rect 83918 173884 83924 173936
rect 83976 173924 83982 173936
rect 87414 173924 87420 173936
rect 83976 173896 87420 173924
rect 83976 173884 83982 173896
rect 87414 173884 87420 173896
rect 87472 173884 87478 173936
rect 1104 173562 5152 173584
rect 1104 173510 3982 173562
rect 4034 173510 4046 173562
rect 4098 173510 4110 173562
rect 4162 173510 4174 173562
rect 4226 173510 5152 173562
rect 1104 173488 5152 173510
rect 84180 173562 90896 173584
rect 84180 173510 87982 173562
rect 88034 173510 88046 173562
rect 88098 173510 88110 173562
rect 88162 173510 88174 173562
rect 88226 173510 90896 173562
rect 84180 173488 90896 173510
rect 1104 173018 5152 173040
rect 1104 172966 1982 173018
rect 2034 172966 2046 173018
rect 2098 172966 2110 173018
rect 2162 172966 2174 173018
rect 2226 172966 5152 173018
rect 1104 172944 5152 172966
rect 84180 173018 90896 173040
rect 84180 172966 85982 173018
rect 86034 172966 86046 173018
rect 86098 172966 86110 173018
rect 86162 172966 86174 173018
rect 86226 172966 89982 173018
rect 90034 172966 90046 173018
rect 90098 172966 90110 173018
rect 90162 172966 90174 173018
rect 90226 172966 90896 173018
rect 84180 172944 90896 172966
rect 1104 172474 5152 172496
rect 1104 172422 3982 172474
rect 4034 172422 4046 172474
rect 4098 172422 4110 172474
rect 4162 172422 4174 172474
rect 4226 172422 5152 172474
rect 1104 172400 5152 172422
rect 84180 172474 90896 172496
rect 84180 172422 87982 172474
rect 88034 172422 88046 172474
rect 88098 172422 88110 172474
rect 88162 172422 88174 172474
rect 88226 172422 90896 172474
rect 84180 172400 90896 172422
rect 1104 171930 5152 171952
rect 1104 171878 1982 171930
rect 2034 171878 2046 171930
rect 2098 171878 2110 171930
rect 2162 171878 2174 171930
rect 2226 171878 5152 171930
rect 1104 171856 5152 171878
rect 84180 171930 90896 171952
rect 84180 171878 85982 171930
rect 86034 171878 86046 171930
rect 86098 171878 86110 171930
rect 86162 171878 86174 171930
rect 86226 171878 89982 171930
rect 90034 171878 90046 171930
rect 90098 171878 90110 171930
rect 90162 171878 90174 171930
rect 90226 171878 90896 171930
rect 84180 171856 90896 171878
rect 1104 171386 5152 171408
rect 1104 171334 3982 171386
rect 4034 171334 4046 171386
rect 4098 171334 4110 171386
rect 4162 171334 4174 171386
rect 4226 171334 5152 171386
rect 1104 171312 5152 171334
rect 84180 171386 90896 171408
rect 84180 171334 87982 171386
rect 88034 171334 88046 171386
rect 88098 171334 88110 171386
rect 88162 171334 88174 171386
rect 88226 171334 90896 171386
rect 84180 171312 90896 171334
rect 1104 170842 5152 170864
rect 1104 170790 1982 170842
rect 2034 170790 2046 170842
rect 2098 170790 2110 170842
rect 2162 170790 2174 170842
rect 2226 170790 5152 170842
rect 1104 170768 5152 170790
rect 84180 170842 90896 170864
rect 84180 170790 85982 170842
rect 86034 170790 86046 170842
rect 86098 170790 86110 170842
rect 86162 170790 86174 170842
rect 86226 170790 89982 170842
rect 90034 170790 90046 170842
rect 90098 170790 90110 170842
rect 90162 170790 90174 170842
rect 90226 170790 90896 170842
rect 84180 170768 90896 170790
rect 1104 170298 5152 170320
rect 1104 170246 3982 170298
rect 4034 170246 4046 170298
rect 4098 170246 4110 170298
rect 4162 170246 4174 170298
rect 4226 170246 5152 170298
rect 1104 170224 5152 170246
rect 84180 170298 90896 170320
rect 84180 170246 87982 170298
rect 88034 170246 88046 170298
rect 88098 170246 88110 170298
rect 88162 170246 88174 170298
rect 88226 170246 90896 170298
rect 84180 170224 90896 170246
rect 1104 169754 5152 169776
rect 1104 169702 1982 169754
rect 2034 169702 2046 169754
rect 2098 169702 2110 169754
rect 2162 169702 2174 169754
rect 2226 169702 5152 169754
rect 1104 169680 5152 169702
rect 84180 169754 90896 169776
rect 84180 169702 85982 169754
rect 86034 169702 86046 169754
rect 86098 169702 86110 169754
rect 86162 169702 86174 169754
rect 86226 169702 89982 169754
rect 90034 169702 90046 169754
rect 90098 169702 90110 169754
rect 90162 169702 90174 169754
rect 90226 169702 90896 169754
rect 84180 169680 90896 169702
rect 1104 169210 5152 169232
rect 1104 169158 3982 169210
rect 4034 169158 4046 169210
rect 4098 169158 4110 169210
rect 4162 169158 4174 169210
rect 4226 169158 5152 169210
rect 1104 169136 5152 169158
rect 84180 169210 90896 169232
rect 84180 169158 87982 169210
rect 88034 169158 88046 169210
rect 88098 169158 88110 169210
rect 88162 169158 88174 169210
rect 88226 169158 90896 169210
rect 84180 169136 90896 169158
rect 1104 168666 5152 168688
rect 1104 168614 1982 168666
rect 2034 168614 2046 168666
rect 2098 168614 2110 168666
rect 2162 168614 2174 168666
rect 2226 168614 5152 168666
rect 1104 168592 5152 168614
rect 84180 168666 90896 168688
rect 84180 168614 85982 168666
rect 86034 168614 86046 168666
rect 86098 168614 86110 168666
rect 86162 168614 86174 168666
rect 86226 168614 89982 168666
rect 90034 168614 90046 168666
rect 90098 168614 90110 168666
rect 90162 168614 90174 168666
rect 90226 168614 90896 168666
rect 84180 168592 90896 168614
rect 84010 168376 84016 168428
rect 84068 168416 84074 168428
rect 87874 168416 87880 168428
rect 84068 168388 87880 168416
rect 84068 168376 84074 168388
rect 87874 168376 87880 168388
rect 87932 168376 87938 168428
rect 1104 168122 5152 168144
rect 1104 168070 3982 168122
rect 4034 168070 4046 168122
rect 4098 168070 4110 168122
rect 4162 168070 4174 168122
rect 4226 168070 5152 168122
rect 1104 168048 5152 168070
rect 84180 168122 90896 168144
rect 84180 168070 87982 168122
rect 88034 168070 88046 168122
rect 88098 168070 88110 168122
rect 88162 168070 88174 168122
rect 88226 168070 90896 168122
rect 84180 168048 90896 168070
rect 1104 167578 5152 167600
rect 1104 167526 1982 167578
rect 2034 167526 2046 167578
rect 2098 167526 2110 167578
rect 2162 167526 2174 167578
rect 2226 167526 5152 167578
rect 1104 167504 5152 167526
rect 84180 167578 90896 167600
rect 84180 167526 85982 167578
rect 86034 167526 86046 167578
rect 86098 167526 86110 167578
rect 86162 167526 86174 167578
rect 86226 167526 89982 167578
rect 90034 167526 90046 167578
rect 90098 167526 90110 167578
rect 90162 167526 90174 167578
rect 90226 167526 90896 167578
rect 84180 167504 90896 167526
rect 84470 167464 84476 167476
rect 84431 167436 84476 167464
rect 84470 167424 84476 167436
rect 84528 167424 84534 167476
rect 83550 167084 83556 167136
rect 83608 167124 83614 167136
rect 87046 167124 87052 167136
rect 83608 167096 87052 167124
rect 83608 167084 83614 167096
rect 87046 167084 87052 167096
rect 87104 167084 87110 167136
rect 1104 167034 5152 167056
rect 1104 166982 3982 167034
rect 4034 166982 4046 167034
rect 4098 166982 4110 167034
rect 4162 166982 4174 167034
rect 4226 166982 5152 167034
rect 1104 166960 5152 166982
rect 84180 167034 90896 167056
rect 84180 166982 87982 167034
rect 88034 166982 88046 167034
rect 88098 166982 88110 167034
rect 88162 166982 88174 167034
rect 88226 166982 90896 167034
rect 84180 166960 90896 166982
rect 1104 166490 5152 166512
rect 1104 166438 1982 166490
rect 2034 166438 2046 166490
rect 2098 166438 2110 166490
rect 2162 166438 2174 166490
rect 2226 166438 5152 166490
rect 1104 166416 5152 166438
rect 84180 166490 90896 166512
rect 84180 166438 85982 166490
rect 86034 166438 86046 166490
rect 86098 166438 86110 166490
rect 86162 166438 86174 166490
rect 86226 166438 89982 166490
rect 90034 166438 90046 166490
rect 90098 166438 90110 166490
rect 90162 166438 90174 166490
rect 90226 166438 90896 166490
rect 84180 166416 90896 166438
rect 1104 165946 5152 165968
rect 1104 165894 3982 165946
rect 4034 165894 4046 165946
rect 4098 165894 4110 165946
rect 4162 165894 4174 165946
rect 4226 165894 5152 165946
rect 1104 165872 5152 165894
rect 84180 165946 90896 165968
rect 84180 165894 87982 165946
rect 88034 165894 88046 165946
rect 88098 165894 88110 165946
rect 88162 165894 88174 165946
rect 88226 165894 90896 165946
rect 84180 165872 90896 165894
rect 1104 165402 5152 165424
rect 1104 165350 1982 165402
rect 2034 165350 2046 165402
rect 2098 165350 2110 165402
rect 2162 165350 2174 165402
rect 2226 165350 5152 165402
rect 1104 165328 5152 165350
rect 84180 165402 90896 165424
rect 84180 165350 85982 165402
rect 86034 165350 86046 165402
rect 86098 165350 86110 165402
rect 86162 165350 86174 165402
rect 86226 165350 89982 165402
rect 90034 165350 90046 165402
rect 90098 165350 90110 165402
rect 90162 165350 90174 165402
rect 90226 165350 90896 165402
rect 84180 165328 90896 165350
rect 1104 164858 5152 164880
rect 1104 164806 3982 164858
rect 4034 164806 4046 164858
rect 4098 164806 4110 164858
rect 4162 164806 4174 164858
rect 4226 164806 5152 164858
rect 1104 164784 5152 164806
rect 84180 164858 90896 164880
rect 84180 164806 87982 164858
rect 88034 164806 88046 164858
rect 88098 164806 88110 164858
rect 88162 164806 88174 164858
rect 88226 164806 90896 164858
rect 84180 164784 90896 164806
rect 83826 164364 83832 164416
rect 83884 164404 83890 164416
rect 87874 164404 87880 164416
rect 83884 164376 87880 164404
rect 83884 164364 83890 164376
rect 87874 164364 87880 164376
rect 87932 164364 87938 164416
rect 1104 164314 5152 164336
rect 1104 164262 1982 164314
rect 2034 164262 2046 164314
rect 2098 164262 2110 164314
rect 2162 164262 2174 164314
rect 2226 164262 5152 164314
rect 1104 164240 5152 164262
rect 84180 164314 90896 164336
rect 84180 164262 85982 164314
rect 86034 164262 86046 164314
rect 86098 164262 86110 164314
rect 86162 164262 86174 164314
rect 86226 164262 89982 164314
rect 90034 164262 90046 164314
rect 90098 164262 90110 164314
rect 90162 164262 90174 164314
rect 90226 164262 90896 164314
rect 84180 164240 90896 164262
rect 1104 163770 5152 163792
rect 1104 163718 3982 163770
rect 4034 163718 4046 163770
rect 4098 163718 4110 163770
rect 4162 163718 4174 163770
rect 4226 163718 5152 163770
rect 1104 163696 5152 163718
rect 84180 163770 90896 163792
rect 84180 163718 87982 163770
rect 88034 163718 88046 163770
rect 88098 163718 88110 163770
rect 88162 163718 88174 163770
rect 88226 163718 90896 163770
rect 84180 163696 90896 163718
rect 1104 163226 5152 163248
rect 1104 163174 1982 163226
rect 2034 163174 2046 163226
rect 2098 163174 2110 163226
rect 2162 163174 2174 163226
rect 2226 163174 5152 163226
rect 1104 163152 5152 163174
rect 84180 163226 90896 163248
rect 84180 163174 85982 163226
rect 86034 163174 86046 163226
rect 86098 163174 86110 163226
rect 86162 163174 86174 163226
rect 86226 163174 89982 163226
rect 90034 163174 90046 163226
rect 90098 163174 90110 163226
rect 90162 163174 90174 163226
rect 90226 163174 90896 163226
rect 84180 163152 90896 163174
rect 82446 162868 82452 162920
rect 82504 162908 82510 162920
rect 87874 162908 87880 162920
rect 82504 162880 87880 162908
rect 82504 162868 82510 162880
rect 87874 162868 87880 162880
rect 87932 162868 87938 162920
rect 1104 162682 5152 162704
rect 1104 162630 3982 162682
rect 4034 162630 4046 162682
rect 4098 162630 4110 162682
rect 4162 162630 4174 162682
rect 4226 162630 5152 162682
rect 1104 162608 5152 162630
rect 84180 162682 90896 162704
rect 84180 162630 87982 162682
rect 88034 162630 88046 162682
rect 88098 162630 88110 162682
rect 88162 162630 88174 162682
rect 88226 162630 90896 162682
rect 84180 162608 90896 162630
rect 84654 162432 84660 162444
rect 84615 162404 84660 162432
rect 84654 162392 84660 162404
rect 84712 162392 84718 162444
rect 85114 162364 85120 162376
rect 85075 162336 85120 162364
rect 85114 162324 85120 162336
rect 85172 162324 85178 162376
rect 1104 162138 5152 162160
rect 1104 162086 1982 162138
rect 2034 162086 2046 162138
rect 2098 162086 2110 162138
rect 2162 162086 2174 162138
rect 2226 162086 5152 162138
rect 1104 162064 5152 162086
rect 84180 162138 90896 162160
rect 84180 162086 85982 162138
rect 86034 162086 86046 162138
rect 86098 162086 86110 162138
rect 86162 162086 86174 162138
rect 86226 162086 89982 162138
rect 90034 162086 90046 162138
rect 90098 162086 90110 162138
rect 90162 162086 90174 162138
rect 90226 162086 90896 162138
rect 84180 162064 90896 162086
rect 84654 162024 84660 162036
rect 84615 161996 84660 162024
rect 84654 161984 84660 161996
rect 84712 161984 84718 162036
rect 1104 161594 5152 161616
rect 1104 161542 3982 161594
rect 4034 161542 4046 161594
rect 4098 161542 4110 161594
rect 4162 161542 4174 161594
rect 4226 161542 5152 161594
rect 1104 161520 5152 161542
rect 84180 161594 90896 161616
rect 84180 161542 87982 161594
rect 88034 161542 88046 161594
rect 88098 161542 88110 161594
rect 88162 161542 88174 161594
rect 88226 161542 90896 161594
rect 84180 161520 90896 161542
rect 1104 161050 5152 161072
rect 1104 160998 1982 161050
rect 2034 160998 2046 161050
rect 2098 160998 2110 161050
rect 2162 160998 2174 161050
rect 2226 160998 5152 161050
rect 1104 160976 5152 160998
rect 84180 161050 90896 161072
rect 84180 160998 85982 161050
rect 86034 160998 86046 161050
rect 86098 160998 86110 161050
rect 86162 160998 86174 161050
rect 86226 160998 89982 161050
rect 90034 160998 90046 161050
rect 90098 160998 90110 161050
rect 90162 160998 90174 161050
rect 90226 160998 90896 161050
rect 84180 160976 90896 160998
rect 1104 160506 5152 160528
rect 1104 160454 3982 160506
rect 4034 160454 4046 160506
rect 4098 160454 4110 160506
rect 4162 160454 4174 160506
rect 4226 160454 5152 160506
rect 1104 160432 5152 160454
rect 84180 160506 90896 160528
rect 84180 160454 87982 160506
rect 88034 160454 88046 160506
rect 88098 160454 88110 160506
rect 88162 160454 88174 160506
rect 88226 160454 90896 160506
rect 84180 160432 90896 160454
rect 84470 160120 84476 160132
rect 84431 160092 84476 160120
rect 84470 160080 84476 160092
rect 84528 160080 84534 160132
rect 1104 159962 5152 159984
rect 1104 159910 1982 159962
rect 2034 159910 2046 159962
rect 2098 159910 2110 159962
rect 2162 159910 2174 159962
rect 2226 159910 5152 159962
rect 1104 159888 5152 159910
rect 84180 159962 90896 159984
rect 84180 159910 85982 159962
rect 86034 159910 86046 159962
rect 86098 159910 86110 159962
rect 86162 159910 86174 159962
rect 86226 159910 89982 159962
rect 90034 159910 90046 159962
rect 90098 159910 90110 159962
rect 90162 159910 90174 159962
rect 90226 159910 90896 159962
rect 84180 159888 90896 159910
rect 1104 159418 5152 159440
rect 1104 159366 3982 159418
rect 4034 159366 4046 159418
rect 4098 159366 4110 159418
rect 4162 159366 4174 159418
rect 4226 159366 5152 159418
rect 1104 159344 5152 159366
rect 84180 159418 90896 159440
rect 84180 159366 87982 159418
rect 88034 159366 88046 159418
rect 88098 159366 88110 159418
rect 88162 159366 88174 159418
rect 88226 159366 90896 159418
rect 84180 159344 90896 159366
rect 1104 158874 5152 158896
rect 1104 158822 1982 158874
rect 2034 158822 2046 158874
rect 2098 158822 2110 158874
rect 2162 158822 2174 158874
rect 2226 158822 5152 158874
rect 1104 158800 5152 158822
rect 84180 158874 90896 158896
rect 84180 158822 85982 158874
rect 86034 158822 86046 158874
rect 86098 158822 86110 158874
rect 86162 158822 86174 158874
rect 86226 158822 89982 158874
rect 90034 158822 90046 158874
rect 90098 158822 90110 158874
rect 90162 158822 90174 158874
rect 90226 158822 90896 158874
rect 84180 158800 90896 158822
rect 1104 158330 5152 158352
rect 1104 158278 3982 158330
rect 4034 158278 4046 158330
rect 4098 158278 4110 158330
rect 4162 158278 4174 158330
rect 4226 158278 5152 158330
rect 1104 158256 5152 158278
rect 84180 158330 90896 158352
rect 84180 158278 87982 158330
rect 88034 158278 88046 158330
rect 88098 158278 88110 158330
rect 88162 158278 88174 158330
rect 88226 158278 90896 158330
rect 84180 158256 90896 158278
rect 1104 157786 5152 157808
rect 1104 157734 1982 157786
rect 2034 157734 2046 157786
rect 2098 157734 2110 157786
rect 2162 157734 2174 157786
rect 2226 157734 5152 157786
rect 1104 157712 5152 157734
rect 84180 157786 90896 157808
rect 84180 157734 85982 157786
rect 86034 157734 86046 157786
rect 86098 157734 86110 157786
rect 86162 157734 86174 157786
rect 86226 157734 89982 157786
rect 90034 157734 90046 157786
rect 90098 157734 90110 157786
rect 90162 157734 90174 157786
rect 90226 157734 90896 157786
rect 84180 157712 90896 157734
rect 1104 157242 5152 157264
rect 1104 157190 3982 157242
rect 4034 157190 4046 157242
rect 4098 157190 4110 157242
rect 4162 157190 4174 157242
rect 4226 157190 5152 157242
rect 1104 157168 5152 157190
rect 84180 157242 90896 157264
rect 84180 157190 87982 157242
rect 88034 157190 88046 157242
rect 88098 157190 88110 157242
rect 88162 157190 88174 157242
rect 88226 157190 90896 157242
rect 84180 157168 90896 157190
rect 1104 156698 5152 156720
rect 1104 156646 1982 156698
rect 2034 156646 2046 156698
rect 2098 156646 2110 156698
rect 2162 156646 2174 156698
rect 2226 156646 5152 156698
rect 1104 156624 5152 156646
rect 84180 156698 90896 156720
rect 84180 156646 85982 156698
rect 86034 156646 86046 156698
rect 86098 156646 86110 156698
rect 86162 156646 86174 156698
rect 86226 156646 89982 156698
rect 90034 156646 90046 156698
rect 90098 156646 90110 156698
rect 90162 156646 90174 156698
rect 90226 156646 90896 156698
rect 84180 156624 90896 156646
rect 1104 156154 5152 156176
rect 1104 156102 3982 156154
rect 4034 156102 4046 156154
rect 4098 156102 4110 156154
rect 4162 156102 4174 156154
rect 4226 156102 5152 156154
rect 1104 156080 5152 156102
rect 84180 156154 90896 156176
rect 84180 156102 87982 156154
rect 88034 156102 88046 156154
rect 88098 156102 88110 156154
rect 88162 156102 88174 156154
rect 88226 156102 90896 156154
rect 84180 156080 90896 156102
rect 1104 155610 5152 155632
rect 1104 155558 1982 155610
rect 2034 155558 2046 155610
rect 2098 155558 2110 155610
rect 2162 155558 2174 155610
rect 2226 155558 5152 155610
rect 1104 155536 5152 155558
rect 84180 155610 90896 155632
rect 84180 155558 85982 155610
rect 86034 155558 86046 155610
rect 86098 155558 86110 155610
rect 86162 155558 86174 155610
rect 86226 155558 89982 155610
rect 90034 155558 90046 155610
rect 90098 155558 90110 155610
rect 90162 155558 90174 155610
rect 90226 155558 90896 155610
rect 84180 155536 90896 155558
rect 1104 155066 5152 155088
rect 1104 155014 3982 155066
rect 4034 155014 4046 155066
rect 4098 155014 4110 155066
rect 4162 155014 4174 155066
rect 4226 155014 5152 155066
rect 1104 154992 5152 155014
rect 84180 155066 90896 155088
rect 84180 155014 87982 155066
rect 88034 155014 88046 155066
rect 88098 155014 88110 155066
rect 88162 155014 88174 155066
rect 88226 155014 90896 155066
rect 84180 154992 90896 155014
rect 1104 154522 5152 154544
rect 1104 154470 1982 154522
rect 2034 154470 2046 154522
rect 2098 154470 2110 154522
rect 2162 154470 2174 154522
rect 2226 154470 5152 154522
rect 1104 154448 5152 154470
rect 84180 154522 90896 154544
rect 84180 154470 85982 154522
rect 86034 154470 86046 154522
rect 86098 154470 86110 154522
rect 86162 154470 86174 154522
rect 86226 154470 89982 154522
rect 90034 154470 90046 154522
rect 90098 154470 90110 154522
rect 90162 154470 90174 154522
rect 90226 154470 90896 154522
rect 84180 154448 90896 154470
rect 1104 153978 5152 154000
rect 1104 153926 3982 153978
rect 4034 153926 4046 153978
rect 4098 153926 4110 153978
rect 4162 153926 4174 153978
rect 4226 153926 5152 153978
rect 1104 153904 5152 153926
rect 84180 153978 90896 154000
rect 84180 153926 87982 153978
rect 88034 153926 88046 153978
rect 88098 153926 88110 153978
rect 88162 153926 88174 153978
rect 88226 153926 90896 153978
rect 84180 153904 90896 153926
rect 84378 153824 84384 153876
rect 84436 153864 84442 153876
rect 84657 153867 84715 153873
rect 84657 153864 84669 153867
rect 84436 153836 84669 153864
rect 84436 153824 84442 153836
rect 84657 153833 84669 153836
rect 84703 153833 84715 153867
rect 84657 153827 84715 153833
rect 1104 153434 5152 153456
rect 1104 153382 1982 153434
rect 2034 153382 2046 153434
rect 2098 153382 2110 153434
rect 2162 153382 2174 153434
rect 2226 153382 5152 153434
rect 1104 153360 5152 153382
rect 84180 153434 90896 153456
rect 84180 153382 85982 153434
rect 86034 153382 86046 153434
rect 86098 153382 86110 153434
rect 86162 153382 86174 153434
rect 86226 153382 89982 153434
rect 90034 153382 90046 153434
rect 90098 153382 90110 153434
rect 90162 153382 90174 153434
rect 90226 153382 90896 153434
rect 84180 153360 90896 153382
rect 1104 152890 5152 152912
rect 1104 152838 3982 152890
rect 4034 152838 4046 152890
rect 4098 152838 4110 152890
rect 4162 152838 4174 152890
rect 4226 152838 5152 152890
rect 1104 152816 5152 152838
rect 84180 152890 90896 152912
rect 84180 152838 87982 152890
rect 88034 152838 88046 152890
rect 88098 152838 88110 152890
rect 88162 152838 88174 152890
rect 88226 152838 90896 152890
rect 84180 152816 90896 152838
rect 1104 152346 5152 152368
rect 1104 152294 1982 152346
rect 2034 152294 2046 152346
rect 2098 152294 2110 152346
rect 2162 152294 2174 152346
rect 2226 152294 5152 152346
rect 1104 152272 5152 152294
rect 84180 152346 90896 152368
rect 84180 152294 85982 152346
rect 86034 152294 86046 152346
rect 86098 152294 86110 152346
rect 86162 152294 86174 152346
rect 86226 152294 89982 152346
rect 90034 152294 90046 152346
rect 90098 152294 90110 152346
rect 90162 152294 90174 152346
rect 90226 152294 90896 152346
rect 84180 152272 90896 152294
rect 1104 151802 5152 151824
rect 1104 151750 3982 151802
rect 4034 151750 4046 151802
rect 4098 151750 4110 151802
rect 4162 151750 4174 151802
rect 4226 151750 5152 151802
rect 1104 151728 5152 151750
rect 84180 151802 90896 151824
rect 84180 151750 87982 151802
rect 88034 151750 88046 151802
rect 88098 151750 88110 151802
rect 88162 151750 88174 151802
rect 88226 151750 90896 151802
rect 84180 151728 90896 151750
rect 1104 151258 5152 151280
rect 1104 151206 1982 151258
rect 2034 151206 2046 151258
rect 2098 151206 2110 151258
rect 2162 151206 2174 151258
rect 2226 151206 5152 151258
rect 1104 151184 5152 151206
rect 84180 151258 90896 151280
rect 84180 151206 85982 151258
rect 86034 151206 86046 151258
rect 86098 151206 86110 151258
rect 86162 151206 86174 151258
rect 86226 151206 89982 151258
rect 90034 151206 90046 151258
rect 90098 151206 90110 151258
rect 90162 151206 90174 151258
rect 90226 151206 90896 151258
rect 84180 151184 90896 151206
rect 1104 150714 5152 150736
rect 1104 150662 3982 150714
rect 4034 150662 4046 150714
rect 4098 150662 4110 150714
rect 4162 150662 4174 150714
rect 4226 150662 5152 150714
rect 1104 150640 5152 150662
rect 84180 150714 90896 150736
rect 84180 150662 87982 150714
rect 88034 150662 88046 150714
rect 88098 150662 88110 150714
rect 88162 150662 88174 150714
rect 88226 150662 90896 150714
rect 84180 150640 90896 150662
rect 1104 150170 5152 150192
rect 1104 150118 1982 150170
rect 2034 150118 2046 150170
rect 2098 150118 2110 150170
rect 2162 150118 2174 150170
rect 2226 150118 5152 150170
rect 1104 150096 5152 150118
rect 84180 150170 90896 150192
rect 84180 150118 85982 150170
rect 86034 150118 86046 150170
rect 86098 150118 86110 150170
rect 86162 150118 86174 150170
rect 86226 150118 89982 150170
rect 90034 150118 90046 150170
rect 90098 150118 90110 150170
rect 90162 150118 90174 150170
rect 90226 150118 90896 150170
rect 84180 150096 90896 150118
rect 1104 149626 5152 149648
rect 1104 149574 3982 149626
rect 4034 149574 4046 149626
rect 4098 149574 4110 149626
rect 4162 149574 4174 149626
rect 4226 149574 5152 149626
rect 1104 149552 5152 149574
rect 84180 149626 90896 149648
rect 84180 149574 87982 149626
rect 88034 149574 88046 149626
rect 88098 149574 88110 149626
rect 88162 149574 88174 149626
rect 88226 149574 90896 149626
rect 84180 149552 90896 149574
rect 1104 149082 5152 149104
rect 1104 149030 1982 149082
rect 2034 149030 2046 149082
rect 2098 149030 2110 149082
rect 2162 149030 2174 149082
rect 2226 149030 5152 149082
rect 1104 149008 5152 149030
rect 84180 149082 90896 149104
rect 84180 149030 85982 149082
rect 86034 149030 86046 149082
rect 86098 149030 86110 149082
rect 86162 149030 86174 149082
rect 86226 149030 89982 149082
rect 90034 149030 90046 149082
rect 90098 149030 90110 149082
rect 90162 149030 90174 149082
rect 90226 149030 90896 149082
rect 84180 149008 90896 149030
rect 1104 148538 5152 148560
rect 1104 148486 3982 148538
rect 4034 148486 4046 148538
rect 4098 148486 4110 148538
rect 4162 148486 4174 148538
rect 4226 148486 5152 148538
rect 1104 148464 5152 148486
rect 84180 148538 90896 148560
rect 84180 148486 87982 148538
rect 88034 148486 88046 148538
rect 88098 148486 88110 148538
rect 88162 148486 88174 148538
rect 88226 148486 90896 148538
rect 84180 148464 90896 148486
rect 1104 147994 5152 148016
rect 1104 147942 1982 147994
rect 2034 147942 2046 147994
rect 2098 147942 2110 147994
rect 2162 147942 2174 147994
rect 2226 147942 5152 147994
rect 1104 147920 5152 147942
rect 84180 147994 90896 148016
rect 84180 147942 85982 147994
rect 86034 147942 86046 147994
rect 86098 147942 86110 147994
rect 86162 147942 86174 147994
rect 86226 147942 89982 147994
rect 90034 147942 90046 147994
rect 90098 147942 90110 147994
rect 90162 147942 90174 147994
rect 90226 147942 90896 147994
rect 84180 147920 90896 147942
rect 1104 147450 5152 147472
rect 1104 147398 3982 147450
rect 4034 147398 4046 147450
rect 4098 147398 4110 147450
rect 4162 147398 4174 147450
rect 4226 147398 5152 147450
rect 1104 147376 5152 147398
rect 84180 147450 90896 147472
rect 84180 147398 87982 147450
rect 88034 147398 88046 147450
rect 88098 147398 88110 147450
rect 88162 147398 88174 147450
rect 88226 147398 90896 147450
rect 84180 147376 90896 147398
rect 1104 146906 5152 146928
rect 1104 146854 1982 146906
rect 2034 146854 2046 146906
rect 2098 146854 2110 146906
rect 2162 146854 2174 146906
rect 2226 146854 5152 146906
rect 1104 146832 5152 146854
rect 84180 146906 90896 146928
rect 84180 146854 85982 146906
rect 86034 146854 86046 146906
rect 86098 146854 86110 146906
rect 86162 146854 86174 146906
rect 86226 146854 89982 146906
rect 90034 146854 90046 146906
rect 90098 146854 90110 146906
rect 90162 146854 90174 146906
rect 90226 146854 90896 146906
rect 84180 146832 90896 146854
rect 1104 146362 5152 146384
rect 1104 146310 3982 146362
rect 4034 146310 4046 146362
rect 4098 146310 4110 146362
rect 4162 146310 4174 146362
rect 4226 146310 5152 146362
rect 1104 146288 5152 146310
rect 84180 146362 90896 146384
rect 84180 146310 87982 146362
rect 88034 146310 88046 146362
rect 88098 146310 88110 146362
rect 88162 146310 88174 146362
rect 88226 146310 90896 146362
rect 84180 146288 90896 146310
rect 1104 145818 5152 145840
rect 1104 145766 1982 145818
rect 2034 145766 2046 145818
rect 2098 145766 2110 145818
rect 2162 145766 2174 145818
rect 2226 145766 5152 145818
rect 1104 145744 5152 145766
rect 84180 145818 90896 145840
rect 84180 145766 85982 145818
rect 86034 145766 86046 145818
rect 86098 145766 86110 145818
rect 86162 145766 86174 145818
rect 86226 145766 89982 145818
rect 90034 145766 90046 145818
rect 90098 145766 90110 145818
rect 90162 145766 90174 145818
rect 90226 145766 90896 145818
rect 84180 145744 90896 145766
rect 1104 145274 5152 145296
rect 1104 145222 3982 145274
rect 4034 145222 4046 145274
rect 4098 145222 4110 145274
rect 4162 145222 4174 145274
rect 4226 145222 5152 145274
rect 1104 145200 5152 145222
rect 84180 145274 90896 145296
rect 84180 145222 87982 145274
rect 88034 145222 88046 145274
rect 88098 145222 88110 145274
rect 88162 145222 88174 145274
rect 88226 145222 90896 145274
rect 84180 145200 90896 145222
rect 84746 144916 84752 144968
rect 84804 144956 84810 144968
rect 87966 144956 87972 144968
rect 84804 144928 87972 144956
rect 84804 144916 84810 144928
rect 87966 144916 87972 144928
rect 88024 144916 88030 144968
rect 1104 144730 5152 144752
rect 1104 144678 1982 144730
rect 2034 144678 2046 144730
rect 2098 144678 2110 144730
rect 2162 144678 2174 144730
rect 2226 144678 5152 144730
rect 1104 144656 5152 144678
rect 84180 144730 90896 144752
rect 84180 144678 85982 144730
rect 86034 144678 86046 144730
rect 86098 144678 86110 144730
rect 86162 144678 86174 144730
rect 86226 144678 89982 144730
rect 90034 144678 90046 144730
rect 90098 144678 90110 144730
rect 90162 144678 90174 144730
rect 90226 144678 90896 144730
rect 84180 144656 90896 144678
rect 1104 144186 5152 144208
rect 1104 144134 3982 144186
rect 4034 144134 4046 144186
rect 4098 144134 4110 144186
rect 4162 144134 4174 144186
rect 4226 144134 5152 144186
rect 1104 144112 5152 144134
rect 84180 144186 90896 144208
rect 84180 144134 87982 144186
rect 88034 144134 88046 144186
rect 88098 144134 88110 144186
rect 88162 144134 88174 144186
rect 88226 144134 90896 144186
rect 84180 144112 90896 144134
rect 85758 143692 85764 143744
rect 85816 143732 85822 143744
rect 88058 143732 88064 143744
rect 85816 143704 88064 143732
rect 85816 143692 85822 143704
rect 88058 143692 88064 143704
rect 88116 143692 88122 143744
rect 1104 143642 5152 143664
rect 1104 143590 1982 143642
rect 2034 143590 2046 143642
rect 2098 143590 2110 143642
rect 2162 143590 2174 143642
rect 2226 143590 5152 143642
rect 1104 143568 5152 143590
rect 84180 143642 90896 143664
rect 84180 143590 85982 143642
rect 86034 143590 86046 143642
rect 86098 143590 86110 143642
rect 86162 143590 86174 143642
rect 86226 143590 89982 143642
rect 90034 143590 90046 143642
rect 90098 143590 90110 143642
rect 90162 143590 90174 143642
rect 90226 143590 90896 143642
rect 84180 143568 90896 143590
rect 1104 143098 5152 143120
rect 1104 143046 3982 143098
rect 4034 143046 4046 143098
rect 4098 143046 4110 143098
rect 4162 143046 4174 143098
rect 4226 143046 5152 143098
rect 1104 143024 5152 143046
rect 84180 143098 90896 143120
rect 84180 143046 87982 143098
rect 88034 143046 88046 143098
rect 88098 143046 88110 143098
rect 88162 143046 88174 143098
rect 88226 143046 90896 143098
rect 84180 143024 90896 143046
rect 1104 142554 5152 142576
rect 1104 142502 1982 142554
rect 2034 142502 2046 142554
rect 2098 142502 2110 142554
rect 2162 142502 2174 142554
rect 2226 142502 5152 142554
rect 1104 142480 5152 142502
rect 84180 142554 90896 142576
rect 84180 142502 85982 142554
rect 86034 142502 86046 142554
rect 86098 142502 86110 142554
rect 86162 142502 86174 142554
rect 86226 142502 89982 142554
rect 90034 142502 90046 142554
rect 90098 142502 90110 142554
rect 90162 142502 90174 142554
rect 90226 142502 90896 142554
rect 84180 142480 90896 142502
rect 85850 142400 85856 142452
rect 85908 142440 85914 142452
rect 87966 142440 87972 142452
rect 85908 142412 87972 142440
rect 85908 142400 85914 142412
rect 87966 142400 87972 142412
rect 88024 142400 88030 142452
rect 1104 142010 5152 142032
rect 1104 141958 3982 142010
rect 4034 141958 4046 142010
rect 4098 141958 4110 142010
rect 4162 141958 4174 142010
rect 4226 141958 5152 142010
rect 1104 141936 5152 141958
rect 84180 142010 90896 142032
rect 84180 141958 87982 142010
rect 88034 141958 88046 142010
rect 88098 141958 88110 142010
rect 88162 141958 88174 142010
rect 88226 141958 90896 142010
rect 84180 141936 90896 141958
rect 1104 141466 5152 141488
rect 1104 141414 1982 141466
rect 2034 141414 2046 141466
rect 2098 141414 2110 141466
rect 2162 141414 2174 141466
rect 2226 141414 5152 141466
rect 1104 141392 5152 141414
rect 84180 141466 90896 141488
rect 84180 141414 85982 141466
rect 86034 141414 86046 141466
rect 86098 141414 86110 141466
rect 86162 141414 86174 141466
rect 86226 141414 89982 141466
rect 90034 141414 90046 141466
rect 90098 141414 90110 141466
rect 90162 141414 90174 141466
rect 90226 141414 90896 141466
rect 84180 141392 90896 141414
rect 84194 141176 84200 141228
rect 84252 141216 84258 141228
rect 87966 141216 87972 141228
rect 84252 141188 87972 141216
rect 84252 141176 84258 141188
rect 87966 141176 87972 141188
rect 88024 141176 88030 141228
rect 84933 141151 84991 141157
rect 84933 141117 84945 141151
rect 84979 141148 84991 141151
rect 84979 141120 85252 141148
rect 84979 141117 84991 141120
rect 84933 141111 84991 141117
rect 84654 141080 84660 141092
rect 84615 141052 84660 141080
rect 84654 141040 84660 141052
rect 84712 141040 84718 141092
rect 85224 141024 85252 141120
rect 85206 141012 85212 141024
rect 85167 140984 85212 141012
rect 85206 140972 85212 140984
rect 85264 140972 85270 141024
rect 1104 140922 5152 140944
rect 1104 140870 3982 140922
rect 4034 140870 4046 140922
rect 4098 140870 4110 140922
rect 4162 140870 4174 140922
rect 4226 140870 5152 140922
rect 1104 140848 5152 140870
rect 84180 140922 90896 140944
rect 84180 140870 87982 140922
rect 88034 140870 88046 140922
rect 88098 140870 88110 140922
rect 88162 140870 88174 140922
rect 88226 140870 90896 140922
rect 84180 140848 90896 140870
rect 1104 140378 5152 140400
rect 1104 140326 1982 140378
rect 2034 140326 2046 140378
rect 2098 140326 2110 140378
rect 2162 140326 2174 140378
rect 2226 140326 5152 140378
rect 1104 140304 5152 140326
rect 84180 140378 90896 140400
rect 84180 140326 85982 140378
rect 86034 140326 86046 140378
rect 86098 140326 86110 140378
rect 86162 140326 86174 140378
rect 86226 140326 89982 140378
rect 90034 140326 90046 140378
rect 90098 140326 90110 140378
rect 90162 140326 90174 140378
rect 90226 140326 90896 140378
rect 84180 140304 90896 140326
rect 85114 139952 85120 140004
rect 85172 139992 85178 140004
rect 88242 139992 88248 140004
rect 85172 139964 88248 139992
rect 85172 139952 85178 139964
rect 88242 139952 88248 139964
rect 88300 139952 88306 140004
rect 1104 139834 5152 139856
rect 1104 139782 3982 139834
rect 4034 139782 4046 139834
rect 4098 139782 4110 139834
rect 4162 139782 4174 139834
rect 4226 139782 5152 139834
rect 1104 139760 5152 139782
rect 84180 139834 90896 139856
rect 84180 139782 87982 139834
rect 88034 139782 88046 139834
rect 88098 139782 88110 139834
rect 88162 139782 88174 139834
rect 88226 139782 90896 139834
rect 84180 139760 90896 139782
rect 1104 139290 5152 139312
rect 1104 139238 1982 139290
rect 2034 139238 2046 139290
rect 2098 139238 2110 139290
rect 2162 139238 2174 139290
rect 2226 139238 5152 139290
rect 1104 139216 5152 139238
rect 84180 139290 90896 139312
rect 84180 139238 85982 139290
rect 86034 139238 86046 139290
rect 86098 139238 86110 139290
rect 86162 139238 86174 139290
rect 86226 139238 89982 139290
rect 90034 139238 90046 139290
rect 90098 139238 90110 139290
rect 90162 139238 90174 139290
rect 90226 139238 90896 139290
rect 84180 139216 90896 139238
rect 84838 138864 84844 138916
rect 84896 138904 84902 138916
rect 88058 138904 88064 138916
rect 84896 138876 88064 138904
rect 84896 138864 84902 138876
rect 88058 138864 88064 138876
rect 88116 138864 88122 138916
rect 1104 138746 5152 138768
rect 1104 138694 3982 138746
rect 4034 138694 4046 138746
rect 4098 138694 4110 138746
rect 4162 138694 4174 138746
rect 4226 138694 5152 138746
rect 1104 138672 5152 138694
rect 84180 138746 90896 138768
rect 84180 138694 87982 138746
rect 88034 138694 88046 138746
rect 88098 138694 88110 138746
rect 88162 138694 88174 138746
rect 88226 138694 90896 138746
rect 84180 138672 90896 138694
rect 1104 138202 5152 138224
rect 1104 138150 1982 138202
rect 2034 138150 2046 138202
rect 2098 138150 2110 138202
rect 2162 138150 2174 138202
rect 2226 138150 5152 138202
rect 1104 138128 5152 138150
rect 84180 138202 90896 138224
rect 84180 138150 85982 138202
rect 86034 138150 86046 138202
rect 86098 138150 86110 138202
rect 86162 138150 86174 138202
rect 86226 138150 89982 138202
rect 90034 138150 90046 138202
rect 90098 138150 90110 138202
rect 90162 138150 90174 138202
rect 90226 138150 90896 138202
rect 84180 138128 90896 138150
rect 1104 137658 5152 137680
rect 1104 137606 3982 137658
rect 4034 137606 4046 137658
rect 4098 137606 4110 137658
rect 4162 137606 4174 137658
rect 4226 137606 5152 137658
rect 1104 137584 5152 137606
rect 84180 137658 90896 137680
rect 84180 137606 87982 137658
rect 88034 137606 88046 137658
rect 88098 137606 88110 137658
rect 88162 137606 88174 137658
rect 88226 137606 90896 137658
rect 84180 137584 90896 137606
rect 1104 137114 5152 137136
rect 1104 137062 1982 137114
rect 2034 137062 2046 137114
rect 2098 137062 2110 137114
rect 2162 137062 2174 137114
rect 2226 137062 5152 137114
rect 1104 137040 5152 137062
rect 84180 137114 90896 137136
rect 84180 137062 85982 137114
rect 86034 137062 86046 137114
rect 86098 137062 86110 137114
rect 86162 137062 86174 137114
rect 86226 137062 89982 137114
rect 90034 137062 90046 137114
rect 90098 137062 90110 137114
rect 90162 137062 90174 137114
rect 90226 137062 90896 137114
rect 84180 137040 90896 137062
rect 1104 136570 5152 136592
rect 1104 136518 3982 136570
rect 4034 136518 4046 136570
rect 4098 136518 4110 136570
rect 4162 136518 4174 136570
rect 4226 136518 5152 136570
rect 1104 136496 5152 136518
rect 84180 136570 90896 136592
rect 84180 136518 87982 136570
rect 88034 136518 88046 136570
rect 88098 136518 88110 136570
rect 88162 136518 88174 136570
rect 88226 136518 90896 136570
rect 84180 136496 90896 136518
rect 1104 136026 5152 136048
rect 1104 135974 1982 136026
rect 2034 135974 2046 136026
rect 2098 135974 2110 136026
rect 2162 135974 2174 136026
rect 2226 135974 5152 136026
rect 1104 135952 5152 135974
rect 84180 136026 90896 136048
rect 84180 135974 85982 136026
rect 86034 135974 86046 136026
rect 86098 135974 86110 136026
rect 86162 135974 86174 136026
rect 86226 135974 89982 136026
rect 90034 135974 90046 136026
rect 90098 135974 90110 136026
rect 90162 135974 90174 136026
rect 90226 135974 90896 136026
rect 84180 135952 90896 135974
rect 1104 135482 5152 135504
rect 1104 135430 3982 135482
rect 4034 135430 4046 135482
rect 4098 135430 4110 135482
rect 4162 135430 4174 135482
rect 4226 135430 5152 135482
rect 1104 135408 5152 135430
rect 84180 135482 90896 135504
rect 84180 135430 87982 135482
rect 88034 135430 88046 135482
rect 88098 135430 88110 135482
rect 88162 135430 88174 135482
rect 88226 135430 90896 135482
rect 84180 135408 90896 135430
rect 1104 134938 5152 134960
rect 1104 134886 1982 134938
rect 2034 134886 2046 134938
rect 2098 134886 2110 134938
rect 2162 134886 2174 134938
rect 2226 134886 5152 134938
rect 1104 134864 5152 134886
rect 84180 134938 90896 134960
rect 84180 134886 85982 134938
rect 86034 134886 86046 134938
rect 86098 134886 86110 134938
rect 86162 134886 86174 134938
rect 86226 134886 89982 134938
rect 90034 134886 90046 134938
rect 90098 134886 90110 134938
rect 90162 134886 90174 134938
rect 90226 134886 90896 134938
rect 84180 134864 90896 134886
rect 1104 134394 5152 134416
rect 1104 134342 3982 134394
rect 4034 134342 4046 134394
rect 4098 134342 4110 134394
rect 4162 134342 4174 134394
rect 4226 134342 5152 134394
rect 1104 134320 5152 134342
rect 84180 134394 90896 134416
rect 84180 134342 87982 134394
rect 88034 134342 88046 134394
rect 88098 134342 88110 134394
rect 88162 134342 88174 134394
rect 88226 134342 90896 134394
rect 84180 134320 90896 134342
rect 1104 133850 5152 133872
rect 1104 133798 1982 133850
rect 2034 133798 2046 133850
rect 2098 133798 2110 133850
rect 2162 133798 2174 133850
rect 2226 133798 5152 133850
rect 1104 133776 5152 133798
rect 84180 133850 90896 133872
rect 84180 133798 85982 133850
rect 86034 133798 86046 133850
rect 86098 133798 86110 133850
rect 86162 133798 86174 133850
rect 86226 133798 89982 133850
rect 90034 133798 90046 133850
rect 90098 133798 90110 133850
rect 90162 133798 90174 133850
rect 90226 133798 90896 133850
rect 84180 133776 90896 133798
rect 1104 133306 5152 133328
rect 1104 133254 3982 133306
rect 4034 133254 4046 133306
rect 4098 133254 4110 133306
rect 4162 133254 4174 133306
rect 4226 133254 5152 133306
rect 1104 133232 5152 133254
rect 84180 133306 90896 133328
rect 84180 133254 87982 133306
rect 88034 133254 88046 133306
rect 88098 133254 88110 133306
rect 88162 133254 88174 133306
rect 88226 133254 90896 133306
rect 84180 133232 90896 133254
rect 1104 132762 5152 132784
rect 1104 132710 1982 132762
rect 2034 132710 2046 132762
rect 2098 132710 2110 132762
rect 2162 132710 2174 132762
rect 2226 132710 5152 132762
rect 1104 132688 5152 132710
rect 84180 132762 90896 132784
rect 84180 132710 85982 132762
rect 86034 132710 86046 132762
rect 86098 132710 86110 132762
rect 86162 132710 86174 132762
rect 86226 132710 89982 132762
rect 90034 132710 90046 132762
rect 90098 132710 90110 132762
rect 90162 132710 90174 132762
rect 90226 132710 90896 132762
rect 84180 132688 90896 132710
rect 1104 132218 5152 132240
rect 1104 132166 3982 132218
rect 4034 132166 4046 132218
rect 4098 132166 4110 132218
rect 4162 132166 4174 132218
rect 4226 132166 5152 132218
rect 1104 132144 5152 132166
rect 84180 132218 90896 132240
rect 84180 132166 87982 132218
rect 88034 132166 88046 132218
rect 88098 132166 88110 132218
rect 88162 132166 88174 132218
rect 88226 132166 90896 132218
rect 84180 132144 90896 132166
rect 1104 131674 5152 131696
rect 1104 131622 1982 131674
rect 2034 131622 2046 131674
rect 2098 131622 2110 131674
rect 2162 131622 2174 131674
rect 2226 131622 5152 131674
rect 1104 131600 5152 131622
rect 84180 131674 90896 131696
rect 84180 131622 85982 131674
rect 86034 131622 86046 131674
rect 86098 131622 86110 131674
rect 86162 131622 86174 131674
rect 86226 131622 89982 131674
rect 90034 131622 90046 131674
rect 90098 131622 90110 131674
rect 90162 131622 90174 131674
rect 90226 131622 90896 131674
rect 84180 131600 90896 131622
rect 85574 131248 85580 131300
rect 85632 131288 85638 131300
rect 88242 131288 88248 131300
rect 85632 131260 88248 131288
rect 85632 131248 85638 131260
rect 88242 131248 88248 131260
rect 88300 131248 88306 131300
rect 84930 131180 84936 131232
rect 84988 131220 84994 131232
rect 85850 131220 85856 131232
rect 84988 131192 85856 131220
rect 84988 131180 84994 131192
rect 85850 131180 85856 131192
rect 85908 131180 85914 131232
rect 1104 131130 5152 131152
rect 1104 131078 3982 131130
rect 4034 131078 4046 131130
rect 4098 131078 4110 131130
rect 4162 131078 4174 131130
rect 4226 131078 5152 131130
rect 1104 131056 5152 131078
rect 84180 131130 90896 131152
rect 84180 131078 87982 131130
rect 88034 131078 88046 131130
rect 88098 131078 88110 131130
rect 88162 131078 88174 131130
rect 88226 131078 90896 131130
rect 84180 131056 90896 131078
rect 1104 130586 5152 130608
rect 1104 130534 1982 130586
rect 2034 130534 2046 130586
rect 2098 130534 2110 130586
rect 2162 130534 2174 130586
rect 2226 130534 5152 130586
rect 1104 130512 5152 130534
rect 84180 130586 90896 130608
rect 84180 130534 85982 130586
rect 86034 130534 86046 130586
rect 86098 130534 86110 130586
rect 86162 130534 86174 130586
rect 86226 130534 89982 130586
rect 90034 130534 90046 130586
rect 90098 130534 90110 130586
rect 90162 130534 90174 130586
rect 90226 130534 90896 130586
rect 84180 130512 90896 130534
rect 1104 130042 5152 130064
rect 1104 129990 3982 130042
rect 4034 129990 4046 130042
rect 4098 129990 4110 130042
rect 4162 129990 4174 130042
rect 4226 129990 5152 130042
rect 1104 129968 5152 129990
rect 84180 130042 90896 130064
rect 84180 129990 87982 130042
rect 88034 129990 88046 130042
rect 88098 129990 88110 130042
rect 88162 129990 88174 130042
rect 88226 129990 90896 130042
rect 84180 129968 90896 129990
rect 1104 129498 5152 129520
rect 1104 129446 1982 129498
rect 2034 129446 2046 129498
rect 2098 129446 2110 129498
rect 2162 129446 2174 129498
rect 2226 129446 5152 129498
rect 1104 129424 5152 129446
rect 84180 129498 90896 129520
rect 84180 129446 85982 129498
rect 86034 129446 86046 129498
rect 86098 129446 86110 129498
rect 86162 129446 86174 129498
rect 86226 129446 89982 129498
rect 90034 129446 90046 129498
rect 90098 129446 90110 129498
rect 90162 129446 90174 129498
rect 90226 129446 90896 129498
rect 84180 129424 90896 129446
rect 1104 128954 5152 128976
rect 1104 128902 3982 128954
rect 4034 128902 4046 128954
rect 4098 128902 4110 128954
rect 4162 128902 4174 128954
rect 4226 128902 5152 128954
rect 1104 128880 5152 128902
rect 84180 128954 90896 128976
rect 84180 128902 87982 128954
rect 88034 128902 88046 128954
rect 88098 128902 88110 128954
rect 88162 128902 88174 128954
rect 88226 128902 90896 128954
rect 84180 128880 90896 128902
rect 84010 128460 84016 128512
rect 84068 128500 84074 128512
rect 88242 128500 88248 128512
rect 84068 128472 88248 128500
rect 84068 128460 84074 128472
rect 88242 128460 88248 128472
rect 88300 128460 88306 128512
rect 1104 128410 5152 128432
rect 1104 128358 1982 128410
rect 2034 128358 2046 128410
rect 2098 128358 2110 128410
rect 2162 128358 2174 128410
rect 2226 128358 5152 128410
rect 1104 128336 5152 128358
rect 84180 128410 90896 128432
rect 84180 128358 85982 128410
rect 86034 128358 86046 128410
rect 86098 128358 86110 128410
rect 86162 128358 86174 128410
rect 86226 128358 89982 128410
rect 90034 128358 90046 128410
rect 90098 128358 90110 128410
rect 90162 128358 90174 128410
rect 90226 128358 90896 128410
rect 84180 128336 90896 128358
rect 1104 127866 5152 127888
rect 1104 127814 3982 127866
rect 4034 127814 4046 127866
rect 4098 127814 4110 127866
rect 4162 127814 4174 127866
rect 4226 127814 5152 127866
rect 1104 127792 5152 127814
rect 84180 127866 90896 127888
rect 84180 127814 87982 127866
rect 88034 127814 88046 127866
rect 88098 127814 88110 127866
rect 88162 127814 88174 127866
rect 88226 127814 90896 127866
rect 84180 127792 90896 127814
rect 1104 127322 5152 127344
rect 1104 127270 1982 127322
rect 2034 127270 2046 127322
rect 2098 127270 2110 127322
rect 2162 127270 2174 127322
rect 2226 127270 5152 127322
rect 1104 127248 5152 127270
rect 84180 127322 90896 127344
rect 84180 127270 85982 127322
rect 86034 127270 86046 127322
rect 86098 127270 86110 127322
rect 86162 127270 86174 127322
rect 86226 127270 89982 127322
rect 90034 127270 90046 127322
rect 90098 127270 90110 127322
rect 90162 127270 90174 127322
rect 90226 127270 90896 127322
rect 84180 127248 90896 127270
rect 83366 126964 83372 127016
rect 83424 127004 83430 127016
rect 88242 127004 88248 127016
rect 83424 126976 88248 127004
rect 83424 126964 83430 126976
rect 88242 126964 88248 126976
rect 88300 126964 88306 127016
rect 1104 126778 5152 126800
rect 1104 126726 3982 126778
rect 4034 126726 4046 126778
rect 4098 126726 4110 126778
rect 4162 126726 4174 126778
rect 4226 126726 5152 126778
rect 1104 126704 5152 126726
rect 84180 126778 90896 126800
rect 84180 126726 87982 126778
rect 88034 126726 88046 126778
rect 88098 126726 88110 126778
rect 88162 126726 88174 126778
rect 88226 126726 90896 126778
rect 84180 126704 90896 126726
rect 1104 126234 5152 126256
rect 1104 126182 1982 126234
rect 2034 126182 2046 126234
rect 2098 126182 2110 126234
rect 2162 126182 2174 126234
rect 2226 126182 5152 126234
rect 1104 126160 5152 126182
rect 84180 126234 90896 126256
rect 84180 126182 85982 126234
rect 86034 126182 86046 126234
rect 86098 126182 86110 126234
rect 86162 126182 86174 126234
rect 86226 126182 89982 126234
rect 90034 126182 90046 126234
rect 90098 126182 90110 126234
rect 90162 126182 90174 126234
rect 90226 126182 90896 126234
rect 84180 126160 90896 126182
rect 83274 125808 83280 125860
rect 83332 125848 83338 125860
rect 87966 125848 87972 125860
rect 83332 125820 87972 125848
rect 83332 125808 83338 125820
rect 87966 125808 87972 125820
rect 88024 125808 88030 125860
rect 84562 125740 84568 125792
rect 84620 125780 84626 125792
rect 84657 125783 84715 125789
rect 84657 125780 84669 125783
rect 84620 125752 84669 125780
rect 84620 125740 84626 125752
rect 84657 125749 84669 125752
rect 84703 125749 84715 125783
rect 84657 125743 84715 125749
rect 1104 125690 5152 125712
rect 1104 125638 3982 125690
rect 4034 125638 4046 125690
rect 4098 125638 4110 125690
rect 4162 125638 4174 125690
rect 4226 125638 5152 125690
rect 1104 125616 5152 125638
rect 84180 125690 90896 125712
rect 84180 125638 87982 125690
rect 88034 125638 88046 125690
rect 88098 125638 88110 125690
rect 88162 125638 88174 125690
rect 88226 125638 90896 125690
rect 84180 125616 90896 125638
rect 1104 125146 5152 125168
rect 1104 125094 1982 125146
rect 2034 125094 2046 125146
rect 2098 125094 2110 125146
rect 2162 125094 2174 125146
rect 2226 125094 5152 125146
rect 1104 125072 5152 125094
rect 84180 125146 90896 125168
rect 84180 125094 85982 125146
rect 86034 125094 86046 125146
rect 86098 125094 86110 125146
rect 86162 125094 86174 125146
rect 86226 125094 89982 125146
rect 90034 125094 90046 125146
rect 90098 125094 90110 125146
rect 90162 125094 90174 125146
rect 90226 125094 90896 125146
rect 84180 125072 90896 125094
rect 1104 124602 5152 124624
rect 1104 124550 3982 124602
rect 4034 124550 4046 124602
rect 4098 124550 4110 124602
rect 4162 124550 4174 124602
rect 4226 124550 5152 124602
rect 1104 124528 5152 124550
rect 84180 124602 90896 124624
rect 84180 124550 87982 124602
rect 88034 124550 88046 124602
rect 88098 124550 88110 124602
rect 88162 124550 88174 124602
rect 88226 124550 90896 124602
rect 84180 124528 90896 124550
rect 84470 124448 84476 124500
rect 84528 124488 84534 124500
rect 84657 124491 84715 124497
rect 84657 124488 84669 124491
rect 84528 124460 84669 124488
rect 84528 124448 84534 124460
rect 84657 124457 84669 124460
rect 84703 124457 84715 124491
rect 84657 124451 84715 124457
rect 1104 124058 5152 124080
rect 1104 124006 1982 124058
rect 2034 124006 2046 124058
rect 2098 124006 2110 124058
rect 2162 124006 2174 124058
rect 2226 124006 5152 124058
rect 1104 123984 5152 124006
rect 84180 124058 90896 124080
rect 84180 124006 85982 124058
rect 86034 124006 86046 124058
rect 86098 124006 86110 124058
rect 86162 124006 86174 124058
rect 86226 124006 89982 124058
rect 90034 124006 90046 124058
rect 90098 124006 90110 124058
rect 90162 124006 90174 124058
rect 90226 124006 90896 124058
rect 84180 123984 90896 124006
rect 1104 123514 5152 123536
rect 1104 123462 3982 123514
rect 4034 123462 4046 123514
rect 4098 123462 4110 123514
rect 4162 123462 4174 123514
rect 4226 123462 5152 123514
rect 1104 123440 5152 123462
rect 84180 123514 90896 123536
rect 84180 123462 87982 123514
rect 88034 123462 88046 123514
rect 88098 123462 88110 123514
rect 88162 123462 88174 123514
rect 88226 123462 90896 123514
rect 84180 123440 90896 123462
rect 84378 123360 84384 123412
rect 84436 123400 84442 123412
rect 84657 123403 84715 123409
rect 84657 123400 84669 123403
rect 84436 123372 84669 123400
rect 84436 123360 84442 123372
rect 84657 123369 84669 123372
rect 84703 123369 84715 123403
rect 84657 123363 84715 123369
rect 1104 122970 5152 122992
rect 1104 122918 1982 122970
rect 2034 122918 2046 122970
rect 2098 122918 2110 122970
rect 2162 122918 2174 122970
rect 2226 122918 5152 122970
rect 1104 122896 5152 122918
rect 84180 122970 90896 122992
rect 84180 122918 85982 122970
rect 86034 122918 86046 122970
rect 86098 122918 86110 122970
rect 86162 122918 86174 122970
rect 86226 122918 89982 122970
rect 90034 122918 90046 122970
rect 90098 122918 90110 122970
rect 90162 122918 90174 122970
rect 90226 122918 90896 122970
rect 84180 122896 90896 122918
rect 83182 122816 83188 122868
rect 83240 122856 83246 122868
rect 87966 122856 87972 122868
rect 83240 122828 87972 122856
rect 83240 122816 83246 122828
rect 87966 122816 87972 122828
rect 88024 122816 88030 122868
rect 1104 122426 5152 122448
rect 1104 122374 3982 122426
rect 4034 122374 4046 122426
rect 4098 122374 4110 122426
rect 4162 122374 4174 122426
rect 4226 122374 5152 122426
rect 1104 122352 5152 122374
rect 84180 122426 90896 122448
rect 84180 122374 87982 122426
rect 88034 122374 88046 122426
rect 88098 122374 88110 122426
rect 88162 122374 88174 122426
rect 88226 122374 90896 122426
rect 84180 122352 90896 122374
rect 87230 122136 87236 122188
rect 87288 122176 87294 122188
rect 87874 122176 87880 122188
rect 87288 122148 87880 122176
rect 87288 122136 87294 122148
rect 87874 122136 87880 122148
rect 87932 122136 87938 122188
rect 1104 121882 5152 121904
rect 1104 121830 1982 121882
rect 2034 121830 2046 121882
rect 2098 121830 2110 121882
rect 2162 121830 2174 121882
rect 2226 121830 5152 121882
rect 1104 121808 5152 121830
rect 84180 121882 90896 121904
rect 84180 121830 85982 121882
rect 86034 121830 86046 121882
rect 86098 121830 86110 121882
rect 86162 121830 86174 121882
rect 86226 121830 89982 121882
rect 90034 121830 90046 121882
rect 90098 121830 90110 121882
rect 90162 121830 90174 121882
rect 90226 121830 90896 121882
rect 84180 121808 90896 121830
rect 83090 121456 83096 121508
rect 83148 121496 83154 121508
rect 87874 121496 87880 121508
rect 83148 121468 87880 121496
rect 83148 121456 83154 121468
rect 87874 121456 87880 121468
rect 87932 121456 87938 121508
rect 1104 121338 5152 121360
rect 1104 121286 3982 121338
rect 4034 121286 4046 121338
rect 4098 121286 4110 121338
rect 4162 121286 4174 121338
rect 4226 121286 5152 121338
rect 1104 121264 5152 121286
rect 84180 121338 90896 121360
rect 84180 121286 87982 121338
rect 88034 121286 88046 121338
rect 88098 121286 88110 121338
rect 88162 121286 88174 121338
rect 88226 121286 90896 121338
rect 84180 121264 90896 121286
rect 84470 120844 84476 120896
rect 84528 120884 84534 120896
rect 84657 120887 84715 120893
rect 84657 120884 84669 120887
rect 84528 120856 84669 120884
rect 84528 120844 84534 120856
rect 84657 120853 84669 120856
rect 84703 120853 84715 120887
rect 84657 120847 84715 120853
rect 1104 120794 5152 120816
rect 1104 120742 1982 120794
rect 2034 120742 2046 120794
rect 2098 120742 2110 120794
rect 2162 120742 2174 120794
rect 2226 120742 5152 120794
rect 1104 120720 5152 120742
rect 84180 120794 90896 120816
rect 84180 120742 85982 120794
rect 86034 120742 86046 120794
rect 86098 120742 86110 120794
rect 86162 120742 86174 120794
rect 86226 120742 89982 120794
rect 90034 120742 90046 120794
rect 90098 120742 90110 120794
rect 90162 120742 90174 120794
rect 90226 120742 90896 120794
rect 84180 120720 90896 120742
rect 1104 120250 5152 120272
rect 1104 120198 3982 120250
rect 4034 120198 4046 120250
rect 4098 120198 4110 120250
rect 4162 120198 4174 120250
rect 4226 120198 5152 120250
rect 1104 120176 5152 120198
rect 84180 120250 90896 120272
rect 84180 120198 87982 120250
rect 88034 120198 88046 120250
rect 88098 120198 88110 120250
rect 88162 120198 88174 120250
rect 88226 120198 90896 120250
rect 84180 120176 90896 120198
rect 82998 120096 83004 120148
rect 83056 120136 83062 120148
rect 87874 120136 87880 120148
rect 83056 120108 87880 120136
rect 83056 120096 83062 120108
rect 87874 120096 87880 120108
rect 87932 120096 87938 120148
rect 84562 120028 84568 120080
rect 84620 120068 84626 120080
rect 84657 120071 84715 120077
rect 84657 120068 84669 120071
rect 84620 120040 84669 120068
rect 84620 120028 84626 120040
rect 84657 120037 84669 120040
rect 84703 120037 84715 120071
rect 84657 120031 84715 120037
rect 1104 119706 5152 119728
rect 1104 119654 1982 119706
rect 2034 119654 2046 119706
rect 2098 119654 2110 119706
rect 2162 119654 2174 119706
rect 2226 119654 5152 119706
rect 1104 119632 5152 119654
rect 84180 119706 90896 119728
rect 84180 119654 85982 119706
rect 86034 119654 86046 119706
rect 86098 119654 86110 119706
rect 86162 119654 86174 119706
rect 86226 119654 89982 119706
rect 90034 119654 90046 119706
rect 90098 119654 90110 119706
rect 90162 119654 90174 119706
rect 90226 119654 90896 119706
rect 84180 119632 90896 119654
rect 1104 119162 5152 119184
rect 1104 119110 3982 119162
rect 4034 119110 4046 119162
rect 4098 119110 4110 119162
rect 4162 119110 4174 119162
rect 4226 119110 5152 119162
rect 1104 119088 5152 119110
rect 84180 119162 90896 119184
rect 84180 119110 87982 119162
rect 88034 119110 88046 119162
rect 88098 119110 88110 119162
rect 88162 119110 88174 119162
rect 88226 119110 90896 119162
rect 84180 119088 90896 119110
rect 82906 118668 82912 118720
rect 82964 118708 82970 118720
rect 87874 118708 87880 118720
rect 82964 118680 87880 118708
rect 82964 118668 82970 118680
rect 87874 118668 87880 118680
rect 87932 118668 87938 118720
rect 1104 118618 5152 118640
rect 1104 118566 1982 118618
rect 2034 118566 2046 118618
rect 2098 118566 2110 118618
rect 2162 118566 2174 118618
rect 2226 118566 5152 118618
rect 1104 118544 5152 118566
rect 84180 118618 90896 118640
rect 84180 118566 85982 118618
rect 86034 118566 86046 118618
rect 86098 118566 86110 118618
rect 86162 118566 86174 118618
rect 86226 118566 89982 118618
rect 90034 118566 90046 118618
rect 90098 118566 90110 118618
rect 90162 118566 90174 118618
rect 90226 118566 90896 118618
rect 84180 118544 90896 118566
rect 84378 118124 84384 118176
rect 84436 118164 84442 118176
rect 84657 118167 84715 118173
rect 84657 118164 84669 118167
rect 84436 118136 84669 118164
rect 84436 118124 84442 118136
rect 84657 118133 84669 118136
rect 84703 118133 84715 118167
rect 84657 118127 84715 118133
rect 1104 118074 5152 118096
rect 1104 118022 3982 118074
rect 4034 118022 4046 118074
rect 4098 118022 4110 118074
rect 4162 118022 4174 118074
rect 4226 118022 5152 118074
rect 1104 118000 5152 118022
rect 84180 118074 90896 118096
rect 84180 118022 87982 118074
rect 88034 118022 88046 118074
rect 88098 118022 88110 118074
rect 88162 118022 88174 118074
rect 88226 118022 90896 118074
rect 84180 118000 90896 118022
rect 1104 117530 5152 117552
rect 1104 117478 1982 117530
rect 2034 117478 2046 117530
rect 2098 117478 2110 117530
rect 2162 117478 2174 117530
rect 2226 117478 5152 117530
rect 1104 117456 5152 117478
rect 84180 117530 90896 117552
rect 84180 117478 85982 117530
rect 86034 117478 86046 117530
rect 86098 117478 86110 117530
rect 86162 117478 86174 117530
rect 86226 117478 89982 117530
rect 90034 117478 90046 117530
rect 90098 117478 90110 117530
rect 90162 117478 90174 117530
rect 90226 117478 90896 117530
rect 84180 117456 90896 117478
rect 84562 117036 84568 117088
rect 84620 117076 84626 117088
rect 84657 117079 84715 117085
rect 84657 117076 84669 117079
rect 84620 117048 84669 117076
rect 84620 117036 84626 117048
rect 84657 117045 84669 117048
rect 84703 117045 84715 117079
rect 84657 117039 84715 117045
rect 1104 116986 5152 117008
rect 1104 116934 3982 116986
rect 4034 116934 4046 116986
rect 4098 116934 4110 116986
rect 4162 116934 4174 116986
rect 4226 116934 5152 116986
rect 1104 116912 5152 116934
rect 84180 116986 90896 117008
rect 84180 116934 87982 116986
rect 88034 116934 88046 116986
rect 88098 116934 88110 116986
rect 88162 116934 88174 116986
rect 88226 116934 90896 116986
rect 84180 116912 90896 116934
rect 4801 116603 4859 116609
rect 4801 116569 4813 116603
rect 4847 116600 4859 116603
rect 5350 116600 5356 116612
rect 4847 116572 5356 116600
rect 4847 116569 4859 116572
rect 4801 116563 4859 116569
rect 5350 116560 5356 116572
rect 5408 116560 5414 116612
rect 1104 116442 5152 116464
rect 1104 116390 1982 116442
rect 2034 116390 2046 116442
rect 2098 116390 2110 116442
rect 2162 116390 2174 116442
rect 2226 116390 5152 116442
rect 1104 116368 5152 116390
rect 84180 116442 90896 116464
rect 84180 116390 85982 116442
rect 86034 116390 86046 116442
rect 86098 116390 86110 116442
rect 86162 116390 86174 116442
rect 86226 116390 89982 116442
rect 90034 116390 90046 116442
rect 90098 116390 90110 116442
rect 90162 116390 90174 116442
rect 90226 116390 90896 116442
rect 84180 116368 90896 116390
rect 1104 115898 5152 115920
rect 1104 115846 3982 115898
rect 4034 115846 4046 115898
rect 4098 115846 4110 115898
rect 4162 115846 4174 115898
rect 4226 115846 5152 115898
rect 1104 115824 5152 115846
rect 84180 115898 90896 115920
rect 84180 115846 87982 115898
rect 88034 115846 88046 115898
rect 88098 115846 88110 115898
rect 88162 115846 88174 115898
rect 88226 115846 90896 115898
rect 84180 115824 90896 115846
rect 1104 115354 5152 115376
rect 1104 115302 1982 115354
rect 2034 115302 2046 115354
rect 2098 115302 2110 115354
rect 2162 115302 2174 115354
rect 2226 115302 5152 115354
rect 1104 115280 5152 115302
rect 84180 115354 90896 115376
rect 84180 115302 85982 115354
rect 86034 115302 86046 115354
rect 86098 115302 86110 115354
rect 86162 115302 86174 115354
rect 86226 115302 89982 115354
rect 90034 115302 90046 115354
rect 90098 115302 90110 115354
rect 90162 115302 90174 115354
rect 90226 115302 90896 115354
rect 84180 115280 90896 115302
rect 4801 114971 4859 114977
rect 4801 114937 4813 114971
rect 4847 114968 4859 114971
rect 5442 114968 5448 114980
rect 4847 114940 5448 114968
rect 4847 114937 4859 114940
rect 4801 114931 4859 114937
rect 5442 114928 5448 114940
rect 5500 114928 5506 114980
rect 1104 114810 5152 114832
rect 1104 114758 3982 114810
rect 4034 114758 4046 114810
rect 4098 114758 4110 114810
rect 4162 114758 4174 114810
rect 4226 114758 5152 114810
rect 1104 114736 5152 114758
rect 84180 114810 90896 114832
rect 84180 114758 87982 114810
rect 88034 114758 88046 114810
rect 88098 114758 88110 114810
rect 88162 114758 88174 114810
rect 88226 114758 90896 114810
rect 84180 114736 90896 114758
rect 85666 114520 85672 114572
rect 85724 114560 85730 114572
rect 87966 114560 87972 114572
rect 85724 114532 87972 114560
rect 85724 114520 85730 114532
rect 87966 114520 87972 114532
rect 88024 114520 88030 114572
rect 1104 114266 5152 114288
rect 1104 114214 1982 114266
rect 2034 114214 2046 114266
rect 2098 114214 2110 114266
rect 2162 114214 2174 114266
rect 2226 114214 5152 114266
rect 1104 114192 5152 114214
rect 84180 114266 90896 114288
rect 84180 114214 85982 114266
rect 86034 114214 86046 114266
rect 86098 114214 86110 114266
rect 86162 114214 86174 114266
rect 86226 114214 89982 114266
rect 90034 114214 90046 114266
rect 90098 114214 90110 114266
rect 90162 114214 90174 114266
rect 90226 114214 90896 114266
rect 84180 114192 90896 114214
rect 85390 113840 85396 113892
rect 85448 113880 85454 113892
rect 86494 113880 86500 113892
rect 85448 113852 86500 113880
rect 85448 113840 85454 113852
rect 86494 113840 86500 113852
rect 86552 113840 86558 113892
rect 1104 113722 5152 113744
rect 1104 113670 3982 113722
rect 4034 113670 4046 113722
rect 4098 113670 4110 113722
rect 4162 113670 4174 113722
rect 4226 113670 5152 113722
rect 1104 113648 5152 113670
rect 84180 113722 90896 113744
rect 84180 113670 87982 113722
rect 88034 113670 88046 113722
rect 88098 113670 88110 113722
rect 88162 113670 88174 113722
rect 88226 113670 90896 113722
rect 84180 113648 90896 113670
rect 1104 113178 5152 113200
rect 1104 113126 1982 113178
rect 2034 113126 2046 113178
rect 2098 113126 2110 113178
rect 2162 113126 2174 113178
rect 2226 113126 5152 113178
rect 1104 113104 5152 113126
rect 84180 113178 90896 113200
rect 84180 113126 85982 113178
rect 86034 113126 86046 113178
rect 86098 113126 86110 113178
rect 86162 113126 86174 113178
rect 86226 113126 89982 113178
rect 90034 113126 90046 113178
rect 90098 113126 90110 113178
rect 90162 113126 90174 113178
rect 90226 113126 90896 113178
rect 84180 113104 90896 113126
rect 1104 112634 5152 112656
rect 1104 112582 3982 112634
rect 4034 112582 4046 112634
rect 4098 112582 4110 112634
rect 4162 112582 4174 112634
rect 4226 112582 5152 112634
rect 1104 112560 5152 112582
rect 84180 112634 90896 112656
rect 84180 112582 87982 112634
rect 88034 112582 88046 112634
rect 88098 112582 88110 112634
rect 88162 112582 88174 112634
rect 88226 112582 90896 112634
rect 84180 112560 90896 112582
rect 1104 112090 5152 112112
rect 1104 112038 1982 112090
rect 2034 112038 2046 112090
rect 2098 112038 2110 112090
rect 2162 112038 2174 112090
rect 2226 112038 5152 112090
rect 1104 112016 5152 112038
rect 84180 112090 90896 112112
rect 84180 112038 85982 112090
rect 86034 112038 86046 112090
rect 86098 112038 86110 112090
rect 86162 112038 86174 112090
rect 86226 112038 89982 112090
rect 90034 112038 90046 112090
rect 90098 112038 90110 112090
rect 90162 112038 90174 112090
rect 90226 112038 90896 112090
rect 84180 112016 90896 112038
rect 85298 111800 85304 111852
rect 85356 111840 85362 111852
rect 87966 111840 87972 111852
rect 85356 111812 87972 111840
rect 85356 111800 85362 111812
rect 87966 111800 87972 111812
rect 88024 111800 88030 111852
rect 1104 111546 5152 111568
rect 1104 111494 3982 111546
rect 4034 111494 4046 111546
rect 4098 111494 4110 111546
rect 4162 111494 4174 111546
rect 4226 111494 5152 111546
rect 1104 111472 5152 111494
rect 84180 111546 90896 111568
rect 84180 111494 87982 111546
rect 88034 111494 88046 111546
rect 88098 111494 88110 111546
rect 88162 111494 88174 111546
rect 88226 111494 90896 111546
rect 84180 111472 90896 111494
rect 1104 111002 5152 111024
rect 1104 110950 1982 111002
rect 2034 110950 2046 111002
rect 2098 110950 2110 111002
rect 2162 110950 2174 111002
rect 2226 110950 5152 111002
rect 1104 110928 5152 110950
rect 84180 111002 90896 111024
rect 84180 110950 85982 111002
rect 86034 110950 86046 111002
rect 86098 110950 86110 111002
rect 86162 110950 86174 111002
rect 86226 110950 89982 111002
rect 90034 110950 90046 111002
rect 90098 110950 90110 111002
rect 90162 110950 90174 111002
rect 90226 110950 90896 111002
rect 84180 110928 90896 110950
rect 1104 110458 5152 110480
rect 1104 110406 3982 110458
rect 4034 110406 4046 110458
rect 4098 110406 4110 110458
rect 4162 110406 4174 110458
rect 4226 110406 5152 110458
rect 1104 110384 5152 110406
rect 84180 110458 90896 110480
rect 84180 110406 87982 110458
rect 88034 110406 88046 110458
rect 88098 110406 88110 110458
rect 88162 110406 88174 110458
rect 88226 110406 90896 110458
rect 84180 110384 90896 110406
rect 82538 110304 82544 110356
rect 82596 110344 82602 110356
rect 85482 110344 85488 110356
rect 82596 110316 85488 110344
rect 82596 110304 82602 110316
rect 85482 110304 85488 110316
rect 85540 110304 85546 110356
rect 1104 109914 5152 109936
rect 1104 109862 1982 109914
rect 2034 109862 2046 109914
rect 2098 109862 2110 109914
rect 2162 109862 2174 109914
rect 2226 109862 5152 109914
rect 1104 109840 5152 109862
rect 84180 109914 90896 109936
rect 84180 109862 85982 109914
rect 86034 109862 86046 109914
rect 86098 109862 86110 109914
rect 86162 109862 86174 109914
rect 86226 109862 89982 109914
rect 90034 109862 90046 109914
rect 90098 109862 90110 109914
rect 90162 109862 90174 109914
rect 90226 109862 90896 109914
rect 84180 109840 90896 109862
rect 85206 109556 85212 109608
rect 85264 109596 85270 109608
rect 85850 109596 85856 109608
rect 85264 109568 85856 109596
rect 85264 109556 85270 109568
rect 85850 109556 85856 109568
rect 85908 109556 85914 109608
rect 1104 109370 5152 109392
rect 1104 109318 3982 109370
rect 4034 109318 4046 109370
rect 4098 109318 4110 109370
rect 4162 109318 4174 109370
rect 4226 109318 5152 109370
rect 1104 109296 5152 109318
rect 84180 109370 90896 109392
rect 84180 109318 87982 109370
rect 88034 109318 88046 109370
rect 88098 109318 88110 109370
rect 88162 109318 88174 109370
rect 88226 109318 90896 109370
rect 84180 109296 90896 109318
rect 84286 108944 84292 108996
rect 84344 108984 84350 108996
rect 85942 108984 85948 108996
rect 84344 108956 85948 108984
rect 84344 108944 84350 108956
rect 85942 108944 85948 108956
rect 86000 108944 86006 108996
rect 1104 108826 5152 108848
rect 1104 108774 1982 108826
rect 2034 108774 2046 108826
rect 2098 108774 2110 108826
rect 2162 108774 2174 108826
rect 2226 108774 5152 108826
rect 1104 108752 5152 108774
rect 84180 108826 90896 108848
rect 84180 108774 85982 108826
rect 86034 108774 86046 108826
rect 86098 108774 86110 108826
rect 86162 108774 86174 108826
rect 86226 108774 89982 108826
rect 90034 108774 90046 108826
rect 90098 108774 90110 108826
rect 90162 108774 90174 108826
rect 90226 108774 90896 108826
rect 84180 108752 90896 108774
rect 85206 108604 85212 108656
rect 85264 108644 85270 108656
rect 87966 108644 87972 108656
rect 85264 108616 87972 108644
rect 85264 108604 85270 108616
rect 87966 108604 87972 108616
rect 88024 108604 88030 108656
rect 87598 108536 87604 108588
rect 87656 108576 87662 108588
rect 88334 108576 88340 108588
rect 87656 108548 88340 108576
rect 87656 108536 87662 108548
rect 88334 108536 88340 108548
rect 88392 108536 88398 108588
rect 87230 108468 87236 108520
rect 87288 108508 87294 108520
rect 88518 108508 88524 108520
rect 87288 108480 88524 108508
rect 87288 108468 87294 108480
rect 88518 108468 88524 108480
rect 88576 108468 88582 108520
rect 87598 108400 87604 108452
rect 87656 108440 87662 108452
rect 88242 108440 88248 108452
rect 87656 108412 88248 108440
rect 87656 108400 87662 108412
rect 88242 108400 88248 108412
rect 88300 108400 88306 108452
rect 1104 108282 5152 108304
rect 1104 108230 3982 108282
rect 4034 108230 4046 108282
rect 4098 108230 4110 108282
rect 4162 108230 4174 108282
rect 4226 108230 5152 108282
rect 1104 108208 5152 108230
rect 84180 108282 90896 108304
rect 84180 108230 87982 108282
rect 88034 108230 88046 108282
rect 88098 108230 88110 108282
rect 88162 108230 88174 108282
rect 88226 108230 90896 108282
rect 84180 108208 90896 108230
rect 1104 107738 5152 107760
rect 1104 107686 1982 107738
rect 2034 107686 2046 107738
rect 2098 107686 2110 107738
rect 2162 107686 2174 107738
rect 2226 107686 5152 107738
rect 1104 107664 5152 107686
rect 84180 107738 90896 107760
rect 84180 107686 85982 107738
rect 86034 107686 86046 107738
rect 86098 107686 86110 107738
rect 86162 107686 86174 107738
rect 86226 107686 89982 107738
rect 90034 107686 90046 107738
rect 90098 107686 90110 107738
rect 90162 107686 90174 107738
rect 90226 107686 90896 107738
rect 84180 107664 90896 107686
rect 83642 107312 83648 107364
rect 83700 107352 83706 107364
rect 87966 107352 87972 107364
rect 83700 107324 87972 107352
rect 83700 107312 83706 107324
rect 87966 107312 87972 107324
rect 88024 107312 88030 107364
rect 1104 107194 5152 107216
rect 1104 107142 3982 107194
rect 4034 107142 4046 107194
rect 4098 107142 4110 107194
rect 4162 107142 4174 107194
rect 4226 107142 5152 107194
rect 1104 107120 5152 107142
rect 84180 107194 90896 107216
rect 84180 107142 87982 107194
rect 88034 107142 88046 107194
rect 88098 107142 88110 107194
rect 88162 107142 88174 107194
rect 88226 107142 90896 107194
rect 84180 107120 90896 107142
rect 1104 106650 5152 106672
rect 1104 106598 1982 106650
rect 2034 106598 2046 106650
rect 2098 106598 2110 106650
rect 2162 106598 2174 106650
rect 2226 106598 5152 106650
rect 1104 106576 5152 106598
rect 84180 106650 90896 106672
rect 84180 106598 85982 106650
rect 86034 106598 86046 106650
rect 86098 106598 86110 106650
rect 86162 106598 86174 106650
rect 86226 106598 89982 106650
rect 90034 106598 90046 106650
rect 90098 106598 90110 106650
rect 90162 106598 90174 106650
rect 90226 106598 90896 106650
rect 84180 106576 90896 106598
rect 86310 106496 86316 106548
rect 86368 106496 86374 106548
rect 86328 106344 86356 106496
rect 86310 106292 86316 106344
rect 86368 106292 86374 106344
rect 1104 106106 5152 106128
rect 1104 106054 3982 106106
rect 4034 106054 4046 106106
rect 4098 106054 4110 106106
rect 4162 106054 4174 106106
rect 4226 106054 5152 106106
rect 1104 106032 5152 106054
rect 84180 106106 90896 106128
rect 84180 106054 87982 106106
rect 88034 106054 88046 106106
rect 88098 106054 88110 106106
rect 88162 106054 88174 106106
rect 88226 106054 90896 106106
rect 84180 106032 90896 106054
rect 4430 105856 4436 105868
rect 4391 105828 4436 105856
rect 4430 105816 4436 105828
rect 4488 105816 4494 105868
rect 84013 105723 84071 105729
rect 84013 105689 84025 105723
rect 84059 105720 84071 105723
rect 86218 105720 86224 105732
rect 84059 105692 86224 105720
rect 84059 105689 84071 105692
rect 84013 105683 84071 105689
rect 86218 105680 86224 105692
rect 86276 105680 86282 105732
rect 1104 105562 5152 105584
rect 1104 105510 1982 105562
rect 2034 105510 2046 105562
rect 2098 105510 2110 105562
rect 2162 105510 2174 105562
rect 2226 105510 5152 105562
rect 1104 105488 5152 105510
rect 84180 105562 90896 105584
rect 84180 105510 85982 105562
rect 86034 105510 86046 105562
rect 86098 105510 86110 105562
rect 86162 105510 86174 105562
rect 86226 105510 89982 105562
rect 90034 105510 90046 105562
rect 90098 105510 90110 105562
rect 90162 105510 90174 105562
rect 90226 105510 90896 105562
rect 84180 105488 90896 105510
rect 1104 105018 5152 105040
rect 1104 104966 3982 105018
rect 4034 104966 4046 105018
rect 4098 104966 4110 105018
rect 4162 104966 4174 105018
rect 4226 104966 5152 105018
rect 1104 104944 5152 104966
rect 84180 105018 90896 105040
rect 84180 104966 87982 105018
rect 88034 104966 88046 105018
rect 88098 104966 88110 105018
rect 88162 104966 88174 105018
rect 88226 104966 90896 105018
rect 84180 104944 90896 104966
rect 85482 104524 85488 104576
rect 85540 104564 85546 104576
rect 86402 104564 86408 104576
rect 85540 104536 86408 104564
rect 85540 104524 85546 104536
rect 86402 104524 86408 104536
rect 86460 104524 86466 104576
rect 86494 104524 86500 104576
rect 86552 104564 86558 104576
rect 86678 104564 86684 104576
rect 86552 104536 86684 104564
rect 86552 104524 86558 104536
rect 86678 104524 86684 104536
rect 86736 104524 86742 104576
rect 1104 104474 5152 104496
rect 1104 104422 1982 104474
rect 2034 104422 2046 104474
rect 2098 104422 2110 104474
rect 2162 104422 2174 104474
rect 2226 104422 5152 104474
rect 1104 104400 5152 104422
rect 84180 104474 90896 104496
rect 84180 104422 85982 104474
rect 86034 104422 86046 104474
rect 86098 104422 86110 104474
rect 86162 104422 86174 104474
rect 86226 104422 89982 104474
rect 90034 104422 90046 104474
rect 90098 104422 90110 104474
rect 90162 104422 90174 104474
rect 90226 104422 90896 104474
rect 84180 104400 90896 104422
rect 83461 104363 83519 104369
rect 83461 104329 83473 104363
rect 83507 104360 83519 104363
rect 86862 104360 86868 104372
rect 83507 104332 86868 104360
rect 83507 104329 83519 104332
rect 83461 104323 83519 104329
rect 86862 104320 86868 104332
rect 86920 104320 86926 104372
rect 87322 104360 87328 104372
rect 87156 104332 87328 104360
rect 82909 104295 82967 104301
rect 82909 104261 82921 104295
rect 82955 104292 82967 104295
rect 85666 104292 85672 104304
rect 82955 104264 85672 104292
rect 82955 104261 82967 104264
rect 82909 104255 82967 104261
rect 85666 104252 85672 104264
rect 85724 104252 85730 104304
rect 86586 104184 86592 104236
rect 86644 104224 86650 104236
rect 86862 104224 86868 104236
rect 86644 104196 86868 104224
rect 86644 104184 86650 104196
rect 86862 104184 86868 104196
rect 86920 104184 86926 104236
rect 87156 104168 87184 104332
rect 87322 104320 87328 104332
rect 87380 104320 87386 104372
rect 87782 104320 87788 104372
rect 87840 104360 87846 104372
rect 88702 104360 88708 104372
rect 87840 104332 88708 104360
rect 87840 104320 87846 104332
rect 88702 104320 88708 104332
rect 88760 104320 88766 104372
rect 87138 104116 87144 104168
rect 87196 104116 87202 104168
rect 1104 103930 5152 103952
rect 1104 103878 3982 103930
rect 4034 103878 4046 103930
rect 4098 103878 4110 103930
rect 4162 103878 4174 103930
rect 4226 103878 5152 103930
rect 1104 103856 5152 103878
rect 84180 103930 90896 103952
rect 84180 103878 87982 103930
rect 88034 103878 88046 103930
rect 88098 103878 88110 103930
rect 88162 103878 88174 103930
rect 88226 103878 90896 103930
rect 84180 103856 90896 103878
rect 1104 103386 5152 103408
rect 1104 103334 1982 103386
rect 2034 103334 2046 103386
rect 2098 103334 2110 103386
rect 2162 103334 2174 103386
rect 2226 103334 5152 103386
rect 1104 103312 5152 103334
rect 84180 103386 90896 103408
rect 84180 103334 85982 103386
rect 86034 103334 86046 103386
rect 86098 103334 86110 103386
rect 86162 103334 86174 103386
rect 86226 103334 89982 103386
rect 90034 103334 90046 103386
rect 90098 103334 90110 103386
rect 90162 103334 90174 103386
rect 90226 103334 90896 103386
rect 84180 103312 90896 103334
rect 1104 102842 5152 102864
rect 1104 102790 3982 102842
rect 4034 102790 4046 102842
rect 4098 102790 4110 102842
rect 4162 102790 4174 102842
rect 4226 102790 5152 102842
rect 1104 102768 5152 102790
rect 84180 102842 90896 102864
rect 84180 102790 87982 102842
rect 88034 102790 88046 102842
rect 88098 102790 88110 102842
rect 88162 102790 88174 102842
rect 88226 102790 90896 102842
rect 84180 102768 90896 102790
rect 1104 102298 5152 102320
rect 1104 102246 1982 102298
rect 2034 102246 2046 102298
rect 2098 102246 2110 102298
rect 2162 102246 2174 102298
rect 2226 102246 5152 102298
rect 1104 102224 5152 102246
rect 84180 102298 90896 102320
rect 84180 102246 85982 102298
rect 86034 102246 86046 102298
rect 86098 102246 86110 102298
rect 86162 102246 86174 102298
rect 86226 102246 89982 102298
rect 90034 102246 90046 102298
rect 90098 102246 90110 102298
rect 90162 102246 90174 102298
rect 90226 102246 90896 102298
rect 84180 102224 90896 102246
rect 1104 101754 5152 101776
rect 1104 101702 3982 101754
rect 4034 101702 4046 101754
rect 4098 101702 4110 101754
rect 4162 101702 4174 101754
rect 4226 101702 5152 101754
rect 1104 101680 5152 101702
rect 84180 101754 90896 101776
rect 84180 101702 87982 101754
rect 88034 101702 88046 101754
rect 88098 101702 88110 101754
rect 88162 101702 88174 101754
rect 88226 101702 90896 101754
rect 84180 101680 90896 101702
rect 1104 101210 5152 101232
rect 1104 101158 1982 101210
rect 2034 101158 2046 101210
rect 2098 101158 2110 101210
rect 2162 101158 2174 101210
rect 2226 101158 5152 101210
rect 1104 101136 5152 101158
rect 84180 101210 90896 101232
rect 84180 101158 85982 101210
rect 86034 101158 86046 101210
rect 86098 101158 86110 101210
rect 86162 101158 86174 101210
rect 86226 101158 89982 101210
rect 90034 101158 90046 101210
rect 90098 101158 90110 101210
rect 90162 101158 90174 101210
rect 90226 101158 90896 101210
rect 84180 101136 90896 101158
rect 87874 101056 87880 101108
rect 87932 101096 87938 101108
rect 88426 101096 88432 101108
rect 87932 101068 88432 101096
rect 87932 101056 87938 101068
rect 88426 101056 88432 101068
rect 88484 101056 88490 101108
rect 1104 100666 5152 100688
rect 1104 100614 3982 100666
rect 4034 100614 4046 100666
rect 4098 100614 4110 100666
rect 4162 100614 4174 100666
rect 4226 100614 5152 100666
rect 1104 100592 5152 100614
rect 84180 100666 90896 100688
rect 84180 100614 87982 100666
rect 88034 100614 88046 100666
rect 88098 100614 88110 100666
rect 88162 100614 88174 100666
rect 88226 100614 90896 100666
rect 84180 100592 90896 100614
rect 1104 100122 5152 100144
rect 1104 100070 1982 100122
rect 2034 100070 2046 100122
rect 2098 100070 2110 100122
rect 2162 100070 2174 100122
rect 2226 100070 5152 100122
rect 1104 100048 5152 100070
rect 84180 100122 90896 100144
rect 84180 100070 85982 100122
rect 86034 100070 86046 100122
rect 86098 100070 86110 100122
rect 86162 100070 86174 100122
rect 86226 100070 89982 100122
rect 90034 100070 90046 100122
rect 90098 100070 90110 100122
rect 90162 100070 90174 100122
rect 90226 100070 90896 100122
rect 84180 100048 90896 100070
rect 85758 99968 85764 100020
rect 85816 100008 85822 100020
rect 86402 100008 86408 100020
rect 85816 99980 86408 100008
rect 85816 99968 85822 99980
rect 86402 99968 86408 99980
rect 86460 99968 86466 100020
rect 86126 99900 86132 99952
rect 86184 99940 86190 99952
rect 86678 99940 86684 99952
rect 86184 99912 86684 99940
rect 86184 99900 86190 99912
rect 86678 99900 86684 99912
rect 86736 99900 86742 99952
rect 87230 99900 87236 99952
rect 87288 99940 87294 99952
rect 88610 99940 88616 99952
rect 87288 99912 88616 99940
rect 87288 99900 87294 99912
rect 88610 99900 88616 99912
rect 88668 99900 88674 99952
rect 85850 99832 85856 99884
rect 85908 99872 85914 99884
rect 86218 99872 86224 99884
rect 85908 99844 86224 99872
rect 85908 99832 85914 99844
rect 86218 99832 86224 99844
rect 86276 99832 86282 99884
rect 87598 99832 87604 99884
rect 87656 99872 87662 99884
rect 88426 99872 88432 99884
rect 87656 99844 88432 99872
rect 87656 99832 87662 99844
rect 88426 99832 88432 99844
rect 88484 99832 88490 99884
rect 88518 99804 88524 99816
rect 86880 99776 88524 99804
rect 86880 99680 86908 99776
rect 88518 99764 88524 99776
rect 88576 99764 88582 99816
rect 87598 99696 87604 99748
rect 87656 99736 87662 99748
rect 87874 99736 87880 99748
rect 87656 99708 87880 99736
rect 87656 99696 87662 99708
rect 87874 99696 87880 99708
rect 87932 99696 87938 99748
rect 85022 99628 85028 99680
rect 85080 99668 85086 99680
rect 85390 99668 85396 99680
rect 85080 99640 85396 99668
rect 85080 99628 85086 99640
rect 85390 99628 85396 99640
rect 85448 99628 85454 99680
rect 85482 99628 85488 99680
rect 85540 99668 85546 99680
rect 85666 99668 85672 99680
rect 85540 99640 85672 99668
rect 85540 99628 85546 99640
rect 85666 99628 85672 99640
rect 85724 99628 85730 99680
rect 86862 99628 86868 99680
rect 86920 99628 86926 99680
rect 1104 99578 5152 99600
rect 1104 99526 3982 99578
rect 4034 99526 4046 99578
rect 4098 99526 4110 99578
rect 4162 99526 4174 99578
rect 4226 99526 5152 99578
rect 1104 99504 5152 99526
rect 84180 99578 90896 99600
rect 84180 99526 87982 99578
rect 88034 99526 88046 99578
rect 88098 99526 88110 99578
rect 88162 99526 88174 99578
rect 88226 99526 90896 99578
rect 84180 99504 90896 99526
rect 85390 99424 85396 99476
rect 85448 99464 85454 99476
rect 86494 99464 86500 99476
rect 85448 99436 86500 99464
rect 85448 99424 85454 99436
rect 86494 99424 86500 99436
rect 86552 99424 86558 99476
rect 85574 99356 85580 99408
rect 85632 99396 85638 99408
rect 86126 99396 86132 99408
rect 85632 99368 86132 99396
rect 85632 99356 85638 99368
rect 86126 99356 86132 99368
rect 86184 99356 86190 99408
rect 82722 99288 82728 99340
rect 82780 99328 82786 99340
rect 87414 99328 87420 99340
rect 82780 99300 87420 99328
rect 82780 99288 82786 99300
rect 87414 99288 87420 99300
rect 87472 99288 87478 99340
rect 85390 99220 85396 99272
rect 85448 99260 85454 99272
rect 85850 99260 85856 99272
rect 85448 99232 85856 99260
rect 85448 99220 85454 99232
rect 85850 99220 85856 99232
rect 85908 99220 85914 99272
rect 87506 99260 87512 99272
rect 85960 99232 87512 99260
rect 82541 99195 82599 99201
rect 82541 99161 82553 99195
rect 82587 99192 82599 99195
rect 85960 99192 85988 99232
rect 87506 99220 87512 99232
rect 87564 99220 87570 99272
rect 82587 99164 85988 99192
rect 82587 99161 82599 99164
rect 82541 99155 82599 99161
rect 87414 99152 87420 99204
rect 87472 99192 87478 99204
rect 88426 99192 88432 99204
rect 87472 99164 88432 99192
rect 87472 99152 87478 99164
rect 88426 99152 88432 99164
rect 88484 99152 88490 99204
rect 87506 99084 87512 99136
rect 87564 99124 87570 99136
rect 88610 99124 88616 99136
rect 87564 99096 88616 99124
rect 87564 99084 87570 99096
rect 88610 99084 88616 99096
rect 88668 99084 88674 99136
rect 1104 99034 5152 99056
rect 1104 98982 1982 99034
rect 2034 98982 2046 99034
rect 2098 98982 2110 99034
rect 2162 98982 2174 99034
rect 2226 98982 5152 99034
rect 1104 98960 5152 98982
rect 84180 99034 90896 99056
rect 84180 98982 85982 99034
rect 86034 98982 86046 99034
rect 86098 98982 86110 99034
rect 86162 98982 86174 99034
rect 86226 98982 89982 99034
rect 90034 98982 90046 99034
rect 90098 98982 90110 99034
rect 90162 98982 90174 99034
rect 90226 98982 90896 99034
rect 84180 98960 90896 98982
rect 83001 98923 83059 98929
rect 83001 98889 83013 98923
rect 83047 98920 83059 98923
rect 87598 98920 87604 98932
rect 83047 98892 87604 98920
rect 83047 98889 83059 98892
rect 83001 98883 83059 98889
rect 87598 98880 87604 98892
rect 87656 98880 87662 98932
rect 87690 98880 87696 98932
rect 87748 98920 87754 98932
rect 87874 98920 87880 98932
rect 87748 98892 87880 98920
rect 87748 98880 87754 98892
rect 87874 98880 87880 98892
rect 87932 98880 87938 98932
rect 87782 98676 87788 98728
rect 87840 98716 87846 98728
rect 88334 98716 88340 98728
rect 87840 98688 88340 98716
rect 87840 98676 87846 98688
rect 88334 98676 88340 98688
rect 88392 98676 88398 98728
rect 4338 98580 4344 98592
rect 4299 98552 4344 98580
rect 4338 98540 4344 98552
rect 4396 98540 4402 98592
rect 4801 98583 4859 98589
rect 4801 98549 4813 98583
rect 4847 98580 4859 98583
rect 6730 98580 6736 98592
rect 4847 98552 6736 98580
rect 4847 98549 4859 98552
rect 4801 98543 4859 98549
rect 6730 98540 6736 98552
rect 6788 98540 6794 98592
rect 1104 98490 5152 98512
rect 1104 98438 3982 98490
rect 4034 98438 4046 98490
rect 4098 98438 4110 98490
rect 4162 98438 4174 98490
rect 4226 98438 5152 98490
rect 1104 98416 5152 98438
rect 84180 98490 90896 98512
rect 84180 98438 87982 98490
rect 88034 98438 88046 98490
rect 88098 98438 88110 98490
rect 88162 98438 88174 98490
rect 88226 98438 90896 98490
rect 84180 98416 90896 98438
rect 82722 98308 82728 98320
rect 82683 98280 82728 98308
rect 82722 98268 82728 98280
rect 82780 98268 82786 98320
rect 82722 98132 82728 98184
rect 82780 98172 82786 98184
rect 87230 98172 87236 98184
rect 82780 98144 87236 98172
rect 82780 98132 82786 98144
rect 87230 98132 87236 98144
rect 87288 98132 87294 98184
rect 3697 98107 3755 98113
rect 3697 98073 3709 98107
rect 3743 98104 3755 98107
rect 6822 98104 6828 98116
rect 3743 98076 6828 98104
rect 3743 98073 3755 98076
rect 3697 98067 3755 98073
rect 6822 98064 6828 98076
rect 6880 98064 6886 98116
rect 83458 98064 83464 98116
rect 83516 98104 83522 98116
rect 86954 98104 86960 98116
rect 83516 98076 86960 98104
rect 83516 98064 83522 98076
rect 86954 98064 86960 98076
rect 87012 98064 87018 98116
rect 4430 98036 4436 98048
rect 4391 98008 4436 98036
rect 4430 97996 4436 98008
rect 4488 97996 4494 98048
rect 4522 97996 4528 98048
rect 4580 98036 4586 98048
rect 4709 98039 4767 98045
rect 4709 98036 4721 98039
rect 4580 98008 4721 98036
rect 4580 97996 4586 98008
rect 4709 98005 4721 98008
rect 4755 98036 4767 98039
rect 5350 98036 5356 98048
rect 4755 98008 5356 98036
rect 4755 98005 4767 98008
rect 4709 97999 4767 98005
rect 5350 97996 5356 98008
rect 5408 97996 5414 98048
rect 83645 98039 83703 98045
rect 83645 98005 83657 98039
rect 83691 98036 83703 98039
rect 84657 98039 84715 98045
rect 84657 98036 84669 98039
rect 83691 98008 84669 98036
rect 83691 98005 83703 98008
rect 83645 97999 83703 98005
rect 84657 98005 84669 98008
rect 84703 98036 84715 98039
rect 84930 98036 84936 98048
rect 84703 98008 84936 98036
rect 84703 98005 84715 98008
rect 84657 97999 84715 98005
rect 84930 97996 84936 98008
rect 84988 97996 84994 98048
rect 1104 97946 5152 97968
rect 1104 97894 1982 97946
rect 2034 97894 2046 97946
rect 2098 97894 2110 97946
rect 2162 97894 2174 97946
rect 2226 97894 5152 97946
rect 1104 97872 5152 97894
rect 84180 97946 90896 97968
rect 84180 97894 85982 97946
rect 86034 97894 86046 97946
rect 86098 97894 86110 97946
rect 86162 97894 86174 97946
rect 86226 97894 89982 97946
rect 90034 97894 90046 97946
rect 90098 97894 90110 97946
rect 90162 97894 90174 97946
rect 90226 97894 90896 97946
rect 84180 97872 90896 97894
rect 2590 97792 2596 97844
rect 2648 97832 2654 97844
rect 6825 97835 6883 97841
rect 6825 97832 6837 97835
rect 2648 97804 6837 97832
rect 2648 97792 2654 97804
rect 6825 97801 6837 97804
rect 6871 97801 6883 97835
rect 84838 97832 84844 97844
rect 84799 97804 84844 97832
rect 6825 97795 6883 97801
rect 84838 97792 84844 97804
rect 84896 97792 84902 97844
rect 85117 97835 85175 97841
rect 85117 97801 85129 97835
rect 85163 97832 85175 97835
rect 85390 97832 85396 97844
rect 85163 97804 85396 97832
rect 85163 97801 85175 97804
rect 85117 97795 85175 97801
rect 85390 97792 85396 97804
rect 85448 97792 85454 97844
rect 3697 97767 3755 97773
rect 3697 97733 3709 97767
rect 3743 97764 3755 97767
rect 5810 97764 5816 97776
rect 3743 97736 5816 97764
rect 3743 97733 3755 97736
rect 3697 97727 3755 97733
rect 5810 97724 5816 97736
rect 5868 97724 5874 97776
rect 4065 97699 4123 97705
rect 4065 97665 4077 97699
rect 4111 97696 4123 97699
rect 5718 97696 5724 97708
rect 4111 97668 5724 97696
rect 4111 97665 4123 97668
rect 4065 97659 4123 97665
rect 5718 97656 5724 97668
rect 5776 97656 5782 97708
rect 87874 97656 87880 97708
rect 87932 97696 87938 97708
rect 90358 97696 90364 97708
rect 87932 97668 90364 97696
rect 87932 97656 87938 97668
rect 90358 97656 90364 97668
rect 90416 97656 90422 97708
rect 4433 97631 4491 97637
rect 4433 97597 4445 97631
rect 4479 97628 4491 97631
rect 5261 97631 5319 97637
rect 5261 97628 5273 97631
rect 4479 97600 5273 97628
rect 4479 97597 4491 97600
rect 4433 97591 4491 97597
rect 5261 97597 5273 97600
rect 5307 97597 5319 97631
rect 5261 97591 5319 97597
rect 82817 97631 82875 97637
rect 82817 97597 82829 97631
rect 82863 97628 82875 97631
rect 87966 97628 87972 97640
rect 82863 97600 87972 97628
rect 82863 97597 82875 97600
rect 82817 97591 82875 97597
rect 87966 97588 87972 97600
rect 88024 97588 88030 97640
rect 2961 97563 3019 97569
rect 2961 97529 2973 97563
rect 3007 97560 3019 97563
rect 82633 97563 82691 97569
rect 3007 97532 6684 97560
rect 3007 97529 3019 97532
rect 2961 97523 3019 97529
rect 3326 97492 3332 97504
rect 3287 97464 3332 97492
rect 3326 97452 3332 97464
rect 3384 97452 3390 97504
rect 4801 97495 4859 97501
rect 4801 97461 4813 97495
rect 4847 97492 4859 97495
rect 5626 97492 5632 97504
rect 4847 97464 5632 97492
rect 4847 97461 4859 97464
rect 4801 97455 4859 97461
rect 5626 97452 5632 97464
rect 5684 97452 5690 97504
rect 1104 97402 5152 97424
rect 1104 97350 3982 97402
rect 4034 97350 4046 97402
rect 4098 97350 4110 97402
rect 4162 97350 4174 97402
rect 4226 97350 5152 97402
rect 1104 97328 5152 97350
rect 2590 97288 2596 97300
rect 2551 97260 2596 97288
rect 2590 97248 2596 97260
rect 2648 97248 2654 97300
rect 3329 97291 3387 97297
rect 3329 97257 3341 97291
rect 3375 97288 3387 97291
rect 5902 97288 5908 97300
rect 3375 97260 5908 97288
rect 3375 97257 3387 97260
rect 3329 97251 3387 97257
rect 5902 97248 5908 97260
rect 5960 97248 5966 97300
rect 3602 97180 3608 97232
rect 3660 97220 3666 97232
rect 3697 97223 3755 97229
rect 3697 97220 3709 97223
rect 3660 97192 3709 97220
rect 3660 97180 3666 97192
rect 3697 97189 3709 97192
rect 3743 97220 3755 97223
rect 6549 97223 6607 97229
rect 6549 97220 6561 97223
rect 3743 97192 6561 97220
rect 3743 97189 3755 97192
rect 3697 97183 3755 97189
rect 6549 97189 6561 97192
rect 6595 97189 6607 97223
rect 6656 97220 6684 97532
rect 82633 97529 82645 97563
rect 82679 97560 82691 97563
rect 87690 97560 87696 97572
rect 82679 97532 87696 97560
rect 82679 97529 82691 97532
rect 82633 97523 82691 97529
rect 87690 97520 87696 97532
rect 87748 97520 87754 97572
rect 84286 97452 84292 97504
rect 84344 97492 84350 97504
rect 84657 97495 84715 97501
rect 84657 97492 84669 97495
rect 84344 97464 84669 97492
rect 84344 97452 84350 97464
rect 84657 97461 84669 97464
rect 84703 97461 84715 97495
rect 84838 97492 84844 97504
rect 84799 97464 84844 97492
rect 84657 97455 84715 97461
rect 84838 97452 84844 97464
rect 84896 97452 84902 97504
rect 82449 97427 82507 97433
rect 82449 97393 82461 97427
rect 82495 97424 82507 97427
rect 82495 97396 83596 97424
rect 82495 97393 82507 97396
rect 82449 97387 82507 97393
rect 6730 97316 6736 97368
rect 6788 97356 6794 97368
rect 15933 97359 15991 97365
rect 6788 97328 15884 97356
rect 6788 97316 6794 97328
rect 7009 97291 7067 97297
rect 7009 97257 7021 97291
rect 7055 97288 7067 97291
rect 15856 97288 15884 97328
rect 15933 97325 15945 97359
rect 15979 97356 15991 97359
rect 83458 97356 83464 97368
rect 15979 97328 83464 97356
rect 15979 97325 15991 97328
rect 15933 97319 15991 97325
rect 83458 97316 83464 97328
rect 83516 97316 83522 97368
rect 83568 97365 83596 97396
rect 84180 97402 90896 97424
rect 83553 97359 83611 97365
rect 83553 97325 83565 97359
rect 83599 97356 83611 97359
rect 83599 97328 84148 97356
rect 84180 97350 87982 97402
rect 88034 97350 88046 97402
rect 88098 97350 88110 97402
rect 88162 97350 88174 97402
rect 88226 97350 90896 97402
rect 84180 97328 90896 97350
rect 83599 97325 83611 97328
rect 83553 97319 83611 97325
rect 22833 97291 22891 97297
rect 22833 97288 22845 97291
rect 7055 97260 15792 97288
rect 15856 97260 22845 97288
rect 7055 97257 7067 97260
rect 7009 97251 7067 97257
rect 15657 97223 15715 97229
rect 15657 97220 15669 97223
rect 6656 97192 15669 97220
rect 6549 97183 6607 97189
rect 15657 97189 15669 97192
rect 15703 97189 15715 97223
rect 15764 97220 15792 97260
rect 22833 97257 22845 97260
rect 22879 97257 22891 97291
rect 22833 97251 22891 97257
rect 22922 97248 22928 97300
rect 22980 97288 22986 97300
rect 83001 97291 83059 97297
rect 83001 97288 83013 97291
rect 22980 97260 83013 97288
rect 22980 97248 22986 97260
rect 83001 97257 83013 97260
rect 83047 97257 83059 97291
rect 84120 97288 84148 97328
rect 84657 97291 84715 97297
rect 84657 97288 84669 97291
rect 84120 97260 84669 97288
rect 83001 97251 83059 97257
rect 84657 97257 84669 97260
rect 84703 97257 84715 97291
rect 84657 97251 84715 97257
rect 84746 97248 84752 97300
rect 84804 97288 84810 97300
rect 86954 97288 86960 97300
rect 84804 97260 86960 97288
rect 84804 97248 84810 97260
rect 86954 97248 86960 97260
rect 87012 97248 87018 97300
rect 21910 97220 21916 97232
rect 15764 97192 21916 97220
rect 15657 97183 15715 97189
rect 21910 97180 21916 97192
rect 21968 97180 21974 97232
rect 22005 97223 22063 97229
rect 22005 97189 22017 97223
rect 22051 97220 22063 97223
rect 86770 97220 86776 97232
rect 22051 97192 86776 97220
rect 22051 97189 22063 97192
rect 22005 97183 22063 97189
rect 86770 97180 86776 97192
rect 86828 97180 86834 97232
rect 5074 97112 5080 97164
rect 5132 97152 5138 97164
rect 86954 97152 86960 97164
rect 5132 97124 86960 97152
rect 5132 97112 5138 97124
rect 86954 97112 86960 97124
rect 87012 97112 87018 97164
rect 4433 97087 4491 97093
rect 4433 97053 4445 97087
rect 4479 97084 4491 97087
rect 5534 97084 5540 97096
rect 4479 97056 5540 97084
rect 4479 97053 4491 97056
rect 4433 97047 4491 97053
rect 5534 97044 5540 97056
rect 5592 97084 5598 97096
rect 18046 97084 18052 97096
rect 5592 97056 18052 97084
rect 5592 97044 5598 97056
rect 18046 97044 18052 97056
rect 18104 97084 18110 97096
rect 83642 97084 83648 97096
rect 18104 97056 83648 97084
rect 18104 97044 18110 97056
rect 83642 97044 83648 97056
rect 83700 97044 83706 97096
rect 84013 97087 84071 97093
rect 84013 97053 84025 97087
rect 84059 97084 84071 97087
rect 85025 97087 85083 97093
rect 85025 97084 85037 97087
rect 84059 97056 85037 97084
rect 84059 97053 84071 97056
rect 84013 97047 84071 97053
rect 85025 97053 85037 97056
rect 85071 97053 85083 97087
rect 85025 97047 85083 97053
rect 85853 97087 85911 97093
rect 85853 97053 85865 97087
rect 85899 97084 85911 97087
rect 86402 97084 86408 97096
rect 85899 97056 86408 97084
rect 85899 97053 85911 97056
rect 85853 97047 85911 97053
rect 86402 97044 86408 97056
rect 86460 97044 86466 97096
rect 86770 97044 86776 97096
rect 86828 97084 86834 97096
rect 87138 97084 87144 97096
rect 86828 97056 87144 97084
rect 86828 97044 86834 97056
rect 87138 97044 87144 97056
rect 87196 97044 87202 97096
rect 2225 97019 2283 97025
rect 2225 96985 2237 97019
rect 2271 97016 2283 97019
rect 14642 97016 14648 97028
rect 2271 96988 14648 97016
rect 2271 96985 2283 96988
rect 2225 96979 2283 96985
rect 14642 96976 14648 96988
rect 14700 97016 14706 97028
rect 15565 97019 15623 97025
rect 15565 97016 15577 97019
rect 14700 96988 15577 97016
rect 14700 96976 14706 96988
rect 15565 96985 15577 96988
rect 15611 96985 15623 97019
rect 15565 96979 15623 96985
rect 15657 97019 15715 97025
rect 15657 96985 15669 97019
rect 15703 97016 15715 97019
rect 17126 97016 17132 97028
rect 15703 96988 17132 97016
rect 15703 96985 15715 96988
rect 15657 96979 15715 96985
rect 17126 96976 17132 96988
rect 17184 97016 17190 97028
rect 22005 97019 22063 97025
rect 22005 97016 22017 97019
rect 17184 96988 22017 97016
rect 17184 96976 17190 96988
rect 22005 96985 22017 96988
rect 22051 96985 22063 97019
rect 22005 96979 22063 96985
rect 22646 96976 22652 97028
rect 22704 97016 22710 97028
rect 85298 97016 85304 97028
rect 22704 96988 85304 97016
rect 22704 96976 22710 96988
rect 85298 96976 85304 96988
rect 85356 96976 85362 97028
rect 2958 96948 2964 96960
rect 2919 96920 2964 96948
rect 2958 96908 2964 96920
rect 3016 96908 3022 96960
rect 4801 96951 4859 96957
rect 4801 96917 4813 96951
rect 4847 96948 4859 96951
rect 6454 96948 6460 96960
rect 4847 96920 6460 96948
rect 4847 96917 4859 96920
rect 4801 96911 4859 96917
rect 6454 96908 6460 96920
rect 6512 96908 6518 96960
rect 6549 96951 6607 96957
rect 6549 96917 6561 96951
rect 6595 96948 6607 96951
rect 33134 96948 33140 96960
rect 6595 96920 33140 96948
rect 6595 96917 6607 96920
rect 6549 96911 6607 96917
rect 33134 96908 33140 96920
rect 33192 96948 33198 96960
rect 83182 96948 83188 96960
rect 33192 96920 83188 96948
rect 33192 96908 33198 96920
rect 83182 96908 83188 96920
rect 83240 96908 83246 96960
rect 83458 96908 83464 96960
rect 83516 96948 83522 96960
rect 84286 96948 84292 96960
rect 83516 96920 84292 96948
rect 83516 96908 83522 96920
rect 84286 96908 84292 96920
rect 84344 96908 84350 96960
rect 84930 96908 84936 96960
rect 84988 96948 84994 96960
rect 85393 96951 85451 96957
rect 85393 96948 85405 96951
rect 84988 96920 85405 96948
rect 84988 96908 84994 96920
rect 85393 96917 85405 96920
rect 85439 96917 85451 96951
rect 85393 96911 85451 96917
rect 1104 96858 5152 96880
rect 1104 96806 1982 96858
rect 2034 96806 2046 96858
rect 2098 96806 2110 96858
rect 2162 96806 2174 96858
rect 2226 96806 5152 96858
rect 5626 96840 5632 96892
rect 5684 96880 5690 96892
rect 30098 96880 30104 96892
rect 5684 96852 30104 96880
rect 5684 96840 5690 96852
rect 30098 96840 30104 96852
rect 30156 96880 30162 96892
rect 82906 96880 82912 96892
rect 30156 96852 82912 96880
rect 30156 96840 30162 96852
rect 82906 96840 82912 96852
rect 82964 96840 82970 96892
rect 83642 96880 83648 96892
rect 83603 96852 83648 96880
rect 83642 96840 83648 96852
rect 83700 96840 83706 96892
rect 84180 96858 90896 96880
rect 1104 96784 5152 96806
rect 5261 96815 5319 96821
rect 5261 96781 5273 96815
rect 5307 96812 5319 96815
rect 6270 96812 6276 96824
rect 5307 96784 6276 96812
rect 5307 96781 5319 96784
rect 5261 96775 5319 96781
rect 6270 96772 6276 96784
rect 6328 96812 6334 96824
rect 32030 96812 32036 96824
rect 6328 96784 32036 96812
rect 6328 96772 6334 96784
rect 32030 96772 32036 96784
rect 32088 96812 32094 96824
rect 83090 96812 83096 96824
rect 32088 96784 83096 96812
rect 32088 96772 32094 96784
rect 83090 96772 83096 96784
rect 83148 96772 83154 96824
rect 83274 96772 83280 96824
rect 83332 96812 83338 96824
rect 84013 96815 84071 96821
rect 84013 96812 84025 96815
rect 83332 96784 84025 96812
rect 83332 96772 83338 96784
rect 84013 96781 84025 96784
rect 84059 96781 84071 96815
rect 84180 96806 85982 96858
rect 86034 96806 86046 96858
rect 86098 96806 86110 96858
rect 86162 96806 86174 96858
rect 86226 96806 89982 96858
rect 90034 96806 90046 96858
rect 90098 96806 90110 96858
rect 90162 96806 90174 96858
rect 90226 96806 90896 96858
rect 84180 96784 90896 96806
rect 84013 96775 84071 96781
rect 3326 96704 3332 96756
rect 3384 96744 3390 96756
rect 6733 96747 6791 96753
rect 6733 96744 6745 96747
rect 3384 96716 6745 96744
rect 3384 96704 3390 96716
rect 6733 96713 6745 96716
rect 6779 96713 6791 96747
rect 6733 96707 6791 96713
rect 6825 96747 6883 96753
rect 6825 96713 6837 96747
rect 6871 96744 6883 96747
rect 24302 96744 24308 96756
rect 6871 96716 24308 96744
rect 6871 96713 6883 96716
rect 6825 96707 6883 96713
rect 24302 96704 24308 96716
rect 24360 96744 24366 96756
rect 24360 96716 76880 96744
rect 24360 96704 24366 96716
rect 2958 96636 2964 96688
rect 3016 96676 3022 96688
rect 3418 96676 3424 96688
rect 3016 96648 3424 96676
rect 3016 96636 3022 96648
rect 3418 96636 3424 96648
rect 3476 96676 3482 96688
rect 22094 96676 22100 96688
rect 3476 96648 22100 96676
rect 3476 96636 3482 96648
rect 22094 96636 22100 96648
rect 22152 96676 22158 96688
rect 22922 96676 22928 96688
rect 22152 96648 22928 96676
rect 22152 96636 22158 96648
rect 22922 96636 22928 96648
rect 22980 96636 22986 96688
rect 23017 96679 23075 96685
rect 23017 96645 23029 96679
rect 23063 96676 23075 96679
rect 25406 96676 25412 96688
rect 23063 96648 25412 96676
rect 23063 96645 23075 96648
rect 23017 96639 23075 96645
rect 25406 96636 25412 96648
rect 25464 96676 25470 96688
rect 76745 96679 76803 96685
rect 76745 96676 76757 96679
rect 25464 96648 76757 96676
rect 25464 96636 25470 96648
rect 76745 96645 76757 96648
rect 76791 96645 76803 96679
rect 76852 96676 76880 96716
rect 76926 96704 76932 96756
rect 76984 96744 76990 96756
rect 80054 96744 80060 96756
rect 76984 96716 80060 96744
rect 76984 96704 76990 96716
rect 80054 96704 80060 96716
rect 80112 96704 80118 96756
rect 80149 96747 80207 96753
rect 80149 96713 80161 96747
rect 80195 96744 80207 96747
rect 82909 96747 82967 96753
rect 82909 96744 82921 96747
rect 80195 96716 82921 96744
rect 80195 96713 80207 96716
rect 80149 96707 80207 96713
rect 82909 96713 82921 96716
rect 82955 96713 82967 96747
rect 82909 96707 82967 96713
rect 85574 96676 85580 96688
rect 76852 96648 85580 96676
rect 76745 96639 76803 96645
rect 85574 96636 85580 96648
rect 85632 96636 85638 96688
rect 85942 96636 85948 96688
rect 86000 96676 86006 96688
rect 86402 96676 86408 96688
rect 86000 96648 86408 96676
rect 86000 96636 86006 96648
rect 86402 96636 86408 96648
rect 86460 96636 86466 96688
rect 5442 96568 5448 96620
rect 5500 96608 5506 96620
rect 87046 96608 87052 96620
rect 5500 96580 87052 96608
rect 5500 96568 5506 96580
rect 87046 96568 87052 96580
rect 87104 96568 87110 96620
rect 4065 96543 4123 96549
rect 4065 96509 4077 96543
rect 4111 96540 4123 96543
rect 4614 96540 4620 96552
rect 4111 96512 4620 96540
rect 4111 96509 4123 96512
rect 4065 96503 4123 96509
rect 4614 96500 4620 96512
rect 4672 96540 4678 96552
rect 39574 96540 39580 96552
rect 4672 96512 39580 96540
rect 4672 96500 4678 96512
rect 39574 96500 39580 96512
rect 39632 96500 39638 96552
rect 39669 96543 39727 96549
rect 39669 96509 39681 96543
rect 39715 96540 39727 96543
rect 62298 96540 62304 96552
rect 39715 96512 62304 96540
rect 39715 96509 39727 96512
rect 39669 96503 39727 96509
rect 62298 96500 62304 96512
rect 62356 96500 62362 96552
rect 85758 96540 85764 96552
rect 70366 96512 85764 96540
rect 4433 96475 4491 96481
rect 4433 96441 4445 96475
rect 4479 96472 4491 96475
rect 5353 96475 5411 96481
rect 5353 96472 5365 96475
rect 4479 96444 5365 96472
rect 4479 96441 4491 96444
rect 4433 96435 4491 96441
rect 5353 96441 5365 96444
rect 5399 96441 5411 96475
rect 5353 96435 5411 96441
rect 16482 96432 16488 96484
rect 16540 96472 16546 96484
rect 70366 96472 70394 96512
rect 85758 96500 85764 96512
rect 85816 96500 85822 96552
rect 16540 96444 70394 96472
rect 74629 96475 74687 96481
rect 16540 96432 16546 96444
rect 74629 96441 74641 96475
rect 74675 96472 74687 96475
rect 76650 96472 76656 96484
rect 74675 96444 76656 96472
rect 74675 96441 74687 96444
rect 74629 96435 74687 96441
rect 76650 96432 76656 96444
rect 76708 96432 76714 96484
rect 76745 96475 76803 96481
rect 76745 96441 76757 96475
rect 76791 96472 76803 96475
rect 80149 96475 80207 96481
rect 80149 96472 80161 96475
rect 76791 96444 80161 96472
rect 76791 96441 76803 96444
rect 76745 96435 76803 96441
rect 80149 96441 80161 96444
rect 80195 96441 80207 96475
rect 80149 96435 80207 96441
rect 80333 96475 80391 96481
rect 80333 96441 80345 96475
rect 80379 96472 80391 96475
rect 82081 96475 82139 96481
rect 82081 96472 82093 96475
rect 80379 96444 82093 96472
rect 80379 96441 80391 96444
rect 80333 96435 80391 96441
rect 82081 96441 82093 96444
rect 82127 96441 82139 96475
rect 82081 96435 82139 96441
rect 82170 96432 82176 96484
rect 82228 96472 82234 96484
rect 82814 96472 82820 96484
rect 82228 96444 82820 96472
rect 82228 96432 82234 96444
rect 82814 96432 82820 96444
rect 82872 96432 82878 96484
rect 88978 96472 88984 96484
rect 84488 96444 88984 96472
rect 3326 96404 3332 96416
rect 3287 96376 3332 96404
rect 3326 96364 3332 96376
rect 3384 96364 3390 96416
rect 3694 96404 3700 96416
rect 3655 96376 3700 96404
rect 3694 96364 3700 96376
rect 3752 96364 3758 96416
rect 4801 96407 4859 96413
rect 4801 96373 4813 96407
rect 4847 96404 4859 96407
rect 5902 96404 5908 96416
rect 4847 96376 5908 96404
rect 4847 96373 4859 96376
rect 4801 96367 4859 96373
rect 5902 96364 5908 96376
rect 5960 96404 5966 96416
rect 8481 96407 8539 96413
rect 8481 96404 8493 96407
rect 5960 96376 8493 96404
rect 5960 96364 5966 96376
rect 8481 96373 8493 96376
rect 8527 96373 8539 96407
rect 8481 96367 8539 96373
rect 29178 96364 29184 96416
rect 29236 96404 29242 96416
rect 84488 96404 84516 96444
rect 88978 96432 88984 96444
rect 89036 96432 89042 96484
rect 29236 96376 84516 96404
rect 84749 96407 84807 96413
rect 29236 96364 29242 96376
rect 84749 96373 84761 96407
rect 84795 96404 84807 96407
rect 84838 96404 84844 96416
rect 84795 96376 84844 96404
rect 84795 96373 84807 96376
rect 84749 96367 84807 96373
rect 84838 96364 84844 96376
rect 84896 96364 84902 96416
rect 85114 96404 85120 96416
rect 85027 96376 85120 96404
rect 85114 96364 85120 96376
rect 85172 96404 85178 96416
rect 85390 96404 85396 96416
rect 85172 96376 85396 96404
rect 85172 96364 85178 96376
rect 85390 96364 85396 96376
rect 85448 96364 85454 96416
rect 1104 96314 5152 96336
rect 1104 96262 3982 96314
rect 4034 96262 4046 96314
rect 4098 96262 4110 96314
rect 4162 96262 4174 96314
rect 4226 96262 5152 96314
rect 15746 96296 15752 96348
rect 15804 96336 15810 96348
rect 82722 96336 82728 96348
rect 15804 96308 82728 96336
rect 15804 96296 15810 96308
rect 82722 96296 82728 96308
rect 82780 96296 82786 96348
rect 84180 96314 90896 96336
rect 1104 96240 5152 96262
rect 37826 96228 37832 96280
rect 37884 96268 37890 96280
rect 39669 96271 39727 96277
rect 39669 96268 39681 96271
rect 37884 96240 39681 96268
rect 37884 96228 37890 96240
rect 39669 96237 39681 96240
rect 39715 96237 39727 96271
rect 39669 96231 39727 96237
rect 41138 96228 41144 96280
rect 41196 96268 41202 96280
rect 59354 96268 59360 96280
rect 41196 96240 59360 96268
rect 41196 96228 41202 96240
rect 59354 96228 59360 96240
rect 59412 96228 59418 96280
rect 60642 96268 60648 96280
rect 59464 96240 60648 96268
rect 3697 96203 3755 96209
rect 3697 96169 3709 96203
rect 3743 96200 3755 96203
rect 9582 96200 9588 96212
rect 3743 96172 9588 96200
rect 3743 96169 3755 96172
rect 3697 96163 3755 96169
rect 9582 96160 9588 96172
rect 9640 96160 9646 96212
rect 50338 96160 50344 96212
rect 50396 96200 50402 96212
rect 51166 96200 51172 96212
rect 50396 96172 51172 96200
rect 50396 96160 50402 96172
rect 51166 96160 51172 96172
rect 51224 96160 51230 96212
rect 57606 96160 57612 96212
rect 57664 96200 57670 96212
rect 59464 96200 59492 96240
rect 60642 96228 60648 96240
rect 60700 96228 60706 96280
rect 61562 96228 61568 96280
rect 61620 96268 61626 96280
rect 74997 96271 75055 96277
rect 74997 96268 75009 96271
rect 61620 96240 75009 96268
rect 61620 96228 61626 96240
rect 74997 96237 75009 96240
rect 75043 96237 75055 96271
rect 76561 96271 76619 96277
rect 76561 96268 76573 96271
rect 74997 96231 75055 96237
rect 75104 96240 76573 96268
rect 57664 96172 59492 96200
rect 57664 96160 57670 96172
rect 59538 96160 59544 96212
rect 59596 96200 59602 96212
rect 75104 96200 75132 96240
rect 76561 96237 76573 96240
rect 76607 96237 76619 96271
rect 76561 96231 76619 96237
rect 76653 96271 76711 96277
rect 76653 96237 76665 96271
rect 76699 96268 76711 96271
rect 82633 96271 82691 96277
rect 82633 96268 82645 96271
rect 76699 96240 82645 96268
rect 76699 96237 76711 96240
rect 76653 96231 76711 96237
rect 82633 96237 82645 96240
rect 82679 96237 82691 96271
rect 84180 96262 87982 96314
rect 88034 96262 88046 96314
rect 88098 96262 88110 96314
rect 88162 96262 88174 96314
rect 88226 96262 90896 96314
rect 84180 96240 90896 96262
rect 82633 96231 82691 96237
rect 59596 96172 75132 96200
rect 59596 96160 59602 96172
rect 75178 96160 75184 96212
rect 75236 96200 75242 96212
rect 84746 96200 84752 96212
rect 75236 96172 84752 96200
rect 75236 96160 75242 96172
rect 84746 96160 84752 96172
rect 84804 96160 84810 96212
rect 3326 96092 3332 96144
rect 3384 96132 3390 96144
rect 6086 96132 6092 96144
rect 3384 96104 6092 96132
rect 3384 96092 3390 96104
rect 6086 96092 6092 96104
rect 6144 96132 6150 96144
rect 27982 96132 27988 96144
rect 6144 96104 27988 96132
rect 6144 96092 6150 96104
rect 27982 96092 27988 96104
rect 28040 96132 28046 96144
rect 28902 96132 28908 96144
rect 28040 96104 28908 96132
rect 28040 96092 28046 96104
rect 28902 96092 28908 96104
rect 28960 96092 28966 96144
rect 59722 96092 59728 96144
rect 59780 96132 59786 96144
rect 74537 96135 74595 96141
rect 74537 96132 74549 96135
rect 59780 96104 74549 96132
rect 59780 96092 59786 96104
rect 74537 96101 74549 96104
rect 74583 96101 74595 96135
rect 74537 96095 74595 96101
rect 74626 96092 74632 96144
rect 74684 96132 74690 96144
rect 80146 96132 80152 96144
rect 74684 96104 80152 96132
rect 74684 96092 74690 96104
rect 80146 96092 80152 96104
rect 80204 96092 80210 96144
rect 80241 96135 80299 96141
rect 80241 96101 80253 96135
rect 80287 96132 80299 96135
rect 82265 96135 82323 96141
rect 82265 96132 82277 96135
rect 80287 96104 82277 96132
rect 80287 96101 80299 96104
rect 80241 96095 80299 96101
rect 82265 96101 82277 96104
rect 82311 96101 82323 96135
rect 82265 96095 82323 96101
rect 82354 96092 82360 96144
rect 82412 96132 82418 96144
rect 82817 96135 82875 96141
rect 82817 96132 82829 96135
rect 82412 96104 82829 96132
rect 82412 96092 82418 96104
rect 82817 96101 82829 96104
rect 82863 96101 82875 96135
rect 82817 96095 82875 96101
rect 57882 96024 57888 96076
rect 57940 96064 57946 96076
rect 79229 96067 79287 96073
rect 79229 96064 79241 96067
rect 57940 96036 79241 96064
rect 57940 96024 57946 96036
rect 79229 96033 79241 96036
rect 79275 96033 79287 96067
rect 79229 96027 79287 96033
rect 79321 96067 79379 96073
rect 79321 96033 79333 96067
rect 79367 96064 79379 96067
rect 85850 96064 85856 96076
rect 79367 96036 85856 96064
rect 79367 96033 79379 96036
rect 79321 96027 79379 96033
rect 85850 96024 85856 96036
rect 85908 96024 85914 96076
rect 4433 95999 4491 96005
rect 4433 95965 4445 95999
rect 4479 95996 4491 95999
rect 6914 95996 6920 96008
rect 4479 95968 6920 95996
rect 4479 95965 4491 95968
rect 4433 95959 4491 95965
rect 6914 95956 6920 95968
rect 6972 95996 6978 96008
rect 41966 95996 41972 96008
rect 6972 95968 41972 95996
rect 6972 95956 6978 95968
rect 41966 95956 41972 95968
rect 42024 95956 42030 96008
rect 54570 95956 54576 96008
rect 54628 95996 54634 96008
rect 76745 95999 76803 96005
rect 76745 95996 76757 95999
rect 54628 95968 76757 95996
rect 54628 95956 54634 95968
rect 76745 95965 76757 95968
rect 76791 95965 76803 95999
rect 76745 95959 76803 95965
rect 76834 95956 76840 96008
rect 76892 95996 76898 96008
rect 79686 95996 79692 96008
rect 76892 95968 79692 95996
rect 76892 95956 76898 95968
rect 79686 95956 79692 95968
rect 79744 95956 79750 96008
rect 79778 95956 79784 96008
rect 79836 95996 79842 96008
rect 80241 95999 80299 96005
rect 80241 95996 80253 95999
rect 79836 95968 80253 95996
rect 79836 95956 79842 95968
rect 80241 95965 80253 95968
rect 80287 95965 80299 95999
rect 80241 95959 80299 95965
rect 80330 95956 80336 96008
rect 80388 95996 80394 96008
rect 87230 95996 87236 96008
rect 80388 95968 87236 95996
rect 80388 95956 80394 95968
rect 87230 95956 87236 95968
rect 87288 95956 87294 96008
rect 4890 95888 4896 95940
rect 4948 95928 4954 95940
rect 5442 95928 5448 95940
rect 4948 95900 5448 95928
rect 4948 95888 4954 95900
rect 5442 95888 5448 95900
rect 5500 95928 5506 95940
rect 86954 95928 86960 95940
rect 5500 95900 86960 95928
rect 5500 95888 5506 95900
rect 86954 95888 86960 95900
rect 87012 95888 87018 95940
rect 4801 95863 4859 95869
rect 4801 95829 4813 95863
rect 4847 95860 4859 95863
rect 5261 95863 5319 95869
rect 5261 95860 5273 95863
rect 4847 95832 5273 95860
rect 4847 95829 4859 95832
rect 4801 95823 4859 95829
rect 5261 95829 5273 95832
rect 5307 95829 5319 95863
rect 5261 95823 5319 95829
rect 5353 95863 5411 95869
rect 5353 95829 5365 95863
rect 5399 95860 5411 95863
rect 5810 95860 5816 95872
rect 5399 95832 5816 95860
rect 5399 95829 5411 95832
rect 5353 95823 5411 95829
rect 5810 95820 5816 95832
rect 5868 95860 5874 95872
rect 8573 95863 8631 95869
rect 8573 95860 8585 95863
rect 5868 95832 8585 95860
rect 5868 95820 5874 95832
rect 8573 95829 8585 95832
rect 8619 95829 8631 95863
rect 8573 95823 8631 95829
rect 52178 95820 52184 95872
rect 52236 95860 52242 95872
rect 82722 95860 82728 95872
rect 52236 95832 82728 95860
rect 52236 95820 52242 95832
rect 82722 95820 82728 95832
rect 82780 95820 82786 95872
rect 84749 95863 84807 95869
rect 84749 95829 84761 95863
rect 84795 95860 84807 95863
rect 85022 95860 85028 95872
rect 84795 95832 85028 95860
rect 84795 95829 84807 95832
rect 84749 95823 84807 95829
rect 85022 95820 85028 95832
rect 85080 95860 85086 95872
rect 85482 95860 85488 95872
rect 85080 95832 85488 95860
rect 85080 95820 85086 95832
rect 85482 95820 85488 95832
rect 85540 95820 85546 95872
rect 15746 95792 15752 95804
rect 1104 95770 5152 95792
rect 1104 95718 1982 95770
rect 2034 95718 2046 95770
rect 2098 95718 2110 95770
rect 2162 95718 2174 95770
rect 2226 95718 5152 95770
rect 1104 95696 5152 95718
rect 8404 95764 15752 95792
rect 4433 95659 4491 95665
rect 4433 95625 4445 95659
rect 4479 95656 4491 95659
rect 8404 95656 8432 95764
rect 15746 95752 15752 95764
rect 15804 95752 15810 95804
rect 24578 95752 24584 95804
rect 24636 95792 24642 95804
rect 62022 95792 62028 95804
rect 24636 95764 62028 95792
rect 24636 95752 24642 95764
rect 62022 95752 62028 95764
rect 62080 95752 62086 95804
rect 62114 95752 62120 95804
rect 62172 95792 62178 95804
rect 79137 95795 79195 95801
rect 79137 95792 79149 95795
rect 62172 95764 79149 95792
rect 62172 95752 62178 95764
rect 79137 95761 79149 95764
rect 79183 95761 79195 95795
rect 79137 95755 79195 95761
rect 79229 95795 79287 95801
rect 79229 95761 79241 95795
rect 79275 95792 79287 95795
rect 79965 95795 80023 95801
rect 79965 95792 79977 95795
rect 79275 95764 79977 95792
rect 79275 95761 79287 95764
rect 79229 95755 79287 95761
rect 79965 95761 79977 95764
rect 80011 95761 80023 95795
rect 79965 95755 80023 95761
rect 80149 95795 80207 95801
rect 80149 95761 80161 95795
rect 80195 95792 80207 95795
rect 80195 95764 83136 95792
rect 80195 95761 80207 95764
rect 80149 95755 80207 95761
rect 8573 95727 8631 95733
rect 8573 95693 8585 95727
rect 8619 95724 8631 95727
rect 34974 95724 34980 95736
rect 8619 95696 34980 95724
rect 8619 95693 8631 95696
rect 8573 95687 8631 95693
rect 34974 95684 34980 95696
rect 35032 95724 35038 95736
rect 76653 95727 76711 95733
rect 76653 95724 76665 95727
rect 35032 95696 76665 95724
rect 35032 95684 35038 95696
rect 76653 95693 76665 95696
rect 76699 95693 76711 95727
rect 76653 95687 76711 95693
rect 76745 95727 76803 95733
rect 76745 95693 76757 95727
rect 76791 95724 76803 95727
rect 79873 95727 79931 95733
rect 79873 95724 79885 95727
rect 76791 95696 79885 95724
rect 76791 95693 76803 95696
rect 76745 95687 76803 95693
rect 79873 95693 79885 95696
rect 79919 95693 79931 95727
rect 79873 95687 79931 95693
rect 80057 95727 80115 95733
rect 80057 95693 80069 95727
rect 80103 95724 80115 95727
rect 82909 95727 82967 95733
rect 82909 95724 82921 95727
rect 80103 95696 82921 95724
rect 80103 95693 80115 95696
rect 80057 95687 80115 95693
rect 82909 95693 82921 95696
rect 82955 95693 82967 95727
rect 82909 95687 82967 95693
rect 4479 95628 8432 95656
rect 8481 95659 8539 95665
rect 4479 95625 4491 95628
rect 4433 95619 4491 95625
rect 8481 95625 8493 95659
rect 8527 95656 8539 95659
rect 31478 95656 31484 95668
rect 8527 95628 31484 95656
rect 8527 95625 8539 95628
rect 8481 95619 8539 95625
rect 31478 95616 31484 95628
rect 31536 95656 31542 95668
rect 82998 95656 83004 95668
rect 31536 95628 83004 95656
rect 31536 95616 31542 95628
rect 82998 95616 83004 95628
rect 83056 95616 83062 95668
rect 83108 95656 83136 95764
rect 84180 95770 90896 95792
rect 84180 95718 85982 95770
rect 86034 95718 86046 95770
rect 86098 95718 86110 95770
rect 86162 95718 86174 95770
rect 86226 95718 89982 95770
rect 90034 95718 90046 95770
rect 90098 95718 90110 95770
rect 90162 95718 90174 95770
rect 90226 95718 90896 95770
rect 84180 95696 90896 95718
rect 87506 95656 87512 95668
rect 83108 95628 87512 95656
rect 87506 95616 87512 95628
rect 87564 95616 87570 95668
rect 6822 95548 6828 95600
rect 6880 95588 6886 95600
rect 16482 95588 16488 95600
rect 6880 95560 16488 95588
rect 6880 95548 6886 95560
rect 16482 95548 16488 95560
rect 16540 95548 16546 95600
rect 27522 95548 27528 95600
rect 27580 95588 27586 95600
rect 79321 95591 79379 95597
rect 79321 95588 79333 95591
rect 27580 95560 79333 95588
rect 27580 95548 27586 95560
rect 79321 95557 79333 95560
rect 79367 95557 79379 95591
rect 79321 95551 79379 95557
rect 79413 95591 79471 95597
rect 79413 95557 79425 95591
rect 79459 95588 79471 95591
rect 83182 95588 83188 95600
rect 79459 95560 83188 95588
rect 79459 95557 79471 95560
rect 79413 95551 79471 95557
rect 83182 95548 83188 95560
rect 83240 95548 83246 95600
rect 5261 95523 5319 95529
rect 5261 95489 5273 95523
rect 5307 95520 5319 95523
rect 6546 95520 6552 95532
rect 5307 95492 6552 95520
rect 5307 95489 5319 95492
rect 5261 95483 5319 95489
rect 6546 95480 6552 95492
rect 6604 95520 6610 95532
rect 38470 95520 38476 95532
rect 6604 95492 38476 95520
rect 6604 95480 6610 95492
rect 38470 95480 38476 95492
rect 38528 95480 38534 95532
rect 58066 95480 58072 95532
rect 58124 95520 58130 95532
rect 83001 95523 83059 95529
rect 83001 95520 83013 95523
rect 58124 95492 83013 95520
rect 58124 95480 58130 95492
rect 83001 95489 83013 95492
rect 83047 95489 83059 95523
rect 83001 95483 83059 95489
rect 28902 95412 28908 95464
rect 28960 95452 28966 95464
rect 80057 95455 80115 95461
rect 80057 95452 80069 95455
rect 28960 95424 80069 95452
rect 28960 95412 28966 95424
rect 80057 95421 80069 95424
rect 80103 95421 80115 95455
rect 80057 95415 80115 95421
rect 80146 95412 80152 95464
rect 80204 95452 80210 95464
rect 83826 95452 83832 95464
rect 80204 95424 83832 95452
rect 80204 95412 80210 95424
rect 83826 95412 83832 95424
rect 83884 95412 83890 95464
rect 3694 95344 3700 95396
rect 3752 95384 3758 95396
rect 3878 95384 3884 95396
rect 3752 95356 3884 95384
rect 3752 95344 3758 95356
rect 3878 95344 3884 95356
rect 3936 95384 3942 95396
rect 20990 95384 20996 95396
rect 3936 95356 20996 95384
rect 3936 95344 3942 95356
rect 20990 95344 20996 95356
rect 21048 95384 21054 95396
rect 80333 95387 80391 95393
rect 21048 95356 80100 95384
rect 21048 95344 21054 95356
rect 4801 95319 4859 95325
rect 4801 95285 4813 95319
rect 4847 95316 4859 95319
rect 5350 95316 5356 95328
rect 4847 95288 5356 95316
rect 4847 95285 4859 95288
rect 4801 95279 4859 95285
rect 5350 95276 5356 95288
rect 5408 95316 5414 95328
rect 26786 95316 26792 95328
rect 5408 95288 26792 95316
rect 5408 95276 5414 95288
rect 26786 95276 26792 95288
rect 26844 95316 26850 95328
rect 27522 95316 27528 95328
rect 26844 95288 27528 95316
rect 26844 95276 26850 95288
rect 27522 95276 27528 95288
rect 27580 95276 27586 95328
rect 64138 95276 64144 95328
rect 64196 95316 64202 95328
rect 79965 95319 80023 95325
rect 79965 95316 79977 95319
rect 64196 95288 79977 95316
rect 64196 95276 64202 95288
rect 79965 95285 79977 95288
rect 80011 95285 80023 95319
rect 79965 95279 80023 95285
rect 1104 95226 5152 95248
rect 1104 95174 3982 95226
rect 4034 95174 4046 95226
rect 4098 95174 4110 95226
rect 4162 95174 4174 95226
rect 4226 95174 5152 95226
rect 45370 95208 45376 95260
rect 45428 95248 45434 95260
rect 49510 95248 49516 95260
rect 45428 95220 49516 95248
rect 45428 95208 45434 95220
rect 49510 95208 49516 95220
rect 49568 95208 49574 95260
rect 49602 95208 49608 95260
rect 49660 95248 49666 95260
rect 64782 95248 64788 95260
rect 49660 95220 64788 95248
rect 49660 95208 49666 95220
rect 64782 95208 64788 95220
rect 64840 95208 64846 95260
rect 74537 95251 74595 95257
rect 74537 95217 74549 95251
rect 74583 95248 74595 95251
rect 79137 95251 79195 95257
rect 74583 95220 78444 95248
rect 74583 95217 74595 95220
rect 74537 95211 74595 95217
rect 1104 95152 5152 95174
rect 24762 95140 24768 95192
rect 24820 95180 24826 95192
rect 78309 95183 78367 95189
rect 78309 95180 78321 95183
rect 24820 95152 78321 95180
rect 24820 95140 24826 95152
rect 78309 95149 78321 95152
rect 78355 95149 78367 95183
rect 78416 95180 78444 95220
rect 79137 95217 79149 95251
rect 79183 95248 79195 95251
rect 79870 95248 79876 95260
rect 79183 95220 79876 95248
rect 79183 95217 79195 95220
rect 79137 95211 79195 95217
rect 79870 95208 79876 95220
rect 79928 95208 79934 95260
rect 80072 95248 80100 95356
rect 80333 95353 80345 95387
rect 80379 95384 80391 95387
rect 82998 95384 83004 95396
rect 80379 95356 83004 95384
rect 80379 95353 80391 95356
rect 80333 95347 80391 95353
rect 82998 95344 83004 95356
rect 83056 95344 83062 95396
rect 80425 95319 80483 95325
rect 80425 95285 80437 95319
rect 80471 95316 80483 95319
rect 83274 95316 83280 95328
rect 80471 95288 83280 95316
rect 80471 95285 80483 95288
rect 80425 95279 80483 95285
rect 83274 95276 83280 95288
rect 83332 95276 83338 95328
rect 87414 95316 87420 95328
rect 83384 95288 87420 95316
rect 80333 95251 80391 95257
rect 80072 95220 80284 95248
rect 79413 95183 79471 95189
rect 79413 95180 79425 95183
rect 78416 95152 79425 95180
rect 78309 95143 78367 95149
rect 79413 95149 79425 95152
rect 79459 95149 79471 95183
rect 79413 95143 79471 95149
rect 79505 95183 79563 95189
rect 79505 95149 79517 95183
rect 79551 95180 79563 95183
rect 80146 95180 80152 95192
rect 79551 95152 80152 95180
rect 79551 95149 79563 95152
rect 79505 95143 79563 95149
rect 80146 95140 80152 95152
rect 80204 95140 80210 95192
rect 80256 95180 80284 95220
rect 80333 95217 80345 95251
rect 80379 95248 80391 95251
rect 83090 95248 83096 95260
rect 80379 95220 83096 95248
rect 80379 95217 80391 95220
rect 80333 95211 80391 95217
rect 83090 95208 83096 95220
rect 83148 95208 83154 95260
rect 83384 95248 83412 95288
rect 87414 95276 87420 95288
rect 87472 95276 87478 95328
rect 83200 95220 83412 95248
rect 84180 95226 90896 95248
rect 83200 95180 83228 95220
rect 80256 95152 83228 95180
rect 83366 95140 83372 95192
rect 83424 95180 83430 95192
rect 83550 95180 83556 95192
rect 83424 95152 83556 95180
rect 83424 95140 83430 95152
rect 83550 95140 83556 95152
rect 83608 95140 83614 95192
rect 84180 95174 87982 95226
rect 88034 95174 88046 95226
rect 88098 95174 88110 95226
rect 88162 95174 88174 95226
rect 88226 95174 90896 95226
rect 84180 95152 90896 95174
rect 19334 95072 19340 95124
rect 19392 95112 19398 95124
rect 85206 95112 85212 95124
rect 19392 95084 85212 95112
rect 19392 95072 19398 95084
rect 85206 95072 85212 95084
rect 85264 95072 85270 95124
rect 25958 95004 25964 95056
rect 26016 95044 26022 95056
rect 82538 95044 82544 95056
rect 26016 95016 82544 95044
rect 26016 95004 26022 95016
rect 82538 95004 82544 95016
rect 82596 95004 82602 95056
rect 4338 94936 4344 94988
rect 4396 94976 4402 94988
rect 29178 94976 29184 94988
rect 4396 94948 29184 94976
rect 4396 94936 4402 94948
rect 29178 94936 29184 94948
rect 29236 94936 29242 94988
rect 30282 94936 30288 94988
rect 30340 94976 30346 94988
rect 76469 94979 76527 94985
rect 76469 94976 76481 94979
rect 30340 94948 76481 94976
rect 30340 94936 30346 94948
rect 76469 94945 76481 94948
rect 76515 94945 76527 94979
rect 76469 94939 76527 94945
rect 76561 94979 76619 94985
rect 76561 94945 76573 94979
rect 76607 94976 76619 94979
rect 80057 94979 80115 94985
rect 80057 94976 80069 94979
rect 76607 94948 80069 94976
rect 76607 94945 76619 94948
rect 76561 94939 76619 94945
rect 80057 94945 80069 94948
rect 80103 94945 80115 94979
rect 80057 94939 80115 94945
rect 80146 94936 80152 94988
rect 80204 94976 80210 94988
rect 80204 94948 80376 94976
rect 80204 94936 80210 94948
rect 31662 94868 31668 94920
rect 31720 94908 31726 94920
rect 74534 94908 74540 94920
rect 31720 94880 74540 94908
rect 31720 94868 31726 94880
rect 74534 94868 74540 94880
rect 74592 94868 74598 94920
rect 74629 94911 74687 94917
rect 74629 94877 74641 94911
rect 74675 94908 74687 94911
rect 80238 94908 80244 94920
rect 74675 94880 80244 94908
rect 74675 94877 74687 94880
rect 74629 94871 74687 94877
rect 80238 94868 80244 94880
rect 80296 94868 80302 94920
rect 80348 94908 80376 94948
rect 80422 94936 80428 94988
rect 80480 94976 80486 94988
rect 82449 94979 82507 94985
rect 82449 94976 82461 94979
rect 80480 94948 82461 94976
rect 80480 94936 80486 94948
rect 82449 94945 82461 94948
rect 82495 94945 82507 94979
rect 82449 94939 82507 94945
rect 85850 94936 85856 94988
rect 85908 94976 85914 94988
rect 86862 94976 86868 94988
rect 85908 94948 86868 94976
rect 85908 94936 85914 94948
rect 86862 94936 86868 94948
rect 86920 94936 86926 94988
rect 82814 94908 82820 94920
rect 80348 94880 82820 94908
rect 82814 94868 82820 94880
rect 82872 94908 82878 94920
rect 83642 94908 83648 94920
rect 82872 94880 83648 94908
rect 82872 94868 82878 94880
rect 83642 94868 83648 94880
rect 83700 94868 83706 94920
rect 20622 94800 20628 94852
rect 20680 94840 20686 94852
rect 44174 94840 44180 94852
rect 20680 94812 44180 94840
rect 20680 94800 20686 94812
rect 44174 94800 44180 94812
rect 44232 94800 44238 94852
rect 45186 94800 45192 94852
rect 45244 94840 45250 94852
rect 78214 94840 78220 94852
rect 45244 94812 78220 94840
rect 45244 94800 45250 94812
rect 78214 94800 78220 94812
rect 78272 94800 78278 94852
rect 78309 94843 78367 94849
rect 78309 94809 78321 94843
rect 78355 94840 78367 94843
rect 82725 94843 82783 94849
rect 82725 94840 82737 94843
rect 78355 94812 82737 94840
rect 78355 94809 78367 94812
rect 78309 94803 78367 94809
rect 82725 94809 82737 94812
rect 82771 94809 82783 94843
rect 82725 94803 82783 94809
rect 86310 94800 86316 94852
rect 86368 94840 86374 94852
rect 86862 94840 86868 94852
rect 86368 94812 86868 94840
rect 86368 94800 86374 94812
rect 86862 94800 86868 94812
rect 86920 94800 86926 94852
rect 4430 94732 4436 94784
rect 4488 94772 4494 94784
rect 19334 94772 19340 94784
rect 4488 94744 19340 94772
rect 4488 94732 4494 94744
rect 19334 94732 19340 94744
rect 19392 94732 19398 94784
rect 45554 94732 45560 94784
rect 45612 94772 45618 94784
rect 74537 94775 74595 94781
rect 74537 94772 74549 94775
rect 45612 94744 74549 94772
rect 45612 94732 45618 94744
rect 74537 94741 74549 94744
rect 74583 94741 74595 94775
rect 74537 94735 74595 94741
rect 74813 94775 74871 94781
rect 74813 94741 74825 94775
rect 74859 94772 74871 94775
rect 76098 94772 76104 94784
rect 74859 94744 76104 94772
rect 74859 94741 74871 94744
rect 74813 94735 74871 94741
rect 76098 94732 76104 94744
rect 76156 94732 76162 94784
rect 76193 94775 76251 94781
rect 76193 94741 76205 94775
rect 76239 94772 76251 94775
rect 80057 94775 80115 94781
rect 80057 94772 80069 94775
rect 76239 94744 80069 94772
rect 76239 94741 76251 94744
rect 76193 94735 76251 94741
rect 80057 94741 80069 94744
rect 80103 94741 80115 94775
rect 80057 94735 80115 94741
rect 80606 94732 80612 94784
rect 80664 94772 80670 94784
rect 82354 94772 82360 94784
rect 80664 94744 82360 94772
rect 80664 94732 80670 94744
rect 82354 94732 82360 94744
rect 82412 94732 82418 94784
rect 82449 94775 82507 94781
rect 82449 94741 82461 94775
rect 82495 94772 82507 94775
rect 85758 94772 85764 94784
rect 82495 94744 85764 94772
rect 82495 94741 82507 94744
rect 82449 94735 82507 94741
rect 85758 94732 85764 94744
rect 85816 94732 85822 94784
rect 1104 94682 5152 94704
rect 1104 94630 1982 94682
rect 2034 94630 2046 94682
rect 2098 94630 2110 94682
rect 2162 94630 2174 94682
rect 2226 94630 5152 94682
rect 38562 94664 38568 94716
rect 38620 94704 38626 94716
rect 46842 94704 46848 94716
rect 38620 94676 46848 94704
rect 38620 94664 38626 94676
rect 46842 94664 46848 94676
rect 46900 94664 46906 94716
rect 47946 94664 47952 94716
rect 48004 94704 48010 94716
rect 74997 94707 75055 94713
rect 48004 94676 74948 94704
rect 48004 94664 48010 94676
rect 1104 94608 5152 94630
rect 6454 94596 6460 94648
rect 6512 94636 6518 94648
rect 12802 94636 12808 94648
rect 6512 94608 12808 94636
rect 6512 94596 6518 94608
rect 12802 94596 12808 94608
rect 12860 94636 12866 94648
rect 13722 94636 13728 94648
rect 12860 94608 13728 94636
rect 12860 94596 12866 94608
rect 13722 94596 13728 94608
rect 13780 94596 13786 94648
rect 23382 94596 23388 94648
rect 23440 94636 23446 94648
rect 48222 94636 48228 94648
rect 23440 94608 48228 94636
rect 23440 94596 23446 94608
rect 48222 94596 48228 94608
rect 48280 94596 48286 94648
rect 49878 94596 49884 94648
rect 49936 94636 49942 94648
rect 50798 94636 50804 94648
rect 49936 94608 50804 94636
rect 49936 94596 49942 94608
rect 50798 94596 50804 94608
rect 50856 94596 50862 94648
rect 52546 94596 52552 94648
rect 52604 94636 52610 94648
rect 74813 94639 74871 94645
rect 74813 94636 74825 94639
rect 52604 94608 74825 94636
rect 52604 94596 52610 94608
rect 74813 94605 74825 94608
rect 74859 94605 74871 94639
rect 74920 94636 74948 94676
rect 74997 94673 75009 94707
rect 75043 94704 75055 94707
rect 80149 94707 80207 94713
rect 80149 94704 80161 94707
rect 75043 94676 80161 94704
rect 75043 94673 75055 94676
rect 74997 94667 75055 94673
rect 80149 94673 80161 94676
rect 80195 94673 80207 94707
rect 80149 94667 80207 94673
rect 80238 94664 80244 94716
rect 80296 94704 80302 94716
rect 80425 94707 80483 94713
rect 80425 94704 80437 94707
rect 80296 94676 80437 94704
rect 80296 94664 80302 94676
rect 80425 94673 80437 94676
rect 80471 94673 80483 94707
rect 80425 94667 80483 94673
rect 80514 94664 80520 94716
rect 80572 94704 80578 94716
rect 83550 94704 83556 94716
rect 80572 94676 83556 94704
rect 80572 94664 80578 94676
rect 83550 94664 83556 94676
rect 83608 94664 83614 94716
rect 84180 94682 90896 94704
rect 76377 94639 76435 94645
rect 76377 94636 76389 94639
rect 74920 94608 76389 94636
rect 74813 94599 74871 94605
rect 76377 94605 76389 94608
rect 76423 94605 76435 94639
rect 76377 94599 76435 94605
rect 76469 94639 76527 94645
rect 76469 94605 76481 94639
rect 76515 94636 76527 94639
rect 83918 94636 83924 94648
rect 76515 94608 83924 94636
rect 76515 94605 76527 94608
rect 76469 94599 76527 94605
rect 83918 94596 83924 94608
rect 83976 94596 83982 94648
rect 84180 94630 85982 94682
rect 86034 94630 86046 94682
rect 86098 94630 86110 94682
rect 86162 94630 86174 94682
rect 86226 94630 89982 94682
rect 90034 94630 90046 94682
rect 90098 94630 90110 94682
rect 90162 94630 90174 94682
rect 90226 94630 90896 94682
rect 84180 94608 90896 94630
rect 4522 94528 4528 94580
rect 4580 94568 4586 94580
rect 37274 94568 37280 94580
rect 4580 94540 37280 94568
rect 4580 94528 4586 94540
rect 37274 94528 37280 94540
rect 37332 94528 37338 94580
rect 46658 94528 46664 94580
rect 46716 94568 46722 94580
rect 74534 94568 74540 94580
rect 46716 94540 74540 94568
rect 46716 94528 46722 94540
rect 74534 94528 74540 94540
rect 74592 94528 74598 94580
rect 74626 94528 74632 94580
rect 74684 94568 74690 94580
rect 80422 94568 80428 94580
rect 74684 94540 80428 94568
rect 74684 94528 74690 94540
rect 80422 94528 80428 94540
rect 80480 94528 80486 94580
rect 80517 94571 80575 94577
rect 80517 94537 80529 94571
rect 80563 94568 80575 94571
rect 82449 94571 82507 94577
rect 82449 94568 82461 94571
rect 80563 94540 82461 94568
rect 80563 94537 80575 94540
rect 80517 94531 80575 94537
rect 82449 94537 82461 94540
rect 82495 94537 82507 94571
rect 82449 94531 82507 94537
rect 82541 94571 82599 94577
rect 82541 94537 82553 94571
rect 82587 94568 82599 94571
rect 85482 94568 85488 94580
rect 82587 94540 85488 94568
rect 82587 94537 82599 94540
rect 82541 94531 82599 94537
rect 85482 94528 85488 94540
rect 85540 94528 85546 94580
rect 4890 94460 4896 94512
rect 4948 94500 4954 94512
rect 86954 94500 86960 94512
rect 4948 94472 86960 94500
rect 4948 94460 4954 94472
rect 86954 94460 86960 94472
rect 87012 94460 87018 94512
rect 49970 94392 49976 94444
rect 50028 94432 50034 94444
rect 50028 94404 74764 94432
rect 50028 94392 50034 94404
rect 51442 94324 51448 94376
rect 51500 94364 51506 94376
rect 74736 94364 74764 94404
rect 74810 94392 74816 94444
rect 74868 94432 74874 94444
rect 79229 94435 79287 94441
rect 79229 94432 79241 94435
rect 74868 94404 79241 94432
rect 74868 94392 74874 94404
rect 79229 94401 79241 94404
rect 79275 94401 79287 94435
rect 79229 94395 79287 94401
rect 79321 94435 79379 94441
rect 79321 94401 79333 94435
rect 79367 94432 79379 94435
rect 85390 94432 85396 94444
rect 79367 94404 85396 94432
rect 79367 94401 79379 94404
rect 79321 94395 79379 94401
rect 85390 94392 85396 94404
rect 85448 94392 85454 94444
rect 85298 94364 85304 94376
rect 51500 94336 74672 94364
rect 74736 94336 85304 94364
rect 51500 94324 51506 94336
rect 45094 94256 45100 94308
rect 45152 94296 45158 94308
rect 53742 94296 53748 94308
rect 45152 94268 53748 94296
rect 45152 94256 45158 94268
rect 53742 94256 53748 94268
rect 53800 94256 53806 94308
rect 54018 94256 54024 94308
rect 54076 94296 54082 94308
rect 74537 94299 74595 94305
rect 74537 94296 74549 94299
rect 54076 94268 74549 94296
rect 54076 94256 54082 94268
rect 74537 94265 74549 94268
rect 74583 94265 74595 94299
rect 74644 94296 74672 94336
rect 85298 94324 85304 94336
rect 85356 94324 85362 94376
rect 79321 94299 79379 94305
rect 79321 94296 79333 94299
rect 74644 94268 79333 94296
rect 74537 94259 74595 94265
rect 79321 94265 79333 94268
rect 79367 94265 79379 94299
rect 79321 94259 79379 94265
rect 79413 94299 79471 94305
rect 79413 94265 79425 94299
rect 79459 94296 79471 94299
rect 83366 94296 83372 94308
rect 79459 94268 83372 94296
rect 79459 94265 79471 94268
rect 79413 94259 79471 94265
rect 83366 94256 83372 94268
rect 83424 94256 83430 94308
rect 83458 94256 83464 94308
rect 83516 94296 83522 94308
rect 84838 94296 84844 94308
rect 83516 94268 84844 94296
rect 83516 94256 83522 94268
rect 84838 94256 84844 94268
rect 84896 94256 84902 94308
rect 4430 94188 4436 94240
rect 4488 94228 4494 94240
rect 5258 94228 5264 94240
rect 4488 94200 5264 94228
rect 4488 94188 4494 94200
rect 5258 94188 5264 94200
rect 5316 94188 5322 94240
rect 44082 94188 44088 94240
rect 44140 94228 44146 94240
rect 54846 94228 54852 94240
rect 44140 94200 54852 94228
rect 44140 94188 44146 94200
rect 54846 94188 54852 94200
rect 54904 94188 54910 94240
rect 54938 94188 54944 94240
rect 54996 94228 55002 94240
rect 76193 94231 76251 94237
rect 76193 94228 76205 94231
rect 54996 94200 76205 94228
rect 54996 94188 55002 94200
rect 76193 94197 76205 94200
rect 76239 94197 76251 94231
rect 87506 94228 87512 94240
rect 76193 94191 76251 94197
rect 76300 94200 87512 94228
rect 1104 94138 5152 94160
rect 1104 94086 3982 94138
rect 4034 94086 4046 94138
rect 4098 94086 4110 94138
rect 4162 94086 4174 94138
rect 4226 94086 5152 94138
rect 42702 94120 42708 94172
rect 42760 94160 42766 94172
rect 42760 94132 45554 94160
rect 42760 94120 42766 94132
rect 1104 94064 5152 94086
rect 45526 94092 45554 94132
rect 48130 94120 48136 94172
rect 48188 94160 48194 94172
rect 50982 94160 50988 94172
rect 48188 94132 50988 94160
rect 48188 94120 48194 94132
rect 50982 94120 50988 94132
rect 51040 94120 51046 94172
rect 53282 94120 53288 94172
rect 53340 94160 53346 94172
rect 59906 94160 59912 94172
rect 53340 94132 59912 94160
rect 53340 94120 53346 94132
rect 59906 94120 59912 94132
rect 59964 94120 59970 94172
rect 62022 94120 62028 94172
rect 62080 94160 62086 94172
rect 76300 94160 76328 94200
rect 87506 94188 87512 94200
rect 87564 94188 87570 94240
rect 62080 94132 76328 94160
rect 76377 94163 76435 94169
rect 62080 94120 62086 94132
rect 76377 94129 76389 94163
rect 76423 94160 76435 94163
rect 79137 94163 79195 94169
rect 79137 94160 79149 94163
rect 76423 94132 79149 94160
rect 76423 94129 76435 94132
rect 76377 94123 76435 94129
rect 79137 94129 79149 94132
rect 79183 94129 79195 94163
rect 79137 94123 79195 94129
rect 79226 94120 79232 94172
rect 79284 94160 79290 94172
rect 81434 94160 81440 94172
rect 79284 94132 81440 94160
rect 79284 94120 79290 94132
rect 81434 94120 81440 94132
rect 81492 94120 81498 94172
rect 83458 94160 83464 94172
rect 82188 94132 83464 94160
rect 61930 94092 61936 94104
rect 45526 94064 61936 94092
rect 61930 94052 61936 94064
rect 61988 94052 61994 94104
rect 62298 94052 62304 94104
rect 62356 94092 62362 94104
rect 76193 94095 76251 94101
rect 76193 94092 76205 94095
rect 62356 94064 76205 94092
rect 62356 94052 62362 94064
rect 76193 94061 76205 94064
rect 76239 94061 76251 94095
rect 82188 94092 82216 94132
rect 83458 94120 83464 94132
rect 83516 94120 83522 94172
rect 84180 94138 90896 94160
rect 76193 94055 76251 94061
rect 76300 94064 82216 94092
rect 84180 94086 87982 94138
rect 88034 94086 88046 94138
rect 88098 94086 88110 94138
rect 88162 94086 88174 94138
rect 88226 94086 90896 94138
rect 84180 94064 90896 94086
rect 49050 93984 49056 94036
rect 49108 94024 49114 94036
rect 76300 94024 76328 94064
rect 49108 93996 76328 94024
rect 76377 94027 76435 94033
rect 49108 93984 49114 93996
rect 76377 93993 76389 94027
rect 76423 94024 76435 94027
rect 87782 94024 87788 94036
rect 76423 93996 87788 94024
rect 76423 93993 76435 93996
rect 76377 93987 76435 93993
rect 87782 93984 87788 93996
rect 87840 93984 87846 94036
rect 13722 93916 13728 93968
rect 13780 93956 13786 93968
rect 84930 93956 84936 93968
rect 13780 93928 84936 93956
rect 13780 93916 13786 93928
rect 84930 93916 84936 93928
rect 84988 93916 84994 93968
rect 86586 93916 86592 93968
rect 86644 93956 86650 93968
rect 87598 93956 87604 93968
rect 86644 93928 87604 93956
rect 86644 93916 86650 93928
rect 87598 93916 87604 93928
rect 87656 93916 87662 93968
rect 4522 93848 4528 93900
rect 4580 93888 4586 93900
rect 5261 93891 5319 93897
rect 5261 93888 5273 93891
rect 4580 93860 5273 93888
rect 4580 93848 4586 93860
rect 5261 93857 5273 93860
rect 5307 93857 5319 93891
rect 5261 93851 5319 93857
rect 9582 93848 9588 93900
rect 9640 93888 9646 93900
rect 85298 93888 85304 93900
rect 9640 93860 85304 93888
rect 9640 93848 9646 93860
rect 85298 93848 85304 93860
rect 85356 93848 85362 93900
rect 50614 93780 50620 93832
rect 50672 93820 50678 93832
rect 87690 93820 87696 93832
rect 50672 93792 87696 93820
rect 50672 93780 50678 93792
rect 87690 93780 87696 93792
rect 87748 93780 87754 93832
rect 49510 93712 49516 93764
rect 49568 93752 49574 93764
rect 86954 93752 86960 93764
rect 49568 93724 86960 93752
rect 49568 93712 49574 93724
rect 86954 93712 86960 93724
rect 87012 93712 87018 93764
rect 4522 93644 4528 93696
rect 4580 93684 4586 93696
rect 79321 93687 79379 93693
rect 79321 93684 79333 93687
rect 4580 93656 79333 93684
rect 4580 93644 4586 93656
rect 79321 93653 79333 93656
rect 79367 93653 79379 93687
rect 79321 93647 79379 93653
rect 79410 93644 79416 93696
rect 79468 93684 79474 93696
rect 82906 93684 82912 93696
rect 79468 93656 82912 93684
rect 79468 93644 79474 93656
rect 82906 93644 82912 93656
rect 82964 93644 82970 93696
rect 87230 93684 87236 93696
rect 83292 93656 87236 93684
rect 1104 93594 5152 93616
rect 1104 93542 1982 93594
rect 2034 93542 2046 93594
rect 2098 93542 2110 93594
rect 2162 93542 2174 93594
rect 2226 93542 5152 93594
rect 48774 93576 48780 93628
rect 48832 93616 48838 93628
rect 54202 93616 54208 93628
rect 48832 93588 54208 93616
rect 48832 93576 48838 93588
rect 54202 93576 54208 93588
rect 54260 93576 54266 93628
rect 64782 93576 64788 93628
rect 64840 93616 64846 93628
rect 83292 93616 83320 93656
rect 87230 93644 87236 93656
rect 87288 93644 87294 93696
rect 83458 93616 83464 93628
rect 64840 93588 83320 93616
rect 83419 93588 83464 93616
rect 64840 93576 64846 93588
rect 83458 93576 83464 93588
rect 83516 93576 83522 93628
rect 84180 93594 90896 93616
rect 1104 93520 5152 93542
rect 59354 93508 59360 93560
rect 59412 93548 59418 93560
rect 78585 93551 78643 93557
rect 59412 93520 78536 93548
rect 59412 93508 59418 93520
rect 51258 93440 51264 93492
rect 51316 93480 51322 93492
rect 78401 93483 78459 93489
rect 78401 93480 78413 93483
rect 51316 93452 78413 93480
rect 51316 93440 51322 93452
rect 78401 93449 78413 93452
rect 78447 93449 78459 93483
rect 78508 93480 78536 93520
rect 78585 93517 78597 93551
rect 78631 93548 78643 93551
rect 84010 93548 84016 93560
rect 78631 93520 84016 93548
rect 78631 93517 78643 93520
rect 78585 93511 78643 93517
rect 84010 93508 84016 93520
rect 84068 93508 84074 93560
rect 84180 93542 85982 93594
rect 86034 93542 86046 93594
rect 86098 93542 86110 93594
rect 86162 93542 86174 93594
rect 86226 93542 89982 93594
rect 90034 93542 90046 93594
rect 90098 93542 90110 93594
rect 90162 93542 90174 93594
rect 90226 93542 90896 93594
rect 84180 93520 90896 93542
rect 87322 93480 87328 93492
rect 78508 93452 87328 93480
rect 78401 93443 78459 93449
rect 87322 93440 87328 93452
rect 87380 93440 87386 93492
rect 53742 93372 53748 93424
rect 53800 93412 53806 93424
rect 77294 93412 77300 93424
rect 53800 93384 77300 93412
rect 53800 93372 53806 93384
rect 77294 93372 77300 93384
rect 77352 93372 77358 93424
rect 77389 93415 77447 93421
rect 77389 93381 77401 93415
rect 77435 93412 77447 93415
rect 78217 93415 78275 93421
rect 78217 93412 78229 93415
rect 77435 93384 78229 93412
rect 77435 93381 77447 93384
rect 77389 93375 77447 93381
rect 78217 93381 78229 93384
rect 78263 93381 78275 93415
rect 79229 93415 79287 93421
rect 79229 93412 79241 93415
rect 78217 93375 78275 93381
rect 78324 93384 79241 93412
rect 47946 93304 47952 93356
rect 48004 93344 48010 93356
rect 78324 93344 78352 93384
rect 79229 93381 79241 93384
rect 79275 93381 79287 93415
rect 79229 93375 79287 93381
rect 79321 93415 79379 93421
rect 79321 93381 79333 93415
rect 79367 93412 79379 93415
rect 84562 93412 84568 93424
rect 79367 93384 84568 93412
rect 79367 93381 79379 93384
rect 79321 93375 79379 93381
rect 84562 93372 84568 93384
rect 84620 93372 84626 93424
rect 84746 93412 84752 93424
rect 84707 93384 84752 93412
rect 84746 93372 84752 93384
rect 84804 93372 84810 93424
rect 85114 93412 85120 93424
rect 85075 93384 85120 93412
rect 85114 93372 85120 93384
rect 85172 93372 85178 93424
rect 48004 93316 78352 93344
rect 78401 93347 78459 93353
rect 48004 93304 48010 93316
rect 78401 93313 78413 93347
rect 78447 93344 78459 93347
rect 82446 93344 82452 93356
rect 78447 93316 82452 93344
rect 78447 93313 78459 93316
rect 78401 93307 78459 93313
rect 82446 93304 82452 93316
rect 82504 93304 82510 93356
rect 82814 93344 82820 93356
rect 82775 93316 82820 93344
rect 82814 93304 82820 93316
rect 82872 93304 82878 93356
rect 46658 93236 46664 93288
rect 46716 93276 46722 93288
rect 77389 93279 77447 93285
rect 77389 93276 77401 93279
rect 46716 93248 77401 93276
rect 46716 93236 46722 93248
rect 77389 93245 77401 93248
rect 77435 93245 77447 93279
rect 77389 93239 77447 93245
rect 77478 93236 77484 93288
rect 77536 93276 77542 93288
rect 79502 93276 79508 93288
rect 77536 93248 79508 93276
rect 77536 93236 77542 93248
rect 79502 93236 79508 93248
rect 79560 93236 79566 93288
rect 79597 93279 79655 93285
rect 79597 93245 79609 93279
rect 79643 93276 79655 93279
rect 84102 93276 84108 93288
rect 79643 93248 84108 93276
rect 79643 93245 79655 93248
rect 79597 93239 79655 93245
rect 84102 93236 84108 93248
rect 84160 93236 84166 93288
rect 44082 93168 44088 93220
rect 44140 93208 44146 93220
rect 78217 93211 78275 93217
rect 78217 93208 78229 93211
rect 44140 93180 78229 93208
rect 44140 93168 44146 93180
rect 78217 93177 78229 93180
rect 78263 93177 78275 93211
rect 78217 93171 78275 93177
rect 78309 93211 78367 93217
rect 78309 93177 78321 93211
rect 78355 93208 78367 93211
rect 83734 93208 83740 93220
rect 78355 93180 83740 93208
rect 78355 93177 78367 93180
rect 78309 93171 78367 93177
rect 83734 93168 83740 93180
rect 83792 93168 83798 93220
rect 42610 93100 42616 93152
rect 42668 93140 42674 93152
rect 84194 93140 84200 93152
rect 42668 93112 84200 93140
rect 42668 93100 42674 93112
rect 84194 93100 84200 93112
rect 84252 93100 84258 93152
rect 1104 93050 5152 93072
rect 1104 92998 3982 93050
rect 4034 92998 4046 93050
rect 4098 92998 4110 93050
rect 4162 92998 4174 93050
rect 4226 92998 5152 93050
rect 39942 93032 39948 93084
rect 40000 93072 40006 93084
rect 78309 93075 78367 93081
rect 78309 93072 78321 93075
rect 40000 93044 78321 93072
rect 40000 93032 40006 93044
rect 78309 93041 78321 93044
rect 78355 93041 78367 93075
rect 78309 93035 78367 93041
rect 78401 93075 78459 93081
rect 78401 93041 78413 93075
rect 78447 93072 78459 93075
rect 82357 93075 82415 93081
rect 82357 93072 82369 93075
rect 78447 93044 82369 93072
rect 78447 93041 78459 93044
rect 78401 93035 78459 93041
rect 82357 93041 82369 93044
rect 82403 93041 82415 93075
rect 82357 93035 82415 93041
rect 84180 93050 90896 93072
rect 1104 92976 5152 92998
rect 38378 92964 38384 93016
rect 38436 93004 38442 93016
rect 78585 93007 78643 93013
rect 38436 92976 78536 93004
rect 38436 92964 38442 92976
rect 35250 92896 35256 92948
rect 35308 92936 35314 92948
rect 78401 92939 78459 92945
rect 78401 92936 78413 92939
rect 35308 92908 78413 92936
rect 35308 92896 35314 92908
rect 78401 92905 78413 92908
rect 78447 92905 78459 92939
rect 78508 92936 78536 92976
rect 78585 92973 78597 93007
rect 78631 93004 78643 93007
rect 83918 93004 83924 93016
rect 78631 92976 83924 93004
rect 78631 92973 78643 92976
rect 78585 92967 78643 92973
rect 83918 92964 83924 92976
rect 83976 92964 83982 93016
rect 84180 92998 87982 93050
rect 88034 92998 88046 93050
rect 88098 92998 88110 93050
rect 88162 92998 88174 93050
rect 88226 92998 90896 93050
rect 84180 92976 90896 92998
rect 84286 92936 84292 92948
rect 78508 92908 84292 92936
rect 78401 92899 78459 92905
rect 84286 92896 84292 92908
rect 84344 92896 84350 92948
rect 36722 92828 36728 92880
rect 36780 92868 36786 92880
rect 82265 92871 82323 92877
rect 82265 92868 82277 92871
rect 36780 92840 82277 92868
rect 36780 92828 36786 92840
rect 82265 92837 82277 92840
rect 82311 92837 82323 92871
rect 82265 92831 82323 92837
rect 82357 92871 82415 92877
rect 82357 92837 82369 92871
rect 82403 92868 82415 92871
rect 84746 92868 84752 92880
rect 82403 92840 84752 92868
rect 82403 92837 82415 92840
rect 82357 92831 82415 92837
rect 84746 92828 84752 92840
rect 84804 92828 84810 92880
rect 32858 92760 32864 92812
rect 32916 92760 32922 92812
rect 34146 92760 34152 92812
rect 34204 92800 34210 92812
rect 34204 92772 85252 92800
rect 34204 92760 34210 92772
rect 32876 92732 32904 92760
rect 85224 92744 85252 92772
rect 84838 92732 84844 92744
rect 32876 92704 84844 92732
rect 84838 92692 84844 92704
rect 84896 92692 84902 92744
rect 85206 92692 85212 92744
rect 85264 92692 85270 92744
rect 82449 92667 82507 92673
rect 82449 92633 82461 92667
rect 82495 92664 82507 92667
rect 87414 92664 87420 92676
rect 82495 92636 87420 92664
rect 82495 92633 82507 92636
rect 82449 92627 82507 92633
rect 87414 92624 87420 92636
rect 87472 92624 87478 92676
rect 1104 92506 5152 92528
rect 1104 92454 1982 92506
rect 2034 92454 2046 92506
rect 2098 92454 2110 92506
rect 2162 92454 2174 92506
rect 2226 92454 5152 92506
rect 1104 92432 5152 92454
rect 84180 92506 90896 92528
rect 84180 92454 85982 92506
rect 86034 92454 86046 92506
rect 86098 92454 86110 92506
rect 86162 92454 86174 92506
rect 86226 92454 89982 92506
rect 90034 92454 90046 92506
rect 90098 92454 90110 92506
rect 90162 92454 90174 92506
rect 90226 92454 90896 92506
rect 84180 92432 90896 92454
rect 83001 92395 83059 92401
rect 83001 92361 83013 92395
rect 83047 92392 83059 92395
rect 87046 92392 87052 92404
rect 83047 92364 87052 92392
rect 83047 92361 83059 92364
rect 83001 92355 83059 92361
rect 87046 92352 87052 92364
rect 87104 92352 87110 92404
rect 82909 92327 82967 92333
rect 82909 92293 82921 92327
rect 82955 92324 82967 92327
rect 87138 92324 87144 92336
rect 82955 92296 87144 92324
rect 82955 92293 82967 92296
rect 82909 92287 82967 92293
rect 87138 92284 87144 92296
rect 87196 92284 87202 92336
rect 82814 92216 82820 92268
rect 82872 92256 82878 92268
rect 87506 92256 87512 92268
rect 82872 92228 87512 92256
rect 82872 92216 82878 92228
rect 87506 92216 87512 92228
rect 87564 92216 87570 92268
rect 82814 92120 82820 92132
rect 82775 92092 82820 92120
rect 82814 92080 82820 92092
rect 82872 92080 82878 92132
rect 84749 92055 84807 92061
rect 84749 92021 84761 92055
rect 84795 92052 84807 92055
rect 85574 92052 85580 92064
rect 84795 92024 85580 92052
rect 84795 92021 84807 92024
rect 84749 92015 84807 92021
rect 85574 92012 85580 92024
rect 85632 92052 85638 92064
rect 86770 92052 86776 92064
rect 85632 92024 86776 92052
rect 85632 92012 85638 92024
rect 86770 92012 86776 92024
rect 86828 92012 86834 92064
rect 1104 91962 5152 91984
rect 1104 91910 3982 91962
rect 4034 91910 4046 91962
rect 4098 91910 4110 91962
rect 4162 91910 4174 91962
rect 4226 91910 5152 91962
rect 1104 91888 5152 91910
rect 84180 91962 90896 91984
rect 84180 91910 87982 91962
rect 88034 91910 88046 91962
rect 88098 91910 88110 91962
rect 88162 91910 88174 91962
rect 88226 91910 90896 91962
rect 84180 91888 90896 91910
rect 82633 91783 82691 91789
rect 82633 91749 82645 91783
rect 82679 91780 82691 91783
rect 88334 91780 88340 91792
rect 82679 91752 88340 91780
rect 82679 91749 82691 91752
rect 82633 91743 82691 91749
rect 88334 91740 88340 91752
rect 88392 91740 88398 91792
rect 1104 91418 5152 91440
rect 1104 91366 1982 91418
rect 2034 91366 2046 91418
rect 2098 91366 2110 91418
rect 2162 91366 2174 91418
rect 2226 91366 5152 91418
rect 1104 91344 5152 91366
rect 84180 91418 90896 91440
rect 84180 91366 85982 91418
rect 86034 91366 86046 91418
rect 86098 91366 86110 91418
rect 86162 91366 86174 91418
rect 86226 91366 89982 91418
rect 90034 91366 90046 91418
rect 90098 91366 90110 91418
rect 90162 91366 90174 91418
rect 90226 91366 90896 91418
rect 84180 91344 90896 91366
rect 1104 90874 5152 90896
rect 1104 90822 3982 90874
rect 4034 90822 4046 90874
rect 4098 90822 4110 90874
rect 4162 90822 4174 90874
rect 4226 90822 5152 90874
rect 1104 90800 5152 90822
rect 84180 90874 90896 90896
rect 84180 90822 87982 90874
rect 88034 90822 88046 90874
rect 88098 90822 88110 90874
rect 88162 90822 88174 90874
rect 88226 90822 90896 90874
rect 84180 90800 90896 90822
rect 86402 90720 86408 90772
rect 86460 90760 86466 90772
rect 86678 90760 86684 90772
rect 86460 90732 86684 90760
rect 86460 90720 86466 90732
rect 86678 90720 86684 90732
rect 86736 90720 86742 90772
rect 4890 90652 4896 90704
rect 4948 90692 4954 90704
rect 5442 90692 5448 90704
rect 4948 90664 5448 90692
rect 4948 90652 4954 90664
rect 5442 90652 5448 90664
rect 5500 90652 5506 90704
rect 4338 90516 4344 90568
rect 4396 90556 4402 90568
rect 5442 90556 5448 90568
rect 4396 90528 5448 90556
rect 4396 90516 4402 90528
rect 5442 90516 5448 90528
rect 5500 90516 5506 90568
rect 4338 90380 4344 90432
rect 4396 90420 4402 90432
rect 5261 90423 5319 90429
rect 5261 90420 5273 90423
rect 4396 90392 5273 90420
rect 4396 90380 4402 90392
rect 5261 90389 5273 90392
rect 5307 90389 5319 90423
rect 5261 90383 5319 90389
rect 1104 90330 5152 90352
rect 1104 90278 1982 90330
rect 2034 90278 2046 90330
rect 2098 90278 2110 90330
rect 2162 90278 2174 90330
rect 2226 90278 5152 90330
rect 1104 90256 5152 90278
rect 84180 90330 90896 90352
rect 84180 90278 85982 90330
rect 86034 90278 86046 90330
rect 86098 90278 86110 90330
rect 86162 90278 86174 90330
rect 86226 90278 89982 90330
rect 90034 90278 90046 90330
rect 90098 90278 90110 90330
rect 90162 90278 90174 90330
rect 90226 90278 90896 90330
rect 84180 90256 90896 90278
rect 86678 90040 86684 90092
rect 86736 90080 86742 90092
rect 86954 90080 86960 90092
rect 86736 90052 86960 90080
rect 86736 90040 86742 90052
rect 86954 90040 86960 90052
rect 87012 90040 87018 90092
rect 1104 89786 5152 89808
rect 1104 89734 3982 89786
rect 4034 89734 4046 89786
rect 4098 89734 4110 89786
rect 4162 89734 4174 89786
rect 4226 89734 5152 89786
rect 1104 89712 5152 89734
rect 84180 89786 90896 89808
rect 84180 89734 87982 89786
rect 88034 89734 88046 89786
rect 88098 89734 88110 89786
rect 88162 89734 88174 89786
rect 88226 89734 90896 89786
rect 84180 89712 90896 89734
rect 86862 89672 86868 89684
rect 86696 89644 86868 89672
rect 86696 89480 86724 89644
rect 86862 89632 86868 89644
rect 86920 89632 86926 89684
rect 87506 89632 87512 89684
rect 87564 89672 87570 89684
rect 88334 89672 88340 89684
rect 87564 89644 88340 89672
rect 87564 89632 87570 89644
rect 88334 89632 88340 89644
rect 88392 89632 88398 89684
rect 86678 89428 86684 89480
rect 86736 89428 86742 89480
rect 5074 89360 5080 89412
rect 5132 89400 5138 89412
rect 5132 89372 5212 89400
rect 5132 89360 5138 89372
rect 1104 89242 5152 89264
rect 1104 89190 1982 89242
rect 2034 89190 2046 89242
rect 2098 89190 2110 89242
rect 2162 89190 2174 89242
rect 2226 89190 5152 89242
rect 1104 89168 5152 89190
rect 4798 89060 4804 89072
rect 4759 89032 4804 89060
rect 4798 89020 4804 89032
rect 4856 89060 4862 89072
rect 5184 89060 5212 89372
rect 84180 89242 90896 89264
rect 84180 89190 85982 89242
rect 86034 89190 86046 89242
rect 86098 89190 86110 89242
rect 86162 89190 86174 89242
rect 86226 89190 89982 89242
rect 90034 89190 90046 89242
rect 90098 89190 90110 89242
rect 90162 89190 90174 89242
rect 90226 89190 90896 89242
rect 84180 89168 90896 89190
rect 4856 89032 5212 89060
rect 4856 89020 4862 89032
rect 4338 88952 4344 89004
rect 4396 88992 4402 89004
rect 4890 88992 4896 89004
rect 4396 88964 4896 88992
rect 4396 88952 4402 88964
rect 4890 88952 4896 88964
rect 4948 88952 4954 89004
rect 4338 88816 4344 88868
rect 4396 88856 4402 88868
rect 5258 88856 5264 88868
rect 4396 88828 5264 88856
rect 4396 88816 4402 88828
rect 5258 88816 5264 88828
rect 5316 88816 5322 88868
rect 1104 88698 5152 88720
rect 1104 88646 3982 88698
rect 4034 88646 4046 88698
rect 4098 88646 4110 88698
rect 4162 88646 4174 88698
rect 4226 88646 5152 88698
rect 1104 88624 5152 88646
rect 84180 88698 90896 88720
rect 84180 88646 87982 88698
rect 88034 88646 88046 88698
rect 88098 88646 88110 88698
rect 88162 88646 88174 88698
rect 88226 88646 90896 88698
rect 84180 88624 90896 88646
rect 84930 88272 84936 88324
rect 84988 88312 84994 88324
rect 87966 88312 87972 88324
rect 84988 88284 87972 88312
rect 84988 88272 84994 88284
rect 87966 88272 87972 88284
rect 88024 88272 88030 88324
rect 1104 88154 5152 88176
rect 1104 88102 1982 88154
rect 2034 88102 2046 88154
rect 2098 88102 2110 88154
rect 2162 88102 2174 88154
rect 2226 88102 5152 88154
rect 1104 88080 5152 88102
rect 84180 88154 90896 88176
rect 84180 88102 85982 88154
rect 86034 88102 86046 88154
rect 86098 88102 86110 88154
rect 86162 88102 86174 88154
rect 86226 88102 89982 88154
rect 90034 88102 90046 88154
rect 90098 88102 90110 88154
rect 90162 88102 90174 88154
rect 90226 88102 90896 88154
rect 84180 88080 90896 88102
rect 4801 88043 4859 88049
rect 4801 88009 4813 88043
rect 4847 88040 4859 88043
rect 4982 88040 4988 88052
rect 4847 88012 4988 88040
rect 4847 88009 4859 88012
rect 4801 88003 4859 88009
rect 4982 88000 4988 88012
rect 5040 88000 5046 88052
rect 1104 87610 5152 87632
rect 1104 87558 3982 87610
rect 4034 87558 4046 87610
rect 4098 87558 4110 87610
rect 4162 87558 4174 87610
rect 4226 87558 5152 87610
rect 1104 87536 5152 87558
rect 84180 87610 90896 87632
rect 84180 87558 87982 87610
rect 88034 87558 88046 87610
rect 88098 87558 88110 87610
rect 88162 87558 88174 87610
rect 88226 87558 90896 87610
rect 84180 87536 90896 87558
rect 1104 87066 5152 87088
rect 1104 87014 1982 87066
rect 2034 87014 2046 87066
rect 2098 87014 2110 87066
rect 2162 87014 2174 87066
rect 2226 87014 5152 87066
rect 1104 86992 5152 87014
rect 84180 87066 90896 87088
rect 84180 87014 85982 87066
rect 86034 87014 86046 87066
rect 86098 87014 86110 87066
rect 86162 87014 86174 87066
rect 86226 87014 89982 87066
rect 90034 87014 90046 87066
rect 90098 87014 90110 87066
rect 90162 87014 90174 87066
rect 90226 87014 90896 87066
rect 84180 86992 90896 87014
rect 1104 86522 5152 86544
rect 1104 86470 3982 86522
rect 4034 86470 4046 86522
rect 4098 86470 4110 86522
rect 4162 86470 4174 86522
rect 4226 86470 5152 86522
rect 1104 86448 5152 86470
rect 84180 86522 90896 86544
rect 84180 86470 87982 86522
rect 88034 86470 88046 86522
rect 88098 86470 88110 86522
rect 88162 86470 88174 86522
rect 88226 86470 90896 86522
rect 84180 86448 90896 86470
rect 4801 86411 4859 86417
rect 4801 86377 4813 86411
rect 4847 86408 4859 86411
rect 5166 86408 5172 86420
rect 4847 86380 5172 86408
rect 4847 86377 4859 86380
rect 4801 86371 4859 86377
rect 5166 86368 5172 86380
rect 5224 86368 5230 86420
rect 82998 86300 83004 86352
rect 83056 86340 83062 86352
rect 87966 86340 87972 86352
rect 83056 86312 87972 86340
rect 83056 86300 83062 86312
rect 87966 86300 87972 86312
rect 88024 86300 88030 86352
rect 1104 85978 5152 86000
rect 1104 85926 1982 85978
rect 2034 85926 2046 85978
rect 2098 85926 2110 85978
rect 2162 85926 2174 85978
rect 2226 85926 5152 85978
rect 1104 85904 5152 85926
rect 84180 85978 90896 86000
rect 84180 85926 85982 85978
rect 86034 85926 86046 85978
rect 86098 85926 86110 85978
rect 86162 85926 86174 85978
rect 86226 85926 89982 85978
rect 90034 85926 90046 85978
rect 90098 85926 90110 85978
rect 90162 85926 90174 85978
rect 90226 85926 90896 85978
rect 84180 85904 90896 85926
rect 1104 85434 5152 85456
rect 1104 85382 3982 85434
rect 4034 85382 4046 85434
rect 4098 85382 4110 85434
rect 4162 85382 4174 85434
rect 4226 85382 5152 85434
rect 1104 85360 5152 85382
rect 84180 85434 90896 85456
rect 84180 85382 87982 85434
rect 88034 85382 88046 85434
rect 88098 85382 88110 85434
rect 88162 85382 88174 85434
rect 88226 85382 90896 85434
rect 84180 85360 90896 85382
rect 4706 85320 4712 85332
rect 4667 85292 4712 85320
rect 4706 85280 4712 85292
rect 4764 85280 4770 85332
rect 83826 85212 83832 85264
rect 83884 85252 83890 85264
rect 87966 85252 87972 85264
rect 83884 85224 87972 85252
rect 83884 85212 83890 85224
rect 87966 85212 87972 85224
rect 88024 85212 88030 85264
rect 84838 85076 84844 85128
rect 84896 85116 84902 85128
rect 85574 85116 85580 85128
rect 84896 85088 85580 85116
rect 84896 85076 84902 85088
rect 85574 85076 85580 85088
rect 85632 85076 85638 85128
rect 84562 84940 84568 84992
rect 84620 84980 84626 84992
rect 84838 84980 84844 84992
rect 84620 84952 84844 84980
rect 84620 84940 84626 84952
rect 84838 84940 84844 84952
rect 84896 84940 84902 84992
rect 1104 84890 5152 84912
rect 1104 84838 1982 84890
rect 2034 84838 2046 84890
rect 2098 84838 2110 84890
rect 2162 84838 2174 84890
rect 2226 84838 5152 84890
rect 1104 84816 5152 84838
rect 84180 84890 90896 84912
rect 84180 84838 85982 84890
rect 86034 84838 86046 84890
rect 86098 84838 86110 84890
rect 86162 84838 86174 84890
rect 86226 84838 89982 84890
rect 90034 84838 90046 84890
rect 90098 84838 90110 84890
rect 90162 84838 90174 84890
rect 90226 84838 90896 84890
rect 84180 84816 90896 84838
rect 85022 84736 85028 84788
rect 85080 84776 85086 84788
rect 85206 84776 85212 84788
rect 85080 84748 85212 84776
rect 85080 84736 85086 84748
rect 85206 84736 85212 84748
rect 85264 84736 85270 84788
rect 86954 84736 86960 84788
rect 87012 84776 87018 84788
rect 87230 84776 87236 84788
rect 87012 84748 87236 84776
rect 87012 84736 87018 84748
rect 87230 84736 87236 84748
rect 87288 84736 87294 84788
rect 82906 84532 82912 84584
rect 82964 84572 82970 84584
rect 84102 84572 84108 84584
rect 82964 84544 84108 84572
rect 82964 84532 82970 84544
rect 84102 84532 84108 84544
rect 84160 84532 84166 84584
rect 1104 84346 5152 84368
rect 1104 84294 3982 84346
rect 4034 84294 4046 84346
rect 4098 84294 4110 84346
rect 4162 84294 4174 84346
rect 4226 84294 5152 84346
rect 1104 84272 5152 84294
rect 84180 84346 90896 84368
rect 84180 84294 87982 84346
rect 88034 84294 88046 84346
rect 88098 84294 88110 84346
rect 88162 84294 88174 84346
rect 88226 84294 90896 84346
rect 84180 84272 90896 84294
rect 83090 84124 83096 84176
rect 83148 84164 83154 84176
rect 87966 84164 87972 84176
rect 83148 84136 87972 84164
rect 83148 84124 83154 84136
rect 87966 84124 87972 84136
rect 88024 84124 88030 84176
rect 1104 83802 5152 83824
rect 1104 83750 1982 83802
rect 2034 83750 2046 83802
rect 2098 83750 2110 83802
rect 2162 83750 2174 83802
rect 2226 83750 5152 83802
rect 1104 83728 5152 83750
rect 84180 83802 90896 83824
rect 84180 83750 85982 83802
rect 86034 83750 86046 83802
rect 86098 83750 86110 83802
rect 86162 83750 86174 83802
rect 86226 83750 89982 83802
rect 90034 83750 90046 83802
rect 90098 83750 90110 83802
rect 90162 83750 90174 83802
rect 90226 83750 90896 83802
rect 84180 83728 90896 83750
rect 4798 83348 4804 83360
rect 4759 83320 4804 83348
rect 4798 83308 4804 83320
rect 4856 83308 4862 83360
rect 1104 83258 5152 83280
rect 1104 83206 3982 83258
rect 4034 83206 4046 83258
rect 4098 83206 4110 83258
rect 4162 83206 4174 83258
rect 4226 83206 5152 83258
rect 1104 83184 5152 83206
rect 84180 83258 90896 83280
rect 84180 83206 87982 83258
rect 88034 83206 88046 83258
rect 88098 83206 88110 83258
rect 88162 83206 88174 83258
rect 88226 83206 90896 83258
rect 84180 83184 90896 83206
rect 1104 82714 5152 82736
rect 1104 82662 1982 82714
rect 2034 82662 2046 82714
rect 2098 82662 2110 82714
rect 2162 82662 2174 82714
rect 2226 82662 5152 82714
rect 1104 82640 5152 82662
rect 84180 82714 90896 82736
rect 84180 82662 85982 82714
rect 86034 82662 86046 82714
rect 86098 82662 86110 82714
rect 86162 82662 86174 82714
rect 86226 82662 89982 82714
rect 90034 82662 90046 82714
rect 90098 82662 90110 82714
rect 90162 82662 90174 82714
rect 90226 82662 90896 82714
rect 84180 82640 90896 82662
rect 4798 82260 4804 82272
rect 4759 82232 4804 82260
rect 4798 82220 4804 82232
rect 4856 82220 4862 82272
rect 1104 82170 5152 82192
rect 1104 82118 3982 82170
rect 4034 82118 4046 82170
rect 4098 82118 4110 82170
rect 4162 82118 4174 82170
rect 4226 82118 5152 82170
rect 1104 82096 5152 82118
rect 84180 82170 90896 82192
rect 84180 82118 87982 82170
rect 88034 82118 88046 82170
rect 88098 82118 88110 82170
rect 88162 82118 88174 82170
rect 88226 82118 90896 82170
rect 84180 82096 90896 82118
rect 83182 81948 83188 82000
rect 83240 81988 83246 82000
rect 87966 81988 87972 82000
rect 83240 81960 87972 81988
rect 83240 81948 83246 81960
rect 87966 81948 87972 81960
rect 88024 81948 88030 82000
rect 1104 81626 5152 81648
rect 1104 81574 1982 81626
rect 2034 81574 2046 81626
rect 2098 81574 2110 81626
rect 2162 81574 2174 81626
rect 2226 81574 5152 81626
rect 1104 81552 5152 81574
rect 84180 81626 90896 81648
rect 84180 81574 85982 81626
rect 86034 81574 86046 81626
rect 86098 81574 86110 81626
rect 86162 81574 86174 81626
rect 86226 81574 89982 81626
rect 90034 81574 90046 81626
rect 90098 81574 90110 81626
rect 90162 81574 90174 81626
rect 90226 81574 90896 81626
rect 84180 81552 90896 81574
rect 1104 81082 5152 81104
rect 1104 81030 3982 81082
rect 4034 81030 4046 81082
rect 4098 81030 4110 81082
rect 4162 81030 4174 81082
rect 4226 81030 5152 81082
rect 1104 81008 5152 81030
rect 84180 81082 90896 81104
rect 84180 81030 87982 81082
rect 88034 81030 88046 81082
rect 88098 81030 88110 81082
rect 88162 81030 88174 81082
rect 88226 81030 90896 81082
rect 84180 81008 90896 81030
rect 83274 80860 83280 80912
rect 83332 80900 83338 80912
rect 87966 80900 87972 80912
rect 83332 80872 87972 80900
rect 83332 80860 83338 80872
rect 87966 80860 87972 80872
rect 88024 80860 88030 80912
rect 1104 80538 5152 80560
rect 1104 80486 1982 80538
rect 2034 80486 2046 80538
rect 2098 80486 2110 80538
rect 2162 80486 2174 80538
rect 2226 80486 5152 80538
rect 1104 80464 5152 80486
rect 84180 80538 90896 80560
rect 84180 80486 85982 80538
rect 86034 80486 86046 80538
rect 86098 80486 86110 80538
rect 86162 80486 86174 80538
rect 86226 80486 89982 80538
rect 90034 80486 90046 80538
rect 90098 80486 90110 80538
rect 90162 80486 90174 80538
rect 90226 80486 90896 80538
rect 84180 80464 90896 80486
rect 4798 80424 4804 80436
rect 4759 80396 4804 80424
rect 4798 80384 4804 80396
rect 4856 80384 4862 80436
rect 86770 80112 86776 80164
rect 86828 80152 86834 80164
rect 87322 80152 87328 80164
rect 86828 80124 87328 80152
rect 86828 80112 86834 80124
rect 87322 80112 87328 80124
rect 87380 80112 87386 80164
rect 87506 80112 87512 80164
rect 87564 80152 87570 80164
rect 88334 80152 88340 80164
rect 87564 80124 88340 80152
rect 87564 80112 87570 80124
rect 88334 80112 88340 80124
rect 88392 80112 88398 80164
rect 1104 79994 5152 80016
rect 1104 79942 3982 79994
rect 4034 79942 4046 79994
rect 4098 79942 4110 79994
rect 4162 79942 4174 79994
rect 4226 79942 5152 79994
rect 1104 79920 5152 79942
rect 84180 79994 90896 80016
rect 84180 79942 87982 79994
rect 88034 79942 88046 79994
rect 88098 79942 88110 79994
rect 88162 79942 88174 79994
rect 88226 79942 90896 79994
rect 84180 79920 90896 79942
rect 1104 79450 5152 79472
rect 1104 79398 1982 79450
rect 2034 79398 2046 79450
rect 2098 79398 2110 79450
rect 2162 79398 2174 79450
rect 2226 79398 5152 79450
rect 1104 79376 5152 79398
rect 84180 79450 90896 79472
rect 84180 79398 85982 79450
rect 86034 79398 86046 79450
rect 86098 79398 86110 79450
rect 86162 79398 86174 79450
rect 86226 79398 89982 79450
rect 90034 79398 90046 79450
rect 90098 79398 90110 79450
rect 90162 79398 90174 79450
rect 90226 79398 90896 79450
rect 84180 79376 90896 79398
rect 1104 78906 5152 78928
rect 1104 78854 3982 78906
rect 4034 78854 4046 78906
rect 4098 78854 4110 78906
rect 4162 78854 4174 78906
rect 4226 78854 5152 78906
rect 1104 78832 5152 78854
rect 84180 78906 90896 78928
rect 84180 78854 87982 78906
rect 88034 78854 88046 78906
rect 88098 78854 88110 78906
rect 88162 78854 88174 78906
rect 88226 78854 90896 78906
rect 84180 78832 90896 78854
rect 1104 78362 5152 78384
rect 1104 78310 1982 78362
rect 2034 78310 2046 78362
rect 2098 78310 2110 78362
rect 2162 78310 2174 78362
rect 2226 78310 5152 78362
rect 1104 78288 5152 78310
rect 84180 78362 90896 78384
rect 84180 78310 85982 78362
rect 86034 78310 86046 78362
rect 86098 78310 86110 78362
rect 86162 78310 86174 78362
rect 86226 78310 89982 78362
rect 90034 78310 90046 78362
rect 90098 78310 90110 78362
rect 90162 78310 90174 78362
rect 90226 78310 90896 78362
rect 84180 78288 90896 78310
rect 1104 77818 5152 77840
rect 1104 77766 3982 77818
rect 4034 77766 4046 77818
rect 4098 77766 4110 77818
rect 4162 77766 4174 77818
rect 4226 77766 5152 77818
rect 1104 77744 5152 77766
rect 84180 77818 90896 77840
rect 84180 77766 87982 77818
rect 88034 77766 88046 77818
rect 88098 77766 88110 77818
rect 88162 77766 88174 77818
rect 88226 77766 90896 77818
rect 84180 77744 90896 77766
rect 1104 77274 5152 77296
rect 1104 77222 1982 77274
rect 2034 77222 2046 77274
rect 2098 77222 2110 77274
rect 2162 77222 2174 77274
rect 2226 77222 5152 77274
rect 1104 77200 5152 77222
rect 84180 77274 90896 77296
rect 84180 77222 85982 77274
rect 86034 77222 86046 77274
rect 86098 77222 86110 77274
rect 86162 77222 86174 77274
rect 86226 77222 89982 77274
rect 90034 77222 90046 77274
rect 90098 77222 90110 77274
rect 90162 77222 90174 77274
rect 90226 77222 90896 77274
rect 84180 77200 90896 77222
rect 84102 77120 84108 77172
rect 84160 77160 84166 77172
rect 87046 77160 87052 77172
rect 84160 77132 87052 77160
rect 84160 77120 84166 77132
rect 87046 77120 87052 77132
rect 87104 77120 87110 77172
rect 1104 76730 5152 76752
rect 1104 76678 3982 76730
rect 4034 76678 4046 76730
rect 4098 76678 4110 76730
rect 4162 76678 4174 76730
rect 4226 76678 5152 76730
rect 1104 76656 5152 76678
rect 84180 76730 90896 76752
rect 84180 76678 87982 76730
rect 88034 76678 88046 76730
rect 88098 76678 88110 76730
rect 88162 76678 88174 76730
rect 88226 76678 90896 76730
rect 84180 76656 90896 76678
rect 1104 76186 5152 76208
rect 1104 76134 1982 76186
rect 2034 76134 2046 76186
rect 2098 76134 2110 76186
rect 2162 76134 2174 76186
rect 2226 76134 5152 76186
rect 1104 76112 5152 76134
rect 84180 76186 90896 76208
rect 84180 76134 85982 76186
rect 86034 76134 86046 76186
rect 86098 76134 86110 76186
rect 86162 76134 86174 76186
rect 86226 76134 89982 76186
rect 90034 76134 90046 76186
rect 90098 76134 90110 76186
rect 90162 76134 90174 76186
rect 90226 76134 90896 76186
rect 84180 76112 90896 76134
rect 1104 75642 5152 75664
rect 1104 75590 3982 75642
rect 4034 75590 4046 75642
rect 4098 75590 4110 75642
rect 4162 75590 4174 75642
rect 4226 75590 5152 75642
rect 1104 75568 5152 75590
rect 84180 75642 90896 75664
rect 84180 75590 87982 75642
rect 88034 75590 88046 75642
rect 88098 75590 88110 75642
rect 88162 75590 88174 75642
rect 88226 75590 90896 75642
rect 84180 75568 90896 75590
rect 87138 75488 87144 75540
rect 87196 75528 87202 75540
rect 87414 75528 87420 75540
rect 87196 75500 87420 75528
rect 87196 75488 87202 75500
rect 87414 75488 87420 75500
rect 87472 75488 87478 75540
rect 87414 75216 87420 75268
rect 87472 75256 87478 75268
rect 87782 75256 87788 75268
rect 87472 75228 87788 75256
rect 87472 75216 87478 75228
rect 87782 75216 87788 75228
rect 87840 75216 87846 75268
rect 1104 75098 5152 75120
rect 1104 75046 1982 75098
rect 2034 75046 2046 75098
rect 2098 75046 2110 75098
rect 2162 75046 2174 75098
rect 2226 75046 5152 75098
rect 1104 75024 5152 75046
rect 84180 75098 90896 75120
rect 84180 75046 85982 75098
rect 86034 75046 86046 75098
rect 86098 75046 86110 75098
rect 86162 75046 86174 75098
rect 86226 75046 89982 75098
rect 90034 75046 90046 75098
rect 90098 75046 90110 75098
rect 90162 75046 90174 75098
rect 90226 75046 90896 75098
rect 84180 75024 90896 75046
rect 1104 74554 5152 74576
rect 1104 74502 3982 74554
rect 4034 74502 4046 74554
rect 4098 74502 4110 74554
rect 4162 74502 4174 74554
rect 4226 74502 5152 74554
rect 1104 74480 5152 74502
rect 84180 74554 90896 74576
rect 84180 74502 87982 74554
rect 88034 74502 88046 74554
rect 88098 74502 88110 74554
rect 88162 74502 88174 74554
rect 88226 74502 90896 74554
rect 84180 74480 90896 74502
rect 82446 74400 82452 74452
rect 82504 74440 82510 74452
rect 86954 74440 86960 74452
rect 82504 74412 86960 74440
rect 82504 74400 82510 74412
rect 86954 74400 86960 74412
rect 87012 74400 87018 74452
rect 1104 74010 5152 74032
rect 1104 73958 1982 74010
rect 2034 73958 2046 74010
rect 2098 73958 2110 74010
rect 2162 73958 2174 74010
rect 2226 73958 5152 74010
rect 1104 73936 5152 73958
rect 84180 74010 90896 74032
rect 84180 73958 85982 74010
rect 86034 73958 86046 74010
rect 86098 73958 86110 74010
rect 86162 73958 86174 74010
rect 86226 73958 89982 74010
rect 90034 73958 90046 74010
rect 90098 73958 90110 74010
rect 90162 73958 90174 74010
rect 90226 73958 90896 74010
rect 84180 73936 90896 73958
rect 1104 73466 5152 73488
rect 1104 73414 3982 73466
rect 4034 73414 4046 73466
rect 4098 73414 4110 73466
rect 4162 73414 4174 73466
rect 4226 73414 5152 73466
rect 1104 73392 5152 73414
rect 84180 73466 90896 73488
rect 84180 73414 87982 73466
rect 88034 73414 88046 73466
rect 88098 73414 88110 73466
rect 88162 73414 88174 73466
rect 88226 73414 90896 73466
rect 84180 73392 90896 73414
rect 1104 72922 5152 72944
rect 1104 72870 1982 72922
rect 2034 72870 2046 72922
rect 2098 72870 2110 72922
rect 2162 72870 2174 72922
rect 2226 72870 5152 72922
rect 1104 72848 5152 72870
rect 84180 72922 90896 72944
rect 84180 72870 85982 72922
rect 86034 72870 86046 72922
rect 86098 72870 86110 72922
rect 86162 72870 86174 72922
rect 86226 72870 89982 72922
rect 90034 72870 90046 72922
rect 90098 72870 90110 72922
rect 90162 72870 90174 72922
rect 90226 72870 90896 72922
rect 84180 72848 90896 72870
rect 1104 72378 5152 72400
rect 1104 72326 3982 72378
rect 4034 72326 4046 72378
rect 4098 72326 4110 72378
rect 4162 72326 4174 72378
rect 4226 72326 5152 72378
rect 1104 72304 5152 72326
rect 84180 72378 90896 72400
rect 84180 72326 87982 72378
rect 88034 72326 88046 72378
rect 88098 72326 88110 72378
rect 88162 72326 88174 72378
rect 88226 72326 90896 72378
rect 84180 72304 90896 72326
rect 1104 71834 5152 71856
rect 1104 71782 1982 71834
rect 2034 71782 2046 71834
rect 2098 71782 2110 71834
rect 2162 71782 2174 71834
rect 2226 71782 5152 71834
rect 1104 71760 5152 71782
rect 84180 71834 90896 71856
rect 84180 71782 85982 71834
rect 86034 71782 86046 71834
rect 86098 71782 86110 71834
rect 86162 71782 86174 71834
rect 86226 71782 89982 71834
rect 90034 71782 90046 71834
rect 90098 71782 90110 71834
rect 90162 71782 90174 71834
rect 90226 71782 90896 71834
rect 84180 71760 90896 71782
rect 1104 71290 5152 71312
rect 1104 71238 3982 71290
rect 4034 71238 4046 71290
rect 4098 71238 4110 71290
rect 4162 71238 4174 71290
rect 4226 71238 5152 71290
rect 1104 71216 5152 71238
rect 84180 71290 90896 71312
rect 84180 71238 87982 71290
rect 88034 71238 88046 71290
rect 88098 71238 88110 71290
rect 88162 71238 88174 71290
rect 88226 71238 90896 71290
rect 84180 71216 90896 71238
rect 1104 70746 5152 70768
rect 1104 70694 1982 70746
rect 2034 70694 2046 70746
rect 2098 70694 2110 70746
rect 2162 70694 2174 70746
rect 2226 70694 5152 70746
rect 1104 70672 5152 70694
rect 84180 70746 90896 70768
rect 84180 70694 85982 70746
rect 86034 70694 86046 70746
rect 86098 70694 86110 70746
rect 86162 70694 86174 70746
rect 86226 70694 89982 70746
rect 90034 70694 90046 70746
rect 90098 70694 90110 70746
rect 90162 70694 90174 70746
rect 90226 70694 90896 70746
rect 84180 70672 90896 70694
rect 84010 70320 84016 70372
rect 84068 70360 84074 70372
rect 87782 70360 87788 70372
rect 84068 70332 87788 70360
rect 84068 70320 84074 70332
rect 87782 70320 87788 70332
rect 87840 70320 87846 70372
rect 1104 70202 5152 70224
rect 1104 70150 3982 70202
rect 4034 70150 4046 70202
rect 4098 70150 4110 70202
rect 4162 70150 4174 70202
rect 4226 70150 5152 70202
rect 1104 70128 5152 70150
rect 84180 70202 90896 70224
rect 84180 70150 87982 70202
rect 88034 70150 88046 70202
rect 88098 70150 88110 70202
rect 88162 70150 88174 70202
rect 88226 70150 90896 70202
rect 84180 70128 90896 70150
rect 1104 69658 5152 69680
rect 1104 69606 1982 69658
rect 2034 69606 2046 69658
rect 2098 69606 2110 69658
rect 2162 69606 2174 69658
rect 2226 69606 5152 69658
rect 1104 69584 5152 69606
rect 84180 69658 90896 69680
rect 84180 69606 85982 69658
rect 86034 69606 86046 69658
rect 86098 69606 86110 69658
rect 86162 69606 86174 69658
rect 86226 69606 89982 69658
rect 90034 69606 90046 69658
rect 90098 69606 90110 69658
rect 90162 69606 90174 69658
rect 90226 69606 90896 69658
rect 84180 69584 90896 69606
rect 1104 69114 5152 69136
rect 1104 69062 3982 69114
rect 4034 69062 4046 69114
rect 4098 69062 4110 69114
rect 4162 69062 4174 69114
rect 4226 69062 5152 69114
rect 1104 69040 5152 69062
rect 84180 69114 90896 69136
rect 84180 69062 87982 69114
rect 88034 69062 88046 69114
rect 88098 69062 88110 69114
rect 88162 69062 88174 69114
rect 88226 69062 90896 69114
rect 84180 69040 90896 69062
rect 83918 68960 83924 69012
rect 83976 69000 83982 69012
rect 87138 69000 87144 69012
rect 83976 68972 87144 69000
rect 83976 68960 83982 68972
rect 87138 68960 87144 68972
rect 87196 68960 87202 69012
rect 1104 68570 5152 68592
rect 1104 68518 1982 68570
rect 2034 68518 2046 68570
rect 2098 68518 2110 68570
rect 2162 68518 2174 68570
rect 2226 68518 5152 68570
rect 1104 68496 5152 68518
rect 84180 68570 90896 68592
rect 84180 68518 85982 68570
rect 86034 68518 86046 68570
rect 86098 68518 86110 68570
rect 86162 68518 86174 68570
rect 86226 68518 89982 68570
rect 90034 68518 90046 68570
rect 90098 68518 90110 68570
rect 90162 68518 90174 68570
rect 90226 68518 90896 68570
rect 84180 68496 90896 68518
rect 1104 68026 5152 68048
rect 1104 67974 3982 68026
rect 4034 67974 4046 68026
rect 4098 67974 4110 68026
rect 4162 67974 4174 68026
rect 4226 67974 5152 68026
rect 1104 67952 5152 67974
rect 84180 68026 90896 68048
rect 84180 67974 87982 68026
rect 88034 67974 88046 68026
rect 88098 67974 88110 68026
rect 88162 67974 88174 68026
rect 88226 67974 90896 68026
rect 84180 67952 90896 67974
rect 1104 67482 5152 67504
rect 1104 67430 1982 67482
rect 2034 67430 2046 67482
rect 2098 67430 2110 67482
rect 2162 67430 2174 67482
rect 2226 67430 5152 67482
rect 1104 67408 5152 67430
rect 84180 67482 90896 67504
rect 84180 67430 85982 67482
rect 86034 67430 86046 67482
rect 86098 67430 86110 67482
rect 86162 67430 86174 67482
rect 86226 67430 89982 67482
rect 90034 67430 90046 67482
rect 90098 67430 90110 67482
rect 90162 67430 90174 67482
rect 90226 67430 90896 67482
rect 84180 67408 90896 67430
rect 1104 66938 5152 66960
rect 1104 66886 3982 66938
rect 4034 66886 4046 66938
rect 4098 66886 4110 66938
rect 4162 66886 4174 66938
rect 4226 66886 5152 66938
rect 1104 66864 5152 66886
rect 84180 66938 90896 66960
rect 84180 66886 87982 66938
rect 88034 66886 88046 66938
rect 88098 66886 88110 66938
rect 88162 66886 88174 66938
rect 88226 66886 90896 66938
rect 84180 66864 90896 66886
rect 1104 66394 5152 66416
rect 1104 66342 1982 66394
rect 2034 66342 2046 66394
rect 2098 66342 2110 66394
rect 2162 66342 2174 66394
rect 2226 66342 5152 66394
rect 1104 66320 5152 66342
rect 84180 66394 90896 66416
rect 84180 66342 85982 66394
rect 86034 66342 86046 66394
rect 86098 66342 86110 66394
rect 86162 66342 86174 66394
rect 86226 66342 89982 66394
rect 90034 66342 90046 66394
rect 90098 66342 90110 66394
rect 90162 66342 90174 66394
rect 90226 66342 90896 66394
rect 84180 66320 90896 66342
rect 83826 66172 83832 66224
rect 83884 66212 83890 66224
rect 87782 66212 87788 66224
rect 83884 66184 87788 66212
rect 83884 66172 83890 66184
rect 87782 66172 87788 66184
rect 87840 66172 87846 66224
rect 84194 66104 84200 66156
rect 84252 66144 84258 66156
rect 87322 66144 87328 66156
rect 84252 66116 87328 66144
rect 84252 66104 84258 66116
rect 87322 66104 87328 66116
rect 87380 66104 87386 66156
rect 1104 65850 5152 65872
rect 1104 65798 3982 65850
rect 4034 65798 4046 65850
rect 4098 65798 4110 65850
rect 4162 65798 4174 65850
rect 4226 65798 5152 65850
rect 1104 65776 5152 65798
rect 84180 65850 90896 65872
rect 84180 65798 87982 65850
rect 88034 65798 88046 65850
rect 88098 65798 88110 65850
rect 88162 65798 88174 65850
rect 88226 65798 90896 65850
rect 84180 65776 90896 65798
rect 1104 65306 5152 65328
rect 1104 65254 1982 65306
rect 2034 65254 2046 65306
rect 2098 65254 2110 65306
rect 2162 65254 2174 65306
rect 2226 65254 5152 65306
rect 1104 65232 5152 65254
rect 84180 65306 90896 65328
rect 84180 65254 85982 65306
rect 86034 65254 86046 65306
rect 86098 65254 86110 65306
rect 86162 65254 86174 65306
rect 86226 65254 89982 65306
rect 90034 65254 90046 65306
rect 90098 65254 90110 65306
rect 90162 65254 90174 65306
rect 90226 65254 90896 65306
rect 84180 65232 90896 65254
rect 1104 64762 5152 64784
rect 1104 64710 3982 64762
rect 4034 64710 4046 64762
rect 4098 64710 4110 64762
rect 4162 64710 4174 64762
rect 4226 64710 5152 64762
rect 1104 64688 5152 64710
rect 84180 64762 90896 64784
rect 84180 64710 87982 64762
rect 88034 64710 88046 64762
rect 88098 64710 88110 64762
rect 88162 64710 88174 64762
rect 88226 64710 90896 64762
rect 84180 64688 90896 64710
rect 1104 64218 5152 64240
rect 1104 64166 1982 64218
rect 2034 64166 2046 64218
rect 2098 64166 2110 64218
rect 2162 64166 2174 64218
rect 2226 64166 5152 64218
rect 1104 64144 5152 64166
rect 84180 64218 90896 64240
rect 84180 64166 85982 64218
rect 86034 64166 86046 64218
rect 86098 64166 86110 64218
rect 86162 64166 86174 64218
rect 86226 64166 89982 64218
rect 90034 64166 90046 64218
rect 90098 64166 90110 64218
rect 90162 64166 90174 64218
rect 90226 64166 90896 64218
rect 84180 64144 90896 64166
rect 1104 63674 5152 63696
rect 1104 63622 3982 63674
rect 4034 63622 4046 63674
rect 4098 63622 4110 63674
rect 4162 63622 4174 63674
rect 4226 63622 5152 63674
rect 1104 63600 5152 63622
rect 84180 63674 90896 63696
rect 84180 63622 87982 63674
rect 88034 63622 88046 63674
rect 88098 63622 88110 63674
rect 88162 63622 88174 63674
rect 88226 63622 90896 63674
rect 84180 63600 90896 63622
rect 83734 63452 83740 63504
rect 83792 63492 83798 63504
rect 87782 63492 87788 63504
rect 83792 63464 87788 63492
rect 83792 63452 83798 63464
rect 87782 63452 87788 63464
rect 87840 63452 87846 63504
rect 1104 63130 5152 63152
rect 1104 63078 1982 63130
rect 2034 63078 2046 63130
rect 2098 63078 2110 63130
rect 2162 63078 2174 63130
rect 2226 63078 5152 63130
rect 1104 63056 5152 63078
rect 84180 63130 90896 63152
rect 84180 63078 85982 63130
rect 86034 63078 86046 63130
rect 86098 63078 86110 63130
rect 86162 63078 86174 63130
rect 86226 63078 89982 63130
rect 90034 63078 90046 63130
rect 90098 63078 90110 63130
rect 90162 63078 90174 63130
rect 90226 63078 90896 63130
rect 84180 63056 90896 63078
rect 1104 62586 5152 62608
rect 1104 62534 3982 62586
rect 4034 62534 4046 62586
rect 4098 62534 4110 62586
rect 4162 62534 4174 62586
rect 4226 62534 5152 62586
rect 1104 62512 5152 62534
rect 84180 62586 90896 62608
rect 84180 62534 87982 62586
rect 88034 62534 88046 62586
rect 88098 62534 88110 62586
rect 88162 62534 88174 62586
rect 88226 62534 90896 62586
rect 84180 62512 90896 62534
rect 1104 62042 5152 62064
rect 1104 61990 1982 62042
rect 2034 61990 2046 62042
rect 2098 61990 2110 62042
rect 2162 61990 2174 62042
rect 2226 61990 5152 62042
rect 1104 61968 5152 61990
rect 84180 62042 90896 62064
rect 84180 61990 85982 62042
rect 86034 61990 86046 62042
rect 86098 61990 86110 62042
rect 86162 61990 86174 62042
rect 86226 61990 89982 62042
rect 90034 61990 90046 62042
rect 90098 61990 90110 62042
rect 90162 61990 90174 62042
rect 90226 61990 90896 62042
rect 84180 61968 90896 61990
rect 84286 61888 84292 61940
rect 84344 61928 84350 61940
rect 87782 61928 87788 61940
rect 84344 61900 87788 61928
rect 84344 61888 84350 61900
rect 87782 61888 87788 61900
rect 87840 61888 87846 61940
rect 1104 61498 5152 61520
rect 1104 61446 3982 61498
rect 4034 61446 4046 61498
rect 4098 61446 4110 61498
rect 4162 61446 4174 61498
rect 4226 61446 5152 61498
rect 1104 61424 5152 61446
rect 84180 61498 90896 61520
rect 84180 61446 87982 61498
rect 88034 61446 88046 61498
rect 88098 61446 88110 61498
rect 88162 61446 88174 61498
rect 88226 61446 90896 61498
rect 84180 61424 90896 61446
rect 1104 60954 5152 60976
rect 1104 60902 1982 60954
rect 2034 60902 2046 60954
rect 2098 60902 2110 60954
rect 2162 60902 2174 60954
rect 2226 60902 5152 60954
rect 1104 60880 5152 60902
rect 84180 60954 90896 60976
rect 84180 60902 85982 60954
rect 86034 60902 86046 60954
rect 86098 60902 86110 60954
rect 86162 60902 86174 60954
rect 86226 60902 89982 60954
rect 90034 60902 90046 60954
rect 90098 60902 90110 60954
rect 90162 60902 90174 60954
rect 90226 60902 90896 60954
rect 84180 60880 90896 60902
rect 1104 60410 5152 60432
rect 1104 60358 3982 60410
rect 4034 60358 4046 60410
rect 4098 60358 4110 60410
rect 4162 60358 4174 60410
rect 4226 60358 5152 60410
rect 1104 60336 5152 60358
rect 84180 60410 90896 60432
rect 84180 60358 87982 60410
rect 88034 60358 88046 60410
rect 88098 60358 88110 60410
rect 88162 60358 88174 60410
rect 88226 60358 90896 60410
rect 84180 60336 90896 60358
rect 1104 59866 5152 59888
rect 1104 59814 1982 59866
rect 2034 59814 2046 59866
rect 2098 59814 2110 59866
rect 2162 59814 2174 59866
rect 2226 59814 5152 59866
rect 1104 59792 5152 59814
rect 84180 59866 90896 59888
rect 84180 59814 85982 59866
rect 86034 59814 86046 59866
rect 86098 59814 86110 59866
rect 86162 59814 86174 59866
rect 86226 59814 89982 59866
rect 90034 59814 90046 59866
rect 90098 59814 90110 59866
rect 90162 59814 90174 59866
rect 90226 59814 90896 59866
rect 84180 59792 90896 59814
rect 1104 59322 5152 59344
rect 1104 59270 3982 59322
rect 4034 59270 4046 59322
rect 4098 59270 4110 59322
rect 4162 59270 4174 59322
rect 4226 59270 5152 59322
rect 1104 59248 5152 59270
rect 84180 59322 90896 59344
rect 84180 59270 87982 59322
rect 88034 59270 88046 59322
rect 88098 59270 88110 59322
rect 88162 59270 88174 59322
rect 88226 59270 90896 59322
rect 84180 59248 90896 59270
rect 1104 58778 5152 58800
rect 1104 58726 1982 58778
rect 2034 58726 2046 58778
rect 2098 58726 2110 58778
rect 2162 58726 2174 58778
rect 2226 58726 5152 58778
rect 1104 58704 5152 58726
rect 84180 58778 90896 58800
rect 84180 58726 85982 58778
rect 86034 58726 86046 58778
rect 86098 58726 86110 58778
rect 86162 58726 86174 58778
rect 86226 58726 89982 58778
rect 90034 58726 90046 58778
rect 90098 58726 90110 58778
rect 90162 58726 90174 58778
rect 90226 58726 90896 58778
rect 84180 58704 90896 58726
rect 1104 58234 5152 58256
rect 1104 58182 3982 58234
rect 4034 58182 4046 58234
rect 4098 58182 4110 58234
rect 4162 58182 4174 58234
rect 4226 58182 5152 58234
rect 1104 58160 5152 58182
rect 84180 58234 90896 58256
rect 84180 58182 87982 58234
rect 88034 58182 88046 58234
rect 88098 58182 88110 58234
rect 88162 58182 88174 58234
rect 88226 58182 90896 58234
rect 84180 58160 90896 58182
rect 4433 57919 4491 57925
rect 4433 57885 4445 57919
rect 4479 57916 4491 57919
rect 4522 57916 4528 57928
rect 4479 57888 4528 57916
rect 4479 57885 4491 57888
rect 4433 57879 4491 57885
rect 4522 57876 4528 57888
rect 4580 57876 4586 57928
rect 84746 57876 84752 57928
rect 84804 57916 84810 57928
rect 86954 57916 86960 57928
rect 84804 57888 86960 57916
rect 84804 57876 84810 57888
rect 86954 57876 86960 57888
rect 87012 57876 87018 57928
rect 1104 57690 5152 57712
rect 1104 57638 1982 57690
rect 2034 57638 2046 57690
rect 2098 57638 2110 57690
rect 2162 57638 2174 57690
rect 2226 57638 5152 57690
rect 1104 57616 5152 57638
rect 84180 57690 90896 57712
rect 84180 57638 85982 57690
rect 86034 57638 86046 57690
rect 86098 57638 86110 57690
rect 86162 57638 86174 57690
rect 86226 57638 89982 57690
rect 90034 57638 90046 57690
rect 90098 57638 90110 57690
rect 90162 57638 90174 57690
rect 90226 57638 90896 57690
rect 84180 57616 90896 57638
rect 1104 57146 5152 57168
rect 1104 57094 3982 57146
rect 4034 57094 4046 57146
rect 4098 57094 4110 57146
rect 4162 57094 4174 57146
rect 4226 57094 5152 57146
rect 1104 57072 5152 57094
rect 84180 57146 90896 57168
rect 84180 57094 87982 57146
rect 88034 57094 88046 57146
rect 88098 57094 88110 57146
rect 88162 57094 88174 57146
rect 88226 57094 90896 57146
rect 84180 57072 90896 57094
rect 1104 56602 5152 56624
rect 1104 56550 1982 56602
rect 2034 56550 2046 56602
rect 2098 56550 2110 56602
rect 2162 56550 2174 56602
rect 2226 56550 5152 56602
rect 1104 56528 5152 56550
rect 84180 56602 90896 56624
rect 84180 56550 85982 56602
rect 86034 56550 86046 56602
rect 86098 56550 86110 56602
rect 86162 56550 86174 56602
rect 86226 56550 89982 56602
rect 90034 56550 90046 56602
rect 90098 56550 90110 56602
rect 90162 56550 90174 56602
rect 90226 56550 90896 56602
rect 84180 56528 90896 56550
rect 85482 56448 85488 56500
rect 85540 56488 85546 56500
rect 86954 56488 86960 56500
rect 85540 56460 86960 56488
rect 85540 56448 85546 56460
rect 86954 56448 86960 56460
rect 87012 56448 87018 56500
rect 85114 56380 85120 56432
rect 85172 56420 85178 56432
rect 87046 56420 87052 56432
rect 85172 56392 87052 56420
rect 85172 56380 85178 56392
rect 87046 56380 87052 56392
rect 87104 56380 87110 56432
rect 1104 56058 5152 56080
rect 1104 56006 3982 56058
rect 4034 56006 4046 56058
rect 4098 56006 4110 56058
rect 4162 56006 4174 56058
rect 4226 56006 5152 56058
rect 1104 55984 5152 56006
rect 84180 56058 90896 56080
rect 84180 56006 87982 56058
rect 88034 56006 88046 56058
rect 88098 56006 88110 56058
rect 88162 56006 88174 56058
rect 88226 56006 90896 56058
rect 84180 55984 90896 56006
rect 1104 55514 5152 55536
rect 1104 55462 1982 55514
rect 2034 55462 2046 55514
rect 2098 55462 2110 55514
rect 2162 55462 2174 55514
rect 2226 55462 5152 55514
rect 1104 55440 5152 55462
rect 84180 55514 90896 55536
rect 84180 55462 85982 55514
rect 86034 55462 86046 55514
rect 86098 55462 86110 55514
rect 86162 55462 86174 55514
rect 86226 55462 89982 55514
rect 90034 55462 90046 55514
rect 90098 55462 90110 55514
rect 90162 55462 90174 55514
rect 90226 55462 90896 55514
rect 84180 55440 90896 55462
rect 1104 54970 5152 54992
rect 1104 54918 3982 54970
rect 4034 54918 4046 54970
rect 4098 54918 4110 54970
rect 4162 54918 4174 54970
rect 4226 54918 5152 54970
rect 1104 54896 5152 54918
rect 84180 54970 90896 54992
rect 84180 54918 87982 54970
rect 88034 54918 88046 54970
rect 88098 54918 88110 54970
rect 88162 54918 88174 54970
rect 88226 54918 90896 54970
rect 84180 54896 90896 54918
rect 85206 54612 85212 54664
rect 85264 54652 85270 54664
rect 86954 54652 86960 54664
rect 85264 54624 86960 54652
rect 85264 54612 85270 54624
rect 86954 54612 86960 54624
rect 87012 54612 87018 54664
rect 1104 54426 5152 54448
rect 1104 54374 1982 54426
rect 2034 54374 2046 54426
rect 2098 54374 2110 54426
rect 2162 54374 2174 54426
rect 2226 54374 5152 54426
rect 1104 54352 5152 54374
rect 84180 54426 90896 54448
rect 84180 54374 85982 54426
rect 86034 54374 86046 54426
rect 86098 54374 86110 54426
rect 86162 54374 86174 54426
rect 86226 54374 89982 54426
rect 90034 54374 90046 54426
rect 90098 54374 90110 54426
rect 90162 54374 90174 54426
rect 90226 54374 90896 54426
rect 84180 54352 90896 54374
rect 1104 53882 5152 53904
rect 1104 53830 3982 53882
rect 4034 53830 4046 53882
rect 4098 53830 4110 53882
rect 4162 53830 4174 53882
rect 4226 53830 5152 53882
rect 1104 53808 5152 53830
rect 84180 53882 90896 53904
rect 84180 53830 87982 53882
rect 88034 53830 88046 53882
rect 88098 53830 88110 53882
rect 88162 53830 88174 53882
rect 88226 53830 90896 53882
rect 84180 53808 90896 53830
rect 84838 53728 84844 53780
rect 84896 53768 84902 53780
rect 86954 53768 86960 53780
rect 84896 53740 86960 53768
rect 84896 53728 84902 53740
rect 86954 53728 86960 53740
rect 87012 53728 87018 53780
rect 1104 53338 5152 53360
rect 1104 53286 1982 53338
rect 2034 53286 2046 53338
rect 2098 53286 2110 53338
rect 2162 53286 2174 53338
rect 2226 53286 5152 53338
rect 1104 53264 5152 53286
rect 84180 53338 90896 53360
rect 84180 53286 85982 53338
rect 86034 53286 86046 53338
rect 86098 53286 86110 53338
rect 86162 53286 86174 53338
rect 86226 53286 89982 53338
rect 90034 53286 90046 53338
rect 90098 53286 90110 53338
rect 90162 53286 90174 53338
rect 90226 53286 90896 53338
rect 84180 53264 90896 53286
rect 1104 52794 5152 52816
rect 1104 52742 3982 52794
rect 4034 52742 4046 52794
rect 4098 52742 4110 52794
rect 4162 52742 4174 52794
rect 4226 52742 5152 52794
rect 1104 52720 5152 52742
rect 84180 52794 90896 52816
rect 84180 52742 87982 52794
rect 88034 52742 88046 52794
rect 88098 52742 88110 52794
rect 88162 52742 88174 52794
rect 88226 52742 90896 52794
rect 84180 52720 90896 52742
rect 1104 52250 5152 52272
rect 1104 52198 1982 52250
rect 2034 52198 2046 52250
rect 2098 52198 2110 52250
rect 2162 52198 2174 52250
rect 2226 52198 5152 52250
rect 1104 52176 5152 52198
rect 84180 52250 90896 52272
rect 84180 52198 85982 52250
rect 86034 52198 86046 52250
rect 86098 52198 86110 52250
rect 86162 52198 86174 52250
rect 86226 52198 89982 52250
rect 90034 52198 90046 52250
rect 90098 52198 90110 52250
rect 90162 52198 90174 52250
rect 90226 52198 90896 52250
rect 84180 52176 90896 52198
rect 1104 51706 5152 51728
rect 1104 51654 3982 51706
rect 4034 51654 4046 51706
rect 4098 51654 4110 51706
rect 4162 51654 4174 51706
rect 4226 51654 5152 51706
rect 1104 51632 5152 51654
rect 84180 51706 90896 51728
rect 84180 51654 87982 51706
rect 88034 51654 88046 51706
rect 88098 51654 88110 51706
rect 88162 51654 88174 51706
rect 88226 51654 90896 51706
rect 84180 51632 90896 51654
rect 1104 51162 5152 51184
rect 1104 51110 1982 51162
rect 2034 51110 2046 51162
rect 2098 51110 2110 51162
rect 2162 51110 2174 51162
rect 2226 51110 5152 51162
rect 1104 51088 5152 51110
rect 84180 51162 90896 51184
rect 84180 51110 85982 51162
rect 86034 51110 86046 51162
rect 86098 51110 86110 51162
rect 86162 51110 86174 51162
rect 86226 51110 89982 51162
rect 90034 51110 90046 51162
rect 90098 51110 90110 51162
rect 90162 51110 90174 51162
rect 90226 51110 90896 51162
rect 84180 51088 90896 51110
rect 1104 50618 5152 50640
rect 1104 50566 3982 50618
rect 4034 50566 4046 50618
rect 4098 50566 4110 50618
rect 4162 50566 4174 50618
rect 4226 50566 5152 50618
rect 1104 50544 5152 50566
rect 84180 50618 90896 50640
rect 84180 50566 87982 50618
rect 88034 50566 88046 50618
rect 88098 50566 88110 50618
rect 88162 50566 88174 50618
rect 88226 50566 90896 50618
rect 84180 50544 90896 50566
rect 1104 50074 5152 50096
rect 1104 50022 1982 50074
rect 2034 50022 2046 50074
rect 2098 50022 2110 50074
rect 2162 50022 2174 50074
rect 2226 50022 5152 50074
rect 1104 50000 5152 50022
rect 84180 50074 90896 50096
rect 84180 50022 85982 50074
rect 86034 50022 86046 50074
rect 86098 50022 86110 50074
rect 86162 50022 86174 50074
rect 86226 50022 89982 50074
rect 90034 50022 90046 50074
rect 90098 50022 90110 50074
rect 90162 50022 90174 50074
rect 90226 50022 90896 50074
rect 84180 50000 90896 50022
rect 4430 49960 4436 49972
rect 4391 49932 4436 49960
rect 4430 49920 4436 49932
rect 4488 49920 4494 49972
rect 82722 49648 82728 49700
rect 82780 49688 82786 49700
rect 87690 49688 87696 49700
rect 82780 49660 87696 49688
rect 82780 49648 82786 49660
rect 87690 49648 87696 49660
rect 87748 49648 87754 49700
rect 1104 49530 5152 49552
rect 1104 49478 3982 49530
rect 4034 49478 4046 49530
rect 4098 49478 4110 49530
rect 4162 49478 4174 49530
rect 4226 49478 5152 49530
rect 1104 49456 5152 49478
rect 84180 49530 90896 49552
rect 84180 49478 87982 49530
rect 88034 49478 88046 49530
rect 88098 49478 88110 49530
rect 88162 49478 88174 49530
rect 88226 49478 90896 49530
rect 84180 49456 90896 49478
rect 1104 48986 5152 49008
rect 1104 48934 1982 48986
rect 2034 48934 2046 48986
rect 2098 48934 2110 48986
rect 2162 48934 2174 48986
rect 2226 48934 5152 48986
rect 1104 48912 5152 48934
rect 84180 48986 90896 49008
rect 84180 48934 85982 48986
rect 86034 48934 86046 48986
rect 86098 48934 86110 48986
rect 86162 48934 86174 48986
rect 86226 48934 89982 48986
rect 90034 48934 90046 48986
rect 90098 48934 90110 48986
rect 90162 48934 90174 48986
rect 90226 48934 90896 48986
rect 84180 48912 90896 48934
rect 1104 48442 5152 48464
rect 1104 48390 3982 48442
rect 4034 48390 4046 48442
rect 4098 48390 4110 48442
rect 4162 48390 4174 48442
rect 4226 48390 5152 48442
rect 1104 48368 5152 48390
rect 84180 48442 90896 48464
rect 84180 48390 87982 48442
rect 88034 48390 88046 48442
rect 88098 48390 88110 48442
rect 88162 48390 88174 48442
rect 88226 48390 90896 48442
rect 84180 48368 90896 48390
rect 1104 47898 5152 47920
rect 1104 47846 1982 47898
rect 2034 47846 2046 47898
rect 2098 47846 2110 47898
rect 2162 47846 2174 47898
rect 2226 47846 5152 47898
rect 1104 47824 5152 47846
rect 84180 47898 90896 47920
rect 84180 47846 85982 47898
rect 86034 47846 86046 47898
rect 86098 47846 86110 47898
rect 86162 47846 86174 47898
rect 86226 47846 89982 47898
rect 90034 47846 90046 47898
rect 90098 47846 90110 47898
rect 90162 47846 90174 47898
rect 90226 47846 90896 47898
rect 84180 47824 90896 47846
rect 1104 47354 5152 47376
rect 1104 47302 3982 47354
rect 4034 47302 4046 47354
rect 4098 47302 4110 47354
rect 4162 47302 4174 47354
rect 4226 47302 5152 47354
rect 1104 47280 5152 47302
rect 84180 47354 90896 47376
rect 84180 47302 87982 47354
rect 88034 47302 88046 47354
rect 88098 47302 88110 47354
rect 88162 47302 88174 47354
rect 88226 47302 90896 47354
rect 84180 47280 90896 47302
rect 1104 46810 5152 46832
rect 1104 46758 1982 46810
rect 2034 46758 2046 46810
rect 2098 46758 2110 46810
rect 2162 46758 2174 46810
rect 2226 46758 5152 46810
rect 1104 46736 5152 46758
rect 84180 46810 90896 46832
rect 84180 46758 85982 46810
rect 86034 46758 86046 46810
rect 86098 46758 86110 46810
rect 86162 46758 86174 46810
rect 86226 46758 89982 46810
rect 90034 46758 90046 46810
rect 90098 46758 90110 46810
rect 90162 46758 90174 46810
rect 90226 46758 90896 46810
rect 84180 46736 90896 46758
rect 1104 46266 5152 46288
rect 1104 46214 3982 46266
rect 4034 46214 4046 46266
rect 4098 46214 4110 46266
rect 4162 46214 4174 46266
rect 4226 46214 5152 46266
rect 1104 46192 5152 46214
rect 84180 46266 90896 46288
rect 84180 46214 87982 46266
rect 88034 46214 88046 46266
rect 88098 46214 88110 46266
rect 88162 46214 88174 46266
rect 88226 46214 90896 46266
rect 84180 46192 90896 46214
rect 1104 45722 5152 45744
rect 1104 45670 1982 45722
rect 2034 45670 2046 45722
rect 2098 45670 2110 45722
rect 2162 45670 2174 45722
rect 2226 45670 5152 45722
rect 1104 45648 5152 45670
rect 84180 45722 90896 45744
rect 84180 45670 85982 45722
rect 86034 45670 86046 45722
rect 86098 45670 86110 45722
rect 86162 45670 86174 45722
rect 86226 45670 89982 45722
rect 90034 45670 90046 45722
rect 90098 45670 90110 45722
rect 90162 45670 90174 45722
rect 90226 45670 90896 45722
rect 84180 45648 90896 45670
rect 83734 45568 83740 45620
rect 83792 45608 83798 45620
rect 87690 45608 87696 45620
rect 83792 45580 87696 45608
rect 83792 45568 83798 45580
rect 87690 45568 87696 45580
rect 87748 45568 87754 45620
rect 1104 45178 5152 45200
rect 1104 45126 3982 45178
rect 4034 45126 4046 45178
rect 4098 45126 4110 45178
rect 4162 45126 4174 45178
rect 4226 45126 5152 45178
rect 1104 45104 5152 45126
rect 84180 45178 90896 45200
rect 84180 45126 87982 45178
rect 88034 45126 88046 45178
rect 88098 45126 88110 45178
rect 88162 45126 88174 45178
rect 88226 45126 90896 45178
rect 84180 45104 90896 45126
rect 1104 44634 5152 44656
rect 1104 44582 1982 44634
rect 2034 44582 2046 44634
rect 2098 44582 2110 44634
rect 2162 44582 2174 44634
rect 2226 44582 5152 44634
rect 1104 44560 5152 44582
rect 84180 44634 90896 44656
rect 84180 44582 85982 44634
rect 86034 44582 86046 44634
rect 86098 44582 86110 44634
rect 86162 44582 86174 44634
rect 86226 44582 89982 44634
rect 90034 44582 90046 44634
rect 90098 44582 90110 44634
rect 90162 44582 90174 44634
rect 90226 44582 90896 44634
rect 84180 44560 90896 44582
rect 83826 44140 83832 44192
rect 83884 44180 83890 44192
rect 87690 44180 87696 44192
rect 83884 44152 87696 44180
rect 83884 44140 83890 44152
rect 87690 44140 87696 44152
rect 87748 44140 87754 44192
rect 1104 44090 5152 44112
rect 1104 44038 3982 44090
rect 4034 44038 4046 44090
rect 4098 44038 4110 44090
rect 4162 44038 4174 44090
rect 4226 44038 5152 44090
rect 1104 44016 5152 44038
rect 84180 44090 90896 44112
rect 84180 44038 87982 44090
rect 88034 44038 88046 44090
rect 88098 44038 88110 44090
rect 88162 44038 88174 44090
rect 88226 44038 90896 44090
rect 84180 44016 90896 44038
rect 1104 43546 5152 43568
rect 1104 43494 1982 43546
rect 2034 43494 2046 43546
rect 2098 43494 2110 43546
rect 2162 43494 2174 43546
rect 2226 43494 5152 43546
rect 1104 43472 5152 43494
rect 84180 43546 90896 43568
rect 84180 43494 85982 43546
rect 86034 43494 86046 43546
rect 86098 43494 86110 43546
rect 86162 43494 86174 43546
rect 86226 43494 89982 43546
rect 90034 43494 90046 43546
rect 90098 43494 90110 43546
rect 90162 43494 90174 43546
rect 90226 43494 90896 43546
rect 84180 43472 90896 43494
rect 1104 43002 5152 43024
rect 1104 42950 3982 43002
rect 4034 42950 4046 43002
rect 4098 42950 4110 43002
rect 4162 42950 4174 43002
rect 4226 42950 5152 43002
rect 1104 42928 5152 42950
rect 84180 43002 90896 43024
rect 84180 42950 87982 43002
rect 88034 42950 88046 43002
rect 88098 42950 88110 43002
rect 88162 42950 88174 43002
rect 88226 42950 90896 43002
rect 84180 42928 90896 42950
rect 1104 42458 5152 42480
rect 1104 42406 1982 42458
rect 2034 42406 2046 42458
rect 2098 42406 2110 42458
rect 2162 42406 2174 42458
rect 2226 42406 5152 42458
rect 1104 42384 5152 42406
rect 84180 42458 90896 42480
rect 84180 42406 85982 42458
rect 86034 42406 86046 42458
rect 86098 42406 86110 42458
rect 86162 42406 86174 42458
rect 86226 42406 89982 42458
rect 90034 42406 90046 42458
rect 90098 42406 90110 42458
rect 90162 42406 90174 42458
rect 90226 42406 90896 42458
rect 84180 42384 90896 42406
rect 1104 41914 5152 41936
rect 1104 41862 3982 41914
rect 4034 41862 4046 41914
rect 4098 41862 4110 41914
rect 4162 41862 4174 41914
rect 4226 41862 5152 41914
rect 1104 41840 5152 41862
rect 84180 41914 90896 41936
rect 84180 41862 87982 41914
rect 88034 41862 88046 41914
rect 88098 41862 88110 41914
rect 88162 41862 88174 41914
rect 88226 41862 90896 41914
rect 84180 41840 90896 41862
rect 1104 41370 5152 41392
rect 1104 41318 1982 41370
rect 2034 41318 2046 41370
rect 2098 41318 2110 41370
rect 2162 41318 2174 41370
rect 2226 41318 5152 41370
rect 1104 41296 5152 41318
rect 84180 41370 90896 41392
rect 84180 41318 85982 41370
rect 86034 41318 86046 41370
rect 86098 41318 86110 41370
rect 86162 41318 86174 41370
rect 86226 41318 89982 41370
rect 90034 41318 90046 41370
rect 90098 41318 90110 41370
rect 90162 41318 90174 41370
rect 90226 41318 90896 41370
rect 84180 41296 90896 41318
rect 1104 40826 5152 40848
rect 1104 40774 3982 40826
rect 4034 40774 4046 40826
rect 4098 40774 4110 40826
rect 4162 40774 4174 40826
rect 4226 40774 5152 40826
rect 1104 40752 5152 40774
rect 84180 40826 90896 40848
rect 84180 40774 87982 40826
rect 88034 40774 88046 40826
rect 88098 40774 88110 40826
rect 88162 40774 88174 40826
rect 88226 40774 90896 40826
rect 84180 40752 90896 40774
rect 87322 40672 87328 40724
rect 87380 40712 87386 40724
rect 87874 40712 87880 40724
rect 87380 40684 87880 40712
rect 87380 40672 87386 40684
rect 87874 40672 87880 40684
rect 87932 40672 87938 40724
rect 1104 40282 5152 40304
rect 1104 40230 1982 40282
rect 2034 40230 2046 40282
rect 2098 40230 2110 40282
rect 2162 40230 2174 40282
rect 2226 40230 5152 40282
rect 1104 40208 5152 40230
rect 84180 40282 90896 40304
rect 84180 40230 85982 40282
rect 86034 40230 86046 40282
rect 86098 40230 86110 40282
rect 86162 40230 86174 40282
rect 86226 40230 89982 40282
rect 90034 40230 90046 40282
rect 90098 40230 90110 40282
rect 90162 40230 90174 40282
rect 90226 40230 90896 40282
rect 84180 40208 90896 40230
rect 84838 40060 84844 40112
rect 84896 40100 84902 40112
rect 87874 40100 87880 40112
rect 84896 40072 87880 40100
rect 84896 40060 84902 40072
rect 87874 40060 87880 40072
rect 87932 40060 87938 40112
rect 1104 39738 5152 39760
rect 1104 39686 3982 39738
rect 4034 39686 4046 39738
rect 4098 39686 4110 39738
rect 4162 39686 4174 39738
rect 4226 39686 5152 39738
rect 1104 39664 5152 39686
rect 84180 39738 90896 39760
rect 84180 39686 87982 39738
rect 88034 39686 88046 39738
rect 88098 39686 88110 39738
rect 88162 39686 88174 39738
rect 88226 39686 90896 39738
rect 84180 39664 90896 39686
rect 1104 39194 5152 39216
rect 1104 39142 1982 39194
rect 2034 39142 2046 39194
rect 2098 39142 2110 39194
rect 2162 39142 2174 39194
rect 2226 39142 5152 39194
rect 1104 39120 5152 39142
rect 84180 39194 90896 39216
rect 84180 39142 85982 39194
rect 86034 39142 86046 39194
rect 86098 39142 86110 39194
rect 86162 39142 86174 39194
rect 86226 39142 89982 39194
rect 90034 39142 90046 39194
rect 90098 39142 90110 39194
rect 90162 39142 90174 39194
rect 90226 39142 90896 39194
rect 84180 39120 90896 39142
rect 84378 39040 84384 39092
rect 84436 39080 84442 39092
rect 84473 39083 84531 39089
rect 84473 39080 84485 39083
rect 84436 39052 84485 39080
rect 84436 39040 84442 39052
rect 84473 39049 84485 39052
rect 84519 39049 84531 39083
rect 84473 39043 84531 39049
rect 1104 38650 5152 38672
rect 1104 38598 3982 38650
rect 4034 38598 4046 38650
rect 4098 38598 4110 38650
rect 4162 38598 4174 38650
rect 4226 38598 5152 38650
rect 1104 38576 5152 38598
rect 84180 38650 90896 38672
rect 84180 38598 87982 38650
rect 88034 38598 88046 38650
rect 88098 38598 88110 38650
rect 88162 38598 88174 38650
rect 88226 38598 90896 38650
rect 84180 38576 90896 38598
rect 1104 38106 5152 38128
rect 1104 38054 1982 38106
rect 2034 38054 2046 38106
rect 2098 38054 2110 38106
rect 2162 38054 2174 38106
rect 2226 38054 5152 38106
rect 1104 38032 5152 38054
rect 84180 38106 90896 38128
rect 84180 38054 85982 38106
rect 86034 38054 86046 38106
rect 86098 38054 86110 38106
rect 86162 38054 86174 38106
rect 86226 38054 89982 38106
rect 90034 38054 90046 38106
rect 90098 38054 90110 38106
rect 90162 38054 90174 38106
rect 90226 38054 90896 38106
rect 84180 38032 90896 38054
rect 1104 37562 5152 37584
rect 1104 37510 3982 37562
rect 4034 37510 4046 37562
rect 4098 37510 4110 37562
rect 4162 37510 4174 37562
rect 4226 37510 5152 37562
rect 1104 37488 5152 37510
rect 84180 37562 90896 37584
rect 84180 37510 87982 37562
rect 88034 37510 88046 37562
rect 88098 37510 88110 37562
rect 88162 37510 88174 37562
rect 88226 37510 90896 37562
rect 84180 37488 90896 37510
rect 1104 37018 5152 37040
rect 1104 36966 1982 37018
rect 2034 36966 2046 37018
rect 2098 36966 2110 37018
rect 2162 36966 2174 37018
rect 2226 36966 5152 37018
rect 1104 36944 5152 36966
rect 84180 37018 90896 37040
rect 84180 36966 85982 37018
rect 86034 36966 86046 37018
rect 86098 36966 86110 37018
rect 86162 36966 86174 37018
rect 86226 36966 89982 37018
rect 90034 36966 90046 37018
rect 90098 36966 90110 37018
rect 90162 36966 90174 37018
rect 90226 36966 90896 37018
rect 84180 36944 90896 36966
rect 1104 36474 5152 36496
rect 1104 36422 3982 36474
rect 4034 36422 4046 36474
rect 4098 36422 4110 36474
rect 4162 36422 4174 36474
rect 4226 36422 5152 36474
rect 1104 36400 5152 36422
rect 84180 36474 90896 36496
rect 84180 36422 87982 36474
rect 88034 36422 88046 36474
rect 88098 36422 88110 36474
rect 88162 36422 88174 36474
rect 88226 36422 90896 36474
rect 84180 36400 90896 36422
rect 85114 36320 85120 36372
rect 85172 36360 85178 36372
rect 86954 36360 86960 36372
rect 85172 36332 86960 36360
rect 85172 36320 85178 36332
rect 86954 36320 86960 36332
rect 87012 36320 87018 36372
rect 1104 35930 5152 35952
rect 1104 35878 1982 35930
rect 2034 35878 2046 35930
rect 2098 35878 2110 35930
rect 2162 35878 2174 35930
rect 2226 35878 5152 35930
rect 1104 35856 5152 35878
rect 84180 35930 90896 35952
rect 84180 35878 85982 35930
rect 86034 35878 86046 35930
rect 86098 35878 86110 35930
rect 86162 35878 86174 35930
rect 86226 35878 89982 35930
rect 90034 35878 90046 35930
rect 90098 35878 90110 35930
rect 90162 35878 90174 35930
rect 90226 35878 90896 35930
rect 84180 35856 90896 35878
rect 1104 35386 5152 35408
rect 1104 35334 3982 35386
rect 4034 35334 4046 35386
rect 4098 35334 4110 35386
rect 4162 35334 4174 35386
rect 4226 35334 5152 35386
rect 1104 35312 5152 35334
rect 84180 35386 90896 35408
rect 84180 35334 87982 35386
rect 88034 35334 88046 35386
rect 88098 35334 88110 35386
rect 88162 35334 88174 35386
rect 88226 35334 90896 35386
rect 84180 35312 90896 35334
rect 1104 34842 5152 34864
rect 1104 34790 1982 34842
rect 2034 34790 2046 34842
rect 2098 34790 2110 34842
rect 2162 34790 2174 34842
rect 2226 34790 5152 34842
rect 1104 34768 5152 34790
rect 84180 34842 90896 34864
rect 84180 34790 85982 34842
rect 86034 34790 86046 34842
rect 86098 34790 86110 34842
rect 86162 34790 86174 34842
rect 86226 34790 89982 34842
rect 90034 34790 90046 34842
rect 90098 34790 90110 34842
rect 90162 34790 90174 34842
rect 90226 34790 90896 34842
rect 84180 34768 90896 34790
rect 85206 34484 85212 34536
rect 85264 34524 85270 34536
rect 86954 34524 86960 34536
rect 85264 34496 86960 34524
rect 85264 34484 85270 34496
rect 86954 34484 86960 34496
rect 87012 34484 87018 34536
rect 1104 34298 5152 34320
rect 1104 34246 3982 34298
rect 4034 34246 4046 34298
rect 4098 34246 4110 34298
rect 4162 34246 4174 34298
rect 4226 34246 5152 34298
rect 1104 34224 5152 34246
rect 84180 34298 90896 34320
rect 84180 34246 87982 34298
rect 88034 34246 88046 34298
rect 88098 34246 88110 34298
rect 88162 34246 88174 34298
rect 88226 34246 90896 34298
rect 84180 34224 90896 34246
rect 1104 33754 5152 33776
rect 1104 33702 1982 33754
rect 2034 33702 2046 33754
rect 2098 33702 2110 33754
rect 2162 33702 2174 33754
rect 2226 33702 5152 33754
rect 1104 33680 5152 33702
rect 84180 33754 90896 33776
rect 84180 33702 85982 33754
rect 86034 33702 86046 33754
rect 86098 33702 86110 33754
rect 86162 33702 86174 33754
rect 86226 33702 89982 33754
rect 90034 33702 90046 33754
rect 90098 33702 90110 33754
rect 90162 33702 90174 33754
rect 90226 33702 90896 33754
rect 84180 33680 90896 33702
rect 1104 33210 5152 33232
rect 1104 33158 3982 33210
rect 4034 33158 4046 33210
rect 4098 33158 4110 33210
rect 4162 33158 4174 33210
rect 4226 33158 5152 33210
rect 1104 33136 5152 33158
rect 84180 33210 90896 33232
rect 84180 33158 87982 33210
rect 88034 33158 88046 33210
rect 88098 33158 88110 33210
rect 88162 33158 88174 33210
rect 88226 33158 90896 33210
rect 84180 33136 90896 33158
rect 1104 32666 5152 32688
rect 1104 32614 1982 32666
rect 2034 32614 2046 32666
rect 2098 32614 2110 32666
rect 2162 32614 2174 32666
rect 2226 32614 5152 32666
rect 1104 32592 5152 32614
rect 84180 32666 90896 32688
rect 84180 32614 85982 32666
rect 86034 32614 86046 32666
rect 86098 32614 86110 32666
rect 86162 32614 86174 32666
rect 86226 32614 89982 32666
rect 90034 32614 90046 32666
rect 90098 32614 90110 32666
rect 90162 32614 90174 32666
rect 90226 32614 90896 32666
rect 84180 32592 90896 32614
rect 1104 32122 5152 32144
rect 1104 32070 3982 32122
rect 4034 32070 4046 32122
rect 4098 32070 4110 32122
rect 4162 32070 4174 32122
rect 4226 32070 5152 32122
rect 1104 32048 5152 32070
rect 84180 32122 90896 32144
rect 84180 32070 87982 32122
rect 88034 32070 88046 32122
rect 88098 32070 88110 32122
rect 88162 32070 88174 32122
rect 88226 32070 90896 32122
rect 84180 32048 90896 32070
rect 84746 32008 84752 32020
rect 84659 31980 84752 32008
rect 84746 31968 84752 31980
rect 84804 32008 84810 32020
rect 86586 32008 86592 32020
rect 84804 31980 86592 32008
rect 84804 31968 84810 31980
rect 86586 31968 86592 31980
rect 86644 31968 86650 32020
rect 85482 31764 85488 31816
rect 85540 31804 85546 31816
rect 86954 31804 86960 31816
rect 85540 31776 86960 31804
rect 85540 31764 85546 31776
rect 86954 31764 86960 31776
rect 87012 31764 87018 31816
rect 1104 31578 5152 31600
rect 1104 31526 1982 31578
rect 2034 31526 2046 31578
rect 2098 31526 2110 31578
rect 2162 31526 2174 31578
rect 2226 31526 5152 31578
rect 1104 31504 5152 31526
rect 84180 31578 90896 31600
rect 84180 31526 85982 31578
rect 86034 31526 86046 31578
rect 86098 31526 86110 31578
rect 86162 31526 86174 31578
rect 86226 31526 89982 31578
rect 90034 31526 90046 31578
rect 90098 31526 90110 31578
rect 90162 31526 90174 31578
rect 90226 31526 90896 31578
rect 84180 31504 90896 31526
rect 1104 31034 5152 31056
rect 1104 30982 3982 31034
rect 4034 30982 4046 31034
rect 4098 30982 4110 31034
rect 4162 30982 4174 31034
rect 4226 30982 5152 31034
rect 1104 30960 5152 30982
rect 84180 31034 90896 31056
rect 84180 30982 87982 31034
rect 88034 30982 88046 31034
rect 88098 30982 88110 31034
rect 88162 30982 88174 31034
rect 88226 30982 90896 31034
rect 84180 30960 90896 30982
rect 1104 30490 5152 30512
rect 1104 30438 1982 30490
rect 2034 30438 2046 30490
rect 2098 30438 2110 30490
rect 2162 30438 2174 30490
rect 2226 30438 5152 30490
rect 1104 30416 5152 30438
rect 84180 30490 90896 30512
rect 84180 30438 85982 30490
rect 86034 30438 86046 30490
rect 86098 30438 86110 30490
rect 86162 30438 86174 30490
rect 86226 30438 89982 30490
rect 90034 30438 90046 30490
rect 90098 30438 90110 30490
rect 90162 30438 90174 30490
rect 90226 30438 90896 30490
rect 84180 30416 90896 30438
rect 84746 30308 84752 30320
rect 84659 30280 84752 30308
rect 84746 30268 84752 30280
rect 84804 30308 84810 30320
rect 87230 30308 87236 30320
rect 84804 30280 87236 30308
rect 84804 30268 84810 30280
rect 87230 30268 87236 30280
rect 87288 30268 87294 30320
rect 1104 29946 5152 29968
rect 1104 29894 3982 29946
rect 4034 29894 4046 29946
rect 4098 29894 4110 29946
rect 4162 29894 4174 29946
rect 4226 29894 5152 29946
rect 1104 29872 5152 29894
rect 84180 29946 90896 29968
rect 84180 29894 87982 29946
rect 88034 29894 88046 29946
rect 88098 29894 88110 29946
rect 88162 29894 88174 29946
rect 88226 29894 90896 29946
rect 84180 29872 90896 29894
rect 1104 29402 5152 29424
rect 1104 29350 1982 29402
rect 2034 29350 2046 29402
rect 2098 29350 2110 29402
rect 2162 29350 2174 29402
rect 2226 29350 5152 29402
rect 1104 29328 5152 29350
rect 84180 29402 90896 29424
rect 84180 29350 85982 29402
rect 86034 29350 86046 29402
rect 86098 29350 86110 29402
rect 86162 29350 86174 29402
rect 86226 29350 89982 29402
rect 90034 29350 90046 29402
rect 90098 29350 90110 29402
rect 90162 29350 90174 29402
rect 90226 29350 90896 29402
rect 84180 29328 90896 29350
rect 84562 29248 84568 29300
rect 84620 29288 84626 29300
rect 84749 29291 84807 29297
rect 84749 29288 84761 29291
rect 84620 29260 84761 29288
rect 84620 29248 84626 29260
rect 84749 29257 84761 29260
rect 84795 29288 84807 29291
rect 86494 29288 86500 29300
rect 84795 29260 86500 29288
rect 84795 29257 84807 29260
rect 84749 29251 84807 29257
rect 86494 29248 86500 29260
rect 86552 29248 86558 29300
rect 84746 28976 84752 29028
rect 84804 29016 84810 29028
rect 86954 29016 86960 29028
rect 84804 28988 86960 29016
rect 84804 28976 84810 28988
rect 86954 28976 86960 28988
rect 87012 28976 87018 29028
rect 1104 28858 5152 28880
rect 1104 28806 3982 28858
rect 4034 28806 4046 28858
rect 4098 28806 4110 28858
rect 4162 28806 4174 28858
rect 4226 28806 5152 28858
rect 1104 28784 5152 28806
rect 84180 28858 90896 28880
rect 84180 28806 87982 28858
rect 88034 28806 88046 28858
rect 88098 28806 88110 28858
rect 88162 28806 88174 28858
rect 88226 28806 90896 28858
rect 84180 28784 90896 28806
rect 1104 28314 5152 28336
rect 1104 28262 1982 28314
rect 2034 28262 2046 28314
rect 2098 28262 2110 28314
rect 2162 28262 2174 28314
rect 2226 28262 5152 28314
rect 1104 28240 5152 28262
rect 84180 28314 90896 28336
rect 84180 28262 85982 28314
rect 86034 28262 86046 28314
rect 86098 28262 86110 28314
rect 86162 28262 86174 28314
rect 86226 28262 89982 28314
rect 90034 28262 90046 28314
rect 90098 28262 90110 28314
rect 90162 28262 90174 28314
rect 90226 28262 90896 28314
rect 84180 28240 90896 28262
rect 1104 27770 5152 27792
rect 1104 27718 3982 27770
rect 4034 27718 4046 27770
rect 4098 27718 4110 27770
rect 4162 27718 4174 27770
rect 4226 27718 5152 27770
rect 1104 27696 5152 27718
rect 84180 27770 90896 27792
rect 84180 27718 87982 27770
rect 88034 27718 88046 27770
rect 88098 27718 88110 27770
rect 88162 27718 88174 27770
rect 88226 27718 90896 27770
rect 84180 27696 90896 27718
rect 83918 27616 83924 27668
rect 83976 27656 83982 27668
rect 86954 27656 86960 27668
rect 83976 27628 86960 27656
rect 83976 27616 83982 27628
rect 86954 27616 86960 27628
rect 87012 27616 87018 27668
rect 84562 27548 84568 27600
rect 84620 27588 84626 27600
rect 84749 27591 84807 27597
rect 84749 27588 84761 27591
rect 84620 27560 84761 27588
rect 84620 27548 84626 27560
rect 84749 27557 84761 27560
rect 84795 27588 84807 27591
rect 86402 27588 86408 27600
rect 84795 27560 86408 27588
rect 84795 27557 84807 27560
rect 84749 27551 84807 27557
rect 86402 27548 86408 27560
rect 86460 27548 86466 27600
rect 1104 27226 5152 27248
rect 1104 27174 1982 27226
rect 2034 27174 2046 27226
rect 2098 27174 2110 27226
rect 2162 27174 2174 27226
rect 2226 27174 5152 27226
rect 1104 27152 5152 27174
rect 84180 27226 90896 27248
rect 84180 27174 85982 27226
rect 86034 27174 86046 27226
rect 86098 27174 86110 27226
rect 86162 27174 86174 27226
rect 86226 27174 89982 27226
rect 90034 27174 90046 27226
rect 90098 27174 90110 27226
rect 90162 27174 90174 27226
rect 90226 27174 90896 27226
rect 84180 27152 90896 27174
rect 1104 26682 5152 26704
rect 1104 26630 3982 26682
rect 4034 26630 4046 26682
rect 4098 26630 4110 26682
rect 4162 26630 4174 26682
rect 4226 26630 5152 26682
rect 1104 26608 5152 26630
rect 84180 26682 90896 26704
rect 84180 26630 87982 26682
rect 88034 26630 88046 26682
rect 88098 26630 88110 26682
rect 88162 26630 88174 26682
rect 88226 26630 90896 26682
rect 84180 26608 90896 26630
rect 84562 26528 84568 26580
rect 84620 26568 84626 26580
rect 84749 26571 84807 26577
rect 84749 26568 84761 26571
rect 84620 26540 84761 26568
rect 84620 26528 84626 26540
rect 84749 26537 84761 26540
rect 84795 26568 84807 26571
rect 86310 26568 86316 26580
rect 84795 26540 86316 26568
rect 84795 26537 84807 26540
rect 84749 26531 84807 26537
rect 86310 26528 86316 26540
rect 86368 26528 86374 26580
rect 84010 26256 84016 26308
rect 84068 26296 84074 26308
rect 86954 26296 86960 26308
rect 84068 26268 86960 26296
rect 84068 26256 84074 26268
rect 86954 26256 86960 26268
rect 87012 26256 87018 26308
rect 1104 26138 5152 26160
rect 1104 26086 1982 26138
rect 2034 26086 2046 26138
rect 2098 26086 2110 26138
rect 2162 26086 2174 26138
rect 2226 26086 5152 26138
rect 1104 26064 5152 26086
rect 84180 26138 90896 26160
rect 84180 26086 85982 26138
rect 86034 26086 86046 26138
rect 86098 26086 86110 26138
rect 86162 26086 86174 26138
rect 86226 26086 89982 26138
rect 90034 26086 90046 26138
rect 90098 26086 90110 26138
rect 90162 26086 90174 26138
rect 90226 26086 90896 26138
rect 84180 26064 90896 26086
rect 1104 25594 5152 25616
rect 1104 25542 3982 25594
rect 4034 25542 4046 25594
rect 4098 25542 4110 25594
rect 4162 25542 4174 25594
rect 4226 25542 5152 25594
rect 1104 25520 5152 25542
rect 84180 25594 90896 25616
rect 84180 25542 87982 25594
rect 88034 25542 88046 25594
rect 88098 25542 88110 25594
rect 88162 25542 88174 25594
rect 88226 25542 90896 25594
rect 84180 25520 90896 25542
rect 1104 25050 5152 25072
rect 1104 24998 1982 25050
rect 2034 24998 2046 25050
rect 2098 24998 2110 25050
rect 2162 24998 2174 25050
rect 2226 24998 5152 25050
rect 1104 24976 5152 24998
rect 84180 25050 90896 25072
rect 84180 24998 85982 25050
rect 86034 24998 86046 25050
rect 86098 24998 86110 25050
rect 86162 24998 86174 25050
rect 86226 24998 89982 25050
rect 90034 24998 90046 25050
rect 90098 24998 90110 25050
rect 90162 24998 90174 25050
rect 90226 24998 90896 25050
rect 84180 24976 90896 24998
rect 1104 24506 5152 24528
rect 1104 24454 3982 24506
rect 4034 24454 4046 24506
rect 4098 24454 4110 24506
rect 4162 24454 4174 24506
rect 4226 24454 5152 24506
rect 1104 24432 5152 24454
rect 84180 24506 90896 24528
rect 84180 24454 87982 24506
rect 88034 24454 88046 24506
rect 88098 24454 88110 24506
rect 88162 24454 88174 24506
rect 88226 24454 90896 24506
rect 84180 24432 90896 24454
rect 84286 24352 84292 24404
rect 84344 24392 84350 24404
rect 84749 24395 84807 24401
rect 84749 24392 84761 24395
rect 84344 24364 84761 24392
rect 84344 24352 84350 24364
rect 84749 24361 84761 24364
rect 84795 24392 84807 24395
rect 85850 24392 85856 24404
rect 84795 24364 85856 24392
rect 84795 24361 84807 24364
rect 84749 24355 84807 24361
rect 85850 24352 85856 24364
rect 85908 24352 85914 24404
rect 1104 23962 5152 23984
rect 1104 23910 1982 23962
rect 2034 23910 2046 23962
rect 2098 23910 2110 23962
rect 2162 23910 2174 23962
rect 2226 23910 5152 23962
rect 1104 23888 5152 23910
rect 84180 23962 90896 23984
rect 84180 23910 85982 23962
rect 86034 23910 86046 23962
rect 86098 23910 86110 23962
rect 86162 23910 86174 23962
rect 86226 23910 89982 23962
rect 90034 23910 90046 23962
rect 90098 23910 90110 23962
rect 90162 23910 90174 23962
rect 90226 23910 90896 23962
rect 84180 23888 90896 23910
rect 83366 23536 83372 23588
rect 83424 23576 83430 23588
rect 87046 23576 87052 23588
rect 83424 23548 87052 23576
rect 83424 23536 83430 23548
rect 87046 23536 87052 23548
rect 87104 23536 87110 23588
rect 84102 23468 84108 23520
rect 84160 23508 84166 23520
rect 86954 23508 86960 23520
rect 84160 23480 86960 23508
rect 84160 23468 84166 23480
rect 86954 23468 86960 23480
rect 87012 23468 87018 23520
rect 1104 23418 5152 23440
rect 1104 23366 3982 23418
rect 4034 23366 4046 23418
rect 4098 23366 4110 23418
rect 4162 23366 4174 23418
rect 4226 23366 5152 23418
rect 1104 23344 5152 23366
rect 84180 23418 90896 23440
rect 84180 23366 87982 23418
rect 88034 23366 88046 23418
rect 88098 23366 88110 23418
rect 88162 23366 88174 23418
rect 88226 23366 90896 23418
rect 84180 23344 90896 23366
rect 84286 23264 84292 23316
rect 84344 23304 84350 23316
rect 84749 23307 84807 23313
rect 84749 23304 84761 23307
rect 84344 23276 84761 23304
rect 84344 23264 84350 23276
rect 84749 23273 84761 23276
rect 84795 23304 84807 23307
rect 85666 23304 85672 23316
rect 84795 23276 85672 23304
rect 84795 23273 84807 23276
rect 84749 23267 84807 23273
rect 85666 23264 85672 23276
rect 85724 23264 85730 23316
rect 1104 22874 5152 22896
rect 1104 22822 1982 22874
rect 2034 22822 2046 22874
rect 2098 22822 2110 22874
rect 2162 22822 2174 22874
rect 2226 22822 5152 22874
rect 1104 22800 5152 22822
rect 84180 22874 90896 22896
rect 84180 22822 85982 22874
rect 86034 22822 86046 22874
rect 86098 22822 86110 22874
rect 86162 22822 86174 22874
rect 86226 22822 89982 22874
rect 90034 22822 90046 22874
rect 90098 22822 90110 22874
rect 90162 22822 90174 22874
rect 90226 22822 90896 22874
rect 84180 22800 90896 22822
rect 4706 22420 4712 22432
rect 4667 22392 4712 22420
rect 4706 22380 4712 22392
rect 4764 22380 4770 22432
rect 1104 22330 5152 22352
rect 1104 22278 3982 22330
rect 4034 22278 4046 22330
rect 4098 22278 4110 22330
rect 4162 22278 4174 22330
rect 4226 22278 5152 22330
rect 1104 22256 5152 22278
rect 84180 22330 90896 22352
rect 84180 22278 87982 22330
rect 88034 22278 88046 22330
rect 88098 22278 88110 22330
rect 88162 22278 88174 22330
rect 88226 22278 90896 22330
rect 84180 22256 90896 22278
rect 84562 22176 84568 22228
rect 84620 22216 84626 22228
rect 87138 22216 87144 22228
rect 84620 22188 87144 22216
rect 84620 22176 84626 22188
rect 87138 22176 87144 22188
rect 87196 22176 87202 22228
rect 1104 21786 5152 21808
rect 1104 21734 1982 21786
rect 2034 21734 2046 21786
rect 2098 21734 2110 21786
rect 2162 21734 2174 21786
rect 2226 21734 5152 21786
rect 1104 21712 5152 21734
rect 84180 21786 90896 21808
rect 84180 21734 85982 21786
rect 86034 21734 86046 21786
rect 86098 21734 86110 21786
rect 86162 21734 86174 21786
rect 86226 21734 89982 21786
rect 90034 21734 90046 21786
rect 90098 21734 90110 21786
rect 90162 21734 90174 21786
rect 90226 21734 90896 21786
rect 84180 21712 90896 21734
rect 1104 21242 5152 21264
rect 1104 21190 3982 21242
rect 4034 21190 4046 21242
rect 4098 21190 4110 21242
rect 4162 21190 4174 21242
rect 4226 21190 5152 21242
rect 1104 21168 5152 21190
rect 84180 21242 90896 21264
rect 84180 21190 87982 21242
rect 88034 21190 88046 21242
rect 88098 21190 88110 21242
rect 88162 21190 88174 21242
rect 88226 21190 90896 21242
rect 84180 21168 90896 21190
rect 4798 20856 4804 20868
rect 4759 20828 4804 20856
rect 4798 20816 4804 20828
rect 4856 20856 4862 20868
rect 4982 20856 4988 20868
rect 4856 20828 4988 20856
rect 4856 20816 4862 20828
rect 4982 20816 4988 20828
rect 5040 20816 5046 20868
rect 83274 20748 83280 20800
rect 83332 20788 83338 20800
rect 87874 20788 87880 20800
rect 83332 20760 87880 20788
rect 83332 20748 83338 20760
rect 87874 20748 87880 20760
rect 87932 20748 87938 20800
rect 1104 20698 5152 20720
rect 1104 20646 1982 20698
rect 2034 20646 2046 20698
rect 2098 20646 2110 20698
rect 2162 20646 2174 20698
rect 2226 20646 5152 20698
rect 1104 20624 5152 20646
rect 84180 20698 90896 20720
rect 84180 20646 85982 20698
rect 86034 20646 86046 20698
rect 86098 20646 86110 20698
rect 86162 20646 86174 20698
rect 86226 20646 89982 20698
rect 90034 20646 90046 20698
rect 90098 20646 90110 20698
rect 90162 20646 90174 20698
rect 90226 20646 90896 20698
rect 84180 20624 90896 20646
rect 87230 20544 87236 20596
rect 87288 20584 87294 20596
rect 87874 20584 87880 20596
rect 87288 20556 87880 20584
rect 87288 20544 87294 20556
rect 87874 20544 87880 20556
rect 87932 20544 87938 20596
rect 1104 20154 5152 20176
rect 1104 20102 3982 20154
rect 4034 20102 4046 20154
rect 4098 20102 4110 20154
rect 4162 20102 4174 20154
rect 4226 20102 5152 20154
rect 1104 20080 5152 20102
rect 84180 20154 90896 20176
rect 84180 20102 87982 20154
rect 88034 20102 88046 20154
rect 88098 20102 88110 20154
rect 88162 20102 88174 20154
rect 88226 20102 90896 20154
rect 84180 20080 90896 20102
rect 1104 19610 5152 19632
rect 1104 19558 1982 19610
rect 2034 19558 2046 19610
rect 2098 19558 2110 19610
rect 2162 19558 2174 19610
rect 2226 19558 5152 19610
rect 1104 19536 5152 19558
rect 84180 19610 90896 19632
rect 84180 19558 85982 19610
rect 86034 19558 86046 19610
rect 86098 19558 86110 19610
rect 86162 19558 86174 19610
rect 86226 19558 89982 19610
rect 90034 19558 90046 19610
rect 90098 19558 90110 19610
rect 90162 19558 90174 19610
rect 90226 19558 90896 19610
rect 84180 19536 90896 19558
rect 1104 19066 5152 19088
rect 1104 19014 3982 19066
rect 4034 19014 4046 19066
rect 4098 19014 4110 19066
rect 4162 19014 4174 19066
rect 4226 19014 5152 19066
rect 1104 18992 5152 19014
rect 84180 19066 90896 19088
rect 84180 19014 87982 19066
rect 88034 19014 88046 19066
rect 88098 19014 88110 19066
rect 88162 19014 88174 19066
rect 88226 19014 90896 19066
rect 84180 18992 90896 19014
rect 1104 18522 5152 18544
rect 1104 18470 1982 18522
rect 2034 18470 2046 18522
rect 2098 18470 2110 18522
rect 2162 18470 2174 18522
rect 2226 18470 5152 18522
rect 1104 18448 5152 18470
rect 84180 18522 90896 18544
rect 84180 18470 85982 18522
rect 86034 18470 86046 18522
rect 86098 18470 86110 18522
rect 86162 18470 86174 18522
rect 86226 18470 89982 18522
rect 90034 18470 90046 18522
rect 90098 18470 90110 18522
rect 90162 18470 90174 18522
rect 90226 18470 90896 18522
rect 84180 18448 90896 18470
rect 1104 17978 5152 18000
rect 1104 17926 3982 17978
rect 4034 17926 4046 17978
rect 4098 17926 4110 17978
rect 4162 17926 4174 17978
rect 4226 17926 5152 17978
rect 1104 17904 5152 17926
rect 84180 17978 90896 18000
rect 84180 17926 87982 17978
rect 88034 17926 88046 17978
rect 88098 17926 88110 17978
rect 88162 17926 88174 17978
rect 88226 17926 90896 17978
rect 84180 17904 90896 17926
rect 84470 17728 84476 17740
rect 84431 17700 84476 17728
rect 84470 17688 84476 17700
rect 84528 17688 84534 17740
rect 1104 17434 5152 17456
rect 1104 17382 1982 17434
rect 2034 17382 2046 17434
rect 2098 17382 2110 17434
rect 2162 17382 2174 17434
rect 2226 17382 5152 17434
rect 1104 17360 5152 17382
rect 84180 17434 90896 17456
rect 84180 17382 85982 17434
rect 86034 17382 86046 17434
rect 86098 17382 86110 17434
rect 86162 17382 86174 17434
rect 86226 17382 89982 17434
rect 90034 17382 90046 17434
rect 90098 17382 90110 17434
rect 90162 17382 90174 17434
rect 90226 17382 90896 17434
rect 84180 17360 90896 17382
rect 1104 16890 5152 16912
rect 1104 16838 3982 16890
rect 4034 16838 4046 16890
rect 4098 16838 4110 16890
rect 4162 16838 4174 16890
rect 4226 16838 5152 16890
rect 1104 16816 5152 16838
rect 84180 16890 90896 16912
rect 84180 16838 87982 16890
rect 88034 16838 88046 16890
rect 88098 16838 88110 16890
rect 88162 16838 88174 16890
rect 88226 16838 90896 16890
rect 84180 16816 90896 16838
rect 87046 16532 87052 16584
rect 87104 16572 87110 16584
rect 87230 16572 87236 16584
rect 87104 16544 87236 16572
rect 87104 16532 87110 16544
rect 87230 16532 87236 16544
rect 87288 16532 87294 16584
rect 1104 16346 5152 16368
rect 1104 16294 1982 16346
rect 2034 16294 2046 16346
rect 2098 16294 2110 16346
rect 2162 16294 2174 16346
rect 2226 16294 5152 16346
rect 1104 16272 5152 16294
rect 84180 16346 90896 16368
rect 84180 16294 85982 16346
rect 86034 16294 86046 16346
rect 86098 16294 86110 16346
rect 86162 16294 86174 16346
rect 86226 16294 89982 16346
rect 90034 16294 90046 16346
rect 90098 16294 90110 16346
rect 90162 16294 90174 16346
rect 90226 16294 90896 16346
rect 84180 16272 90896 16294
rect 1104 15802 5152 15824
rect 1104 15750 3982 15802
rect 4034 15750 4046 15802
rect 4098 15750 4110 15802
rect 4162 15750 4174 15802
rect 4226 15750 5152 15802
rect 1104 15728 5152 15750
rect 84180 15802 90896 15824
rect 84180 15750 87982 15802
rect 88034 15750 88046 15802
rect 88098 15750 88110 15802
rect 88162 15750 88174 15802
rect 88226 15750 90896 15802
rect 84180 15728 90896 15750
rect 84470 15308 84476 15360
rect 84528 15348 84534 15360
rect 87138 15348 87144 15360
rect 84528 15320 87144 15348
rect 84528 15308 84534 15320
rect 87138 15308 87144 15320
rect 87196 15308 87202 15360
rect 1104 15258 5152 15280
rect 1104 15206 1982 15258
rect 2034 15206 2046 15258
rect 2098 15206 2110 15258
rect 2162 15206 2174 15258
rect 2226 15206 5152 15258
rect 1104 15184 5152 15206
rect 84180 15258 90896 15280
rect 84180 15206 85982 15258
rect 86034 15206 86046 15258
rect 86098 15206 86110 15258
rect 86162 15206 86174 15258
rect 86226 15206 89982 15258
rect 90034 15206 90046 15258
rect 90098 15206 90110 15258
rect 90162 15206 90174 15258
rect 90226 15206 90896 15258
rect 84180 15184 90896 15206
rect 1104 14714 5152 14736
rect 1104 14662 3982 14714
rect 4034 14662 4046 14714
rect 4098 14662 4110 14714
rect 4162 14662 4174 14714
rect 4226 14662 5152 14714
rect 1104 14640 5152 14662
rect 84180 14714 90896 14736
rect 84180 14662 87982 14714
rect 88034 14662 88046 14714
rect 88098 14662 88110 14714
rect 88162 14662 88174 14714
rect 88226 14662 90896 14714
rect 84180 14640 90896 14662
rect 84654 14600 84660 14612
rect 84615 14572 84660 14600
rect 84654 14560 84660 14572
rect 84712 14560 84718 14612
rect 1104 14170 5152 14192
rect 1104 14118 1982 14170
rect 2034 14118 2046 14170
rect 2098 14118 2110 14170
rect 2162 14118 2174 14170
rect 2226 14118 5152 14170
rect 1104 14096 5152 14118
rect 84180 14170 90896 14192
rect 84180 14118 85982 14170
rect 86034 14118 86046 14170
rect 86098 14118 86110 14170
rect 86162 14118 86174 14170
rect 86226 14118 89982 14170
rect 90034 14118 90046 14170
rect 90098 14118 90110 14170
rect 90162 14118 90174 14170
rect 90226 14118 90896 14170
rect 84180 14096 90896 14118
rect 85298 13920 85304 13932
rect 85259 13892 85304 13920
rect 85298 13880 85304 13892
rect 85356 13880 85362 13932
rect 84654 13852 84660 13864
rect 84615 13824 84660 13852
rect 84654 13812 84660 13824
rect 84712 13812 84718 13864
rect 1104 13626 5152 13648
rect 1104 13574 3982 13626
rect 4034 13574 4046 13626
rect 4098 13574 4110 13626
rect 4162 13574 4174 13626
rect 4226 13574 5152 13626
rect 1104 13552 5152 13574
rect 84180 13626 90896 13648
rect 84180 13574 87982 13626
rect 88034 13574 88046 13626
rect 88098 13574 88110 13626
rect 88162 13574 88174 13626
rect 88226 13574 90896 13626
rect 84180 13552 90896 13574
rect 1104 13082 5152 13104
rect 1104 13030 1982 13082
rect 2034 13030 2046 13082
rect 2098 13030 2110 13082
rect 2162 13030 2174 13082
rect 2226 13030 5152 13082
rect 1104 13008 5152 13030
rect 84180 13082 90896 13104
rect 84180 13030 85982 13082
rect 86034 13030 86046 13082
rect 86098 13030 86110 13082
rect 86162 13030 86174 13082
rect 86226 13030 89982 13082
rect 90034 13030 90046 13082
rect 90098 13030 90110 13082
rect 90162 13030 90174 13082
rect 90226 13030 90896 13082
rect 84180 13008 90896 13030
rect 85298 12588 85304 12640
rect 85356 12628 85362 12640
rect 86954 12628 86960 12640
rect 85356 12600 86960 12628
rect 85356 12588 85362 12600
rect 86954 12588 86960 12600
rect 87012 12588 87018 12640
rect 1104 12538 5152 12560
rect 1104 12486 3982 12538
rect 4034 12486 4046 12538
rect 4098 12486 4110 12538
rect 4162 12486 4174 12538
rect 4226 12486 5152 12538
rect 1104 12464 5152 12486
rect 84180 12538 90896 12560
rect 84180 12486 87982 12538
rect 88034 12486 88046 12538
rect 88098 12486 88110 12538
rect 88162 12486 88174 12538
rect 88226 12486 90896 12538
rect 84180 12464 90896 12486
rect 1104 11994 5152 12016
rect 1104 11942 1982 11994
rect 2034 11942 2046 11994
rect 2098 11942 2110 11994
rect 2162 11942 2174 11994
rect 2226 11942 5152 11994
rect 1104 11920 5152 11942
rect 84180 11994 90896 12016
rect 84180 11942 85982 11994
rect 86034 11942 86046 11994
rect 86098 11942 86110 11994
rect 86162 11942 86174 11994
rect 86226 11942 89982 11994
rect 90034 11942 90046 11994
rect 90098 11942 90110 11994
rect 90162 11942 90174 11994
rect 90226 11942 90896 11994
rect 84180 11920 90896 11942
rect 1104 11450 5152 11472
rect 1104 11398 3982 11450
rect 4034 11398 4046 11450
rect 4098 11398 4110 11450
rect 4162 11398 4174 11450
rect 4226 11398 5152 11450
rect 1104 11376 5152 11398
rect 84180 11450 90896 11472
rect 84180 11398 87982 11450
rect 88034 11398 88046 11450
rect 88098 11398 88110 11450
rect 88162 11398 88174 11450
rect 88226 11398 90896 11450
rect 84180 11376 90896 11398
rect 82906 11024 82912 11076
rect 82964 11064 82970 11076
rect 86954 11064 86960 11076
rect 82964 11036 86960 11064
rect 82964 11024 82970 11036
rect 86954 11024 86960 11036
rect 87012 11024 87018 11076
rect 1104 10906 5152 10928
rect 1104 10854 1982 10906
rect 2034 10854 2046 10906
rect 2098 10854 2110 10906
rect 2162 10854 2174 10906
rect 2226 10854 5152 10906
rect 1104 10832 5152 10854
rect 84180 10906 90896 10928
rect 84180 10854 85982 10906
rect 86034 10854 86046 10906
rect 86098 10854 86110 10906
rect 86162 10854 86174 10906
rect 86226 10854 89982 10906
rect 90034 10854 90046 10906
rect 90098 10854 90110 10906
rect 90162 10854 90174 10906
rect 90226 10854 90896 10906
rect 84180 10832 90896 10854
rect 1104 10362 5152 10384
rect 1104 10310 3982 10362
rect 4034 10310 4046 10362
rect 4098 10310 4110 10362
rect 4162 10310 4174 10362
rect 4226 10310 5152 10362
rect 1104 10288 5152 10310
rect 84180 10362 90896 10384
rect 84180 10310 87982 10362
rect 88034 10310 88046 10362
rect 88098 10310 88110 10362
rect 88162 10310 88174 10362
rect 88226 10310 90896 10362
rect 84180 10288 90896 10310
rect 4430 10112 4436 10124
rect 4391 10084 4436 10112
rect 4430 10072 4436 10084
rect 4488 10072 4494 10124
rect 1104 9818 5152 9840
rect 1104 9766 1982 9818
rect 2034 9766 2046 9818
rect 2098 9766 2110 9818
rect 2162 9766 2174 9818
rect 2226 9766 5152 9818
rect 1104 9744 5152 9766
rect 84180 9818 90896 9840
rect 84180 9766 85982 9818
rect 86034 9766 86046 9818
rect 86098 9766 86110 9818
rect 86162 9766 86174 9818
rect 86226 9766 89982 9818
rect 90034 9766 90046 9818
rect 90098 9766 90110 9818
rect 90162 9766 90174 9818
rect 90226 9766 90896 9818
rect 84180 9744 90896 9766
rect 1104 9274 5152 9296
rect 1104 9222 3982 9274
rect 4034 9222 4046 9274
rect 4098 9222 4110 9274
rect 4162 9222 4174 9274
rect 4226 9222 5152 9274
rect 1104 9200 5152 9222
rect 84180 9274 90896 9296
rect 84180 9222 87982 9274
rect 88034 9222 88046 9274
rect 88098 9222 88110 9274
rect 88162 9222 88174 9274
rect 88226 9222 90896 9274
rect 84180 9200 90896 9222
rect 1104 8730 5152 8752
rect 1104 8678 1982 8730
rect 2034 8678 2046 8730
rect 2098 8678 2110 8730
rect 2162 8678 2174 8730
rect 2226 8678 5152 8730
rect 1104 8656 5152 8678
rect 84180 8730 90896 8752
rect 84180 8678 85982 8730
rect 86034 8678 86046 8730
rect 86098 8678 86110 8730
rect 86162 8678 86174 8730
rect 86226 8678 89982 8730
rect 90034 8678 90046 8730
rect 90098 8678 90110 8730
rect 90162 8678 90174 8730
rect 90226 8678 90896 8730
rect 84180 8656 90896 8678
rect 83090 8304 83096 8356
rect 83148 8344 83154 8356
rect 86954 8344 86960 8356
rect 83148 8316 86960 8344
rect 83148 8304 83154 8316
rect 86954 8304 86960 8316
rect 87012 8304 87018 8356
rect 87046 8236 87052 8288
rect 87104 8276 87110 8288
rect 87598 8276 87604 8288
rect 87104 8248 87604 8276
rect 87104 8236 87110 8248
rect 87598 8236 87604 8248
rect 87656 8236 87662 8288
rect 1104 8186 5152 8208
rect 1104 8134 3982 8186
rect 4034 8134 4046 8186
rect 4098 8134 4110 8186
rect 4162 8134 4174 8186
rect 4226 8134 5152 8186
rect 1104 8112 5152 8134
rect 84180 8186 90896 8208
rect 84180 8134 87982 8186
rect 88034 8134 88046 8186
rect 88098 8134 88110 8186
rect 88162 8134 88174 8186
rect 88226 8134 90896 8186
rect 84180 8112 90896 8134
rect 87782 8032 87788 8084
rect 87840 8072 87846 8084
rect 87840 8044 88012 8072
rect 87840 8032 87846 8044
rect 87984 8016 88012 8044
rect 87966 7964 87972 8016
rect 88024 7964 88030 8016
rect 5350 7760 5356 7812
rect 5408 7760 5414 7812
rect 1104 7642 5152 7664
rect 1104 7590 1982 7642
rect 2034 7590 2046 7642
rect 2098 7590 2110 7642
rect 2162 7590 2174 7642
rect 2226 7590 5152 7642
rect 5368 7608 5396 7760
rect 84180 7642 90896 7664
rect 1104 7568 5152 7590
rect 5350 7556 5356 7608
rect 5408 7556 5414 7608
rect 84180 7590 85982 7642
rect 86034 7590 86046 7642
rect 86098 7590 86110 7642
rect 86162 7590 86174 7642
rect 86226 7590 89982 7642
rect 90034 7590 90046 7642
rect 90098 7590 90110 7642
rect 90162 7590 90174 7642
rect 90226 7590 90896 7642
rect 84180 7568 90896 7590
rect 86954 7488 86960 7540
rect 87012 7528 87018 7540
rect 87230 7528 87236 7540
rect 87012 7500 87236 7528
rect 87012 7488 87018 7500
rect 87230 7488 87236 7500
rect 87288 7488 87294 7540
rect 87322 7488 87328 7540
rect 87380 7528 87386 7540
rect 87782 7528 87788 7540
rect 87380 7500 87788 7528
rect 87380 7488 87386 7500
rect 87782 7488 87788 7500
rect 87840 7488 87846 7540
rect 87230 7352 87236 7404
rect 87288 7392 87294 7404
rect 87690 7392 87696 7404
rect 87288 7364 87696 7392
rect 87288 7352 87294 7364
rect 87690 7352 87696 7364
rect 87748 7352 87754 7404
rect 87690 7216 87696 7268
rect 87748 7256 87754 7268
rect 87966 7256 87972 7268
rect 87748 7228 87972 7256
rect 87748 7216 87754 7228
rect 87966 7216 87972 7228
rect 88024 7216 88030 7268
rect 1104 7098 5152 7120
rect 1104 7046 3982 7098
rect 4034 7046 4046 7098
rect 4098 7046 4110 7098
rect 4162 7046 4174 7098
rect 4226 7046 5152 7098
rect 1104 7024 5152 7046
rect 84180 7098 90896 7120
rect 84180 7046 87982 7098
rect 88034 7046 88046 7098
rect 88098 7046 88110 7098
rect 88162 7046 88174 7098
rect 88226 7046 90896 7098
rect 84180 7024 90896 7046
rect 1104 6554 5152 6576
rect 1104 6502 1982 6554
rect 2034 6502 2046 6554
rect 2098 6502 2110 6554
rect 2162 6502 2174 6554
rect 2226 6502 5152 6554
rect 1104 6480 5152 6502
rect 84180 6554 90896 6576
rect 84180 6502 85982 6554
rect 86034 6502 86046 6554
rect 86098 6502 86110 6554
rect 86162 6502 86174 6554
rect 86226 6502 89982 6554
rect 90034 6502 90046 6554
rect 90098 6502 90110 6554
rect 90162 6502 90174 6554
rect 90226 6502 90896 6554
rect 84180 6480 90896 6502
rect 1104 6010 5152 6032
rect 1104 5958 3982 6010
rect 4034 5958 4046 6010
rect 4098 5958 4110 6010
rect 4162 5958 4174 6010
rect 4226 5958 5152 6010
rect 1104 5936 5152 5958
rect 84180 6010 90896 6032
rect 84180 5958 87982 6010
rect 88034 5958 88046 6010
rect 88098 5958 88110 6010
rect 88162 5958 88174 6010
rect 88226 5958 90896 6010
rect 84180 5936 90896 5958
rect 1104 5466 5152 5488
rect 1104 5414 1982 5466
rect 2034 5414 2046 5466
rect 2098 5414 2110 5466
rect 2162 5414 2174 5466
rect 2226 5414 5152 5466
rect 1104 5392 5152 5414
rect 84180 5466 90896 5488
rect 84180 5414 85982 5466
rect 86034 5414 86046 5466
rect 86098 5414 86110 5466
rect 86162 5414 86174 5466
rect 86226 5414 89982 5466
rect 90034 5414 90046 5466
rect 90098 5414 90110 5466
rect 90162 5414 90174 5466
rect 90226 5414 90896 5466
rect 84180 5392 90896 5414
rect 85850 5312 85856 5364
rect 85908 5352 85914 5364
rect 87046 5352 87052 5364
rect 85908 5324 87052 5352
rect 85908 5312 85914 5324
rect 87046 5312 87052 5324
rect 87104 5312 87110 5364
rect 4801 5015 4859 5021
rect 4801 4981 4813 5015
rect 4847 5012 4859 5015
rect 5442 5012 5448 5024
rect 4847 4984 5448 5012
rect 4847 4981 4859 4984
rect 4801 4975 4859 4981
rect 5442 4972 5448 4984
rect 5500 4972 5506 5024
rect 1104 4922 5152 4944
rect 1104 4870 3982 4922
rect 4034 4870 4046 4922
rect 4098 4870 4110 4922
rect 4162 4870 4174 4922
rect 4226 4870 5152 4922
rect 1104 4848 5152 4870
rect 84180 4922 90896 4944
rect 84180 4870 87982 4922
rect 88034 4870 88046 4922
rect 88098 4870 88110 4922
rect 88162 4870 88174 4922
rect 88226 4870 90896 4922
rect 84180 4848 90896 4870
rect 4801 4811 4859 4817
rect 4801 4777 4813 4811
rect 4847 4808 4859 4811
rect 5074 4808 5080 4820
rect 4847 4780 5080 4808
rect 4847 4777 4859 4780
rect 4801 4771 4859 4777
rect 5074 4768 5080 4780
rect 5132 4808 5138 4820
rect 5718 4808 5724 4820
rect 5132 4780 5724 4808
rect 5132 4768 5138 4780
rect 5718 4768 5724 4780
rect 5776 4768 5782 4820
rect 4433 4743 4491 4749
rect 4433 4709 4445 4743
rect 4479 4740 4491 4743
rect 5166 4740 5172 4752
rect 4479 4712 5172 4740
rect 4479 4709 4491 4712
rect 4433 4703 4491 4709
rect 5166 4700 5172 4712
rect 5224 4740 5230 4752
rect 5994 4740 6000 4752
rect 5224 4712 6000 4740
rect 5224 4700 5230 4712
rect 5994 4700 6000 4712
rect 6052 4700 6058 4752
rect 87690 4700 87696 4752
rect 87748 4740 87754 4752
rect 87966 4740 87972 4752
rect 87748 4712 87972 4740
rect 87748 4700 87754 4712
rect 87966 4700 87972 4712
rect 88024 4700 88030 4752
rect 1104 4378 5152 4400
rect 1104 4326 1982 4378
rect 2034 4326 2046 4378
rect 2098 4326 2110 4378
rect 2162 4326 2174 4378
rect 2226 4326 5152 4378
rect 83182 4360 83188 4412
rect 83240 4400 83246 4412
rect 83458 4400 83464 4412
rect 83240 4372 83464 4400
rect 83240 4360 83246 4372
rect 83458 4360 83464 4372
rect 83516 4360 83522 4412
rect 84180 4378 90896 4400
rect 83642 4332 83648 4344
rect 1104 4304 5152 4326
rect 83603 4304 83648 4332
rect 83642 4292 83648 4304
rect 83700 4292 83706 4344
rect 84180 4326 85982 4378
rect 86034 4326 86046 4378
rect 86098 4326 86110 4378
rect 86162 4326 86174 4378
rect 86226 4326 89982 4378
rect 90034 4326 90046 4378
rect 90098 4326 90110 4378
rect 90162 4326 90174 4378
rect 90226 4326 90896 4378
rect 84180 4304 90896 4326
rect 83642 4156 83648 4208
rect 83700 4196 83706 4208
rect 87046 4196 87052 4208
rect 83700 4168 87052 4196
rect 83700 4156 83706 4168
rect 87046 4156 87052 4168
rect 87104 4156 87110 4208
rect 3878 4088 3884 4140
rect 3936 4128 3942 4140
rect 3973 4131 4031 4137
rect 3973 4128 3985 4131
rect 3936 4100 3985 4128
rect 3936 4088 3942 4100
rect 3973 4097 3985 4100
rect 4019 4097 4031 4131
rect 3973 4091 4031 4097
rect 4522 4088 4528 4140
rect 4580 4128 4586 4140
rect 5902 4128 5908 4140
rect 4580 4100 5908 4128
rect 4580 4088 4586 4100
rect 5902 4088 5908 4100
rect 5960 4088 5966 4140
rect 82814 4088 82820 4140
rect 82872 4128 82878 4140
rect 84657 4131 84715 4137
rect 84657 4128 84669 4131
rect 82872 4100 84669 4128
rect 82872 4088 82878 4100
rect 84657 4097 84669 4100
rect 84703 4097 84715 4131
rect 84657 4091 84715 4097
rect 4433 4063 4491 4069
rect 4433 4029 4445 4063
rect 4479 4060 4491 4063
rect 5718 4060 5724 4072
rect 4479 4032 5724 4060
rect 4479 4029 4491 4032
rect 4433 4023 4491 4029
rect 5718 4020 5724 4032
rect 5776 4060 5782 4072
rect 6362 4060 6368 4072
rect 5776 4032 6368 4060
rect 5776 4020 5782 4032
rect 6362 4020 6368 4032
rect 6420 4020 6426 4072
rect 82722 4020 82728 4072
rect 82780 4060 82786 4072
rect 87690 4060 87696 4072
rect 82780 4032 87696 4060
rect 82780 4020 82786 4032
rect 87690 4020 87696 4032
rect 87748 4020 87754 4072
rect 3329 3995 3387 4001
rect 3329 3961 3341 3995
rect 3375 3992 3387 3995
rect 3375 3964 6960 3992
rect 3375 3961 3387 3964
rect 3329 3955 3387 3961
rect 3697 3927 3755 3933
rect 3697 3893 3709 3927
rect 3743 3924 3755 3927
rect 3786 3924 3792 3936
rect 3743 3896 3792 3924
rect 3743 3893 3755 3896
rect 3697 3887 3755 3893
rect 3786 3884 3792 3896
rect 3844 3884 3850 3936
rect 4798 3924 4804 3936
rect 4759 3896 4804 3924
rect 4798 3884 4804 3896
rect 4856 3884 4862 3936
rect 1104 3834 5152 3856
rect 1104 3782 3982 3834
rect 4034 3782 4046 3834
rect 4098 3782 4110 3834
rect 4162 3782 4174 3834
rect 4226 3782 5152 3834
rect 1104 3760 5152 3782
rect 3326 3720 3332 3732
rect 3287 3692 3332 3720
rect 3326 3680 3332 3692
rect 3384 3680 3390 3732
rect 4798 3720 4804 3732
rect 4711 3692 4804 3720
rect 4798 3680 4804 3692
rect 4856 3720 4862 3732
rect 5626 3720 5632 3732
rect 4856 3692 5632 3720
rect 4856 3680 4862 3692
rect 5626 3680 5632 3692
rect 5684 3680 5690 3732
rect 3344 3584 3372 3680
rect 4430 3652 4436 3664
rect 4343 3624 4436 3652
rect 4430 3612 4436 3624
rect 4488 3652 4494 3664
rect 5810 3652 5816 3664
rect 4488 3624 5816 3652
rect 4488 3612 4494 3624
rect 5810 3612 5816 3624
rect 5868 3612 5874 3664
rect 6825 3587 6883 3593
rect 6825 3584 6837 3587
rect 3344 3556 6837 3584
rect 6825 3553 6837 3556
rect 6871 3553 6883 3587
rect 6825 3547 6883 3553
rect 3697 3519 3755 3525
rect 3697 3485 3709 3519
rect 3743 3516 3755 3519
rect 5626 3516 5632 3528
rect 3743 3488 5632 3516
rect 3743 3485 3755 3488
rect 3697 3479 3755 3485
rect 5626 3476 5632 3488
rect 5684 3476 5690 3528
rect 2593 3451 2651 3457
rect 2593 3417 2605 3451
rect 2639 3448 2651 3451
rect 6733 3451 6791 3457
rect 6733 3448 6745 3451
rect 2639 3420 6745 3448
rect 2639 3417 2651 3420
rect 2593 3411 2651 3417
rect 6733 3417 6745 3420
rect 6779 3417 6791 3451
rect 6733 3411 6791 3417
rect 2961 3383 3019 3389
rect 2961 3349 2973 3383
rect 3007 3380 3019 3383
rect 3602 3380 3608 3392
rect 3007 3352 3608 3380
rect 3007 3349 3019 3352
rect 2961 3343 3019 3349
rect 3602 3340 3608 3352
rect 3660 3340 3666 3392
rect 3786 3340 3792 3392
rect 3844 3380 3850 3392
rect 3844 3352 5212 3380
rect 3844 3340 3850 3352
rect 1104 3290 5152 3312
rect 1104 3238 1982 3290
rect 2034 3238 2046 3290
rect 2098 3238 2110 3290
rect 2162 3238 2174 3290
rect 2226 3238 5152 3290
rect 1104 3216 5152 3238
rect 5184 3244 5212 3352
rect 6932 3312 6960 3964
rect 82630 3952 82636 4004
rect 82688 3992 82694 4004
rect 87966 3992 87972 4004
rect 82688 3964 87972 3992
rect 82688 3952 82694 3964
rect 87966 3952 87972 3964
rect 88024 3952 88030 4004
rect 84180 3834 90896 3856
rect 84180 3782 87982 3834
rect 88034 3782 88046 3834
rect 88098 3782 88110 3834
rect 88162 3782 88174 3834
rect 88226 3782 90896 3834
rect 84180 3760 90896 3782
rect 83458 3680 83464 3732
rect 83516 3720 83522 3732
rect 83645 3723 83703 3729
rect 83645 3720 83657 3723
rect 83516 3692 83657 3720
rect 83516 3680 83522 3692
rect 83645 3689 83657 3692
rect 83691 3720 83703 3723
rect 84657 3723 84715 3729
rect 84657 3720 84669 3723
rect 83691 3692 84669 3720
rect 83691 3689 83703 3692
rect 83645 3683 83703 3689
rect 84657 3689 84669 3692
rect 84703 3689 84715 3723
rect 84657 3683 84715 3689
rect 84930 3680 84936 3732
rect 84988 3720 84994 3732
rect 85025 3723 85083 3729
rect 85025 3720 85037 3723
rect 84988 3692 85037 3720
rect 84988 3680 84994 3692
rect 85025 3689 85037 3692
rect 85071 3689 85083 3723
rect 85390 3720 85396 3732
rect 85351 3692 85396 3720
rect 85025 3683 85083 3689
rect 85390 3680 85396 3692
rect 85448 3680 85454 3732
rect 82541 3655 82599 3661
rect 82541 3621 82553 3655
rect 82587 3652 82599 3655
rect 85408 3652 85436 3680
rect 82587 3624 85436 3652
rect 82587 3621 82599 3624
rect 82541 3615 82599 3621
rect 82449 3587 82507 3593
rect 82449 3553 82461 3587
rect 82495 3584 82507 3587
rect 85850 3584 85856 3596
rect 82495 3556 85856 3584
rect 82495 3553 82507 3556
rect 82449 3547 82507 3553
rect 85850 3544 85856 3556
rect 85908 3544 85914 3596
rect 83093 3519 83151 3525
rect 83093 3485 83105 3519
rect 83139 3516 83151 3519
rect 85758 3516 85764 3528
rect 83139 3488 85764 3516
rect 83139 3485 83151 3488
rect 83093 3479 83151 3485
rect 85758 3476 85764 3488
rect 85816 3476 85822 3528
rect 82538 3408 82544 3460
rect 82596 3448 82602 3460
rect 87046 3448 87052 3460
rect 82596 3420 87052 3448
rect 82596 3408 82602 3420
rect 87046 3408 87052 3420
rect 87104 3408 87110 3460
rect 83642 3312 83648 3324
rect 6932 3284 83648 3312
rect 15304 3256 15332 3284
rect 83642 3272 83648 3284
rect 83700 3272 83706 3324
rect 84180 3290 90896 3312
rect 6730 3244 6736 3256
rect 5184 3216 6736 3244
rect 6730 3204 6736 3216
rect 6788 3244 6794 3256
rect 15105 3247 15163 3253
rect 15105 3244 15117 3247
rect 6788 3216 15117 3244
rect 6788 3204 6794 3216
rect 15105 3213 15117 3216
rect 15151 3213 15163 3247
rect 15105 3207 15163 3213
rect 15286 3204 15292 3256
rect 15344 3204 15350 3256
rect 15381 3247 15439 3253
rect 15381 3213 15393 3247
rect 15427 3244 15439 3247
rect 25038 3244 25044 3256
rect 15427 3216 25044 3244
rect 15427 3213 15439 3216
rect 15381 3207 15439 3213
rect 25038 3204 25044 3216
rect 25096 3204 25102 3256
rect 52546 3204 52552 3256
rect 52604 3244 52610 3256
rect 82814 3244 82820 3256
rect 52604 3216 82820 3244
rect 52604 3204 52610 3216
rect 82814 3204 82820 3216
rect 82872 3204 82878 3256
rect 83550 3244 83556 3256
rect 83511 3216 83556 3244
rect 83550 3204 83556 3216
rect 83608 3204 83614 3256
rect 84180 3238 85982 3290
rect 86034 3238 86046 3290
rect 86098 3238 86110 3290
rect 86162 3238 86174 3290
rect 86226 3238 89982 3290
rect 90034 3238 90046 3290
rect 90098 3238 90110 3290
rect 90162 3238 90174 3290
rect 90226 3238 90896 3290
rect 84180 3216 90896 3238
rect 2225 3179 2283 3185
rect 2225 3145 2237 3179
rect 2271 3176 2283 3179
rect 3510 3176 3516 3188
rect 2271 3148 3516 3176
rect 2271 3145 2283 3148
rect 2225 3139 2283 3145
rect 3510 3136 3516 3148
rect 3568 3136 3574 3188
rect 3694 3176 3700 3188
rect 3655 3148 3700 3176
rect 3694 3136 3700 3148
rect 3752 3136 3758 3188
rect 4433 3179 4491 3185
rect 4433 3145 4445 3179
rect 4479 3176 4491 3179
rect 5534 3176 5540 3188
rect 4479 3148 5540 3176
rect 4479 3145 4491 3148
rect 4433 3139 4491 3145
rect 5534 3136 5540 3148
rect 5592 3136 5598 3188
rect 6917 3179 6975 3185
rect 6917 3145 6929 3179
rect 6963 3176 6975 3179
rect 15013 3179 15071 3185
rect 15013 3176 15025 3179
rect 6963 3148 15025 3176
rect 6963 3145 6975 3148
rect 6917 3139 6975 3145
rect 15013 3145 15025 3148
rect 15059 3145 15071 3179
rect 15013 3139 15071 3145
rect 15473 3179 15531 3185
rect 15473 3145 15485 3179
rect 15519 3176 15531 3179
rect 22094 3176 22100 3188
rect 15519 3148 22100 3176
rect 15519 3145 15531 3148
rect 15473 3139 15531 3145
rect 22094 3136 22100 3148
rect 22152 3136 22158 3188
rect 49970 3136 49976 3188
rect 50028 3176 50034 3188
rect 84930 3176 84936 3188
rect 50028 3148 84936 3176
rect 50028 3136 50034 3148
rect 84930 3136 84936 3148
rect 84988 3136 84994 3188
rect 85758 3176 85764 3188
rect 85719 3148 85764 3176
rect 85758 3136 85764 3148
rect 85816 3136 85822 3188
rect 2498 3108 2504 3120
rect 2459 3080 2504 3108
rect 2498 3068 2504 3080
rect 2556 3068 2562 3120
rect 4065 3111 4123 3117
rect 4065 3077 4077 3111
rect 4111 3108 4123 3111
rect 4522 3108 4528 3120
rect 4111 3080 4528 3108
rect 4111 3077 4123 3080
rect 4065 3071 4123 3077
rect 4522 3068 4528 3080
rect 4580 3068 4586 3120
rect 6733 3111 6791 3117
rect 6733 3077 6745 3111
rect 6779 3108 6791 3111
rect 15105 3111 15163 3117
rect 15105 3108 15117 3111
rect 6779 3080 15117 3108
rect 6779 3077 6791 3080
rect 6733 3071 6791 3077
rect 15105 3077 15117 3080
rect 15151 3077 15163 3111
rect 15105 3071 15163 3077
rect 15381 3111 15439 3117
rect 15381 3077 15393 3111
rect 15427 3108 15439 3111
rect 16298 3108 16304 3120
rect 15427 3080 16304 3108
rect 15427 3077 15439 3080
rect 15381 3071 15439 3077
rect 16298 3068 16304 3080
rect 16356 3108 16362 3120
rect 87322 3108 87328 3120
rect 16356 3080 87328 3108
rect 16356 3068 16362 3080
rect 87322 3068 87328 3080
rect 87380 3068 87386 3120
rect 2516 3040 2544 3068
rect 2516 3012 2774 3040
rect 2746 2904 2774 3012
rect 5902 3000 5908 3052
rect 5960 3040 5966 3052
rect 13906 3040 13912 3052
rect 5960 3012 13912 3040
rect 5960 3000 5966 3012
rect 13906 3000 13912 3012
rect 13964 3000 13970 3052
rect 53466 3000 53472 3052
rect 53524 3040 53530 3052
rect 83093 3043 83151 3049
rect 83093 3040 83105 3043
rect 53524 3012 83105 3040
rect 53524 3000 53530 3012
rect 83093 3009 83105 3012
rect 83139 3009 83151 3043
rect 83093 3003 83151 3009
rect 83182 3000 83188 3052
rect 83240 3040 83246 3052
rect 84657 3043 84715 3049
rect 84657 3040 84669 3043
rect 83240 3012 84669 3040
rect 83240 3000 83246 3012
rect 84657 3009 84669 3012
rect 84703 3009 84715 3043
rect 84657 3003 84715 3009
rect 2961 2975 3019 2981
rect 2961 2941 2973 2975
rect 3007 2972 3019 2975
rect 3786 2972 3792 2984
rect 3007 2944 3792 2972
rect 3007 2941 3019 2944
rect 2961 2935 3019 2941
rect 3786 2932 3792 2944
rect 3844 2932 3850 2984
rect 3878 2932 3884 2984
rect 3936 2972 3942 2984
rect 20714 2972 20720 2984
rect 3936 2944 20720 2972
rect 3936 2932 3942 2944
rect 20714 2932 20720 2944
rect 20772 2932 20778 2984
rect 87598 2972 87604 2984
rect 26206 2944 87604 2972
rect 24118 2904 24124 2916
rect 2746 2876 24124 2904
rect 24118 2864 24124 2876
rect 24176 2864 24182 2916
rect 3329 2839 3387 2845
rect 3329 2805 3341 2839
rect 3375 2836 3387 2839
rect 4338 2836 4344 2848
rect 3375 2808 4344 2836
rect 3375 2805 3387 2808
rect 3329 2799 3387 2805
rect 4338 2796 4344 2808
rect 4396 2796 4402 2848
rect 4614 2796 4620 2848
rect 4672 2836 4678 2848
rect 4709 2839 4767 2845
rect 4709 2836 4721 2839
rect 4672 2808 4721 2836
rect 4672 2796 4678 2808
rect 4709 2805 4721 2808
rect 4755 2805 4767 2839
rect 4709 2799 4767 2805
rect 4890 2796 4896 2848
rect 4948 2836 4954 2848
rect 6914 2836 6920 2848
rect 4948 2808 6920 2836
rect 4948 2796 4954 2808
rect 6914 2796 6920 2808
rect 6972 2836 6978 2848
rect 8110 2836 8116 2848
rect 6972 2808 8116 2836
rect 6972 2796 6978 2808
rect 8110 2796 8116 2808
rect 8168 2796 8174 2848
rect 13906 2796 13912 2848
rect 13964 2836 13970 2848
rect 26206 2836 26234 2944
rect 87598 2932 87604 2944
rect 87656 2932 87662 2984
rect 47762 2864 47768 2916
rect 47820 2904 47826 2916
rect 82446 2904 82452 2916
rect 47820 2876 64874 2904
rect 47820 2864 47826 2876
rect 13964 2808 26234 2836
rect 64846 2836 64874 2876
rect 80026 2876 82452 2904
rect 80026 2836 80054 2876
rect 82446 2864 82452 2876
rect 82504 2864 82510 2916
rect 82998 2864 83004 2916
rect 83056 2904 83062 2916
rect 85025 2907 85083 2913
rect 85025 2904 85037 2907
rect 83056 2876 85037 2904
rect 83056 2864 83062 2876
rect 85025 2873 85037 2876
rect 85071 2873 85083 2907
rect 85025 2867 85083 2873
rect 87322 2864 87328 2916
rect 87380 2904 87386 2916
rect 87506 2904 87512 2916
rect 87380 2876 87512 2904
rect 87380 2864 87386 2876
rect 87506 2864 87512 2876
rect 87564 2864 87570 2916
rect 64846 2808 80054 2836
rect 13964 2796 13970 2808
rect 81434 2796 81440 2848
rect 81492 2836 81498 2848
rect 82357 2839 82415 2845
rect 82357 2836 82369 2839
rect 81492 2808 82369 2836
rect 81492 2796 81498 2808
rect 82357 2805 82369 2808
rect 82403 2805 82415 2839
rect 82464 2836 82492 2864
rect 85393 2839 85451 2845
rect 85393 2836 85405 2839
rect 82464 2808 85405 2836
rect 82357 2799 82415 2805
rect 85393 2805 85405 2808
rect 85439 2805 85451 2839
rect 85393 2799 85451 2805
rect 82446 2768 82452 2780
rect 1104 2746 5152 2768
rect 1104 2694 3982 2746
rect 4034 2694 4046 2746
rect 4098 2694 4110 2746
rect 4162 2694 4174 2746
rect 4226 2694 5152 2746
rect 1104 2672 5152 2694
rect 12406 2740 82452 2768
rect 3697 2635 3755 2641
rect 3697 2601 3709 2635
rect 3743 2632 3755 2635
rect 3878 2632 3884 2644
rect 3743 2604 3884 2632
rect 3743 2601 3755 2604
rect 3697 2595 3755 2601
rect 3878 2592 3884 2604
rect 3936 2592 3942 2644
rect 4706 2592 4712 2644
rect 4764 2632 4770 2644
rect 12406 2632 12434 2740
rect 82446 2728 82452 2740
rect 82504 2728 82510 2780
rect 83550 2768 83556 2780
rect 83511 2740 83556 2768
rect 83550 2728 83556 2740
rect 83608 2728 83614 2780
rect 84180 2746 90896 2768
rect 81342 2660 81348 2712
rect 81400 2700 81406 2712
rect 82541 2703 82599 2709
rect 82541 2700 82553 2703
rect 81400 2672 82553 2700
rect 81400 2660 81406 2672
rect 82541 2669 82553 2672
rect 82587 2669 82599 2703
rect 84180 2694 87982 2746
rect 88034 2694 88046 2746
rect 88098 2694 88110 2746
rect 88162 2694 88174 2746
rect 88226 2694 90896 2746
rect 84180 2672 90896 2694
rect 82541 2663 82599 2669
rect 4764 2604 12434 2632
rect 4764 2592 4770 2604
rect 53834 2592 53840 2644
rect 53892 2632 53898 2644
rect 87322 2632 87328 2644
rect 53892 2604 87328 2632
rect 53892 2592 53898 2604
rect 87322 2592 87328 2604
rect 87380 2592 87386 2644
rect 3234 2524 3240 2576
rect 3292 2564 3298 2576
rect 3329 2567 3387 2573
rect 3329 2564 3341 2567
rect 3292 2536 3341 2564
rect 3292 2524 3298 2536
rect 3329 2533 3341 2536
rect 3375 2564 3387 2567
rect 3375 2536 12434 2564
rect 3375 2533 3387 2536
rect 3329 2527 3387 2533
rect 4433 2499 4491 2505
rect 4433 2465 4445 2499
rect 4479 2496 4491 2499
rect 6178 2496 6184 2508
rect 4479 2468 6184 2496
rect 4479 2465 4491 2468
rect 4433 2459 4491 2465
rect 6178 2456 6184 2468
rect 6236 2456 6242 2508
rect 12406 2496 12434 2536
rect 50338 2524 50344 2576
rect 50396 2564 50402 2576
rect 83093 2567 83151 2573
rect 83093 2564 83105 2567
rect 50396 2536 83105 2564
rect 50396 2524 50402 2536
rect 83093 2533 83105 2536
rect 83139 2533 83151 2567
rect 83093 2527 83151 2533
rect 83185 2567 83243 2573
rect 83185 2533 83197 2567
rect 83231 2564 83243 2567
rect 87138 2564 87144 2576
rect 83231 2536 87144 2564
rect 83231 2533 83243 2536
rect 83185 2527 83243 2533
rect 87138 2524 87144 2536
rect 87196 2524 87202 2576
rect 22646 2496 22652 2508
rect 12406 2468 22652 2496
rect 22646 2456 22652 2468
rect 22704 2456 22710 2508
rect 45922 2456 45928 2508
rect 45980 2496 45986 2508
rect 87230 2496 87236 2508
rect 45980 2468 87236 2496
rect 45980 2456 45986 2468
rect 87230 2456 87236 2468
rect 87288 2456 87294 2508
rect 2961 2431 3019 2437
rect 2961 2397 2973 2431
rect 3007 2428 3019 2431
rect 4154 2428 4160 2440
rect 3007 2400 4160 2428
rect 3007 2397 3019 2400
rect 2961 2391 3019 2397
rect 4154 2388 4160 2400
rect 4212 2388 4218 2440
rect 4982 2388 4988 2440
rect 5040 2428 5046 2440
rect 5040 2400 12434 2428
rect 5040 2388 5046 2400
rect 2593 2363 2651 2369
rect 2593 2329 2605 2363
rect 2639 2360 2651 2363
rect 9766 2360 9772 2372
rect 2639 2332 9772 2360
rect 2639 2329 2651 2332
rect 2593 2323 2651 2329
rect 9766 2320 9772 2332
rect 9824 2320 9830 2372
rect 12406 2360 12434 2400
rect 41414 2388 41420 2440
rect 41472 2428 41478 2440
rect 83185 2431 83243 2437
rect 83185 2428 83197 2431
rect 41472 2400 83197 2428
rect 41472 2388 41478 2400
rect 83185 2397 83197 2400
rect 83231 2397 83243 2431
rect 86954 2428 86960 2440
rect 83185 2391 83243 2397
rect 83292 2400 86960 2428
rect 83292 2360 83320 2400
rect 86954 2388 86960 2400
rect 87012 2388 87018 2440
rect 85022 2360 85028 2372
rect 12406 2332 83320 2360
rect 83384 2332 85028 2360
rect 4801 2295 4859 2301
rect 4801 2261 4813 2295
rect 4847 2292 4859 2295
rect 6270 2292 6276 2304
rect 4847 2264 6276 2292
rect 4847 2261 4859 2264
rect 4801 2255 4859 2261
rect 6270 2252 6276 2264
rect 6328 2252 6334 2304
rect 51350 2252 51356 2304
rect 51408 2292 51414 2304
rect 83384 2292 83412 2332
rect 85022 2320 85028 2332
rect 85080 2320 85086 2372
rect 51408 2264 83412 2292
rect 51408 2252 51414 2264
rect 83550 2252 83556 2304
rect 83608 2292 83614 2304
rect 84657 2295 84715 2301
rect 84657 2292 84669 2295
rect 83608 2264 84669 2292
rect 83608 2252 83614 2264
rect 84657 2261 84669 2264
rect 84703 2261 84715 2295
rect 84657 2255 84715 2261
rect 1104 2202 5152 2224
rect 1104 2150 1982 2202
rect 2034 2150 2046 2202
rect 2098 2150 2110 2202
rect 2162 2150 2174 2202
rect 2226 2150 5152 2202
rect 37458 2184 37464 2236
rect 37516 2224 37522 2236
rect 83918 2224 83924 2236
rect 37516 2196 83924 2224
rect 37516 2184 37522 2196
rect 83918 2184 83924 2196
rect 83976 2184 83982 2236
rect 84180 2202 90896 2224
rect 1104 2128 5152 2150
rect 6178 2116 6184 2168
rect 6236 2156 6242 2168
rect 36170 2156 36176 2168
rect 6236 2128 36176 2156
rect 6236 2116 6242 2128
rect 36170 2116 36176 2128
rect 36228 2116 36234 2168
rect 36262 2116 36268 2168
rect 36320 2156 36326 2168
rect 84010 2156 84016 2168
rect 36320 2128 84016 2156
rect 36320 2116 36326 2128
rect 84010 2116 84016 2128
rect 84068 2116 84074 2168
rect 84180 2150 85982 2202
rect 86034 2150 86046 2202
rect 86098 2150 86110 2202
rect 86162 2150 86174 2202
rect 86226 2150 89982 2202
rect 90034 2150 90046 2202
rect 90098 2150 90110 2202
rect 90162 2150 90174 2202
rect 90226 2150 90896 2202
rect 84180 2128 90896 2150
rect 33962 2048 33968 2100
rect 34020 2088 34026 2100
rect 84102 2088 84108 2100
rect 34020 2060 84108 2088
rect 34020 2048 34026 2060
rect 84102 2048 84108 2060
rect 84160 2048 84166 2100
rect 6270 1980 6276 2032
rect 6328 2020 6334 2032
rect 32674 2020 32680 2032
rect 6328 1992 32680 2020
rect 6328 1980 6334 1992
rect 32674 1980 32680 1992
rect 32732 1980 32738 2032
rect 32766 1980 32772 2032
rect 32824 2020 32830 2032
rect 83366 2020 83372 2032
rect 32824 1992 83372 2020
rect 32824 1980 32830 1992
rect 83366 1980 83372 1992
rect 83424 1980 83430 2032
rect 4154 1912 4160 1964
rect 4212 1952 4218 1964
rect 5258 1952 5264 1964
rect 4212 1924 5264 1952
rect 4212 1912 4218 1924
rect 5258 1912 5264 1924
rect 5316 1952 5322 1964
rect 29086 1952 29092 1964
rect 5316 1924 29092 1952
rect 5316 1912 5322 1924
rect 29086 1912 29092 1924
rect 29144 1912 29150 1964
rect 30466 1912 30472 1964
rect 30524 1952 30530 1964
rect 83274 1952 83280 1964
rect 30524 1924 83280 1952
rect 30524 1912 30530 1924
rect 83274 1912 83280 1924
rect 83332 1912 83338 1964
rect 31662 1844 31668 1896
rect 31720 1884 31726 1896
rect 84562 1884 84568 1896
rect 31720 1856 84568 1884
rect 31720 1844 31726 1856
rect 84562 1844 84568 1856
rect 84620 1844 84626 1896
rect 25774 1776 25780 1828
rect 25832 1816 25838 1828
rect 84470 1816 84476 1828
rect 25832 1788 84476 1816
rect 25832 1776 25838 1788
rect 84470 1776 84476 1788
rect 84528 1776 84534 1828
rect 28166 1708 28172 1760
rect 28224 1748 28230 1760
rect 83001 1751 83059 1757
rect 83001 1748 83013 1751
rect 28224 1720 83013 1748
rect 28224 1708 28230 1720
rect 83001 1717 83013 1720
rect 83047 1717 83059 1751
rect 83001 1711 83059 1717
rect 83093 1751 83151 1757
rect 83093 1717 83105 1751
rect 83139 1748 83151 1751
rect 87414 1748 87420 1760
rect 83139 1720 87420 1748
rect 83139 1717 83151 1720
rect 83093 1711 83151 1717
rect 87414 1708 87420 1720
rect 87472 1708 87478 1760
rect 26970 1640 26976 1692
rect 27028 1680 27034 1692
rect 87046 1680 87052 1692
rect 27028 1652 87052 1680
rect 27028 1640 27034 1652
rect 87046 1640 87052 1652
rect 87104 1640 87110 1692
rect 21082 1572 21088 1624
rect 21140 1612 21146 1624
rect 83182 1612 83188 1624
rect 21140 1584 83188 1612
rect 21140 1572 21146 1584
rect 83182 1572 83188 1584
rect 83240 1572 83246 1624
rect 83277 1615 83335 1621
rect 83277 1581 83289 1615
rect 83323 1612 83335 1615
rect 87874 1612 87880 1624
rect 83323 1584 87880 1612
rect 83323 1581 83335 1584
rect 83277 1575 83335 1581
rect 87874 1572 87880 1584
rect 87932 1572 87938 1624
rect 22278 1504 22284 1556
rect 22336 1544 22342 1556
rect 85298 1544 85304 1556
rect 22336 1516 85304 1544
rect 22336 1504 22342 1516
rect 85298 1504 85304 1516
rect 85356 1504 85362 1556
rect 19242 1436 19248 1488
rect 19300 1476 19306 1488
rect 83090 1476 83096 1488
rect 19300 1448 83096 1476
rect 19300 1436 19306 1448
rect 83090 1436 83096 1448
rect 83148 1436 83154 1488
rect 88242 1476 88248 1488
rect 83200 1448 88248 1476
rect 5442 1368 5448 1420
rect 5500 1408 5506 1420
rect 17494 1408 17500 1420
rect 5500 1380 17500 1408
rect 5500 1368 5506 1380
rect 17494 1368 17500 1380
rect 17552 1408 17558 1420
rect 17552 1380 82952 1408
rect 17552 1368 17558 1380
rect 4614 1300 4620 1352
rect 4672 1340 4678 1352
rect 6454 1340 6460 1352
rect 4672 1312 6460 1340
rect 4672 1300 4678 1312
rect 6454 1300 6460 1312
rect 6512 1340 6518 1352
rect 12434 1340 12440 1352
rect 6512 1312 12440 1340
rect 6512 1300 6518 1312
rect 12434 1300 12440 1312
rect 12492 1300 12498 1352
rect 35526 1300 35532 1352
rect 35584 1340 35590 1352
rect 45922 1340 45928 1352
rect 35584 1312 45928 1340
rect 35584 1300 35590 1312
rect 45922 1300 45928 1312
rect 45980 1300 45986 1352
rect 48222 1300 48228 1352
rect 48280 1340 48286 1352
rect 53834 1340 53840 1352
rect 48280 1312 53840 1340
rect 48280 1300 48286 1312
rect 53834 1300 53840 1312
rect 53892 1300 53898 1352
rect 82924 1340 82952 1380
rect 83200 1340 83228 1448
rect 88242 1436 88248 1448
rect 88300 1436 88306 1488
rect 82924 1312 83228 1340
rect 4798 1232 4804 1284
rect 4856 1272 4862 1284
rect 28994 1272 29000 1284
rect 4856 1244 29000 1272
rect 4856 1232 4862 1244
rect 28994 1232 29000 1244
rect 29052 1232 29058 1284
rect 44910 1232 44916 1284
rect 44968 1272 44974 1284
rect 50338 1272 50344 1284
rect 44968 1244 50344 1272
rect 44968 1232 44974 1244
rect 50338 1232 50344 1244
rect 50396 1232 50402 1284
rect 30282 1164 30288 1216
rect 30340 1204 30346 1216
rect 86310 1204 86316 1216
rect 30340 1176 86316 1204
rect 30340 1164 30346 1176
rect 86310 1164 86316 1176
rect 86368 1164 86374 1216
rect 39942 1096 39948 1148
rect 40000 1136 40006 1148
rect 86586 1136 86592 1148
rect 40000 1108 86592 1136
rect 40000 1096 40006 1108
rect 86586 1096 86592 1108
rect 86644 1096 86650 1148
rect 4430 1028 4436 1080
rect 4488 1068 4494 1080
rect 34514 1068 34520 1080
rect 4488 1040 34520 1068
rect 4488 1028 4494 1040
rect 34514 1028 34520 1040
rect 34572 1028 34578 1080
rect 39850 1028 39856 1080
rect 39908 1068 39914 1080
rect 84746 1068 84752 1080
rect 39908 1040 84752 1068
rect 39908 1028 39914 1040
rect 84746 1028 84752 1040
rect 84804 1028 84810 1080
rect 4522 960 4528 1012
rect 4580 1000 4586 1012
rect 30374 1000 30380 1012
rect 4580 972 30380 1000
rect 4580 960 4586 972
rect 30374 960 30380 972
rect 30432 960 30438 1012
rect 41322 960 41328 1012
rect 41380 1000 41386 1012
rect 85482 1000 85488 1012
rect 41380 972 85488 1000
rect 41380 960 41386 972
rect 85482 960 85488 972
rect 85540 960 85546 1012
rect 3878 892 3884 944
rect 3936 932 3942 944
rect 19334 932 19340 944
rect 3936 904 19340 932
rect 3936 892 3942 904
rect 19334 892 19340 904
rect 19392 892 19398 944
rect 24762 892 24768 944
rect 24820 932 24826 944
rect 41414 932 41420 944
rect 24820 904 41420 932
rect 24820 892 24826 904
rect 41414 892 41420 904
rect 41472 892 41478 944
rect 42702 892 42708 944
rect 42760 932 42766 944
rect 86770 932 86776 944
rect 42760 904 86776 932
rect 42760 892 42766 904
rect 86770 892 86776 904
rect 86828 892 86834 944
rect 5626 824 5632 876
rect 5684 864 5690 876
rect 17954 864 17960 876
rect 5684 836 17960 864
rect 5684 824 5690 836
rect 17954 824 17960 836
rect 18012 824 18018 876
rect 44082 824 44088 876
rect 44140 864 44146 876
rect 85206 864 85212 876
rect 44140 836 85212 864
rect 44140 824 44146 836
rect 85206 824 85212 836
rect 85264 824 85270 876
rect 5166 756 5172 808
rect 5224 796 5230 808
rect 27614 796 27620 808
rect 5224 768 27620 796
rect 5224 756 5230 768
rect 27614 756 27620 768
rect 27672 756 27678 808
rect 46842 756 46848 808
rect 46900 796 46906 808
rect 86678 796 86684 808
rect 46900 768 86684 796
rect 46900 756 46906 768
rect 86678 756 86684 768
rect 86736 756 86742 808
rect 3694 688 3700 740
rect 3752 728 3758 740
rect 33134 728 33140 740
rect 3752 700 33140 728
rect 3752 688 3758 700
rect 33134 688 33140 700
rect 33192 688 33198 740
rect 46750 688 46756 740
rect 46808 728 46814 740
rect 85114 728 85120 740
rect 46808 700 85120 728
rect 46808 688 46814 700
rect 85114 688 85120 700
rect 85172 688 85178 740
rect 5074 620 5080 672
rect 5132 660 5138 672
rect 42794 660 42800 672
rect 5132 632 42800 660
rect 5132 620 5138 632
rect 42794 620 42800 632
rect 42852 620 42858 672
rect 49602 620 49608 672
rect 49660 660 49666 672
rect 84838 660 84844 672
rect 49660 632 84844 660
rect 49660 620 49666 632
rect 84838 620 84844 632
rect 84896 620 84902 672
rect 50982 552 50988 604
rect 51040 592 51046 604
rect 82630 592 82636 604
rect 51040 564 82636 592
rect 51040 552 51046 564
rect 82630 552 82636 564
rect 82688 552 82694 604
rect 52362 484 52368 536
rect 52420 524 52426 536
rect 82722 524 82728 536
rect 52420 496 82728 524
rect 52420 484 52426 496
rect 82722 484 82728 496
rect 82780 484 82786 536
rect 53742 416 53748 468
rect 53800 456 53806 468
rect 83826 456 83832 468
rect 53800 428 83832 456
rect 53800 416 53806 428
rect 83826 416 83832 428
rect 83884 416 83890 468
rect 55122 348 55128 400
rect 55180 388 55186 400
rect 83734 388 83740 400
rect 55180 360 83740 388
rect 55180 348 55186 360
rect 83734 348 83740 360
rect 83792 348 83798 400
rect 54662 280 54668 332
rect 54720 320 54726 332
rect 81434 320 81440 332
rect 54720 292 81440 320
rect 54720 280 54726 292
rect 81434 280 81440 292
rect 81492 280 81498 332
rect 55030 212 55036 264
rect 55088 252 55094 264
rect 81342 252 81348 264
rect 55088 224 81348 252
rect 55088 212 55094 224
rect 81342 212 81348 224
rect 81400 212 81406 264
rect 20622 144 20628 196
rect 20680 184 20686 196
rect 86494 184 86500 196
rect 20680 156 86500 184
rect 20680 144 20686 156
rect 86494 144 86500 156
rect 86552 144 86558 196
rect 24762 76 24768 128
rect 24820 116 24826 128
rect 86402 116 86408 128
rect 24820 88 86408 116
rect 24820 76 24826 88
rect 86402 76 86408 88
rect 86460 76 86466 128
<< via1 >>
rect 1982 189286 2034 189338
rect 2046 189286 2098 189338
rect 2110 189286 2162 189338
rect 2174 189286 2226 189338
rect 85982 189286 86034 189338
rect 86046 189286 86098 189338
rect 86110 189286 86162 189338
rect 86174 189286 86226 189338
rect 89982 189286 90034 189338
rect 90046 189286 90098 189338
rect 90110 189286 90162 189338
rect 90174 189286 90226 189338
rect 75828 189048 75880 189100
rect 84476 189048 84528 189100
rect 3982 188742 4034 188794
rect 4046 188742 4098 188794
rect 4110 188742 4162 188794
rect 4174 188742 4226 188794
rect 87982 188742 88034 188794
rect 88046 188742 88098 188794
rect 88110 188742 88162 188794
rect 88174 188742 88226 188794
rect 1982 188198 2034 188250
rect 2046 188198 2098 188250
rect 2110 188198 2162 188250
rect 2174 188198 2226 188250
rect 85982 188198 86034 188250
rect 86046 188198 86098 188250
rect 86110 188198 86162 188250
rect 86174 188198 86226 188250
rect 89982 188198 90034 188250
rect 90046 188198 90098 188250
rect 90110 188198 90162 188250
rect 90174 188198 90226 188250
rect 3982 187654 4034 187706
rect 4046 187654 4098 187706
rect 4110 187654 4162 187706
rect 4174 187654 4226 187706
rect 87982 187654 88034 187706
rect 88046 187654 88098 187706
rect 88110 187654 88162 187706
rect 88174 187654 88226 187706
rect 79324 187348 79376 187400
rect 84476 187212 84528 187264
rect 1982 187110 2034 187162
rect 2046 187110 2098 187162
rect 2110 187110 2162 187162
rect 2174 187110 2226 187162
rect 85982 187110 86034 187162
rect 86046 187110 86098 187162
rect 86110 187110 86162 187162
rect 86174 187110 86226 187162
rect 89982 187110 90034 187162
rect 90046 187110 90098 187162
rect 90110 187110 90162 187162
rect 90174 187110 90226 187162
rect 4436 186736 4488 186788
rect 79324 186804 79376 186856
rect 3982 186566 4034 186618
rect 4046 186566 4098 186618
rect 4110 186566 4162 186618
rect 4174 186566 4226 186618
rect 87982 186566 88034 186618
rect 88046 186566 88098 186618
rect 88110 186566 88162 186618
rect 88174 186566 88226 186618
rect 84384 186328 84436 186380
rect 1982 186022 2034 186074
rect 2046 186022 2098 186074
rect 2110 186022 2162 186074
rect 2174 186022 2226 186074
rect 85982 186022 86034 186074
rect 86046 186022 86098 186074
rect 86110 186022 86162 186074
rect 86174 186022 86226 186074
rect 89982 186022 90034 186074
rect 90046 186022 90098 186074
rect 90110 186022 90162 186074
rect 90174 186022 90226 186074
rect 3982 185478 4034 185530
rect 4046 185478 4098 185530
rect 4110 185478 4162 185530
rect 4174 185478 4226 185530
rect 87982 185478 88034 185530
rect 88046 185478 88098 185530
rect 88110 185478 88162 185530
rect 88174 185478 88226 185530
rect 1982 184934 2034 184986
rect 2046 184934 2098 184986
rect 2110 184934 2162 184986
rect 2174 184934 2226 184986
rect 85982 184934 86034 184986
rect 86046 184934 86098 184986
rect 86110 184934 86162 184986
rect 86174 184934 86226 184986
rect 89982 184934 90034 184986
rect 90046 184934 90098 184986
rect 90110 184934 90162 184986
rect 90174 184934 90226 184986
rect 3982 184390 4034 184442
rect 4046 184390 4098 184442
rect 4110 184390 4162 184442
rect 4174 184390 4226 184442
rect 87982 184390 88034 184442
rect 88046 184390 88098 184442
rect 88110 184390 88162 184442
rect 88174 184390 88226 184442
rect 1982 183846 2034 183898
rect 2046 183846 2098 183898
rect 2110 183846 2162 183898
rect 2174 183846 2226 183898
rect 85982 183846 86034 183898
rect 86046 183846 86098 183898
rect 86110 183846 86162 183898
rect 86174 183846 86226 183898
rect 89982 183846 90034 183898
rect 90046 183846 90098 183898
rect 90110 183846 90162 183898
rect 90174 183846 90226 183898
rect 3982 183302 4034 183354
rect 4046 183302 4098 183354
rect 4110 183302 4162 183354
rect 4174 183302 4226 183354
rect 87982 183302 88034 183354
rect 88046 183302 88098 183354
rect 88110 183302 88162 183354
rect 88174 183302 88226 183354
rect 4804 182971 4856 182980
rect 4804 182937 4813 182971
rect 4813 182937 4847 182971
rect 4847 182937 4856 182971
rect 4804 182928 4856 182937
rect 1982 182758 2034 182810
rect 2046 182758 2098 182810
rect 2110 182758 2162 182810
rect 2174 182758 2226 182810
rect 85982 182758 86034 182810
rect 86046 182758 86098 182810
rect 86110 182758 86162 182810
rect 86174 182758 86226 182810
rect 89982 182758 90034 182810
rect 90046 182758 90098 182810
rect 90110 182758 90162 182810
rect 90174 182758 90226 182810
rect 3982 182214 4034 182266
rect 4046 182214 4098 182266
rect 4110 182214 4162 182266
rect 4174 182214 4226 182266
rect 87982 182214 88034 182266
rect 88046 182214 88098 182266
rect 88110 182214 88162 182266
rect 88174 182214 88226 182266
rect 4804 181883 4856 181892
rect 4804 181849 4813 181883
rect 4813 181849 4847 181883
rect 4847 181849 4856 181883
rect 4804 181840 4856 181849
rect 1982 181670 2034 181722
rect 2046 181670 2098 181722
rect 2110 181670 2162 181722
rect 2174 181670 2226 181722
rect 85982 181670 86034 181722
rect 86046 181670 86098 181722
rect 86110 181670 86162 181722
rect 86174 181670 86226 181722
rect 89982 181670 90034 181722
rect 90046 181670 90098 181722
rect 90110 181670 90162 181722
rect 90174 181670 90226 181722
rect 3982 181126 4034 181178
rect 4046 181126 4098 181178
rect 4110 181126 4162 181178
rect 4174 181126 4226 181178
rect 87982 181126 88034 181178
rect 88046 181126 88098 181178
rect 88110 181126 88162 181178
rect 88174 181126 88226 181178
rect 83740 180820 83792 180872
rect 87696 180820 87748 180872
rect 1982 180582 2034 180634
rect 2046 180582 2098 180634
rect 2110 180582 2162 180634
rect 2174 180582 2226 180634
rect 85982 180582 86034 180634
rect 86046 180582 86098 180634
rect 86110 180582 86162 180634
rect 86174 180582 86226 180634
rect 89982 180582 90034 180634
rect 90046 180582 90098 180634
rect 90110 180582 90162 180634
rect 90174 180582 90226 180634
rect 4620 180140 4672 180192
rect 3982 180038 4034 180090
rect 4046 180038 4098 180090
rect 4110 180038 4162 180090
rect 4174 180038 4226 180090
rect 87982 180038 88034 180090
rect 88046 180038 88098 180090
rect 88110 180038 88162 180090
rect 88174 180038 88226 180090
rect 84568 179596 84620 179648
rect 1982 179494 2034 179546
rect 2046 179494 2098 179546
rect 2110 179494 2162 179546
rect 2174 179494 2226 179546
rect 85982 179494 86034 179546
rect 86046 179494 86098 179546
rect 86110 179494 86162 179546
rect 86174 179494 86226 179546
rect 89982 179494 90034 179546
rect 90046 179494 90098 179546
rect 90110 179494 90162 179546
rect 90174 179494 90226 179546
rect 4528 179052 4580 179104
rect 3982 178950 4034 179002
rect 4046 178950 4098 179002
rect 4110 178950 4162 179002
rect 4174 178950 4226 179002
rect 87982 178950 88034 179002
rect 88046 178950 88098 179002
rect 88110 178950 88162 179002
rect 88174 178950 88226 179002
rect 1982 178406 2034 178458
rect 2046 178406 2098 178458
rect 2110 178406 2162 178458
rect 2174 178406 2226 178458
rect 85982 178406 86034 178458
rect 86046 178406 86098 178458
rect 86110 178406 86162 178458
rect 86174 178406 86226 178458
rect 89982 178406 90034 178458
rect 90046 178406 90098 178458
rect 90110 178406 90162 178458
rect 90174 178406 90226 178458
rect 3982 177862 4034 177914
rect 4046 177862 4098 177914
rect 4110 177862 4162 177914
rect 4174 177862 4226 177914
rect 87982 177862 88034 177914
rect 88046 177862 88098 177914
rect 88110 177862 88162 177914
rect 88174 177862 88226 177914
rect 1982 177318 2034 177370
rect 2046 177318 2098 177370
rect 2110 177318 2162 177370
rect 2174 177318 2226 177370
rect 85982 177318 86034 177370
rect 86046 177318 86098 177370
rect 86110 177318 86162 177370
rect 86174 177318 86226 177370
rect 89982 177318 90034 177370
rect 90046 177318 90098 177370
rect 90110 177318 90162 177370
rect 90174 177318 90226 177370
rect 4712 176919 4764 176928
rect 4712 176885 4721 176919
rect 4721 176885 4755 176919
rect 4755 176885 4764 176919
rect 4712 176876 4764 176885
rect 3982 176774 4034 176826
rect 4046 176774 4098 176826
rect 4110 176774 4162 176826
rect 4174 176774 4226 176826
rect 87982 176774 88034 176826
rect 88046 176774 88098 176826
rect 88110 176774 88162 176826
rect 88174 176774 88226 176826
rect 1982 176230 2034 176282
rect 2046 176230 2098 176282
rect 2110 176230 2162 176282
rect 2174 176230 2226 176282
rect 85982 176230 86034 176282
rect 86046 176230 86098 176282
rect 86110 176230 86162 176282
rect 86174 176230 86226 176282
rect 89982 176230 90034 176282
rect 90046 176230 90098 176282
rect 90110 176230 90162 176282
rect 90174 176230 90226 176282
rect 4804 176171 4856 176180
rect 4804 176137 4813 176171
rect 4813 176137 4847 176171
rect 4847 176137 4856 176171
rect 4804 176128 4856 176137
rect 3982 175686 4034 175738
rect 4046 175686 4098 175738
rect 4110 175686 4162 175738
rect 4174 175686 4226 175738
rect 87982 175686 88034 175738
rect 88046 175686 88098 175738
rect 88110 175686 88162 175738
rect 88174 175686 88226 175738
rect 1982 175142 2034 175194
rect 2046 175142 2098 175194
rect 2110 175142 2162 175194
rect 2174 175142 2226 175194
rect 85982 175142 86034 175194
rect 86046 175142 86098 175194
rect 86110 175142 86162 175194
rect 86174 175142 86226 175194
rect 89982 175142 90034 175194
rect 90046 175142 90098 175194
rect 90110 175142 90162 175194
rect 90174 175142 90226 175194
rect 3982 174598 4034 174650
rect 4046 174598 4098 174650
rect 4110 174598 4162 174650
rect 4174 174598 4226 174650
rect 87982 174598 88034 174650
rect 88046 174598 88098 174650
rect 88110 174598 88162 174650
rect 88174 174598 88226 174650
rect 4804 174539 4856 174548
rect 4804 174505 4813 174539
rect 4813 174505 4847 174539
rect 4847 174505 4856 174539
rect 4804 174496 4856 174505
rect 4528 174360 4580 174412
rect 4804 174360 4856 174412
rect 4620 174292 4672 174344
rect 4988 174292 5040 174344
rect 1982 174054 2034 174106
rect 2046 174054 2098 174106
rect 2110 174054 2162 174106
rect 2174 174054 2226 174106
rect 85982 174054 86034 174106
rect 86046 174054 86098 174106
rect 86110 174054 86162 174106
rect 86174 174054 86226 174106
rect 89982 174054 90034 174106
rect 90046 174054 90098 174106
rect 90110 174054 90162 174106
rect 90174 174054 90226 174106
rect 83924 173884 83976 173936
rect 87420 173884 87472 173936
rect 3982 173510 4034 173562
rect 4046 173510 4098 173562
rect 4110 173510 4162 173562
rect 4174 173510 4226 173562
rect 87982 173510 88034 173562
rect 88046 173510 88098 173562
rect 88110 173510 88162 173562
rect 88174 173510 88226 173562
rect 1982 172966 2034 173018
rect 2046 172966 2098 173018
rect 2110 172966 2162 173018
rect 2174 172966 2226 173018
rect 85982 172966 86034 173018
rect 86046 172966 86098 173018
rect 86110 172966 86162 173018
rect 86174 172966 86226 173018
rect 89982 172966 90034 173018
rect 90046 172966 90098 173018
rect 90110 172966 90162 173018
rect 90174 172966 90226 173018
rect 3982 172422 4034 172474
rect 4046 172422 4098 172474
rect 4110 172422 4162 172474
rect 4174 172422 4226 172474
rect 87982 172422 88034 172474
rect 88046 172422 88098 172474
rect 88110 172422 88162 172474
rect 88174 172422 88226 172474
rect 1982 171878 2034 171930
rect 2046 171878 2098 171930
rect 2110 171878 2162 171930
rect 2174 171878 2226 171930
rect 85982 171878 86034 171930
rect 86046 171878 86098 171930
rect 86110 171878 86162 171930
rect 86174 171878 86226 171930
rect 89982 171878 90034 171930
rect 90046 171878 90098 171930
rect 90110 171878 90162 171930
rect 90174 171878 90226 171930
rect 3982 171334 4034 171386
rect 4046 171334 4098 171386
rect 4110 171334 4162 171386
rect 4174 171334 4226 171386
rect 87982 171334 88034 171386
rect 88046 171334 88098 171386
rect 88110 171334 88162 171386
rect 88174 171334 88226 171386
rect 1982 170790 2034 170842
rect 2046 170790 2098 170842
rect 2110 170790 2162 170842
rect 2174 170790 2226 170842
rect 85982 170790 86034 170842
rect 86046 170790 86098 170842
rect 86110 170790 86162 170842
rect 86174 170790 86226 170842
rect 89982 170790 90034 170842
rect 90046 170790 90098 170842
rect 90110 170790 90162 170842
rect 90174 170790 90226 170842
rect 3982 170246 4034 170298
rect 4046 170246 4098 170298
rect 4110 170246 4162 170298
rect 4174 170246 4226 170298
rect 87982 170246 88034 170298
rect 88046 170246 88098 170298
rect 88110 170246 88162 170298
rect 88174 170246 88226 170298
rect 1982 169702 2034 169754
rect 2046 169702 2098 169754
rect 2110 169702 2162 169754
rect 2174 169702 2226 169754
rect 85982 169702 86034 169754
rect 86046 169702 86098 169754
rect 86110 169702 86162 169754
rect 86174 169702 86226 169754
rect 89982 169702 90034 169754
rect 90046 169702 90098 169754
rect 90110 169702 90162 169754
rect 90174 169702 90226 169754
rect 3982 169158 4034 169210
rect 4046 169158 4098 169210
rect 4110 169158 4162 169210
rect 4174 169158 4226 169210
rect 87982 169158 88034 169210
rect 88046 169158 88098 169210
rect 88110 169158 88162 169210
rect 88174 169158 88226 169210
rect 1982 168614 2034 168666
rect 2046 168614 2098 168666
rect 2110 168614 2162 168666
rect 2174 168614 2226 168666
rect 85982 168614 86034 168666
rect 86046 168614 86098 168666
rect 86110 168614 86162 168666
rect 86174 168614 86226 168666
rect 89982 168614 90034 168666
rect 90046 168614 90098 168666
rect 90110 168614 90162 168666
rect 90174 168614 90226 168666
rect 84016 168376 84068 168428
rect 87880 168376 87932 168428
rect 3982 168070 4034 168122
rect 4046 168070 4098 168122
rect 4110 168070 4162 168122
rect 4174 168070 4226 168122
rect 87982 168070 88034 168122
rect 88046 168070 88098 168122
rect 88110 168070 88162 168122
rect 88174 168070 88226 168122
rect 1982 167526 2034 167578
rect 2046 167526 2098 167578
rect 2110 167526 2162 167578
rect 2174 167526 2226 167578
rect 85982 167526 86034 167578
rect 86046 167526 86098 167578
rect 86110 167526 86162 167578
rect 86174 167526 86226 167578
rect 89982 167526 90034 167578
rect 90046 167526 90098 167578
rect 90110 167526 90162 167578
rect 90174 167526 90226 167578
rect 84476 167467 84528 167476
rect 84476 167433 84485 167467
rect 84485 167433 84519 167467
rect 84519 167433 84528 167467
rect 84476 167424 84528 167433
rect 83556 167084 83608 167136
rect 87052 167084 87104 167136
rect 3982 166982 4034 167034
rect 4046 166982 4098 167034
rect 4110 166982 4162 167034
rect 4174 166982 4226 167034
rect 87982 166982 88034 167034
rect 88046 166982 88098 167034
rect 88110 166982 88162 167034
rect 88174 166982 88226 167034
rect 1982 166438 2034 166490
rect 2046 166438 2098 166490
rect 2110 166438 2162 166490
rect 2174 166438 2226 166490
rect 85982 166438 86034 166490
rect 86046 166438 86098 166490
rect 86110 166438 86162 166490
rect 86174 166438 86226 166490
rect 89982 166438 90034 166490
rect 90046 166438 90098 166490
rect 90110 166438 90162 166490
rect 90174 166438 90226 166490
rect 3982 165894 4034 165946
rect 4046 165894 4098 165946
rect 4110 165894 4162 165946
rect 4174 165894 4226 165946
rect 87982 165894 88034 165946
rect 88046 165894 88098 165946
rect 88110 165894 88162 165946
rect 88174 165894 88226 165946
rect 1982 165350 2034 165402
rect 2046 165350 2098 165402
rect 2110 165350 2162 165402
rect 2174 165350 2226 165402
rect 85982 165350 86034 165402
rect 86046 165350 86098 165402
rect 86110 165350 86162 165402
rect 86174 165350 86226 165402
rect 89982 165350 90034 165402
rect 90046 165350 90098 165402
rect 90110 165350 90162 165402
rect 90174 165350 90226 165402
rect 3982 164806 4034 164858
rect 4046 164806 4098 164858
rect 4110 164806 4162 164858
rect 4174 164806 4226 164858
rect 87982 164806 88034 164858
rect 88046 164806 88098 164858
rect 88110 164806 88162 164858
rect 88174 164806 88226 164858
rect 83832 164364 83884 164416
rect 87880 164364 87932 164416
rect 1982 164262 2034 164314
rect 2046 164262 2098 164314
rect 2110 164262 2162 164314
rect 2174 164262 2226 164314
rect 85982 164262 86034 164314
rect 86046 164262 86098 164314
rect 86110 164262 86162 164314
rect 86174 164262 86226 164314
rect 89982 164262 90034 164314
rect 90046 164262 90098 164314
rect 90110 164262 90162 164314
rect 90174 164262 90226 164314
rect 3982 163718 4034 163770
rect 4046 163718 4098 163770
rect 4110 163718 4162 163770
rect 4174 163718 4226 163770
rect 87982 163718 88034 163770
rect 88046 163718 88098 163770
rect 88110 163718 88162 163770
rect 88174 163718 88226 163770
rect 1982 163174 2034 163226
rect 2046 163174 2098 163226
rect 2110 163174 2162 163226
rect 2174 163174 2226 163226
rect 85982 163174 86034 163226
rect 86046 163174 86098 163226
rect 86110 163174 86162 163226
rect 86174 163174 86226 163226
rect 89982 163174 90034 163226
rect 90046 163174 90098 163226
rect 90110 163174 90162 163226
rect 90174 163174 90226 163226
rect 82452 162868 82504 162920
rect 87880 162868 87932 162920
rect 3982 162630 4034 162682
rect 4046 162630 4098 162682
rect 4110 162630 4162 162682
rect 4174 162630 4226 162682
rect 87982 162630 88034 162682
rect 88046 162630 88098 162682
rect 88110 162630 88162 162682
rect 88174 162630 88226 162682
rect 84660 162435 84712 162444
rect 84660 162401 84669 162435
rect 84669 162401 84703 162435
rect 84703 162401 84712 162435
rect 84660 162392 84712 162401
rect 85120 162367 85172 162376
rect 85120 162333 85129 162367
rect 85129 162333 85163 162367
rect 85163 162333 85172 162367
rect 85120 162324 85172 162333
rect 1982 162086 2034 162138
rect 2046 162086 2098 162138
rect 2110 162086 2162 162138
rect 2174 162086 2226 162138
rect 85982 162086 86034 162138
rect 86046 162086 86098 162138
rect 86110 162086 86162 162138
rect 86174 162086 86226 162138
rect 89982 162086 90034 162138
rect 90046 162086 90098 162138
rect 90110 162086 90162 162138
rect 90174 162086 90226 162138
rect 84660 162027 84712 162036
rect 84660 161993 84669 162027
rect 84669 161993 84703 162027
rect 84703 161993 84712 162027
rect 84660 161984 84712 161993
rect 3982 161542 4034 161594
rect 4046 161542 4098 161594
rect 4110 161542 4162 161594
rect 4174 161542 4226 161594
rect 87982 161542 88034 161594
rect 88046 161542 88098 161594
rect 88110 161542 88162 161594
rect 88174 161542 88226 161594
rect 1982 160998 2034 161050
rect 2046 160998 2098 161050
rect 2110 160998 2162 161050
rect 2174 160998 2226 161050
rect 85982 160998 86034 161050
rect 86046 160998 86098 161050
rect 86110 160998 86162 161050
rect 86174 160998 86226 161050
rect 89982 160998 90034 161050
rect 90046 160998 90098 161050
rect 90110 160998 90162 161050
rect 90174 160998 90226 161050
rect 3982 160454 4034 160506
rect 4046 160454 4098 160506
rect 4110 160454 4162 160506
rect 4174 160454 4226 160506
rect 87982 160454 88034 160506
rect 88046 160454 88098 160506
rect 88110 160454 88162 160506
rect 88174 160454 88226 160506
rect 84476 160123 84528 160132
rect 84476 160089 84485 160123
rect 84485 160089 84519 160123
rect 84519 160089 84528 160123
rect 84476 160080 84528 160089
rect 1982 159910 2034 159962
rect 2046 159910 2098 159962
rect 2110 159910 2162 159962
rect 2174 159910 2226 159962
rect 85982 159910 86034 159962
rect 86046 159910 86098 159962
rect 86110 159910 86162 159962
rect 86174 159910 86226 159962
rect 89982 159910 90034 159962
rect 90046 159910 90098 159962
rect 90110 159910 90162 159962
rect 90174 159910 90226 159962
rect 3982 159366 4034 159418
rect 4046 159366 4098 159418
rect 4110 159366 4162 159418
rect 4174 159366 4226 159418
rect 87982 159366 88034 159418
rect 88046 159366 88098 159418
rect 88110 159366 88162 159418
rect 88174 159366 88226 159418
rect 1982 158822 2034 158874
rect 2046 158822 2098 158874
rect 2110 158822 2162 158874
rect 2174 158822 2226 158874
rect 85982 158822 86034 158874
rect 86046 158822 86098 158874
rect 86110 158822 86162 158874
rect 86174 158822 86226 158874
rect 89982 158822 90034 158874
rect 90046 158822 90098 158874
rect 90110 158822 90162 158874
rect 90174 158822 90226 158874
rect 3982 158278 4034 158330
rect 4046 158278 4098 158330
rect 4110 158278 4162 158330
rect 4174 158278 4226 158330
rect 87982 158278 88034 158330
rect 88046 158278 88098 158330
rect 88110 158278 88162 158330
rect 88174 158278 88226 158330
rect 1982 157734 2034 157786
rect 2046 157734 2098 157786
rect 2110 157734 2162 157786
rect 2174 157734 2226 157786
rect 85982 157734 86034 157786
rect 86046 157734 86098 157786
rect 86110 157734 86162 157786
rect 86174 157734 86226 157786
rect 89982 157734 90034 157786
rect 90046 157734 90098 157786
rect 90110 157734 90162 157786
rect 90174 157734 90226 157786
rect 3982 157190 4034 157242
rect 4046 157190 4098 157242
rect 4110 157190 4162 157242
rect 4174 157190 4226 157242
rect 87982 157190 88034 157242
rect 88046 157190 88098 157242
rect 88110 157190 88162 157242
rect 88174 157190 88226 157242
rect 1982 156646 2034 156698
rect 2046 156646 2098 156698
rect 2110 156646 2162 156698
rect 2174 156646 2226 156698
rect 85982 156646 86034 156698
rect 86046 156646 86098 156698
rect 86110 156646 86162 156698
rect 86174 156646 86226 156698
rect 89982 156646 90034 156698
rect 90046 156646 90098 156698
rect 90110 156646 90162 156698
rect 90174 156646 90226 156698
rect 3982 156102 4034 156154
rect 4046 156102 4098 156154
rect 4110 156102 4162 156154
rect 4174 156102 4226 156154
rect 87982 156102 88034 156154
rect 88046 156102 88098 156154
rect 88110 156102 88162 156154
rect 88174 156102 88226 156154
rect 1982 155558 2034 155610
rect 2046 155558 2098 155610
rect 2110 155558 2162 155610
rect 2174 155558 2226 155610
rect 85982 155558 86034 155610
rect 86046 155558 86098 155610
rect 86110 155558 86162 155610
rect 86174 155558 86226 155610
rect 89982 155558 90034 155610
rect 90046 155558 90098 155610
rect 90110 155558 90162 155610
rect 90174 155558 90226 155610
rect 3982 155014 4034 155066
rect 4046 155014 4098 155066
rect 4110 155014 4162 155066
rect 4174 155014 4226 155066
rect 87982 155014 88034 155066
rect 88046 155014 88098 155066
rect 88110 155014 88162 155066
rect 88174 155014 88226 155066
rect 1982 154470 2034 154522
rect 2046 154470 2098 154522
rect 2110 154470 2162 154522
rect 2174 154470 2226 154522
rect 85982 154470 86034 154522
rect 86046 154470 86098 154522
rect 86110 154470 86162 154522
rect 86174 154470 86226 154522
rect 89982 154470 90034 154522
rect 90046 154470 90098 154522
rect 90110 154470 90162 154522
rect 90174 154470 90226 154522
rect 3982 153926 4034 153978
rect 4046 153926 4098 153978
rect 4110 153926 4162 153978
rect 4174 153926 4226 153978
rect 87982 153926 88034 153978
rect 88046 153926 88098 153978
rect 88110 153926 88162 153978
rect 88174 153926 88226 153978
rect 84384 153824 84436 153876
rect 1982 153382 2034 153434
rect 2046 153382 2098 153434
rect 2110 153382 2162 153434
rect 2174 153382 2226 153434
rect 85982 153382 86034 153434
rect 86046 153382 86098 153434
rect 86110 153382 86162 153434
rect 86174 153382 86226 153434
rect 89982 153382 90034 153434
rect 90046 153382 90098 153434
rect 90110 153382 90162 153434
rect 90174 153382 90226 153434
rect 3982 152838 4034 152890
rect 4046 152838 4098 152890
rect 4110 152838 4162 152890
rect 4174 152838 4226 152890
rect 87982 152838 88034 152890
rect 88046 152838 88098 152890
rect 88110 152838 88162 152890
rect 88174 152838 88226 152890
rect 1982 152294 2034 152346
rect 2046 152294 2098 152346
rect 2110 152294 2162 152346
rect 2174 152294 2226 152346
rect 85982 152294 86034 152346
rect 86046 152294 86098 152346
rect 86110 152294 86162 152346
rect 86174 152294 86226 152346
rect 89982 152294 90034 152346
rect 90046 152294 90098 152346
rect 90110 152294 90162 152346
rect 90174 152294 90226 152346
rect 3982 151750 4034 151802
rect 4046 151750 4098 151802
rect 4110 151750 4162 151802
rect 4174 151750 4226 151802
rect 87982 151750 88034 151802
rect 88046 151750 88098 151802
rect 88110 151750 88162 151802
rect 88174 151750 88226 151802
rect 1982 151206 2034 151258
rect 2046 151206 2098 151258
rect 2110 151206 2162 151258
rect 2174 151206 2226 151258
rect 85982 151206 86034 151258
rect 86046 151206 86098 151258
rect 86110 151206 86162 151258
rect 86174 151206 86226 151258
rect 89982 151206 90034 151258
rect 90046 151206 90098 151258
rect 90110 151206 90162 151258
rect 90174 151206 90226 151258
rect 3982 150662 4034 150714
rect 4046 150662 4098 150714
rect 4110 150662 4162 150714
rect 4174 150662 4226 150714
rect 87982 150662 88034 150714
rect 88046 150662 88098 150714
rect 88110 150662 88162 150714
rect 88174 150662 88226 150714
rect 1982 150118 2034 150170
rect 2046 150118 2098 150170
rect 2110 150118 2162 150170
rect 2174 150118 2226 150170
rect 85982 150118 86034 150170
rect 86046 150118 86098 150170
rect 86110 150118 86162 150170
rect 86174 150118 86226 150170
rect 89982 150118 90034 150170
rect 90046 150118 90098 150170
rect 90110 150118 90162 150170
rect 90174 150118 90226 150170
rect 3982 149574 4034 149626
rect 4046 149574 4098 149626
rect 4110 149574 4162 149626
rect 4174 149574 4226 149626
rect 87982 149574 88034 149626
rect 88046 149574 88098 149626
rect 88110 149574 88162 149626
rect 88174 149574 88226 149626
rect 1982 149030 2034 149082
rect 2046 149030 2098 149082
rect 2110 149030 2162 149082
rect 2174 149030 2226 149082
rect 85982 149030 86034 149082
rect 86046 149030 86098 149082
rect 86110 149030 86162 149082
rect 86174 149030 86226 149082
rect 89982 149030 90034 149082
rect 90046 149030 90098 149082
rect 90110 149030 90162 149082
rect 90174 149030 90226 149082
rect 3982 148486 4034 148538
rect 4046 148486 4098 148538
rect 4110 148486 4162 148538
rect 4174 148486 4226 148538
rect 87982 148486 88034 148538
rect 88046 148486 88098 148538
rect 88110 148486 88162 148538
rect 88174 148486 88226 148538
rect 1982 147942 2034 147994
rect 2046 147942 2098 147994
rect 2110 147942 2162 147994
rect 2174 147942 2226 147994
rect 85982 147942 86034 147994
rect 86046 147942 86098 147994
rect 86110 147942 86162 147994
rect 86174 147942 86226 147994
rect 89982 147942 90034 147994
rect 90046 147942 90098 147994
rect 90110 147942 90162 147994
rect 90174 147942 90226 147994
rect 3982 147398 4034 147450
rect 4046 147398 4098 147450
rect 4110 147398 4162 147450
rect 4174 147398 4226 147450
rect 87982 147398 88034 147450
rect 88046 147398 88098 147450
rect 88110 147398 88162 147450
rect 88174 147398 88226 147450
rect 1982 146854 2034 146906
rect 2046 146854 2098 146906
rect 2110 146854 2162 146906
rect 2174 146854 2226 146906
rect 85982 146854 86034 146906
rect 86046 146854 86098 146906
rect 86110 146854 86162 146906
rect 86174 146854 86226 146906
rect 89982 146854 90034 146906
rect 90046 146854 90098 146906
rect 90110 146854 90162 146906
rect 90174 146854 90226 146906
rect 3982 146310 4034 146362
rect 4046 146310 4098 146362
rect 4110 146310 4162 146362
rect 4174 146310 4226 146362
rect 87982 146310 88034 146362
rect 88046 146310 88098 146362
rect 88110 146310 88162 146362
rect 88174 146310 88226 146362
rect 1982 145766 2034 145818
rect 2046 145766 2098 145818
rect 2110 145766 2162 145818
rect 2174 145766 2226 145818
rect 85982 145766 86034 145818
rect 86046 145766 86098 145818
rect 86110 145766 86162 145818
rect 86174 145766 86226 145818
rect 89982 145766 90034 145818
rect 90046 145766 90098 145818
rect 90110 145766 90162 145818
rect 90174 145766 90226 145818
rect 3982 145222 4034 145274
rect 4046 145222 4098 145274
rect 4110 145222 4162 145274
rect 4174 145222 4226 145274
rect 87982 145222 88034 145274
rect 88046 145222 88098 145274
rect 88110 145222 88162 145274
rect 88174 145222 88226 145274
rect 84752 144916 84804 144968
rect 87972 144916 88024 144968
rect 1982 144678 2034 144730
rect 2046 144678 2098 144730
rect 2110 144678 2162 144730
rect 2174 144678 2226 144730
rect 85982 144678 86034 144730
rect 86046 144678 86098 144730
rect 86110 144678 86162 144730
rect 86174 144678 86226 144730
rect 89982 144678 90034 144730
rect 90046 144678 90098 144730
rect 90110 144678 90162 144730
rect 90174 144678 90226 144730
rect 3982 144134 4034 144186
rect 4046 144134 4098 144186
rect 4110 144134 4162 144186
rect 4174 144134 4226 144186
rect 87982 144134 88034 144186
rect 88046 144134 88098 144186
rect 88110 144134 88162 144186
rect 88174 144134 88226 144186
rect 85764 143692 85816 143744
rect 88064 143692 88116 143744
rect 1982 143590 2034 143642
rect 2046 143590 2098 143642
rect 2110 143590 2162 143642
rect 2174 143590 2226 143642
rect 85982 143590 86034 143642
rect 86046 143590 86098 143642
rect 86110 143590 86162 143642
rect 86174 143590 86226 143642
rect 89982 143590 90034 143642
rect 90046 143590 90098 143642
rect 90110 143590 90162 143642
rect 90174 143590 90226 143642
rect 3982 143046 4034 143098
rect 4046 143046 4098 143098
rect 4110 143046 4162 143098
rect 4174 143046 4226 143098
rect 87982 143046 88034 143098
rect 88046 143046 88098 143098
rect 88110 143046 88162 143098
rect 88174 143046 88226 143098
rect 1982 142502 2034 142554
rect 2046 142502 2098 142554
rect 2110 142502 2162 142554
rect 2174 142502 2226 142554
rect 85982 142502 86034 142554
rect 86046 142502 86098 142554
rect 86110 142502 86162 142554
rect 86174 142502 86226 142554
rect 89982 142502 90034 142554
rect 90046 142502 90098 142554
rect 90110 142502 90162 142554
rect 90174 142502 90226 142554
rect 85856 142400 85908 142452
rect 87972 142400 88024 142452
rect 3982 141958 4034 142010
rect 4046 141958 4098 142010
rect 4110 141958 4162 142010
rect 4174 141958 4226 142010
rect 87982 141958 88034 142010
rect 88046 141958 88098 142010
rect 88110 141958 88162 142010
rect 88174 141958 88226 142010
rect 1982 141414 2034 141466
rect 2046 141414 2098 141466
rect 2110 141414 2162 141466
rect 2174 141414 2226 141466
rect 85982 141414 86034 141466
rect 86046 141414 86098 141466
rect 86110 141414 86162 141466
rect 86174 141414 86226 141466
rect 89982 141414 90034 141466
rect 90046 141414 90098 141466
rect 90110 141414 90162 141466
rect 90174 141414 90226 141466
rect 84200 141176 84252 141228
rect 87972 141176 88024 141228
rect 84660 141083 84712 141092
rect 84660 141049 84669 141083
rect 84669 141049 84703 141083
rect 84703 141049 84712 141083
rect 84660 141040 84712 141049
rect 85212 141015 85264 141024
rect 85212 140981 85221 141015
rect 85221 140981 85255 141015
rect 85255 140981 85264 141015
rect 85212 140972 85264 140981
rect 3982 140870 4034 140922
rect 4046 140870 4098 140922
rect 4110 140870 4162 140922
rect 4174 140870 4226 140922
rect 87982 140870 88034 140922
rect 88046 140870 88098 140922
rect 88110 140870 88162 140922
rect 88174 140870 88226 140922
rect 1982 140326 2034 140378
rect 2046 140326 2098 140378
rect 2110 140326 2162 140378
rect 2174 140326 2226 140378
rect 85982 140326 86034 140378
rect 86046 140326 86098 140378
rect 86110 140326 86162 140378
rect 86174 140326 86226 140378
rect 89982 140326 90034 140378
rect 90046 140326 90098 140378
rect 90110 140326 90162 140378
rect 90174 140326 90226 140378
rect 85120 139952 85172 140004
rect 88248 139952 88300 140004
rect 3982 139782 4034 139834
rect 4046 139782 4098 139834
rect 4110 139782 4162 139834
rect 4174 139782 4226 139834
rect 87982 139782 88034 139834
rect 88046 139782 88098 139834
rect 88110 139782 88162 139834
rect 88174 139782 88226 139834
rect 1982 139238 2034 139290
rect 2046 139238 2098 139290
rect 2110 139238 2162 139290
rect 2174 139238 2226 139290
rect 85982 139238 86034 139290
rect 86046 139238 86098 139290
rect 86110 139238 86162 139290
rect 86174 139238 86226 139290
rect 89982 139238 90034 139290
rect 90046 139238 90098 139290
rect 90110 139238 90162 139290
rect 90174 139238 90226 139290
rect 84844 138864 84896 138916
rect 88064 138864 88116 138916
rect 3982 138694 4034 138746
rect 4046 138694 4098 138746
rect 4110 138694 4162 138746
rect 4174 138694 4226 138746
rect 87982 138694 88034 138746
rect 88046 138694 88098 138746
rect 88110 138694 88162 138746
rect 88174 138694 88226 138746
rect 1982 138150 2034 138202
rect 2046 138150 2098 138202
rect 2110 138150 2162 138202
rect 2174 138150 2226 138202
rect 85982 138150 86034 138202
rect 86046 138150 86098 138202
rect 86110 138150 86162 138202
rect 86174 138150 86226 138202
rect 89982 138150 90034 138202
rect 90046 138150 90098 138202
rect 90110 138150 90162 138202
rect 90174 138150 90226 138202
rect 3982 137606 4034 137658
rect 4046 137606 4098 137658
rect 4110 137606 4162 137658
rect 4174 137606 4226 137658
rect 87982 137606 88034 137658
rect 88046 137606 88098 137658
rect 88110 137606 88162 137658
rect 88174 137606 88226 137658
rect 1982 137062 2034 137114
rect 2046 137062 2098 137114
rect 2110 137062 2162 137114
rect 2174 137062 2226 137114
rect 85982 137062 86034 137114
rect 86046 137062 86098 137114
rect 86110 137062 86162 137114
rect 86174 137062 86226 137114
rect 89982 137062 90034 137114
rect 90046 137062 90098 137114
rect 90110 137062 90162 137114
rect 90174 137062 90226 137114
rect 3982 136518 4034 136570
rect 4046 136518 4098 136570
rect 4110 136518 4162 136570
rect 4174 136518 4226 136570
rect 87982 136518 88034 136570
rect 88046 136518 88098 136570
rect 88110 136518 88162 136570
rect 88174 136518 88226 136570
rect 1982 135974 2034 136026
rect 2046 135974 2098 136026
rect 2110 135974 2162 136026
rect 2174 135974 2226 136026
rect 85982 135974 86034 136026
rect 86046 135974 86098 136026
rect 86110 135974 86162 136026
rect 86174 135974 86226 136026
rect 89982 135974 90034 136026
rect 90046 135974 90098 136026
rect 90110 135974 90162 136026
rect 90174 135974 90226 136026
rect 3982 135430 4034 135482
rect 4046 135430 4098 135482
rect 4110 135430 4162 135482
rect 4174 135430 4226 135482
rect 87982 135430 88034 135482
rect 88046 135430 88098 135482
rect 88110 135430 88162 135482
rect 88174 135430 88226 135482
rect 1982 134886 2034 134938
rect 2046 134886 2098 134938
rect 2110 134886 2162 134938
rect 2174 134886 2226 134938
rect 85982 134886 86034 134938
rect 86046 134886 86098 134938
rect 86110 134886 86162 134938
rect 86174 134886 86226 134938
rect 89982 134886 90034 134938
rect 90046 134886 90098 134938
rect 90110 134886 90162 134938
rect 90174 134886 90226 134938
rect 3982 134342 4034 134394
rect 4046 134342 4098 134394
rect 4110 134342 4162 134394
rect 4174 134342 4226 134394
rect 87982 134342 88034 134394
rect 88046 134342 88098 134394
rect 88110 134342 88162 134394
rect 88174 134342 88226 134394
rect 1982 133798 2034 133850
rect 2046 133798 2098 133850
rect 2110 133798 2162 133850
rect 2174 133798 2226 133850
rect 85982 133798 86034 133850
rect 86046 133798 86098 133850
rect 86110 133798 86162 133850
rect 86174 133798 86226 133850
rect 89982 133798 90034 133850
rect 90046 133798 90098 133850
rect 90110 133798 90162 133850
rect 90174 133798 90226 133850
rect 3982 133254 4034 133306
rect 4046 133254 4098 133306
rect 4110 133254 4162 133306
rect 4174 133254 4226 133306
rect 87982 133254 88034 133306
rect 88046 133254 88098 133306
rect 88110 133254 88162 133306
rect 88174 133254 88226 133306
rect 1982 132710 2034 132762
rect 2046 132710 2098 132762
rect 2110 132710 2162 132762
rect 2174 132710 2226 132762
rect 85982 132710 86034 132762
rect 86046 132710 86098 132762
rect 86110 132710 86162 132762
rect 86174 132710 86226 132762
rect 89982 132710 90034 132762
rect 90046 132710 90098 132762
rect 90110 132710 90162 132762
rect 90174 132710 90226 132762
rect 3982 132166 4034 132218
rect 4046 132166 4098 132218
rect 4110 132166 4162 132218
rect 4174 132166 4226 132218
rect 87982 132166 88034 132218
rect 88046 132166 88098 132218
rect 88110 132166 88162 132218
rect 88174 132166 88226 132218
rect 1982 131622 2034 131674
rect 2046 131622 2098 131674
rect 2110 131622 2162 131674
rect 2174 131622 2226 131674
rect 85982 131622 86034 131674
rect 86046 131622 86098 131674
rect 86110 131622 86162 131674
rect 86174 131622 86226 131674
rect 89982 131622 90034 131674
rect 90046 131622 90098 131674
rect 90110 131622 90162 131674
rect 90174 131622 90226 131674
rect 85580 131248 85632 131300
rect 88248 131248 88300 131300
rect 84936 131180 84988 131232
rect 85856 131180 85908 131232
rect 3982 131078 4034 131130
rect 4046 131078 4098 131130
rect 4110 131078 4162 131130
rect 4174 131078 4226 131130
rect 87982 131078 88034 131130
rect 88046 131078 88098 131130
rect 88110 131078 88162 131130
rect 88174 131078 88226 131130
rect 1982 130534 2034 130586
rect 2046 130534 2098 130586
rect 2110 130534 2162 130586
rect 2174 130534 2226 130586
rect 85982 130534 86034 130586
rect 86046 130534 86098 130586
rect 86110 130534 86162 130586
rect 86174 130534 86226 130586
rect 89982 130534 90034 130586
rect 90046 130534 90098 130586
rect 90110 130534 90162 130586
rect 90174 130534 90226 130586
rect 3982 129990 4034 130042
rect 4046 129990 4098 130042
rect 4110 129990 4162 130042
rect 4174 129990 4226 130042
rect 87982 129990 88034 130042
rect 88046 129990 88098 130042
rect 88110 129990 88162 130042
rect 88174 129990 88226 130042
rect 1982 129446 2034 129498
rect 2046 129446 2098 129498
rect 2110 129446 2162 129498
rect 2174 129446 2226 129498
rect 85982 129446 86034 129498
rect 86046 129446 86098 129498
rect 86110 129446 86162 129498
rect 86174 129446 86226 129498
rect 89982 129446 90034 129498
rect 90046 129446 90098 129498
rect 90110 129446 90162 129498
rect 90174 129446 90226 129498
rect 3982 128902 4034 128954
rect 4046 128902 4098 128954
rect 4110 128902 4162 128954
rect 4174 128902 4226 128954
rect 87982 128902 88034 128954
rect 88046 128902 88098 128954
rect 88110 128902 88162 128954
rect 88174 128902 88226 128954
rect 84016 128460 84068 128512
rect 88248 128460 88300 128512
rect 1982 128358 2034 128410
rect 2046 128358 2098 128410
rect 2110 128358 2162 128410
rect 2174 128358 2226 128410
rect 85982 128358 86034 128410
rect 86046 128358 86098 128410
rect 86110 128358 86162 128410
rect 86174 128358 86226 128410
rect 89982 128358 90034 128410
rect 90046 128358 90098 128410
rect 90110 128358 90162 128410
rect 90174 128358 90226 128410
rect 3982 127814 4034 127866
rect 4046 127814 4098 127866
rect 4110 127814 4162 127866
rect 4174 127814 4226 127866
rect 87982 127814 88034 127866
rect 88046 127814 88098 127866
rect 88110 127814 88162 127866
rect 88174 127814 88226 127866
rect 1982 127270 2034 127322
rect 2046 127270 2098 127322
rect 2110 127270 2162 127322
rect 2174 127270 2226 127322
rect 85982 127270 86034 127322
rect 86046 127270 86098 127322
rect 86110 127270 86162 127322
rect 86174 127270 86226 127322
rect 89982 127270 90034 127322
rect 90046 127270 90098 127322
rect 90110 127270 90162 127322
rect 90174 127270 90226 127322
rect 83372 126964 83424 127016
rect 88248 126964 88300 127016
rect 3982 126726 4034 126778
rect 4046 126726 4098 126778
rect 4110 126726 4162 126778
rect 4174 126726 4226 126778
rect 87982 126726 88034 126778
rect 88046 126726 88098 126778
rect 88110 126726 88162 126778
rect 88174 126726 88226 126778
rect 1982 126182 2034 126234
rect 2046 126182 2098 126234
rect 2110 126182 2162 126234
rect 2174 126182 2226 126234
rect 85982 126182 86034 126234
rect 86046 126182 86098 126234
rect 86110 126182 86162 126234
rect 86174 126182 86226 126234
rect 89982 126182 90034 126234
rect 90046 126182 90098 126234
rect 90110 126182 90162 126234
rect 90174 126182 90226 126234
rect 83280 125808 83332 125860
rect 87972 125808 88024 125860
rect 84568 125740 84620 125792
rect 3982 125638 4034 125690
rect 4046 125638 4098 125690
rect 4110 125638 4162 125690
rect 4174 125638 4226 125690
rect 87982 125638 88034 125690
rect 88046 125638 88098 125690
rect 88110 125638 88162 125690
rect 88174 125638 88226 125690
rect 1982 125094 2034 125146
rect 2046 125094 2098 125146
rect 2110 125094 2162 125146
rect 2174 125094 2226 125146
rect 85982 125094 86034 125146
rect 86046 125094 86098 125146
rect 86110 125094 86162 125146
rect 86174 125094 86226 125146
rect 89982 125094 90034 125146
rect 90046 125094 90098 125146
rect 90110 125094 90162 125146
rect 90174 125094 90226 125146
rect 3982 124550 4034 124602
rect 4046 124550 4098 124602
rect 4110 124550 4162 124602
rect 4174 124550 4226 124602
rect 87982 124550 88034 124602
rect 88046 124550 88098 124602
rect 88110 124550 88162 124602
rect 88174 124550 88226 124602
rect 84476 124448 84528 124500
rect 1982 124006 2034 124058
rect 2046 124006 2098 124058
rect 2110 124006 2162 124058
rect 2174 124006 2226 124058
rect 85982 124006 86034 124058
rect 86046 124006 86098 124058
rect 86110 124006 86162 124058
rect 86174 124006 86226 124058
rect 89982 124006 90034 124058
rect 90046 124006 90098 124058
rect 90110 124006 90162 124058
rect 90174 124006 90226 124058
rect 3982 123462 4034 123514
rect 4046 123462 4098 123514
rect 4110 123462 4162 123514
rect 4174 123462 4226 123514
rect 87982 123462 88034 123514
rect 88046 123462 88098 123514
rect 88110 123462 88162 123514
rect 88174 123462 88226 123514
rect 84384 123360 84436 123412
rect 1982 122918 2034 122970
rect 2046 122918 2098 122970
rect 2110 122918 2162 122970
rect 2174 122918 2226 122970
rect 85982 122918 86034 122970
rect 86046 122918 86098 122970
rect 86110 122918 86162 122970
rect 86174 122918 86226 122970
rect 89982 122918 90034 122970
rect 90046 122918 90098 122970
rect 90110 122918 90162 122970
rect 90174 122918 90226 122970
rect 83188 122816 83240 122868
rect 87972 122816 88024 122868
rect 3982 122374 4034 122426
rect 4046 122374 4098 122426
rect 4110 122374 4162 122426
rect 4174 122374 4226 122426
rect 87982 122374 88034 122426
rect 88046 122374 88098 122426
rect 88110 122374 88162 122426
rect 88174 122374 88226 122426
rect 87236 122136 87288 122188
rect 87880 122136 87932 122188
rect 1982 121830 2034 121882
rect 2046 121830 2098 121882
rect 2110 121830 2162 121882
rect 2174 121830 2226 121882
rect 85982 121830 86034 121882
rect 86046 121830 86098 121882
rect 86110 121830 86162 121882
rect 86174 121830 86226 121882
rect 89982 121830 90034 121882
rect 90046 121830 90098 121882
rect 90110 121830 90162 121882
rect 90174 121830 90226 121882
rect 83096 121456 83148 121508
rect 87880 121456 87932 121508
rect 3982 121286 4034 121338
rect 4046 121286 4098 121338
rect 4110 121286 4162 121338
rect 4174 121286 4226 121338
rect 87982 121286 88034 121338
rect 88046 121286 88098 121338
rect 88110 121286 88162 121338
rect 88174 121286 88226 121338
rect 84476 120844 84528 120896
rect 1982 120742 2034 120794
rect 2046 120742 2098 120794
rect 2110 120742 2162 120794
rect 2174 120742 2226 120794
rect 85982 120742 86034 120794
rect 86046 120742 86098 120794
rect 86110 120742 86162 120794
rect 86174 120742 86226 120794
rect 89982 120742 90034 120794
rect 90046 120742 90098 120794
rect 90110 120742 90162 120794
rect 90174 120742 90226 120794
rect 3982 120198 4034 120250
rect 4046 120198 4098 120250
rect 4110 120198 4162 120250
rect 4174 120198 4226 120250
rect 87982 120198 88034 120250
rect 88046 120198 88098 120250
rect 88110 120198 88162 120250
rect 88174 120198 88226 120250
rect 83004 120096 83056 120148
rect 87880 120096 87932 120148
rect 84568 120028 84620 120080
rect 1982 119654 2034 119706
rect 2046 119654 2098 119706
rect 2110 119654 2162 119706
rect 2174 119654 2226 119706
rect 85982 119654 86034 119706
rect 86046 119654 86098 119706
rect 86110 119654 86162 119706
rect 86174 119654 86226 119706
rect 89982 119654 90034 119706
rect 90046 119654 90098 119706
rect 90110 119654 90162 119706
rect 90174 119654 90226 119706
rect 3982 119110 4034 119162
rect 4046 119110 4098 119162
rect 4110 119110 4162 119162
rect 4174 119110 4226 119162
rect 87982 119110 88034 119162
rect 88046 119110 88098 119162
rect 88110 119110 88162 119162
rect 88174 119110 88226 119162
rect 82912 118668 82964 118720
rect 87880 118668 87932 118720
rect 1982 118566 2034 118618
rect 2046 118566 2098 118618
rect 2110 118566 2162 118618
rect 2174 118566 2226 118618
rect 85982 118566 86034 118618
rect 86046 118566 86098 118618
rect 86110 118566 86162 118618
rect 86174 118566 86226 118618
rect 89982 118566 90034 118618
rect 90046 118566 90098 118618
rect 90110 118566 90162 118618
rect 90174 118566 90226 118618
rect 84384 118124 84436 118176
rect 3982 118022 4034 118074
rect 4046 118022 4098 118074
rect 4110 118022 4162 118074
rect 4174 118022 4226 118074
rect 87982 118022 88034 118074
rect 88046 118022 88098 118074
rect 88110 118022 88162 118074
rect 88174 118022 88226 118074
rect 1982 117478 2034 117530
rect 2046 117478 2098 117530
rect 2110 117478 2162 117530
rect 2174 117478 2226 117530
rect 85982 117478 86034 117530
rect 86046 117478 86098 117530
rect 86110 117478 86162 117530
rect 86174 117478 86226 117530
rect 89982 117478 90034 117530
rect 90046 117478 90098 117530
rect 90110 117478 90162 117530
rect 90174 117478 90226 117530
rect 84568 117036 84620 117088
rect 3982 116934 4034 116986
rect 4046 116934 4098 116986
rect 4110 116934 4162 116986
rect 4174 116934 4226 116986
rect 87982 116934 88034 116986
rect 88046 116934 88098 116986
rect 88110 116934 88162 116986
rect 88174 116934 88226 116986
rect 5356 116560 5408 116612
rect 1982 116390 2034 116442
rect 2046 116390 2098 116442
rect 2110 116390 2162 116442
rect 2174 116390 2226 116442
rect 85982 116390 86034 116442
rect 86046 116390 86098 116442
rect 86110 116390 86162 116442
rect 86174 116390 86226 116442
rect 89982 116390 90034 116442
rect 90046 116390 90098 116442
rect 90110 116390 90162 116442
rect 90174 116390 90226 116442
rect 3982 115846 4034 115898
rect 4046 115846 4098 115898
rect 4110 115846 4162 115898
rect 4174 115846 4226 115898
rect 87982 115846 88034 115898
rect 88046 115846 88098 115898
rect 88110 115846 88162 115898
rect 88174 115846 88226 115898
rect 1982 115302 2034 115354
rect 2046 115302 2098 115354
rect 2110 115302 2162 115354
rect 2174 115302 2226 115354
rect 85982 115302 86034 115354
rect 86046 115302 86098 115354
rect 86110 115302 86162 115354
rect 86174 115302 86226 115354
rect 89982 115302 90034 115354
rect 90046 115302 90098 115354
rect 90110 115302 90162 115354
rect 90174 115302 90226 115354
rect 5448 114928 5500 114980
rect 3982 114758 4034 114810
rect 4046 114758 4098 114810
rect 4110 114758 4162 114810
rect 4174 114758 4226 114810
rect 87982 114758 88034 114810
rect 88046 114758 88098 114810
rect 88110 114758 88162 114810
rect 88174 114758 88226 114810
rect 85672 114520 85724 114572
rect 87972 114520 88024 114572
rect 1982 114214 2034 114266
rect 2046 114214 2098 114266
rect 2110 114214 2162 114266
rect 2174 114214 2226 114266
rect 85982 114214 86034 114266
rect 86046 114214 86098 114266
rect 86110 114214 86162 114266
rect 86174 114214 86226 114266
rect 89982 114214 90034 114266
rect 90046 114214 90098 114266
rect 90110 114214 90162 114266
rect 90174 114214 90226 114266
rect 85396 113840 85448 113892
rect 86500 113840 86552 113892
rect 3982 113670 4034 113722
rect 4046 113670 4098 113722
rect 4110 113670 4162 113722
rect 4174 113670 4226 113722
rect 87982 113670 88034 113722
rect 88046 113670 88098 113722
rect 88110 113670 88162 113722
rect 88174 113670 88226 113722
rect 1982 113126 2034 113178
rect 2046 113126 2098 113178
rect 2110 113126 2162 113178
rect 2174 113126 2226 113178
rect 85982 113126 86034 113178
rect 86046 113126 86098 113178
rect 86110 113126 86162 113178
rect 86174 113126 86226 113178
rect 89982 113126 90034 113178
rect 90046 113126 90098 113178
rect 90110 113126 90162 113178
rect 90174 113126 90226 113178
rect 3982 112582 4034 112634
rect 4046 112582 4098 112634
rect 4110 112582 4162 112634
rect 4174 112582 4226 112634
rect 87982 112582 88034 112634
rect 88046 112582 88098 112634
rect 88110 112582 88162 112634
rect 88174 112582 88226 112634
rect 1982 112038 2034 112090
rect 2046 112038 2098 112090
rect 2110 112038 2162 112090
rect 2174 112038 2226 112090
rect 85982 112038 86034 112090
rect 86046 112038 86098 112090
rect 86110 112038 86162 112090
rect 86174 112038 86226 112090
rect 89982 112038 90034 112090
rect 90046 112038 90098 112090
rect 90110 112038 90162 112090
rect 90174 112038 90226 112090
rect 85304 111800 85356 111852
rect 87972 111800 88024 111852
rect 3982 111494 4034 111546
rect 4046 111494 4098 111546
rect 4110 111494 4162 111546
rect 4174 111494 4226 111546
rect 87982 111494 88034 111546
rect 88046 111494 88098 111546
rect 88110 111494 88162 111546
rect 88174 111494 88226 111546
rect 1982 110950 2034 111002
rect 2046 110950 2098 111002
rect 2110 110950 2162 111002
rect 2174 110950 2226 111002
rect 85982 110950 86034 111002
rect 86046 110950 86098 111002
rect 86110 110950 86162 111002
rect 86174 110950 86226 111002
rect 89982 110950 90034 111002
rect 90046 110950 90098 111002
rect 90110 110950 90162 111002
rect 90174 110950 90226 111002
rect 3982 110406 4034 110458
rect 4046 110406 4098 110458
rect 4110 110406 4162 110458
rect 4174 110406 4226 110458
rect 87982 110406 88034 110458
rect 88046 110406 88098 110458
rect 88110 110406 88162 110458
rect 88174 110406 88226 110458
rect 82544 110304 82596 110356
rect 85488 110304 85540 110356
rect 1982 109862 2034 109914
rect 2046 109862 2098 109914
rect 2110 109862 2162 109914
rect 2174 109862 2226 109914
rect 85982 109862 86034 109914
rect 86046 109862 86098 109914
rect 86110 109862 86162 109914
rect 86174 109862 86226 109914
rect 89982 109862 90034 109914
rect 90046 109862 90098 109914
rect 90110 109862 90162 109914
rect 90174 109862 90226 109914
rect 85212 109556 85264 109608
rect 85856 109556 85908 109608
rect 3982 109318 4034 109370
rect 4046 109318 4098 109370
rect 4110 109318 4162 109370
rect 4174 109318 4226 109370
rect 87982 109318 88034 109370
rect 88046 109318 88098 109370
rect 88110 109318 88162 109370
rect 88174 109318 88226 109370
rect 84292 108944 84344 108996
rect 85948 108944 86000 108996
rect 1982 108774 2034 108826
rect 2046 108774 2098 108826
rect 2110 108774 2162 108826
rect 2174 108774 2226 108826
rect 85982 108774 86034 108826
rect 86046 108774 86098 108826
rect 86110 108774 86162 108826
rect 86174 108774 86226 108826
rect 89982 108774 90034 108826
rect 90046 108774 90098 108826
rect 90110 108774 90162 108826
rect 90174 108774 90226 108826
rect 85212 108604 85264 108656
rect 87972 108604 88024 108656
rect 87604 108536 87656 108588
rect 88340 108536 88392 108588
rect 87236 108468 87288 108520
rect 88524 108468 88576 108520
rect 87604 108400 87656 108452
rect 88248 108400 88300 108452
rect 3982 108230 4034 108282
rect 4046 108230 4098 108282
rect 4110 108230 4162 108282
rect 4174 108230 4226 108282
rect 87982 108230 88034 108282
rect 88046 108230 88098 108282
rect 88110 108230 88162 108282
rect 88174 108230 88226 108282
rect 1982 107686 2034 107738
rect 2046 107686 2098 107738
rect 2110 107686 2162 107738
rect 2174 107686 2226 107738
rect 85982 107686 86034 107738
rect 86046 107686 86098 107738
rect 86110 107686 86162 107738
rect 86174 107686 86226 107738
rect 89982 107686 90034 107738
rect 90046 107686 90098 107738
rect 90110 107686 90162 107738
rect 90174 107686 90226 107738
rect 83648 107312 83700 107364
rect 87972 107312 88024 107364
rect 3982 107142 4034 107194
rect 4046 107142 4098 107194
rect 4110 107142 4162 107194
rect 4174 107142 4226 107194
rect 87982 107142 88034 107194
rect 88046 107142 88098 107194
rect 88110 107142 88162 107194
rect 88174 107142 88226 107194
rect 1982 106598 2034 106650
rect 2046 106598 2098 106650
rect 2110 106598 2162 106650
rect 2174 106598 2226 106650
rect 85982 106598 86034 106650
rect 86046 106598 86098 106650
rect 86110 106598 86162 106650
rect 86174 106598 86226 106650
rect 89982 106598 90034 106650
rect 90046 106598 90098 106650
rect 90110 106598 90162 106650
rect 90174 106598 90226 106650
rect 86316 106496 86368 106548
rect 86316 106292 86368 106344
rect 3982 106054 4034 106106
rect 4046 106054 4098 106106
rect 4110 106054 4162 106106
rect 4174 106054 4226 106106
rect 87982 106054 88034 106106
rect 88046 106054 88098 106106
rect 88110 106054 88162 106106
rect 88174 106054 88226 106106
rect 4436 105859 4488 105868
rect 4436 105825 4445 105859
rect 4445 105825 4479 105859
rect 4479 105825 4488 105859
rect 4436 105816 4488 105825
rect 86224 105680 86276 105732
rect 1982 105510 2034 105562
rect 2046 105510 2098 105562
rect 2110 105510 2162 105562
rect 2174 105510 2226 105562
rect 85982 105510 86034 105562
rect 86046 105510 86098 105562
rect 86110 105510 86162 105562
rect 86174 105510 86226 105562
rect 89982 105510 90034 105562
rect 90046 105510 90098 105562
rect 90110 105510 90162 105562
rect 90174 105510 90226 105562
rect 3982 104966 4034 105018
rect 4046 104966 4098 105018
rect 4110 104966 4162 105018
rect 4174 104966 4226 105018
rect 87982 104966 88034 105018
rect 88046 104966 88098 105018
rect 88110 104966 88162 105018
rect 88174 104966 88226 105018
rect 85488 104524 85540 104576
rect 86408 104524 86460 104576
rect 86500 104524 86552 104576
rect 86684 104524 86736 104576
rect 1982 104422 2034 104474
rect 2046 104422 2098 104474
rect 2110 104422 2162 104474
rect 2174 104422 2226 104474
rect 85982 104422 86034 104474
rect 86046 104422 86098 104474
rect 86110 104422 86162 104474
rect 86174 104422 86226 104474
rect 89982 104422 90034 104474
rect 90046 104422 90098 104474
rect 90110 104422 90162 104474
rect 90174 104422 90226 104474
rect 86868 104320 86920 104372
rect 85672 104252 85724 104304
rect 86592 104184 86644 104236
rect 86868 104184 86920 104236
rect 87328 104320 87380 104372
rect 87788 104320 87840 104372
rect 88708 104320 88760 104372
rect 87144 104116 87196 104168
rect 3982 103878 4034 103930
rect 4046 103878 4098 103930
rect 4110 103878 4162 103930
rect 4174 103878 4226 103930
rect 87982 103878 88034 103930
rect 88046 103878 88098 103930
rect 88110 103878 88162 103930
rect 88174 103878 88226 103930
rect 1982 103334 2034 103386
rect 2046 103334 2098 103386
rect 2110 103334 2162 103386
rect 2174 103334 2226 103386
rect 85982 103334 86034 103386
rect 86046 103334 86098 103386
rect 86110 103334 86162 103386
rect 86174 103334 86226 103386
rect 89982 103334 90034 103386
rect 90046 103334 90098 103386
rect 90110 103334 90162 103386
rect 90174 103334 90226 103386
rect 3982 102790 4034 102842
rect 4046 102790 4098 102842
rect 4110 102790 4162 102842
rect 4174 102790 4226 102842
rect 87982 102790 88034 102842
rect 88046 102790 88098 102842
rect 88110 102790 88162 102842
rect 88174 102790 88226 102842
rect 1982 102246 2034 102298
rect 2046 102246 2098 102298
rect 2110 102246 2162 102298
rect 2174 102246 2226 102298
rect 85982 102246 86034 102298
rect 86046 102246 86098 102298
rect 86110 102246 86162 102298
rect 86174 102246 86226 102298
rect 89982 102246 90034 102298
rect 90046 102246 90098 102298
rect 90110 102246 90162 102298
rect 90174 102246 90226 102298
rect 3982 101702 4034 101754
rect 4046 101702 4098 101754
rect 4110 101702 4162 101754
rect 4174 101702 4226 101754
rect 87982 101702 88034 101754
rect 88046 101702 88098 101754
rect 88110 101702 88162 101754
rect 88174 101702 88226 101754
rect 1982 101158 2034 101210
rect 2046 101158 2098 101210
rect 2110 101158 2162 101210
rect 2174 101158 2226 101210
rect 85982 101158 86034 101210
rect 86046 101158 86098 101210
rect 86110 101158 86162 101210
rect 86174 101158 86226 101210
rect 89982 101158 90034 101210
rect 90046 101158 90098 101210
rect 90110 101158 90162 101210
rect 90174 101158 90226 101210
rect 87880 101056 87932 101108
rect 88432 101056 88484 101108
rect 3982 100614 4034 100666
rect 4046 100614 4098 100666
rect 4110 100614 4162 100666
rect 4174 100614 4226 100666
rect 87982 100614 88034 100666
rect 88046 100614 88098 100666
rect 88110 100614 88162 100666
rect 88174 100614 88226 100666
rect 1982 100070 2034 100122
rect 2046 100070 2098 100122
rect 2110 100070 2162 100122
rect 2174 100070 2226 100122
rect 85982 100070 86034 100122
rect 86046 100070 86098 100122
rect 86110 100070 86162 100122
rect 86174 100070 86226 100122
rect 89982 100070 90034 100122
rect 90046 100070 90098 100122
rect 90110 100070 90162 100122
rect 90174 100070 90226 100122
rect 85764 99968 85816 100020
rect 86408 99968 86460 100020
rect 86132 99900 86184 99952
rect 86684 99900 86736 99952
rect 87236 99900 87288 99952
rect 88616 99900 88668 99952
rect 85856 99832 85908 99884
rect 86224 99832 86276 99884
rect 87604 99832 87656 99884
rect 88432 99832 88484 99884
rect 88524 99764 88576 99816
rect 87604 99696 87656 99748
rect 87880 99696 87932 99748
rect 85028 99628 85080 99680
rect 85396 99628 85448 99680
rect 85488 99628 85540 99680
rect 85672 99628 85724 99680
rect 86868 99628 86920 99680
rect 3982 99526 4034 99578
rect 4046 99526 4098 99578
rect 4110 99526 4162 99578
rect 4174 99526 4226 99578
rect 87982 99526 88034 99578
rect 88046 99526 88098 99578
rect 88110 99526 88162 99578
rect 88174 99526 88226 99578
rect 85396 99424 85448 99476
rect 86500 99424 86552 99476
rect 85580 99356 85632 99408
rect 86132 99356 86184 99408
rect 82728 99288 82780 99340
rect 87420 99288 87472 99340
rect 85396 99220 85448 99272
rect 85856 99220 85908 99272
rect 87512 99220 87564 99272
rect 87420 99152 87472 99204
rect 88432 99152 88484 99204
rect 87512 99084 87564 99136
rect 88616 99084 88668 99136
rect 1982 98982 2034 99034
rect 2046 98982 2098 99034
rect 2110 98982 2162 99034
rect 2174 98982 2226 99034
rect 85982 98982 86034 99034
rect 86046 98982 86098 99034
rect 86110 98982 86162 99034
rect 86174 98982 86226 99034
rect 89982 98982 90034 99034
rect 90046 98982 90098 99034
rect 90110 98982 90162 99034
rect 90174 98982 90226 99034
rect 87604 98880 87656 98932
rect 87696 98880 87748 98932
rect 87880 98880 87932 98932
rect 87788 98676 87840 98728
rect 88340 98676 88392 98728
rect 4344 98583 4396 98592
rect 4344 98549 4353 98583
rect 4353 98549 4387 98583
rect 4387 98549 4396 98583
rect 4344 98540 4396 98549
rect 6736 98540 6788 98592
rect 3982 98438 4034 98490
rect 4046 98438 4098 98490
rect 4110 98438 4162 98490
rect 4174 98438 4226 98490
rect 87982 98438 88034 98490
rect 88046 98438 88098 98490
rect 88110 98438 88162 98490
rect 88174 98438 88226 98490
rect 82728 98311 82780 98320
rect 82728 98277 82737 98311
rect 82737 98277 82771 98311
rect 82771 98277 82780 98311
rect 82728 98268 82780 98277
rect 82728 98132 82780 98184
rect 87236 98132 87288 98184
rect 6828 98064 6880 98116
rect 83464 98064 83516 98116
rect 86960 98064 87012 98116
rect 4436 98039 4488 98048
rect 4436 98005 4445 98039
rect 4445 98005 4479 98039
rect 4479 98005 4488 98039
rect 4436 97996 4488 98005
rect 4528 97996 4580 98048
rect 5356 97996 5408 98048
rect 84936 97996 84988 98048
rect 1982 97894 2034 97946
rect 2046 97894 2098 97946
rect 2110 97894 2162 97946
rect 2174 97894 2226 97946
rect 85982 97894 86034 97946
rect 86046 97894 86098 97946
rect 86110 97894 86162 97946
rect 86174 97894 86226 97946
rect 89982 97894 90034 97946
rect 90046 97894 90098 97946
rect 90110 97894 90162 97946
rect 90174 97894 90226 97946
rect 2596 97792 2648 97844
rect 84844 97835 84896 97844
rect 84844 97801 84853 97835
rect 84853 97801 84887 97835
rect 84887 97801 84896 97835
rect 84844 97792 84896 97801
rect 85396 97792 85448 97844
rect 5816 97724 5868 97776
rect 5724 97656 5776 97708
rect 87880 97656 87932 97708
rect 90364 97656 90416 97708
rect 87972 97588 88024 97640
rect 3332 97495 3384 97504
rect 3332 97461 3341 97495
rect 3341 97461 3375 97495
rect 3375 97461 3384 97495
rect 3332 97452 3384 97461
rect 5632 97452 5684 97504
rect 3982 97350 4034 97402
rect 4046 97350 4098 97402
rect 4110 97350 4162 97402
rect 4174 97350 4226 97402
rect 2596 97291 2648 97300
rect 2596 97257 2605 97291
rect 2605 97257 2639 97291
rect 2639 97257 2648 97291
rect 2596 97248 2648 97257
rect 5908 97248 5960 97300
rect 3608 97180 3660 97232
rect 87696 97520 87748 97572
rect 84292 97452 84344 97504
rect 84844 97495 84896 97504
rect 84844 97461 84853 97495
rect 84853 97461 84887 97495
rect 84887 97461 84896 97495
rect 84844 97452 84896 97461
rect 6736 97316 6788 97368
rect 83464 97316 83516 97368
rect 87982 97350 88034 97402
rect 88046 97350 88098 97402
rect 88110 97350 88162 97402
rect 88174 97350 88226 97402
rect 22928 97248 22980 97300
rect 84752 97248 84804 97300
rect 86960 97248 87012 97300
rect 21916 97180 21968 97232
rect 86776 97180 86828 97232
rect 5080 97112 5132 97164
rect 86960 97112 87012 97164
rect 5540 97044 5592 97096
rect 18052 97044 18104 97096
rect 83648 97044 83700 97096
rect 86408 97044 86460 97096
rect 86776 97044 86828 97096
rect 87144 97044 87196 97096
rect 14648 96976 14700 97028
rect 17132 96976 17184 97028
rect 22652 96976 22704 97028
rect 85304 96976 85356 97028
rect 2964 96951 3016 96960
rect 2964 96917 2973 96951
rect 2973 96917 3007 96951
rect 3007 96917 3016 96951
rect 2964 96908 3016 96917
rect 6460 96908 6512 96960
rect 33140 96908 33192 96960
rect 83188 96908 83240 96960
rect 83464 96908 83516 96960
rect 84292 96908 84344 96960
rect 84936 96908 84988 96960
rect 1982 96806 2034 96858
rect 2046 96806 2098 96858
rect 2110 96806 2162 96858
rect 2174 96806 2226 96858
rect 5632 96840 5684 96892
rect 30104 96840 30156 96892
rect 82912 96840 82964 96892
rect 83648 96883 83700 96892
rect 83648 96849 83657 96883
rect 83657 96849 83691 96883
rect 83691 96849 83700 96883
rect 83648 96840 83700 96849
rect 6276 96772 6328 96824
rect 32036 96772 32088 96824
rect 83096 96772 83148 96824
rect 83280 96772 83332 96824
rect 85982 96806 86034 96858
rect 86046 96806 86098 96858
rect 86110 96806 86162 96858
rect 86174 96806 86226 96858
rect 89982 96806 90034 96858
rect 90046 96806 90098 96858
rect 90110 96806 90162 96858
rect 90174 96806 90226 96858
rect 3332 96704 3384 96756
rect 24308 96704 24360 96756
rect 2964 96636 3016 96688
rect 3424 96636 3476 96688
rect 22100 96636 22152 96688
rect 22928 96636 22980 96688
rect 25412 96636 25464 96688
rect 76932 96704 76984 96756
rect 80060 96704 80112 96756
rect 85580 96636 85632 96688
rect 85948 96636 86000 96688
rect 86408 96636 86460 96688
rect 5448 96568 5500 96620
rect 87052 96568 87104 96620
rect 4620 96500 4672 96552
rect 39580 96500 39632 96552
rect 62304 96500 62356 96552
rect 16488 96432 16540 96484
rect 85764 96500 85816 96552
rect 76656 96432 76708 96484
rect 82176 96432 82228 96484
rect 82820 96432 82872 96484
rect 3332 96407 3384 96416
rect 3332 96373 3341 96407
rect 3341 96373 3375 96407
rect 3375 96373 3384 96407
rect 3332 96364 3384 96373
rect 3700 96407 3752 96416
rect 3700 96373 3709 96407
rect 3709 96373 3743 96407
rect 3743 96373 3752 96407
rect 3700 96364 3752 96373
rect 5908 96364 5960 96416
rect 29184 96364 29236 96416
rect 88984 96432 89036 96484
rect 84844 96364 84896 96416
rect 85120 96407 85172 96416
rect 85120 96373 85129 96407
rect 85129 96373 85163 96407
rect 85163 96373 85172 96407
rect 85120 96364 85172 96373
rect 85396 96364 85448 96416
rect 3982 96262 4034 96314
rect 4046 96262 4098 96314
rect 4110 96262 4162 96314
rect 4174 96262 4226 96314
rect 15752 96296 15804 96348
rect 82728 96296 82780 96348
rect 37832 96228 37884 96280
rect 41144 96228 41196 96280
rect 59360 96228 59412 96280
rect 9588 96160 9640 96212
rect 50344 96160 50396 96212
rect 51172 96160 51224 96212
rect 57612 96160 57664 96212
rect 60648 96228 60700 96280
rect 61568 96228 61620 96280
rect 59544 96160 59596 96212
rect 87982 96262 88034 96314
rect 88046 96262 88098 96314
rect 88110 96262 88162 96314
rect 88174 96262 88226 96314
rect 75184 96160 75236 96212
rect 84752 96160 84804 96212
rect 3332 96092 3384 96144
rect 6092 96092 6144 96144
rect 27988 96092 28040 96144
rect 28908 96092 28960 96144
rect 59728 96092 59780 96144
rect 74632 96092 74684 96144
rect 80152 96092 80204 96144
rect 82360 96092 82412 96144
rect 57888 96024 57940 96076
rect 85856 96024 85908 96076
rect 6920 95956 6972 96008
rect 41972 95956 42024 96008
rect 54576 95956 54628 96008
rect 76840 95956 76892 96008
rect 79692 95956 79744 96008
rect 79784 95956 79836 96008
rect 80336 95956 80388 96008
rect 87236 95956 87288 96008
rect 4896 95888 4948 95940
rect 5448 95888 5500 95940
rect 86960 95888 87012 95940
rect 5816 95820 5868 95872
rect 52184 95820 52236 95872
rect 82728 95820 82780 95872
rect 85028 95820 85080 95872
rect 85488 95820 85540 95872
rect 1982 95718 2034 95770
rect 2046 95718 2098 95770
rect 2110 95718 2162 95770
rect 2174 95718 2226 95770
rect 15752 95752 15804 95804
rect 24584 95752 24636 95804
rect 62028 95752 62080 95804
rect 62120 95752 62172 95804
rect 34980 95684 35032 95736
rect 31484 95616 31536 95668
rect 83004 95616 83056 95668
rect 85982 95718 86034 95770
rect 86046 95718 86098 95770
rect 86110 95718 86162 95770
rect 86174 95718 86226 95770
rect 89982 95718 90034 95770
rect 90046 95718 90098 95770
rect 90110 95718 90162 95770
rect 90174 95718 90226 95770
rect 87512 95616 87564 95668
rect 6828 95548 6880 95600
rect 16488 95548 16540 95600
rect 27528 95548 27580 95600
rect 83188 95548 83240 95600
rect 6552 95480 6604 95532
rect 38476 95480 38528 95532
rect 58072 95480 58124 95532
rect 28908 95412 28960 95464
rect 80152 95412 80204 95464
rect 83832 95412 83884 95464
rect 3700 95344 3752 95396
rect 3884 95344 3936 95396
rect 20996 95344 21048 95396
rect 5356 95276 5408 95328
rect 26792 95276 26844 95328
rect 27528 95276 27580 95328
rect 64144 95276 64196 95328
rect 3982 95174 4034 95226
rect 4046 95174 4098 95226
rect 4110 95174 4162 95226
rect 4174 95174 4226 95226
rect 45376 95208 45428 95260
rect 49516 95208 49568 95260
rect 49608 95208 49660 95260
rect 64788 95208 64840 95260
rect 24768 95140 24820 95192
rect 79876 95208 79928 95260
rect 83004 95344 83056 95396
rect 83280 95276 83332 95328
rect 80152 95140 80204 95192
rect 83096 95208 83148 95260
rect 87420 95276 87472 95328
rect 83372 95140 83424 95192
rect 83556 95140 83608 95192
rect 87982 95174 88034 95226
rect 88046 95174 88098 95226
rect 88110 95174 88162 95226
rect 88174 95174 88226 95226
rect 19340 95072 19392 95124
rect 85212 95072 85264 95124
rect 25964 95004 26016 95056
rect 82544 95004 82596 95056
rect 4344 94936 4396 94988
rect 29184 94936 29236 94988
rect 30288 94936 30340 94988
rect 80152 94936 80204 94988
rect 31668 94868 31720 94920
rect 74540 94868 74592 94920
rect 80244 94868 80296 94920
rect 80428 94936 80480 94988
rect 85856 94936 85908 94988
rect 86868 94936 86920 94988
rect 82820 94868 82872 94920
rect 83648 94868 83700 94920
rect 20628 94800 20680 94852
rect 44180 94800 44232 94852
rect 45192 94800 45244 94852
rect 78220 94800 78272 94852
rect 86316 94800 86368 94852
rect 86868 94800 86920 94852
rect 4436 94732 4488 94784
rect 19340 94732 19392 94784
rect 45560 94732 45612 94784
rect 76104 94732 76156 94784
rect 80612 94732 80664 94784
rect 82360 94732 82412 94784
rect 85764 94732 85816 94784
rect 1982 94630 2034 94682
rect 2046 94630 2098 94682
rect 2110 94630 2162 94682
rect 2174 94630 2226 94682
rect 38568 94664 38620 94716
rect 46848 94664 46900 94716
rect 47952 94664 48004 94716
rect 6460 94596 6512 94648
rect 12808 94596 12860 94648
rect 13728 94596 13780 94648
rect 23388 94596 23440 94648
rect 48228 94596 48280 94648
rect 49884 94596 49936 94648
rect 50804 94596 50856 94648
rect 52552 94596 52604 94648
rect 80244 94664 80296 94716
rect 80520 94664 80572 94716
rect 83556 94664 83608 94716
rect 83924 94596 83976 94648
rect 85982 94630 86034 94682
rect 86046 94630 86098 94682
rect 86110 94630 86162 94682
rect 86174 94630 86226 94682
rect 89982 94630 90034 94682
rect 90046 94630 90098 94682
rect 90110 94630 90162 94682
rect 90174 94630 90226 94682
rect 4528 94528 4580 94580
rect 37280 94528 37332 94580
rect 46664 94528 46716 94580
rect 74540 94528 74592 94580
rect 74632 94528 74684 94580
rect 80428 94528 80480 94580
rect 85488 94528 85540 94580
rect 4896 94460 4948 94512
rect 86960 94460 87012 94512
rect 49976 94392 50028 94444
rect 51448 94324 51500 94376
rect 74816 94392 74868 94444
rect 85396 94392 85448 94444
rect 45100 94256 45152 94308
rect 53748 94256 53800 94308
rect 54024 94256 54076 94308
rect 85304 94324 85356 94376
rect 83372 94256 83424 94308
rect 83464 94256 83516 94308
rect 84844 94256 84896 94308
rect 4436 94188 4488 94240
rect 5264 94188 5316 94240
rect 44088 94188 44140 94240
rect 54852 94188 54904 94240
rect 54944 94188 54996 94240
rect 3982 94086 4034 94138
rect 4046 94086 4098 94138
rect 4110 94086 4162 94138
rect 4174 94086 4226 94138
rect 42708 94120 42760 94172
rect 48136 94120 48188 94172
rect 50988 94120 51040 94172
rect 53288 94120 53340 94172
rect 59912 94120 59964 94172
rect 62028 94120 62080 94172
rect 87512 94188 87564 94240
rect 79232 94120 79284 94172
rect 81440 94120 81492 94172
rect 61936 94052 61988 94104
rect 62304 94052 62356 94104
rect 83464 94120 83516 94172
rect 87982 94086 88034 94138
rect 88046 94086 88098 94138
rect 88110 94086 88162 94138
rect 88174 94086 88226 94138
rect 49056 93984 49108 94036
rect 87788 93984 87840 94036
rect 13728 93916 13780 93968
rect 84936 93916 84988 93968
rect 86592 93916 86644 93968
rect 87604 93916 87656 93968
rect 4528 93848 4580 93900
rect 9588 93848 9640 93900
rect 85304 93848 85356 93900
rect 50620 93780 50672 93832
rect 87696 93780 87748 93832
rect 49516 93712 49568 93764
rect 86960 93712 87012 93764
rect 4528 93644 4580 93696
rect 79416 93644 79468 93696
rect 82912 93644 82964 93696
rect 1982 93542 2034 93594
rect 2046 93542 2098 93594
rect 2110 93542 2162 93594
rect 2174 93542 2226 93594
rect 48780 93576 48832 93628
rect 54208 93576 54260 93628
rect 64788 93576 64840 93628
rect 87236 93644 87288 93696
rect 83464 93619 83516 93628
rect 83464 93585 83473 93619
rect 83473 93585 83507 93619
rect 83507 93585 83516 93619
rect 83464 93576 83516 93585
rect 59360 93508 59412 93560
rect 51264 93440 51316 93492
rect 84016 93508 84068 93560
rect 85982 93542 86034 93594
rect 86046 93542 86098 93594
rect 86110 93542 86162 93594
rect 86174 93542 86226 93594
rect 89982 93542 90034 93594
rect 90046 93542 90098 93594
rect 90110 93542 90162 93594
rect 90174 93542 90226 93594
rect 87328 93440 87380 93492
rect 53748 93372 53800 93424
rect 77300 93372 77352 93424
rect 47952 93304 48004 93356
rect 84568 93372 84620 93424
rect 84752 93415 84804 93424
rect 84752 93381 84761 93415
rect 84761 93381 84795 93415
rect 84795 93381 84804 93415
rect 84752 93372 84804 93381
rect 85120 93415 85172 93424
rect 85120 93381 85129 93415
rect 85129 93381 85163 93415
rect 85163 93381 85172 93415
rect 85120 93372 85172 93381
rect 82452 93304 82504 93356
rect 82820 93347 82872 93356
rect 82820 93313 82829 93347
rect 82829 93313 82863 93347
rect 82863 93313 82872 93347
rect 82820 93304 82872 93313
rect 46664 93236 46716 93288
rect 77484 93236 77536 93288
rect 79508 93236 79560 93288
rect 84108 93236 84160 93288
rect 44088 93168 44140 93220
rect 83740 93168 83792 93220
rect 42616 93100 42668 93152
rect 84200 93100 84252 93152
rect 3982 92998 4034 93050
rect 4046 92998 4098 93050
rect 4110 92998 4162 93050
rect 4174 92998 4226 93050
rect 39948 93032 40000 93084
rect 38384 92964 38436 93016
rect 35256 92896 35308 92948
rect 83924 92964 83976 93016
rect 87982 92998 88034 93050
rect 88046 92998 88098 93050
rect 88110 92998 88162 93050
rect 88174 92998 88226 93050
rect 84292 92896 84344 92948
rect 36728 92828 36780 92880
rect 84752 92828 84804 92880
rect 32864 92760 32916 92812
rect 34152 92760 34204 92812
rect 84844 92692 84896 92744
rect 85212 92692 85264 92744
rect 87420 92624 87472 92676
rect 1982 92454 2034 92506
rect 2046 92454 2098 92506
rect 2110 92454 2162 92506
rect 2174 92454 2226 92506
rect 85982 92454 86034 92506
rect 86046 92454 86098 92506
rect 86110 92454 86162 92506
rect 86174 92454 86226 92506
rect 89982 92454 90034 92506
rect 90046 92454 90098 92506
rect 90110 92454 90162 92506
rect 90174 92454 90226 92506
rect 87052 92352 87104 92404
rect 87144 92284 87196 92336
rect 82820 92216 82872 92268
rect 87512 92216 87564 92268
rect 82820 92123 82872 92132
rect 82820 92089 82829 92123
rect 82829 92089 82863 92123
rect 82863 92089 82872 92123
rect 82820 92080 82872 92089
rect 85580 92012 85632 92064
rect 86776 92012 86828 92064
rect 3982 91910 4034 91962
rect 4046 91910 4098 91962
rect 4110 91910 4162 91962
rect 4174 91910 4226 91962
rect 87982 91910 88034 91962
rect 88046 91910 88098 91962
rect 88110 91910 88162 91962
rect 88174 91910 88226 91962
rect 88340 91740 88392 91792
rect 1982 91366 2034 91418
rect 2046 91366 2098 91418
rect 2110 91366 2162 91418
rect 2174 91366 2226 91418
rect 85982 91366 86034 91418
rect 86046 91366 86098 91418
rect 86110 91366 86162 91418
rect 86174 91366 86226 91418
rect 89982 91366 90034 91418
rect 90046 91366 90098 91418
rect 90110 91366 90162 91418
rect 90174 91366 90226 91418
rect 3982 90822 4034 90874
rect 4046 90822 4098 90874
rect 4110 90822 4162 90874
rect 4174 90822 4226 90874
rect 87982 90822 88034 90874
rect 88046 90822 88098 90874
rect 88110 90822 88162 90874
rect 88174 90822 88226 90874
rect 86408 90720 86460 90772
rect 86684 90720 86736 90772
rect 4896 90652 4948 90704
rect 5448 90652 5500 90704
rect 4344 90516 4396 90568
rect 5448 90516 5500 90568
rect 4344 90380 4396 90432
rect 1982 90278 2034 90330
rect 2046 90278 2098 90330
rect 2110 90278 2162 90330
rect 2174 90278 2226 90330
rect 85982 90278 86034 90330
rect 86046 90278 86098 90330
rect 86110 90278 86162 90330
rect 86174 90278 86226 90330
rect 89982 90278 90034 90330
rect 90046 90278 90098 90330
rect 90110 90278 90162 90330
rect 90174 90278 90226 90330
rect 86684 90040 86736 90092
rect 86960 90040 87012 90092
rect 3982 89734 4034 89786
rect 4046 89734 4098 89786
rect 4110 89734 4162 89786
rect 4174 89734 4226 89786
rect 87982 89734 88034 89786
rect 88046 89734 88098 89786
rect 88110 89734 88162 89786
rect 88174 89734 88226 89786
rect 86868 89632 86920 89684
rect 87512 89632 87564 89684
rect 88340 89632 88392 89684
rect 86684 89428 86736 89480
rect 5080 89360 5132 89412
rect 1982 89190 2034 89242
rect 2046 89190 2098 89242
rect 2110 89190 2162 89242
rect 2174 89190 2226 89242
rect 4804 89063 4856 89072
rect 4804 89029 4813 89063
rect 4813 89029 4847 89063
rect 4847 89029 4856 89063
rect 85982 89190 86034 89242
rect 86046 89190 86098 89242
rect 86110 89190 86162 89242
rect 86174 89190 86226 89242
rect 89982 89190 90034 89242
rect 90046 89190 90098 89242
rect 90110 89190 90162 89242
rect 90174 89190 90226 89242
rect 4804 89020 4856 89029
rect 4344 88952 4396 89004
rect 4896 88952 4948 89004
rect 4344 88816 4396 88868
rect 5264 88816 5316 88868
rect 3982 88646 4034 88698
rect 4046 88646 4098 88698
rect 4110 88646 4162 88698
rect 4174 88646 4226 88698
rect 87982 88646 88034 88698
rect 88046 88646 88098 88698
rect 88110 88646 88162 88698
rect 88174 88646 88226 88698
rect 84936 88272 84988 88324
rect 87972 88272 88024 88324
rect 1982 88102 2034 88154
rect 2046 88102 2098 88154
rect 2110 88102 2162 88154
rect 2174 88102 2226 88154
rect 85982 88102 86034 88154
rect 86046 88102 86098 88154
rect 86110 88102 86162 88154
rect 86174 88102 86226 88154
rect 89982 88102 90034 88154
rect 90046 88102 90098 88154
rect 90110 88102 90162 88154
rect 90174 88102 90226 88154
rect 4988 88000 5040 88052
rect 3982 87558 4034 87610
rect 4046 87558 4098 87610
rect 4110 87558 4162 87610
rect 4174 87558 4226 87610
rect 87982 87558 88034 87610
rect 88046 87558 88098 87610
rect 88110 87558 88162 87610
rect 88174 87558 88226 87610
rect 1982 87014 2034 87066
rect 2046 87014 2098 87066
rect 2110 87014 2162 87066
rect 2174 87014 2226 87066
rect 85982 87014 86034 87066
rect 86046 87014 86098 87066
rect 86110 87014 86162 87066
rect 86174 87014 86226 87066
rect 89982 87014 90034 87066
rect 90046 87014 90098 87066
rect 90110 87014 90162 87066
rect 90174 87014 90226 87066
rect 3982 86470 4034 86522
rect 4046 86470 4098 86522
rect 4110 86470 4162 86522
rect 4174 86470 4226 86522
rect 87982 86470 88034 86522
rect 88046 86470 88098 86522
rect 88110 86470 88162 86522
rect 88174 86470 88226 86522
rect 5172 86368 5224 86420
rect 83004 86300 83056 86352
rect 87972 86300 88024 86352
rect 1982 85926 2034 85978
rect 2046 85926 2098 85978
rect 2110 85926 2162 85978
rect 2174 85926 2226 85978
rect 85982 85926 86034 85978
rect 86046 85926 86098 85978
rect 86110 85926 86162 85978
rect 86174 85926 86226 85978
rect 89982 85926 90034 85978
rect 90046 85926 90098 85978
rect 90110 85926 90162 85978
rect 90174 85926 90226 85978
rect 3982 85382 4034 85434
rect 4046 85382 4098 85434
rect 4110 85382 4162 85434
rect 4174 85382 4226 85434
rect 87982 85382 88034 85434
rect 88046 85382 88098 85434
rect 88110 85382 88162 85434
rect 88174 85382 88226 85434
rect 4712 85323 4764 85332
rect 4712 85289 4721 85323
rect 4721 85289 4755 85323
rect 4755 85289 4764 85323
rect 4712 85280 4764 85289
rect 83832 85212 83884 85264
rect 87972 85212 88024 85264
rect 84844 85076 84896 85128
rect 85580 85076 85632 85128
rect 84568 84940 84620 84992
rect 84844 84940 84896 84992
rect 1982 84838 2034 84890
rect 2046 84838 2098 84890
rect 2110 84838 2162 84890
rect 2174 84838 2226 84890
rect 85982 84838 86034 84890
rect 86046 84838 86098 84890
rect 86110 84838 86162 84890
rect 86174 84838 86226 84890
rect 89982 84838 90034 84890
rect 90046 84838 90098 84890
rect 90110 84838 90162 84890
rect 90174 84838 90226 84890
rect 85028 84736 85080 84788
rect 85212 84736 85264 84788
rect 86960 84736 87012 84788
rect 87236 84736 87288 84788
rect 82912 84532 82964 84584
rect 84108 84532 84160 84584
rect 3982 84294 4034 84346
rect 4046 84294 4098 84346
rect 4110 84294 4162 84346
rect 4174 84294 4226 84346
rect 87982 84294 88034 84346
rect 88046 84294 88098 84346
rect 88110 84294 88162 84346
rect 88174 84294 88226 84346
rect 83096 84124 83148 84176
rect 87972 84124 88024 84176
rect 1982 83750 2034 83802
rect 2046 83750 2098 83802
rect 2110 83750 2162 83802
rect 2174 83750 2226 83802
rect 85982 83750 86034 83802
rect 86046 83750 86098 83802
rect 86110 83750 86162 83802
rect 86174 83750 86226 83802
rect 89982 83750 90034 83802
rect 90046 83750 90098 83802
rect 90110 83750 90162 83802
rect 90174 83750 90226 83802
rect 4804 83351 4856 83360
rect 4804 83317 4813 83351
rect 4813 83317 4847 83351
rect 4847 83317 4856 83351
rect 4804 83308 4856 83317
rect 3982 83206 4034 83258
rect 4046 83206 4098 83258
rect 4110 83206 4162 83258
rect 4174 83206 4226 83258
rect 87982 83206 88034 83258
rect 88046 83206 88098 83258
rect 88110 83206 88162 83258
rect 88174 83206 88226 83258
rect 1982 82662 2034 82714
rect 2046 82662 2098 82714
rect 2110 82662 2162 82714
rect 2174 82662 2226 82714
rect 85982 82662 86034 82714
rect 86046 82662 86098 82714
rect 86110 82662 86162 82714
rect 86174 82662 86226 82714
rect 89982 82662 90034 82714
rect 90046 82662 90098 82714
rect 90110 82662 90162 82714
rect 90174 82662 90226 82714
rect 4804 82263 4856 82272
rect 4804 82229 4813 82263
rect 4813 82229 4847 82263
rect 4847 82229 4856 82263
rect 4804 82220 4856 82229
rect 3982 82118 4034 82170
rect 4046 82118 4098 82170
rect 4110 82118 4162 82170
rect 4174 82118 4226 82170
rect 87982 82118 88034 82170
rect 88046 82118 88098 82170
rect 88110 82118 88162 82170
rect 88174 82118 88226 82170
rect 83188 81948 83240 82000
rect 87972 81948 88024 82000
rect 1982 81574 2034 81626
rect 2046 81574 2098 81626
rect 2110 81574 2162 81626
rect 2174 81574 2226 81626
rect 85982 81574 86034 81626
rect 86046 81574 86098 81626
rect 86110 81574 86162 81626
rect 86174 81574 86226 81626
rect 89982 81574 90034 81626
rect 90046 81574 90098 81626
rect 90110 81574 90162 81626
rect 90174 81574 90226 81626
rect 3982 81030 4034 81082
rect 4046 81030 4098 81082
rect 4110 81030 4162 81082
rect 4174 81030 4226 81082
rect 87982 81030 88034 81082
rect 88046 81030 88098 81082
rect 88110 81030 88162 81082
rect 88174 81030 88226 81082
rect 83280 80860 83332 80912
rect 87972 80860 88024 80912
rect 1982 80486 2034 80538
rect 2046 80486 2098 80538
rect 2110 80486 2162 80538
rect 2174 80486 2226 80538
rect 85982 80486 86034 80538
rect 86046 80486 86098 80538
rect 86110 80486 86162 80538
rect 86174 80486 86226 80538
rect 89982 80486 90034 80538
rect 90046 80486 90098 80538
rect 90110 80486 90162 80538
rect 90174 80486 90226 80538
rect 4804 80427 4856 80436
rect 4804 80393 4813 80427
rect 4813 80393 4847 80427
rect 4847 80393 4856 80427
rect 4804 80384 4856 80393
rect 86776 80112 86828 80164
rect 87328 80112 87380 80164
rect 87512 80112 87564 80164
rect 88340 80112 88392 80164
rect 3982 79942 4034 79994
rect 4046 79942 4098 79994
rect 4110 79942 4162 79994
rect 4174 79942 4226 79994
rect 87982 79942 88034 79994
rect 88046 79942 88098 79994
rect 88110 79942 88162 79994
rect 88174 79942 88226 79994
rect 1982 79398 2034 79450
rect 2046 79398 2098 79450
rect 2110 79398 2162 79450
rect 2174 79398 2226 79450
rect 85982 79398 86034 79450
rect 86046 79398 86098 79450
rect 86110 79398 86162 79450
rect 86174 79398 86226 79450
rect 89982 79398 90034 79450
rect 90046 79398 90098 79450
rect 90110 79398 90162 79450
rect 90174 79398 90226 79450
rect 3982 78854 4034 78906
rect 4046 78854 4098 78906
rect 4110 78854 4162 78906
rect 4174 78854 4226 78906
rect 87982 78854 88034 78906
rect 88046 78854 88098 78906
rect 88110 78854 88162 78906
rect 88174 78854 88226 78906
rect 1982 78310 2034 78362
rect 2046 78310 2098 78362
rect 2110 78310 2162 78362
rect 2174 78310 2226 78362
rect 85982 78310 86034 78362
rect 86046 78310 86098 78362
rect 86110 78310 86162 78362
rect 86174 78310 86226 78362
rect 89982 78310 90034 78362
rect 90046 78310 90098 78362
rect 90110 78310 90162 78362
rect 90174 78310 90226 78362
rect 3982 77766 4034 77818
rect 4046 77766 4098 77818
rect 4110 77766 4162 77818
rect 4174 77766 4226 77818
rect 87982 77766 88034 77818
rect 88046 77766 88098 77818
rect 88110 77766 88162 77818
rect 88174 77766 88226 77818
rect 1982 77222 2034 77274
rect 2046 77222 2098 77274
rect 2110 77222 2162 77274
rect 2174 77222 2226 77274
rect 85982 77222 86034 77274
rect 86046 77222 86098 77274
rect 86110 77222 86162 77274
rect 86174 77222 86226 77274
rect 89982 77222 90034 77274
rect 90046 77222 90098 77274
rect 90110 77222 90162 77274
rect 90174 77222 90226 77274
rect 84108 77120 84160 77172
rect 87052 77120 87104 77172
rect 3982 76678 4034 76730
rect 4046 76678 4098 76730
rect 4110 76678 4162 76730
rect 4174 76678 4226 76730
rect 87982 76678 88034 76730
rect 88046 76678 88098 76730
rect 88110 76678 88162 76730
rect 88174 76678 88226 76730
rect 1982 76134 2034 76186
rect 2046 76134 2098 76186
rect 2110 76134 2162 76186
rect 2174 76134 2226 76186
rect 85982 76134 86034 76186
rect 86046 76134 86098 76186
rect 86110 76134 86162 76186
rect 86174 76134 86226 76186
rect 89982 76134 90034 76186
rect 90046 76134 90098 76186
rect 90110 76134 90162 76186
rect 90174 76134 90226 76186
rect 3982 75590 4034 75642
rect 4046 75590 4098 75642
rect 4110 75590 4162 75642
rect 4174 75590 4226 75642
rect 87982 75590 88034 75642
rect 88046 75590 88098 75642
rect 88110 75590 88162 75642
rect 88174 75590 88226 75642
rect 87144 75488 87196 75540
rect 87420 75488 87472 75540
rect 87420 75216 87472 75268
rect 87788 75216 87840 75268
rect 1982 75046 2034 75098
rect 2046 75046 2098 75098
rect 2110 75046 2162 75098
rect 2174 75046 2226 75098
rect 85982 75046 86034 75098
rect 86046 75046 86098 75098
rect 86110 75046 86162 75098
rect 86174 75046 86226 75098
rect 89982 75046 90034 75098
rect 90046 75046 90098 75098
rect 90110 75046 90162 75098
rect 90174 75046 90226 75098
rect 3982 74502 4034 74554
rect 4046 74502 4098 74554
rect 4110 74502 4162 74554
rect 4174 74502 4226 74554
rect 87982 74502 88034 74554
rect 88046 74502 88098 74554
rect 88110 74502 88162 74554
rect 88174 74502 88226 74554
rect 82452 74400 82504 74452
rect 86960 74400 87012 74452
rect 1982 73958 2034 74010
rect 2046 73958 2098 74010
rect 2110 73958 2162 74010
rect 2174 73958 2226 74010
rect 85982 73958 86034 74010
rect 86046 73958 86098 74010
rect 86110 73958 86162 74010
rect 86174 73958 86226 74010
rect 89982 73958 90034 74010
rect 90046 73958 90098 74010
rect 90110 73958 90162 74010
rect 90174 73958 90226 74010
rect 3982 73414 4034 73466
rect 4046 73414 4098 73466
rect 4110 73414 4162 73466
rect 4174 73414 4226 73466
rect 87982 73414 88034 73466
rect 88046 73414 88098 73466
rect 88110 73414 88162 73466
rect 88174 73414 88226 73466
rect 1982 72870 2034 72922
rect 2046 72870 2098 72922
rect 2110 72870 2162 72922
rect 2174 72870 2226 72922
rect 85982 72870 86034 72922
rect 86046 72870 86098 72922
rect 86110 72870 86162 72922
rect 86174 72870 86226 72922
rect 89982 72870 90034 72922
rect 90046 72870 90098 72922
rect 90110 72870 90162 72922
rect 90174 72870 90226 72922
rect 3982 72326 4034 72378
rect 4046 72326 4098 72378
rect 4110 72326 4162 72378
rect 4174 72326 4226 72378
rect 87982 72326 88034 72378
rect 88046 72326 88098 72378
rect 88110 72326 88162 72378
rect 88174 72326 88226 72378
rect 1982 71782 2034 71834
rect 2046 71782 2098 71834
rect 2110 71782 2162 71834
rect 2174 71782 2226 71834
rect 85982 71782 86034 71834
rect 86046 71782 86098 71834
rect 86110 71782 86162 71834
rect 86174 71782 86226 71834
rect 89982 71782 90034 71834
rect 90046 71782 90098 71834
rect 90110 71782 90162 71834
rect 90174 71782 90226 71834
rect 3982 71238 4034 71290
rect 4046 71238 4098 71290
rect 4110 71238 4162 71290
rect 4174 71238 4226 71290
rect 87982 71238 88034 71290
rect 88046 71238 88098 71290
rect 88110 71238 88162 71290
rect 88174 71238 88226 71290
rect 1982 70694 2034 70746
rect 2046 70694 2098 70746
rect 2110 70694 2162 70746
rect 2174 70694 2226 70746
rect 85982 70694 86034 70746
rect 86046 70694 86098 70746
rect 86110 70694 86162 70746
rect 86174 70694 86226 70746
rect 89982 70694 90034 70746
rect 90046 70694 90098 70746
rect 90110 70694 90162 70746
rect 90174 70694 90226 70746
rect 84016 70320 84068 70372
rect 87788 70320 87840 70372
rect 3982 70150 4034 70202
rect 4046 70150 4098 70202
rect 4110 70150 4162 70202
rect 4174 70150 4226 70202
rect 87982 70150 88034 70202
rect 88046 70150 88098 70202
rect 88110 70150 88162 70202
rect 88174 70150 88226 70202
rect 1982 69606 2034 69658
rect 2046 69606 2098 69658
rect 2110 69606 2162 69658
rect 2174 69606 2226 69658
rect 85982 69606 86034 69658
rect 86046 69606 86098 69658
rect 86110 69606 86162 69658
rect 86174 69606 86226 69658
rect 89982 69606 90034 69658
rect 90046 69606 90098 69658
rect 90110 69606 90162 69658
rect 90174 69606 90226 69658
rect 3982 69062 4034 69114
rect 4046 69062 4098 69114
rect 4110 69062 4162 69114
rect 4174 69062 4226 69114
rect 87982 69062 88034 69114
rect 88046 69062 88098 69114
rect 88110 69062 88162 69114
rect 88174 69062 88226 69114
rect 83924 68960 83976 69012
rect 87144 68960 87196 69012
rect 1982 68518 2034 68570
rect 2046 68518 2098 68570
rect 2110 68518 2162 68570
rect 2174 68518 2226 68570
rect 85982 68518 86034 68570
rect 86046 68518 86098 68570
rect 86110 68518 86162 68570
rect 86174 68518 86226 68570
rect 89982 68518 90034 68570
rect 90046 68518 90098 68570
rect 90110 68518 90162 68570
rect 90174 68518 90226 68570
rect 3982 67974 4034 68026
rect 4046 67974 4098 68026
rect 4110 67974 4162 68026
rect 4174 67974 4226 68026
rect 87982 67974 88034 68026
rect 88046 67974 88098 68026
rect 88110 67974 88162 68026
rect 88174 67974 88226 68026
rect 1982 67430 2034 67482
rect 2046 67430 2098 67482
rect 2110 67430 2162 67482
rect 2174 67430 2226 67482
rect 85982 67430 86034 67482
rect 86046 67430 86098 67482
rect 86110 67430 86162 67482
rect 86174 67430 86226 67482
rect 89982 67430 90034 67482
rect 90046 67430 90098 67482
rect 90110 67430 90162 67482
rect 90174 67430 90226 67482
rect 3982 66886 4034 66938
rect 4046 66886 4098 66938
rect 4110 66886 4162 66938
rect 4174 66886 4226 66938
rect 87982 66886 88034 66938
rect 88046 66886 88098 66938
rect 88110 66886 88162 66938
rect 88174 66886 88226 66938
rect 1982 66342 2034 66394
rect 2046 66342 2098 66394
rect 2110 66342 2162 66394
rect 2174 66342 2226 66394
rect 85982 66342 86034 66394
rect 86046 66342 86098 66394
rect 86110 66342 86162 66394
rect 86174 66342 86226 66394
rect 89982 66342 90034 66394
rect 90046 66342 90098 66394
rect 90110 66342 90162 66394
rect 90174 66342 90226 66394
rect 83832 66172 83884 66224
rect 87788 66172 87840 66224
rect 84200 66104 84252 66156
rect 87328 66104 87380 66156
rect 3982 65798 4034 65850
rect 4046 65798 4098 65850
rect 4110 65798 4162 65850
rect 4174 65798 4226 65850
rect 87982 65798 88034 65850
rect 88046 65798 88098 65850
rect 88110 65798 88162 65850
rect 88174 65798 88226 65850
rect 1982 65254 2034 65306
rect 2046 65254 2098 65306
rect 2110 65254 2162 65306
rect 2174 65254 2226 65306
rect 85982 65254 86034 65306
rect 86046 65254 86098 65306
rect 86110 65254 86162 65306
rect 86174 65254 86226 65306
rect 89982 65254 90034 65306
rect 90046 65254 90098 65306
rect 90110 65254 90162 65306
rect 90174 65254 90226 65306
rect 3982 64710 4034 64762
rect 4046 64710 4098 64762
rect 4110 64710 4162 64762
rect 4174 64710 4226 64762
rect 87982 64710 88034 64762
rect 88046 64710 88098 64762
rect 88110 64710 88162 64762
rect 88174 64710 88226 64762
rect 1982 64166 2034 64218
rect 2046 64166 2098 64218
rect 2110 64166 2162 64218
rect 2174 64166 2226 64218
rect 85982 64166 86034 64218
rect 86046 64166 86098 64218
rect 86110 64166 86162 64218
rect 86174 64166 86226 64218
rect 89982 64166 90034 64218
rect 90046 64166 90098 64218
rect 90110 64166 90162 64218
rect 90174 64166 90226 64218
rect 3982 63622 4034 63674
rect 4046 63622 4098 63674
rect 4110 63622 4162 63674
rect 4174 63622 4226 63674
rect 87982 63622 88034 63674
rect 88046 63622 88098 63674
rect 88110 63622 88162 63674
rect 88174 63622 88226 63674
rect 83740 63452 83792 63504
rect 87788 63452 87840 63504
rect 1982 63078 2034 63130
rect 2046 63078 2098 63130
rect 2110 63078 2162 63130
rect 2174 63078 2226 63130
rect 85982 63078 86034 63130
rect 86046 63078 86098 63130
rect 86110 63078 86162 63130
rect 86174 63078 86226 63130
rect 89982 63078 90034 63130
rect 90046 63078 90098 63130
rect 90110 63078 90162 63130
rect 90174 63078 90226 63130
rect 3982 62534 4034 62586
rect 4046 62534 4098 62586
rect 4110 62534 4162 62586
rect 4174 62534 4226 62586
rect 87982 62534 88034 62586
rect 88046 62534 88098 62586
rect 88110 62534 88162 62586
rect 88174 62534 88226 62586
rect 1982 61990 2034 62042
rect 2046 61990 2098 62042
rect 2110 61990 2162 62042
rect 2174 61990 2226 62042
rect 85982 61990 86034 62042
rect 86046 61990 86098 62042
rect 86110 61990 86162 62042
rect 86174 61990 86226 62042
rect 89982 61990 90034 62042
rect 90046 61990 90098 62042
rect 90110 61990 90162 62042
rect 90174 61990 90226 62042
rect 84292 61888 84344 61940
rect 87788 61888 87840 61940
rect 3982 61446 4034 61498
rect 4046 61446 4098 61498
rect 4110 61446 4162 61498
rect 4174 61446 4226 61498
rect 87982 61446 88034 61498
rect 88046 61446 88098 61498
rect 88110 61446 88162 61498
rect 88174 61446 88226 61498
rect 1982 60902 2034 60954
rect 2046 60902 2098 60954
rect 2110 60902 2162 60954
rect 2174 60902 2226 60954
rect 85982 60902 86034 60954
rect 86046 60902 86098 60954
rect 86110 60902 86162 60954
rect 86174 60902 86226 60954
rect 89982 60902 90034 60954
rect 90046 60902 90098 60954
rect 90110 60902 90162 60954
rect 90174 60902 90226 60954
rect 3982 60358 4034 60410
rect 4046 60358 4098 60410
rect 4110 60358 4162 60410
rect 4174 60358 4226 60410
rect 87982 60358 88034 60410
rect 88046 60358 88098 60410
rect 88110 60358 88162 60410
rect 88174 60358 88226 60410
rect 1982 59814 2034 59866
rect 2046 59814 2098 59866
rect 2110 59814 2162 59866
rect 2174 59814 2226 59866
rect 85982 59814 86034 59866
rect 86046 59814 86098 59866
rect 86110 59814 86162 59866
rect 86174 59814 86226 59866
rect 89982 59814 90034 59866
rect 90046 59814 90098 59866
rect 90110 59814 90162 59866
rect 90174 59814 90226 59866
rect 3982 59270 4034 59322
rect 4046 59270 4098 59322
rect 4110 59270 4162 59322
rect 4174 59270 4226 59322
rect 87982 59270 88034 59322
rect 88046 59270 88098 59322
rect 88110 59270 88162 59322
rect 88174 59270 88226 59322
rect 1982 58726 2034 58778
rect 2046 58726 2098 58778
rect 2110 58726 2162 58778
rect 2174 58726 2226 58778
rect 85982 58726 86034 58778
rect 86046 58726 86098 58778
rect 86110 58726 86162 58778
rect 86174 58726 86226 58778
rect 89982 58726 90034 58778
rect 90046 58726 90098 58778
rect 90110 58726 90162 58778
rect 90174 58726 90226 58778
rect 3982 58182 4034 58234
rect 4046 58182 4098 58234
rect 4110 58182 4162 58234
rect 4174 58182 4226 58234
rect 87982 58182 88034 58234
rect 88046 58182 88098 58234
rect 88110 58182 88162 58234
rect 88174 58182 88226 58234
rect 4528 57876 4580 57928
rect 84752 57876 84804 57928
rect 86960 57876 87012 57928
rect 1982 57638 2034 57690
rect 2046 57638 2098 57690
rect 2110 57638 2162 57690
rect 2174 57638 2226 57690
rect 85982 57638 86034 57690
rect 86046 57638 86098 57690
rect 86110 57638 86162 57690
rect 86174 57638 86226 57690
rect 89982 57638 90034 57690
rect 90046 57638 90098 57690
rect 90110 57638 90162 57690
rect 90174 57638 90226 57690
rect 3982 57094 4034 57146
rect 4046 57094 4098 57146
rect 4110 57094 4162 57146
rect 4174 57094 4226 57146
rect 87982 57094 88034 57146
rect 88046 57094 88098 57146
rect 88110 57094 88162 57146
rect 88174 57094 88226 57146
rect 1982 56550 2034 56602
rect 2046 56550 2098 56602
rect 2110 56550 2162 56602
rect 2174 56550 2226 56602
rect 85982 56550 86034 56602
rect 86046 56550 86098 56602
rect 86110 56550 86162 56602
rect 86174 56550 86226 56602
rect 89982 56550 90034 56602
rect 90046 56550 90098 56602
rect 90110 56550 90162 56602
rect 90174 56550 90226 56602
rect 85488 56448 85540 56500
rect 86960 56448 87012 56500
rect 85120 56380 85172 56432
rect 87052 56380 87104 56432
rect 3982 56006 4034 56058
rect 4046 56006 4098 56058
rect 4110 56006 4162 56058
rect 4174 56006 4226 56058
rect 87982 56006 88034 56058
rect 88046 56006 88098 56058
rect 88110 56006 88162 56058
rect 88174 56006 88226 56058
rect 1982 55462 2034 55514
rect 2046 55462 2098 55514
rect 2110 55462 2162 55514
rect 2174 55462 2226 55514
rect 85982 55462 86034 55514
rect 86046 55462 86098 55514
rect 86110 55462 86162 55514
rect 86174 55462 86226 55514
rect 89982 55462 90034 55514
rect 90046 55462 90098 55514
rect 90110 55462 90162 55514
rect 90174 55462 90226 55514
rect 3982 54918 4034 54970
rect 4046 54918 4098 54970
rect 4110 54918 4162 54970
rect 4174 54918 4226 54970
rect 87982 54918 88034 54970
rect 88046 54918 88098 54970
rect 88110 54918 88162 54970
rect 88174 54918 88226 54970
rect 85212 54612 85264 54664
rect 86960 54612 87012 54664
rect 1982 54374 2034 54426
rect 2046 54374 2098 54426
rect 2110 54374 2162 54426
rect 2174 54374 2226 54426
rect 85982 54374 86034 54426
rect 86046 54374 86098 54426
rect 86110 54374 86162 54426
rect 86174 54374 86226 54426
rect 89982 54374 90034 54426
rect 90046 54374 90098 54426
rect 90110 54374 90162 54426
rect 90174 54374 90226 54426
rect 3982 53830 4034 53882
rect 4046 53830 4098 53882
rect 4110 53830 4162 53882
rect 4174 53830 4226 53882
rect 87982 53830 88034 53882
rect 88046 53830 88098 53882
rect 88110 53830 88162 53882
rect 88174 53830 88226 53882
rect 84844 53728 84896 53780
rect 86960 53728 87012 53780
rect 1982 53286 2034 53338
rect 2046 53286 2098 53338
rect 2110 53286 2162 53338
rect 2174 53286 2226 53338
rect 85982 53286 86034 53338
rect 86046 53286 86098 53338
rect 86110 53286 86162 53338
rect 86174 53286 86226 53338
rect 89982 53286 90034 53338
rect 90046 53286 90098 53338
rect 90110 53286 90162 53338
rect 90174 53286 90226 53338
rect 3982 52742 4034 52794
rect 4046 52742 4098 52794
rect 4110 52742 4162 52794
rect 4174 52742 4226 52794
rect 87982 52742 88034 52794
rect 88046 52742 88098 52794
rect 88110 52742 88162 52794
rect 88174 52742 88226 52794
rect 1982 52198 2034 52250
rect 2046 52198 2098 52250
rect 2110 52198 2162 52250
rect 2174 52198 2226 52250
rect 85982 52198 86034 52250
rect 86046 52198 86098 52250
rect 86110 52198 86162 52250
rect 86174 52198 86226 52250
rect 89982 52198 90034 52250
rect 90046 52198 90098 52250
rect 90110 52198 90162 52250
rect 90174 52198 90226 52250
rect 3982 51654 4034 51706
rect 4046 51654 4098 51706
rect 4110 51654 4162 51706
rect 4174 51654 4226 51706
rect 87982 51654 88034 51706
rect 88046 51654 88098 51706
rect 88110 51654 88162 51706
rect 88174 51654 88226 51706
rect 1982 51110 2034 51162
rect 2046 51110 2098 51162
rect 2110 51110 2162 51162
rect 2174 51110 2226 51162
rect 85982 51110 86034 51162
rect 86046 51110 86098 51162
rect 86110 51110 86162 51162
rect 86174 51110 86226 51162
rect 89982 51110 90034 51162
rect 90046 51110 90098 51162
rect 90110 51110 90162 51162
rect 90174 51110 90226 51162
rect 3982 50566 4034 50618
rect 4046 50566 4098 50618
rect 4110 50566 4162 50618
rect 4174 50566 4226 50618
rect 87982 50566 88034 50618
rect 88046 50566 88098 50618
rect 88110 50566 88162 50618
rect 88174 50566 88226 50618
rect 1982 50022 2034 50074
rect 2046 50022 2098 50074
rect 2110 50022 2162 50074
rect 2174 50022 2226 50074
rect 85982 50022 86034 50074
rect 86046 50022 86098 50074
rect 86110 50022 86162 50074
rect 86174 50022 86226 50074
rect 89982 50022 90034 50074
rect 90046 50022 90098 50074
rect 90110 50022 90162 50074
rect 90174 50022 90226 50074
rect 4436 49963 4488 49972
rect 4436 49929 4445 49963
rect 4445 49929 4479 49963
rect 4479 49929 4488 49963
rect 4436 49920 4488 49929
rect 82728 49648 82780 49700
rect 87696 49648 87748 49700
rect 3982 49478 4034 49530
rect 4046 49478 4098 49530
rect 4110 49478 4162 49530
rect 4174 49478 4226 49530
rect 87982 49478 88034 49530
rect 88046 49478 88098 49530
rect 88110 49478 88162 49530
rect 88174 49478 88226 49530
rect 1982 48934 2034 48986
rect 2046 48934 2098 48986
rect 2110 48934 2162 48986
rect 2174 48934 2226 48986
rect 85982 48934 86034 48986
rect 86046 48934 86098 48986
rect 86110 48934 86162 48986
rect 86174 48934 86226 48986
rect 89982 48934 90034 48986
rect 90046 48934 90098 48986
rect 90110 48934 90162 48986
rect 90174 48934 90226 48986
rect 3982 48390 4034 48442
rect 4046 48390 4098 48442
rect 4110 48390 4162 48442
rect 4174 48390 4226 48442
rect 87982 48390 88034 48442
rect 88046 48390 88098 48442
rect 88110 48390 88162 48442
rect 88174 48390 88226 48442
rect 1982 47846 2034 47898
rect 2046 47846 2098 47898
rect 2110 47846 2162 47898
rect 2174 47846 2226 47898
rect 85982 47846 86034 47898
rect 86046 47846 86098 47898
rect 86110 47846 86162 47898
rect 86174 47846 86226 47898
rect 89982 47846 90034 47898
rect 90046 47846 90098 47898
rect 90110 47846 90162 47898
rect 90174 47846 90226 47898
rect 3982 47302 4034 47354
rect 4046 47302 4098 47354
rect 4110 47302 4162 47354
rect 4174 47302 4226 47354
rect 87982 47302 88034 47354
rect 88046 47302 88098 47354
rect 88110 47302 88162 47354
rect 88174 47302 88226 47354
rect 1982 46758 2034 46810
rect 2046 46758 2098 46810
rect 2110 46758 2162 46810
rect 2174 46758 2226 46810
rect 85982 46758 86034 46810
rect 86046 46758 86098 46810
rect 86110 46758 86162 46810
rect 86174 46758 86226 46810
rect 89982 46758 90034 46810
rect 90046 46758 90098 46810
rect 90110 46758 90162 46810
rect 90174 46758 90226 46810
rect 3982 46214 4034 46266
rect 4046 46214 4098 46266
rect 4110 46214 4162 46266
rect 4174 46214 4226 46266
rect 87982 46214 88034 46266
rect 88046 46214 88098 46266
rect 88110 46214 88162 46266
rect 88174 46214 88226 46266
rect 1982 45670 2034 45722
rect 2046 45670 2098 45722
rect 2110 45670 2162 45722
rect 2174 45670 2226 45722
rect 85982 45670 86034 45722
rect 86046 45670 86098 45722
rect 86110 45670 86162 45722
rect 86174 45670 86226 45722
rect 89982 45670 90034 45722
rect 90046 45670 90098 45722
rect 90110 45670 90162 45722
rect 90174 45670 90226 45722
rect 83740 45568 83792 45620
rect 87696 45568 87748 45620
rect 3982 45126 4034 45178
rect 4046 45126 4098 45178
rect 4110 45126 4162 45178
rect 4174 45126 4226 45178
rect 87982 45126 88034 45178
rect 88046 45126 88098 45178
rect 88110 45126 88162 45178
rect 88174 45126 88226 45178
rect 1982 44582 2034 44634
rect 2046 44582 2098 44634
rect 2110 44582 2162 44634
rect 2174 44582 2226 44634
rect 85982 44582 86034 44634
rect 86046 44582 86098 44634
rect 86110 44582 86162 44634
rect 86174 44582 86226 44634
rect 89982 44582 90034 44634
rect 90046 44582 90098 44634
rect 90110 44582 90162 44634
rect 90174 44582 90226 44634
rect 83832 44140 83884 44192
rect 87696 44140 87748 44192
rect 3982 44038 4034 44090
rect 4046 44038 4098 44090
rect 4110 44038 4162 44090
rect 4174 44038 4226 44090
rect 87982 44038 88034 44090
rect 88046 44038 88098 44090
rect 88110 44038 88162 44090
rect 88174 44038 88226 44090
rect 1982 43494 2034 43546
rect 2046 43494 2098 43546
rect 2110 43494 2162 43546
rect 2174 43494 2226 43546
rect 85982 43494 86034 43546
rect 86046 43494 86098 43546
rect 86110 43494 86162 43546
rect 86174 43494 86226 43546
rect 89982 43494 90034 43546
rect 90046 43494 90098 43546
rect 90110 43494 90162 43546
rect 90174 43494 90226 43546
rect 3982 42950 4034 43002
rect 4046 42950 4098 43002
rect 4110 42950 4162 43002
rect 4174 42950 4226 43002
rect 87982 42950 88034 43002
rect 88046 42950 88098 43002
rect 88110 42950 88162 43002
rect 88174 42950 88226 43002
rect 1982 42406 2034 42458
rect 2046 42406 2098 42458
rect 2110 42406 2162 42458
rect 2174 42406 2226 42458
rect 85982 42406 86034 42458
rect 86046 42406 86098 42458
rect 86110 42406 86162 42458
rect 86174 42406 86226 42458
rect 89982 42406 90034 42458
rect 90046 42406 90098 42458
rect 90110 42406 90162 42458
rect 90174 42406 90226 42458
rect 3982 41862 4034 41914
rect 4046 41862 4098 41914
rect 4110 41862 4162 41914
rect 4174 41862 4226 41914
rect 87982 41862 88034 41914
rect 88046 41862 88098 41914
rect 88110 41862 88162 41914
rect 88174 41862 88226 41914
rect 1982 41318 2034 41370
rect 2046 41318 2098 41370
rect 2110 41318 2162 41370
rect 2174 41318 2226 41370
rect 85982 41318 86034 41370
rect 86046 41318 86098 41370
rect 86110 41318 86162 41370
rect 86174 41318 86226 41370
rect 89982 41318 90034 41370
rect 90046 41318 90098 41370
rect 90110 41318 90162 41370
rect 90174 41318 90226 41370
rect 3982 40774 4034 40826
rect 4046 40774 4098 40826
rect 4110 40774 4162 40826
rect 4174 40774 4226 40826
rect 87982 40774 88034 40826
rect 88046 40774 88098 40826
rect 88110 40774 88162 40826
rect 88174 40774 88226 40826
rect 87328 40672 87380 40724
rect 87880 40672 87932 40724
rect 1982 40230 2034 40282
rect 2046 40230 2098 40282
rect 2110 40230 2162 40282
rect 2174 40230 2226 40282
rect 85982 40230 86034 40282
rect 86046 40230 86098 40282
rect 86110 40230 86162 40282
rect 86174 40230 86226 40282
rect 89982 40230 90034 40282
rect 90046 40230 90098 40282
rect 90110 40230 90162 40282
rect 90174 40230 90226 40282
rect 84844 40060 84896 40112
rect 87880 40060 87932 40112
rect 3982 39686 4034 39738
rect 4046 39686 4098 39738
rect 4110 39686 4162 39738
rect 4174 39686 4226 39738
rect 87982 39686 88034 39738
rect 88046 39686 88098 39738
rect 88110 39686 88162 39738
rect 88174 39686 88226 39738
rect 1982 39142 2034 39194
rect 2046 39142 2098 39194
rect 2110 39142 2162 39194
rect 2174 39142 2226 39194
rect 85982 39142 86034 39194
rect 86046 39142 86098 39194
rect 86110 39142 86162 39194
rect 86174 39142 86226 39194
rect 89982 39142 90034 39194
rect 90046 39142 90098 39194
rect 90110 39142 90162 39194
rect 90174 39142 90226 39194
rect 84384 39040 84436 39092
rect 3982 38598 4034 38650
rect 4046 38598 4098 38650
rect 4110 38598 4162 38650
rect 4174 38598 4226 38650
rect 87982 38598 88034 38650
rect 88046 38598 88098 38650
rect 88110 38598 88162 38650
rect 88174 38598 88226 38650
rect 1982 38054 2034 38106
rect 2046 38054 2098 38106
rect 2110 38054 2162 38106
rect 2174 38054 2226 38106
rect 85982 38054 86034 38106
rect 86046 38054 86098 38106
rect 86110 38054 86162 38106
rect 86174 38054 86226 38106
rect 89982 38054 90034 38106
rect 90046 38054 90098 38106
rect 90110 38054 90162 38106
rect 90174 38054 90226 38106
rect 3982 37510 4034 37562
rect 4046 37510 4098 37562
rect 4110 37510 4162 37562
rect 4174 37510 4226 37562
rect 87982 37510 88034 37562
rect 88046 37510 88098 37562
rect 88110 37510 88162 37562
rect 88174 37510 88226 37562
rect 1982 36966 2034 37018
rect 2046 36966 2098 37018
rect 2110 36966 2162 37018
rect 2174 36966 2226 37018
rect 85982 36966 86034 37018
rect 86046 36966 86098 37018
rect 86110 36966 86162 37018
rect 86174 36966 86226 37018
rect 89982 36966 90034 37018
rect 90046 36966 90098 37018
rect 90110 36966 90162 37018
rect 90174 36966 90226 37018
rect 3982 36422 4034 36474
rect 4046 36422 4098 36474
rect 4110 36422 4162 36474
rect 4174 36422 4226 36474
rect 87982 36422 88034 36474
rect 88046 36422 88098 36474
rect 88110 36422 88162 36474
rect 88174 36422 88226 36474
rect 85120 36320 85172 36372
rect 86960 36320 87012 36372
rect 1982 35878 2034 35930
rect 2046 35878 2098 35930
rect 2110 35878 2162 35930
rect 2174 35878 2226 35930
rect 85982 35878 86034 35930
rect 86046 35878 86098 35930
rect 86110 35878 86162 35930
rect 86174 35878 86226 35930
rect 89982 35878 90034 35930
rect 90046 35878 90098 35930
rect 90110 35878 90162 35930
rect 90174 35878 90226 35930
rect 3982 35334 4034 35386
rect 4046 35334 4098 35386
rect 4110 35334 4162 35386
rect 4174 35334 4226 35386
rect 87982 35334 88034 35386
rect 88046 35334 88098 35386
rect 88110 35334 88162 35386
rect 88174 35334 88226 35386
rect 1982 34790 2034 34842
rect 2046 34790 2098 34842
rect 2110 34790 2162 34842
rect 2174 34790 2226 34842
rect 85982 34790 86034 34842
rect 86046 34790 86098 34842
rect 86110 34790 86162 34842
rect 86174 34790 86226 34842
rect 89982 34790 90034 34842
rect 90046 34790 90098 34842
rect 90110 34790 90162 34842
rect 90174 34790 90226 34842
rect 85212 34484 85264 34536
rect 86960 34484 87012 34536
rect 3982 34246 4034 34298
rect 4046 34246 4098 34298
rect 4110 34246 4162 34298
rect 4174 34246 4226 34298
rect 87982 34246 88034 34298
rect 88046 34246 88098 34298
rect 88110 34246 88162 34298
rect 88174 34246 88226 34298
rect 1982 33702 2034 33754
rect 2046 33702 2098 33754
rect 2110 33702 2162 33754
rect 2174 33702 2226 33754
rect 85982 33702 86034 33754
rect 86046 33702 86098 33754
rect 86110 33702 86162 33754
rect 86174 33702 86226 33754
rect 89982 33702 90034 33754
rect 90046 33702 90098 33754
rect 90110 33702 90162 33754
rect 90174 33702 90226 33754
rect 3982 33158 4034 33210
rect 4046 33158 4098 33210
rect 4110 33158 4162 33210
rect 4174 33158 4226 33210
rect 87982 33158 88034 33210
rect 88046 33158 88098 33210
rect 88110 33158 88162 33210
rect 88174 33158 88226 33210
rect 1982 32614 2034 32666
rect 2046 32614 2098 32666
rect 2110 32614 2162 32666
rect 2174 32614 2226 32666
rect 85982 32614 86034 32666
rect 86046 32614 86098 32666
rect 86110 32614 86162 32666
rect 86174 32614 86226 32666
rect 89982 32614 90034 32666
rect 90046 32614 90098 32666
rect 90110 32614 90162 32666
rect 90174 32614 90226 32666
rect 3982 32070 4034 32122
rect 4046 32070 4098 32122
rect 4110 32070 4162 32122
rect 4174 32070 4226 32122
rect 87982 32070 88034 32122
rect 88046 32070 88098 32122
rect 88110 32070 88162 32122
rect 88174 32070 88226 32122
rect 84752 32011 84804 32020
rect 84752 31977 84761 32011
rect 84761 31977 84795 32011
rect 84795 31977 84804 32011
rect 84752 31968 84804 31977
rect 86592 31968 86644 32020
rect 85488 31764 85540 31816
rect 86960 31764 87012 31816
rect 1982 31526 2034 31578
rect 2046 31526 2098 31578
rect 2110 31526 2162 31578
rect 2174 31526 2226 31578
rect 85982 31526 86034 31578
rect 86046 31526 86098 31578
rect 86110 31526 86162 31578
rect 86174 31526 86226 31578
rect 89982 31526 90034 31578
rect 90046 31526 90098 31578
rect 90110 31526 90162 31578
rect 90174 31526 90226 31578
rect 3982 30982 4034 31034
rect 4046 30982 4098 31034
rect 4110 30982 4162 31034
rect 4174 30982 4226 31034
rect 87982 30982 88034 31034
rect 88046 30982 88098 31034
rect 88110 30982 88162 31034
rect 88174 30982 88226 31034
rect 1982 30438 2034 30490
rect 2046 30438 2098 30490
rect 2110 30438 2162 30490
rect 2174 30438 2226 30490
rect 85982 30438 86034 30490
rect 86046 30438 86098 30490
rect 86110 30438 86162 30490
rect 86174 30438 86226 30490
rect 89982 30438 90034 30490
rect 90046 30438 90098 30490
rect 90110 30438 90162 30490
rect 90174 30438 90226 30490
rect 84752 30311 84804 30320
rect 84752 30277 84761 30311
rect 84761 30277 84795 30311
rect 84795 30277 84804 30311
rect 84752 30268 84804 30277
rect 87236 30268 87288 30320
rect 3982 29894 4034 29946
rect 4046 29894 4098 29946
rect 4110 29894 4162 29946
rect 4174 29894 4226 29946
rect 87982 29894 88034 29946
rect 88046 29894 88098 29946
rect 88110 29894 88162 29946
rect 88174 29894 88226 29946
rect 1982 29350 2034 29402
rect 2046 29350 2098 29402
rect 2110 29350 2162 29402
rect 2174 29350 2226 29402
rect 85982 29350 86034 29402
rect 86046 29350 86098 29402
rect 86110 29350 86162 29402
rect 86174 29350 86226 29402
rect 89982 29350 90034 29402
rect 90046 29350 90098 29402
rect 90110 29350 90162 29402
rect 90174 29350 90226 29402
rect 84568 29248 84620 29300
rect 86500 29248 86552 29300
rect 84752 28976 84804 29028
rect 86960 28976 87012 29028
rect 3982 28806 4034 28858
rect 4046 28806 4098 28858
rect 4110 28806 4162 28858
rect 4174 28806 4226 28858
rect 87982 28806 88034 28858
rect 88046 28806 88098 28858
rect 88110 28806 88162 28858
rect 88174 28806 88226 28858
rect 1982 28262 2034 28314
rect 2046 28262 2098 28314
rect 2110 28262 2162 28314
rect 2174 28262 2226 28314
rect 85982 28262 86034 28314
rect 86046 28262 86098 28314
rect 86110 28262 86162 28314
rect 86174 28262 86226 28314
rect 89982 28262 90034 28314
rect 90046 28262 90098 28314
rect 90110 28262 90162 28314
rect 90174 28262 90226 28314
rect 3982 27718 4034 27770
rect 4046 27718 4098 27770
rect 4110 27718 4162 27770
rect 4174 27718 4226 27770
rect 87982 27718 88034 27770
rect 88046 27718 88098 27770
rect 88110 27718 88162 27770
rect 88174 27718 88226 27770
rect 83924 27616 83976 27668
rect 86960 27616 87012 27668
rect 84568 27548 84620 27600
rect 86408 27548 86460 27600
rect 1982 27174 2034 27226
rect 2046 27174 2098 27226
rect 2110 27174 2162 27226
rect 2174 27174 2226 27226
rect 85982 27174 86034 27226
rect 86046 27174 86098 27226
rect 86110 27174 86162 27226
rect 86174 27174 86226 27226
rect 89982 27174 90034 27226
rect 90046 27174 90098 27226
rect 90110 27174 90162 27226
rect 90174 27174 90226 27226
rect 3982 26630 4034 26682
rect 4046 26630 4098 26682
rect 4110 26630 4162 26682
rect 4174 26630 4226 26682
rect 87982 26630 88034 26682
rect 88046 26630 88098 26682
rect 88110 26630 88162 26682
rect 88174 26630 88226 26682
rect 84568 26528 84620 26580
rect 86316 26528 86368 26580
rect 84016 26256 84068 26308
rect 86960 26256 87012 26308
rect 1982 26086 2034 26138
rect 2046 26086 2098 26138
rect 2110 26086 2162 26138
rect 2174 26086 2226 26138
rect 85982 26086 86034 26138
rect 86046 26086 86098 26138
rect 86110 26086 86162 26138
rect 86174 26086 86226 26138
rect 89982 26086 90034 26138
rect 90046 26086 90098 26138
rect 90110 26086 90162 26138
rect 90174 26086 90226 26138
rect 3982 25542 4034 25594
rect 4046 25542 4098 25594
rect 4110 25542 4162 25594
rect 4174 25542 4226 25594
rect 87982 25542 88034 25594
rect 88046 25542 88098 25594
rect 88110 25542 88162 25594
rect 88174 25542 88226 25594
rect 1982 24998 2034 25050
rect 2046 24998 2098 25050
rect 2110 24998 2162 25050
rect 2174 24998 2226 25050
rect 85982 24998 86034 25050
rect 86046 24998 86098 25050
rect 86110 24998 86162 25050
rect 86174 24998 86226 25050
rect 89982 24998 90034 25050
rect 90046 24998 90098 25050
rect 90110 24998 90162 25050
rect 90174 24998 90226 25050
rect 3982 24454 4034 24506
rect 4046 24454 4098 24506
rect 4110 24454 4162 24506
rect 4174 24454 4226 24506
rect 87982 24454 88034 24506
rect 88046 24454 88098 24506
rect 88110 24454 88162 24506
rect 88174 24454 88226 24506
rect 84292 24352 84344 24404
rect 85856 24352 85908 24404
rect 1982 23910 2034 23962
rect 2046 23910 2098 23962
rect 2110 23910 2162 23962
rect 2174 23910 2226 23962
rect 85982 23910 86034 23962
rect 86046 23910 86098 23962
rect 86110 23910 86162 23962
rect 86174 23910 86226 23962
rect 89982 23910 90034 23962
rect 90046 23910 90098 23962
rect 90110 23910 90162 23962
rect 90174 23910 90226 23962
rect 83372 23536 83424 23588
rect 87052 23536 87104 23588
rect 84108 23468 84160 23520
rect 86960 23468 87012 23520
rect 3982 23366 4034 23418
rect 4046 23366 4098 23418
rect 4110 23366 4162 23418
rect 4174 23366 4226 23418
rect 87982 23366 88034 23418
rect 88046 23366 88098 23418
rect 88110 23366 88162 23418
rect 88174 23366 88226 23418
rect 84292 23264 84344 23316
rect 85672 23264 85724 23316
rect 1982 22822 2034 22874
rect 2046 22822 2098 22874
rect 2110 22822 2162 22874
rect 2174 22822 2226 22874
rect 85982 22822 86034 22874
rect 86046 22822 86098 22874
rect 86110 22822 86162 22874
rect 86174 22822 86226 22874
rect 89982 22822 90034 22874
rect 90046 22822 90098 22874
rect 90110 22822 90162 22874
rect 90174 22822 90226 22874
rect 4712 22423 4764 22432
rect 4712 22389 4721 22423
rect 4721 22389 4755 22423
rect 4755 22389 4764 22423
rect 4712 22380 4764 22389
rect 3982 22278 4034 22330
rect 4046 22278 4098 22330
rect 4110 22278 4162 22330
rect 4174 22278 4226 22330
rect 87982 22278 88034 22330
rect 88046 22278 88098 22330
rect 88110 22278 88162 22330
rect 88174 22278 88226 22330
rect 84568 22176 84620 22228
rect 87144 22176 87196 22228
rect 1982 21734 2034 21786
rect 2046 21734 2098 21786
rect 2110 21734 2162 21786
rect 2174 21734 2226 21786
rect 85982 21734 86034 21786
rect 86046 21734 86098 21786
rect 86110 21734 86162 21786
rect 86174 21734 86226 21786
rect 89982 21734 90034 21786
rect 90046 21734 90098 21786
rect 90110 21734 90162 21786
rect 90174 21734 90226 21786
rect 3982 21190 4034 21242
rect 4046 21190 4098 21242
rect 4110 21190 4162 21242
rect 4174 21190 4226 21242
rect 87982 21190 88034 21242
rect 88046 21190 88098 21242
rect 88110 21190 88162 21242
rect 88174 21190 88226 21242
rect 4804 20859 4856 20868
rect 4804 20825 4813 20859
rect 4813 20825 4847 20859
rect 4847 20825 4856 20859
rect 4804 20816 4856 20825
rect 4988 20816 5040 20868
rect 83280 20748 83332 20800
rect 87880 20748 87932 20800
rect 1982 20646 2034 20698
rect 2046 20646 2098 20698
rect 2110 20646 2162 20698
rect 2174 20646 2226 20698
rect 85982 20646 86034 20698
rect 86046 20646 86098 20698
rect 86110 20646 86162 20698
rect 86174 20646 86226 20698
rect 89982 20646 90034 20698
rect 90046 20646 90098 20698
rect 90110 20646 90162 20698
rect 90174 20646 90226 20698
rect 87236 20544 87288 20596
rect 87880 20544 87932 20596
rect 3982 20102 4034 20154
rect 4046 20102 4098 20154
rect 4110 20102 4162 20154
rect 4174 20102 4226 20154
rect 87982 20102 88034 20154
rect 88046 20102 88098 20154
rect 88110 20102 88162 20154
rect 88174 20102 88226 20154
rect 1982 19558 2034 19610
rect 2046 19558 2098 19610
rect 2110 19558 2162 19610
rect 2174 19558 2226 19610
rect 85982 19558 86034 19610
rect 86046 19558 86098 19610
rect 86110 19558 86162 19610
rect 86174 19558 86226 19610
rect 89982 19558 90034 19610
rect 90046 19558 90098 19610
rect 90110 19558 90162 19610
rect 90174 19558 90226 19610
rect 3982 19014 4034 19066
rect 4046 19014 4098 19066
rect 4110 19014 4162 19066
rect 4174 19014 4226 19066
rect 87982 19014 88034 19066
rect 88046 19014 88098 19066
rect 88110 19014 88162 19066
rect 88174 19014 88226 19066
rect 1982 18470 2034 18522
rect 2046 18470 2098 18522
rect 2110 18470 2162 18522
rect 2174 18470 2226 18522
rect 85982 18470 86034 18522
rect 86046 18470 86098 18522
rect 86110 18470 86162 18522
rect 86174 18470 86226 18522
rect 89982 18470 90034 18522
rect 90046 18470 90098 18522
rect 90110 18470 90162 18522
rect 90174 18470 90226 18522
rect 3982 17926 4034 17978
rect 4046 17926 4098 17978
rect 4110 17926 4162 17978
rect 4174 17926 4226 17978
rect 87982 17926 88034 17978
rect 88046 17926 88098 17978
rect 88110 17926 88162 17978
rect 88174 17926 88226 17978
rect 84476 17731 84528 17740
rect 84476 17697 84485 17731
rect 84485 17697 84519 17731
rect 84519 17697 84528 17731
rect 84476 17688 84528 17697
rect 1982 17382 2034 17434
rect 2046 17382 2098 17434
rect 2110 17382 2162 17434
rect 2174 17382 2226 17434
rect 85982 17382 86034 17434
rect 86046 17382 86098 17434
rect 86110 17382 86162 17434
rect 86174 17382 86226 17434
rect 89982 17382 90034 17434
rect 90046 17382 90098 17434
rect 90110 17382 90162 17434
rect 90174 17382 90226 17434
rect 3982 16838 4034 16890
rect 4046 16838 4098 16890
rect 4110 16838 4162 16890
rect 4174 16838 4226 16890
rect 87982 16838 88034 16890
rect 88046 16838 88098 16890
rect 88110 16838 88162 16890
rect 88174 16838 88226 16890
rect 87052 16532 87104 16584
rect 87236 16532 87288 16584
rect 1982 16294 2034 16346
rect 2046 16294 2098 16346
rect 2110 16294 2162 16346
rect 2174 16294 2226 16346
rect 85982 16294 86034 16346
rect 86046 16294 86098 16346
rect 86110 16294 86162 16346
rect 86174 16294 86226 16346
rect 89982 16294 90034 16346
rect 90046 16294 90098 16346
rect 90110 16294 90162 16346
rect 90174 16294 90226 16346
rect 3982 15750 4034 15802
rect 4046 15750 4098 15802
rect 4110 15750 4162 15802
rect 4174 15750 4226 15802
rect 87982 15750 88034 15802
rect 88046 15750 88098 15802
rect 88110 15750 88162 15802
rect 88174 15750 88226 15802
rect 84476 15308 84528 15360
rect 87144 15308 87196 15360
rect 1982 15206 2034 15258
rect 2046 15206 2098 15258
rect 2110 15206 2162 15258
rect 2174 15206 2226 15258
rect 85982 15206 86034 15258
rect 86046 15206 86098 15258
rect 86110 15206 86162 15258
rect 86174 15206 86226 15258
rect 89982 15206 90034 15258
rect 90046 15206 90098 15258
rect 90110 15206 90162 15258
rect 90174 15206 90226 15258
rect 3982 14662 4034 14714
rect 4046 14662 4098 14714
rect 4110 14662 4162 14714
rect 4174 14662 4226 14714
rect 87982 14662 88034 14714
rect 88046 14662 88098 14714
rect 88110 14662 88162 14714
rect 88174 14662 88226 14714
rect 84660 14603 84712 14612
rect 84660 14569 84669 14603
rect 84669 14569 84703 14603
rect 84703 14569 84712 14603
rect 84660 14560 84712 14569
rect 1982 14118 2034 14170
rect 2046 14118 2098 14170
rect 2110 14118 2162 14170
rect 2174 14118 2226 14170
rect 85982 14118 86034 14170
rect 86046 14118 86098 14170
rect 86110 14118 86162 14170
rect 86174 14118 86226 14170
rect 89982 14118 90034 14170
rect 90046 14118 90098 14170
rect 90110 14118 90162 14170
rect 90174 14118 90226 14170
rect 85304 13923 85356 13932
rect 85304 13889 85313 13923
rect 85313 13889 85347 13923
rect 85347 13889 85356 13923
rect 85304 13880 85356 13889
rect 84660 13855 84712 13864
rect 84660 13821 84669 13855
rect 84669 13821 84703 13855
rect 84703 13821 84712 13855
rect 84660 13812 84712 13821
rect 3982 13574 4034 13626
rect 4046 13574 4098 13626
rect 4110 13574 4162 13626
rect 4174 13574 4226 13626
rect 87982 13574 88034 13626
rect 88046 13574 88098 13626
rect 88110 13574 88162 13626
rect 88174 13574 88226 13626
rect 1982 13030 2034 13082
rect 2046 13030 2098 13082
rect 2110 13030 2162 13082
rect 2174 13030 2226 13082
rect 85982 13030 86034 13082
rect 86046 13030 86098 13082
rect 86110 13030 86162 13082
rect 86174 13030 86226 13082
rect 89982 13030 90034 13082
rect 90046 13030 90098 13082
rect 90110 13030 90162 13082
rect 90174 13030 90226 13082
rect 85304 12588 85356 12640
rect 86960 12588 87012 12640
rect 3982 12486 4034 12538
rect 4046 12486 4098 12538
rect 4110 12486 4162 12538
rect 4174 12486 4226 12538
rect 87982 12486 88034 12538
rect 88046 12486 88098 12538
rect 88110 12486 88162 12538
rect 88174 12486 88226 12538
rect 1982 11942 2034 11994
rect 2046 11942 2098 11994
rect 2110 11942 2162 11994
rect 2174 11942 2226 11994
rect 85982 11942 86034 11994
rect 86046 11942 86098 11994
rect 86110 11942 86162 11994
rect 86174 11942 86226 11994
rect 89982 11942 90034 11994
rect 90046 11942 90098 11994
rect 90110 11942 90162 11994
rect 90174 11942 90226 11994
rect 3982 11398 4034 11450
rect 4046 11398 4098 11450
rect 4110 11398 4162 11450
rect 4174 11398 4226 11450
rect 87982 11398 88034 11450
rect 88046 11398 88098 11450
rect 88110 11398 88162 11450
rect 88174 11398 88226 11450
rect 82912 11024 82964 11076
rect 86960 11024 87012 11076
rect 1982 10854 2034 10906
rect 2046 10854 2098 10906
rect 2110 10854 2162 10906
rect 2174 10854 2226 10906
rect 85982 10854 86034 10906
rect 86046 10854 86098 10906
rect 86110 10854 86162 10906
rect 86174 10854 86226 10906
rect 89982 10854 90034 10906
rect 90046 10854 90098 10906
rect 90110 10854 90162 10906
rect 90174 10854 90226 10906
rect 3982 10310 4034 10362
rect 4046 10310 4098 10362
rect 4110 10310 4162 10362
rect 4174 10310 4226 10362
rect 87982 10310 88034 10362
rect 88046 10310 88098 10362
rect 88110 10310 88162 10362
rect 88174 10310 88226 10362
rect 4436 10115 4488 10124
rect 4436 10081 4445 10115
rect 4445 10081 4479 10115
rect 4479 10081 4488 10115
rect 4436 10072 4488 10081
rect 1982 9766 2034 9818
rect 2046 9766 2098 9818
rect 2110 9766 2162 9818
rect 2174 9766 2226 9818
rect 85982 9766 86034 9818
rect 86046 9766 86098 9818
rect 86110 9766 86162 9818
rect 86174 9766 86226 9818
rect 89982 9766 90034 9818
rect 90046 9766 90098 9818
rect 90110 9766 90162 9818
rect 90174 9766 90226 9818
rect 3982 9222 4034 9274
rect 4046 9222 4098 9274
rect 4110 9222 4162 9274
rect 4174 9222 4226 9274
rect 87982 9222 88034 9274
rect 88046 9222 88098 9274
rect 88110 9222 88162 9274
rect 88174 9222 88226 9274
rect 1982 8678 2034 8730
rect 2046 8678 2098 8730
rect 2110 8678 2162 8730
rect 2174 8678 2226 8730
rect 85982 8678 86034 8730
rect 86046 8678 86098 8730
rect 86110 8678 86162 8730
rect 86174 8678 86226 8730
rect 89982 8678 90034 8730
rect 90046 8678 90098 8730
rect 90110 8678 90162 8730
rect 90174 8678 90226 8730
rect 83096 8304 83148 8356
rect 86960 8304 87012 8356
rect 87052 8236 87104 8288
rect 87604 8236 87656 8288
rect 3982 8134 4034 8186
rect 4046 8134 4098 8186
rect 4110 8134 4162 8186
rect 4174 8134 4226 8186
rect 87982 8134 88034 8186
rect 88046 8134 88098 8186
rect 88110 8134 88162 8186
rect 88174 8134 88226 8186
rect 87788 8032 87840 8084
rect 87972 7964 88024 8016
rect 5356 7760 5408 7812
rect 1982 7590 2034 7642
rect 2046 7590 2098 7642
rect 2110 7590 2162 7642
rect 2174 7590 2226 7642
rect 5356 7556 5408 7608
rect 85982 7590 86034 7642
rect 86046 7590 86098 7642
rect 86110 7590 86162 7642
rect 86174 7590 86226 7642
rect 89982 7590 90034 7642
rect 90046 7590 90098 7642
rect 90110 7590 90162 7642
rect 90174 7590 90226 7642
rect 86960 7488 87012 7540
rect 87236 7488 87288 7540
rect 87328 7488 87380 7540
rect 87788 7488 87840 7540
rect 87236 7352 87288 7404
rect 87696 7352 87748 7404
rect 87696 7216 87748 7268
rect 87972 7216 88024 7268
rect 3982 7046 4034 7098
rect 4046 7046 4098 7098
rect 4110 7046 4162 7098
rect 4174 7046 4226 7098
rect 87982 7046 88034 7098
rect 88046 7046 88098 7098
rect 88110 7046 88162 7098
rect 88174 7046 88226 7098
rect 1982 6502 2034 6554
rect 2046 6502 2098 6554
rect 2110 6502 2162 6554
rect 2174 6502 2226 6554
rect 85982 6502 86034 6554
rect 86046 6502 86098 6554
rect 86110 6502 86162 6554
rect 86174 6502 86226 6554
rect 89982 6502 90034 6554
rect 90046 6502 90098 6554
rect 90110 6502 90162 6554
rect 90174 6502 90226 6554
rect 3982 5958 4034 6010
rect 4046 5958 4098 6010
rect 4110 5958 4162 6010
rect 4174 5958 4226 6010
rect 87982 5958 88034 6010
rect 88046 5958 88098 6010
rect 88110 5958 88162 6010
rect 88174 5958 88226 6010
rect 1982 5414 2034 5466
rect 2046 5414 2098 5466
rect 2110 5414 2162 5466
rect 2174 5414 2226 5466
rect 85982 5414 86034 5466
rect 86046 5414 86098 5466
rect 86110 5414 86162 5466
rect 86174 5414 86226 5466
rect 89982 5414 90034 5466
rect 90046 5414 90098 5466
rect 90110 5414 90162 5466
rect 90174 5414 90226 5466
rect 85856 5312 85908 5364
rect 87052 5312 87104 5364
rect 5448 4972 5500 5024
rect 3982 4870 4034 4922
rect 4046 4870 4098 4922
rect 4110 4870 4162 4922
rect 4174 4870 4226 4922
rect 87982 4870 88034 4922
rect 88046 4870 88098 4922
rect 88110 4870 88162 4922
rect 88174 4870 88226 4922
rect 5080 4768 5132 4820
rect 5724 4768 5776 4820
rect 5172 4700 5224 4752
rect 6000 4700 6052 4752
rect 87696 4700 87748 4752
rect 87972 4700 88024 4752
rect 1982 4326 2034 4378
rect 2046 4326 2098 4378
rect 2110 4326 2162 4378
rect 2174 4326 2226 4378
rect 83188 4360 83240 4412
rect 83464 4360 83516 4412
rect 83648 4335 83700 4344
rect 83648 4301 83657 4335
rect 83657 4301 83691 4335
rect 83691 4301 83700 4335
rect 83648 4292 83700 4301
rect 85982 4326 86034 4378
rect 86046 4326 86098 4378
rect 86110 4326 86162 4378
rect 86174 4326 86226 4378
rect 89982 4326 90034 4378
rect 90046 4326 90098 4378
rect 90110 4326 90162 4378
rect 90174 4326 90226 4378
rect 83648 4156 83700 4208
rect 87052 4156 87104 4208
rect 3884 4088 3936 4140
rect 4528 4088 4580 4140
rect 5908 4088 5960 4140
rect 82820 4088 82872 4140
rect 5724 4020 5776 4072
rect 6368 4020 6420 4072
rect 82728 4020 82780 4072
rect 87696 4020 87748 4072
rect 3792 3884 3844 3936
rect 4804 3927 4856 3936
rect 4804 3893 4813 3927
rect 4813 3893 4847 3927
rect 4847 3893 4856 3927
rect 4804 3884 4856 3893
rect 3982 3782 4034 3834
rect 4046 3782 4098 3834
rect 4110 3782 4162 3834
rect 4174 3782 4226 3834
rect 3332 3723 3384 3732
rect 3332 3689 3341 3723
rect 3341 3689 3375 3723
rect 3375 3689 3384 3723
rect 3332 3680 3384 3689
rect 4804 3723 4856 3732
rect 4804 3689 4813 3723
rect 4813 3689 4847 3723
rect 4847 3689 4856 3723
rect 4804 3680 4856 3689
rect 5632 3680 5684 3732
rect 4436 3655 4488 3664
rect 4436 3621 4445 3655
rect 4445 3621 4479 3655
rect 4479 3621 4488 3655
rect 4436 3612 4488 3621
rect 5816 3612 5868 3664
rect 5632 3476 5684 3528
rect 3608 3340 3660 3392
rect 3792 3340 3844 3392
rect 1982 3238 2034 3290
rect 2046 3238 2098 3290
rect 2110 3238 2162 3290
rect 2174 3238 2226 3290
rect 82636 3952 82688 4004
rect 87972 3952 88024 4004
rect 87982 3782 88034 3834
rect 88046 3782 88098 3834
rect 88110 3782 88162 3834
rect 88174 3782 88226 3834
rect 83464 3680 83516 3732
rect 84936 3680 84988 3732
rect 85396 3723 85448 3732
rect 85396 3689 85405 3723
rect 85405 3689 85439 3723
rect 85439 3689 85448 3723
rect 85396 3680 85448 3689
rect 85856 3544 85908 3596
rect 85764 3476 85816 3528
rect 82544 3408 82596 3460
rect 87052 3408 87104 3460
rect 83648 3272 83700 3324
rect 6736 3204 6788 3256
rect 15292 3204 15344 3256
rect 25044 3204 25096 3256
rect 52552 3204 52604 3256
rect 82820 3204 82872 3256
rect 83556 3247 83608 3256
rect 83556 3213 83565 3247
rect 83565 3213 83599 3247
rect 83599 3213 83608 3247
rect 83556 3204 83608 3213
rect 85982 3238 86034 3290
rect 86046 3238 86098 3290
rect 86110 3238 86162 3290
rect 86174 3238 86226 3290
rect 89982 3238 90034 3290
rect 90046 3238 90098 3290
rect 90110 3238 90162 3290
rect 90174 3238 90226 3290
rect 3516 3136 3568 3188
rect 3700 3179 3752 3188
rect 3700 3145 3709 3179
rect 3709 3145 3743 3179
rect 3743 3145 3752 3179
rect 3700 3136 3752 3145
rect 5540 3136 5592 3188
rect 22100 3136 22152 3188
rect 49976 3136 50028 3188
rect 84936 3136 84988 3188
rect 85764 3179 85816 3188
rect 85764 3145 85773 3179
rect 85773 3145 85807 3179
rect 85807 3145 85816 3179
rect 85764 3136 85816 3145
rect 2504 3111 2556 3120
rect 2504 3077 2513 3111
rect 2513 3077 2547 3111
rect 2547 3077 2556 3111
rect 2504 3068 2556 3077
rect 4528 3068 4580 3120
rect 16304 3068 16356 3120
rect 87328 3068 87380 3120
rect 5908 3000 5960 3052
rect 13912 3000 13964 3052
rect 53472 3000 53524 3052
rect 83188 3000 83240 3052
rect 3792 2932 3844 2984
rect 3884 2932 3936 2984
rect 20720 2932 20772 2984
rect 24124 2864 24176 2916
rect 4344 2796 4396 2848
rect 4620 2796 4672 2848
rect 4896 2796 4948 2848
rect 6920 2796 6972 2848
rect 8116 2796 8168 2848
rect 13912 2796 13964 2848
rect 87604 2932 87656 2984
rect 47768 2864 47820 2916
rect 82452 2864 82504 2916
rect 83004 2864 83056 2916
rect 87328 2864 87380 2916
rect 87512 2864 87564 2916
rect 81440 2796 81492 2848
rect 3982 2694 4034 2746
rect 4046 2694 4098 2746
rect 4110 2694 4162 2746
rect 4174 2694 4226 2746
rect 3884 2592 3936 2644
rect 4712 2592 4764 2644
rect 82452 2728 82504 2780
rect 83556 2771 83608 2780
rect 83556 2737 83565 2771
rect 83565 2737 83599 2771
rect 83599 2737 83608 2771
rect 83556 2728 83608 2737
rect 81348 2660 81400 2712
rect 87982 2694 88034 2746
rect 88046 2694 88098 2746
rect 88110 2694 88162 2746
rect 88174 2694 88226 2746
rect 53840 2592 53892 2644
rect 87328 2592 87380 2644
rect 3240 2524 3292 2576
rect 6184 2456 6236 2508
rect 50344 2524 50396 2576
rect 87144 2524 87196 2576
rect 22652 2456 22704 2508
rect 45928 2456 45980 2508
rect 87236 2456 87288 2508
rect 4160 2388 4212 2440
rect 4988 2388 5040 2440
rect 9772 2320 9824 2372
rect 41420 2388 41472 2440
rect 86960 2388 87012 2440
rect 85028 2363 85080 2372
rect 6276 2252 6328 2304
rect 51356 2252 51408 2304
rect 85028 2329 85037 2363
rect 85037 2329 85071 2363
rect 85071 2329 85080 2363
rect 85028 2320 85080 2329
rect 83556 2252 83608 2304
rect 1982 2150 2034 2202
rect 2046 2150 2098 2202
rect 2110 2150 2162 2202
rect 2174 2150 2226 2202
rect 37464 2184 37516 2236
rect 83924 2184 83976 2236
rect 6184 2116 6236 2168
rect 36176 2116 36228 2168
rect 36268 2116 36320 2168
rect 84016 2116 84068 2168
rect 85982 2150 86034 2202
rect 86046 2150 86098 2202
rect 86110 2150 86162 2202
rect 86174 2150 86226 2202
rect 89982 2150 90034 2202
rect 90046 2150 90098 2202
rect 90110 2150 90162 2202
rect 90174 2150 90226 2202
rect 33968 2048 34020 2100
rect 84108 2048 84160 2100
rect 6276 1980 6328 2032
rect 32680 1980 32732 2032
rect 32772 1980 32824 2032
rect 83372 1980 83424 2032
rect 4160 1912 4212 1964
rect 5264 1912 5316 1964
rect 29092 1912 29144 1964
rect 30472 1912 30524 1964
rect 83280 1912 83332 1964
rect 31668 1844 31720 1896
rect 84568 1844 84620 1896
rect 25780 1776 25832 1828
rect 84476 1776 84528 1828
rect 28172 1708 28224 1760
rect 87420 1708 87472 1760
rect 26976 1640 27028 1692
rect 87052 1640 87104 1692
rect 21088 1572 21140 1624
rect 83188 1572 83240 1624
rect 87880 1572 87932 1624
rect 22284 1504 22336 1556
rect 85304 1504 85356 1556
rect 19248 1436 19300 1488
rect 83096 1436 83148 1488
rect 5448 1368 5500 1420
rect 17500 1368 17552 1420
rect 4620 1300 4672 1352
rect 6460 1300 6512 1352
rect 12440 1300 12492 1352
rect 35532 1300 35584 1352
rect 45928 1300 45980 1352
rect 48228 1300 48280 1352
rect 53840 1300 53892 1352
rect 88248 1436 88300 1488
rect 4804 1232 4856 1284
rect 29000 1232 29052 1284
rect 44916 1232 44968 1284
rect 50344 1232 50396 1284
rect 30288 1164 30340 1216
rect 86316 1164 86368 1216
rect 39948 1096 40000 1148
rect 86592 1096 86644 1148
rect 4436 1028 4488 1080
rect 34520 1028 34572 1080
rect 39856 1028 39908 1080
rect 84752 1028 84804 1080
rect 4528 960 4580 1012
rect 30380 960 30432 1012
rect 41328 960 41380 1012
rect 85488 960 85540 1012
rect 3884 892 3936 944
rect 19340 892 19392 944
rect 24768 892 24820 944
rect 41420 892 41472 944
rect 42708 892 42760 944
rect 86776 892 86828 944
rect 5632 824 5684 876
rect 17960 824 18012 876
rect 44088 824 44140 876
rect 85212 824 85264 876
rect 5172 756 5224 808
rect 27620 756 27672 808
rect 46848 756 46900 808
rect 86684 756 86736 808
rect 3700 688 3752 740
rect 33140 688 33192 740
rect 46756 688 46808 740
rect 85120 688 85172 740
rect 5080 620 5132 672
rect 42800 620 42852 672
rect 49608 620 49660 672
rect 84844 620 84896 672
rect 50988 552 51040 604
rect 82636 552 82688 604
rect 52368 484 52420 536
rect 82728 484 82780 536
rect 53748 416 53800 468
rect 83832 416 83884 468
rect 55128 348 55180 400
rect 83740 348 83792 400
rect 54668 280 54720 332
rect 81440 280 81492 332
rect 55036 212 55088 264
rect 81348 212 81400 264
rect 20628 144 20680 196
rect 86500 144 86552 196
rect 24768 76 24820 128
rect 86408 76 86460 128
<< metal2 >>
rect 1956 189340 2252 189360
rect 2012 189338 2036 189340
rect 2092 189338 2116 189340
rect 2172 189338 2196 189340
rect 2034 189286 2036 189338
rect 2098 189286 2110 189338
rect 2172 189286 2174 189338
rect 2012 189284 2036 189286
rect 2092 189284 2116 189286
rect 2172 189284 2196 189286
rect 1956 189264 2252 189284
rect 85956 189340 86252 189360
rect 86012 189338 86036 189340
rect 86092 189338 86116 189340
rect 86172 189338 86196 189340
rect 86034 189286 86036 189338
rect 86098 189286 86110 189338
rect 86172 189286 86174 189338
rect 86012 189284 86036 189286
rect 86092 189284 86116 189286
rect 86172 189284 86196 189286
rect 85956 189264 86252 189284
rect 89956 189340 90252 189360
rect 90012 189338 90036 189340
rect 90092 189338 90116 189340
rect 90172 189338 90196 189340
rect 90034 189286 90036 189338
rect 90098 189286 90110 189338
rect 90172 189286 90174 189338
rect 90012 189284 90036 189286
rect 90092 189284 90116 189286
rect 90172 189284 90196 189286
rect 89956 189264 90252 189284
rect 75826 189136 75882 189145
rect 75826 189071 75828 189080
rect 75880 189071 75882 189080
rect 84476 189100 84528 189106
rect 75828 189042 75880 189048
rect 84476 189042 84528 189048
rect 3956 188796 4252 188816
rect 4012 188794 4036 188796
rect 4092 188794 4116 188796
rect 4172 188794 4196 188796
rect 4034 188742 4036 188794
rect 4098 188742 4110 188794
rect 4172 188742 4174 188794
rect 4012 188740 4036 188742
rect 4092 188740 4116 188742
rect 4172 188740 4196 188742
rect 3956 188720 4252 188740
rect 1956 188252 2252 188272
rect 2012 188250 2036 188252
rect 2092 188250 2116 188252
rect 2172 188250 2196 188252
rect 2034 188198 2036 188250
rect 2098 188198 2110 188250
rect 2172 188198 2174 188250
rect 2012 188196 2036 188198
rect 2092 188196 2116 188198
rect 2172 188196 2196 188198
rect 1956 188176 2252 188196
rect 3956 187708 4252 187728
rect 4012 187706 4036 187708
rect 4092 187706 4116 187708
rect 4172 187706 4196 187708
rect 4034 187654 4036 187706
rect 4098 187654 4110 187706
rect 4172 187654 4174 187706
rect 4012 187652 4036 187654
rect 4092 187652 4116 187654
rect 4172 187652 4196 187654
rect 3956 187632 4252 187652
rect 79324 187400 79376 187406
rect 79324 187342 79376 187348
rect 1956 187164 2252 187184
rect 2012 187162 2036 187164
rect 2092 187162 2116 187164
rect 2172 187162 2196 187164
rect 2034 187110 2036 187162
rect 2098 187110 2110 187162
rect 2172 187110 2174 187162
rect 2012 187108 2036 187110
rect 2092 187108 2116 187110
rect 2172 187108 2196 187110
rect 1956 187088 2252 187108
rect 79336 187105 79364 187342
rect 84488 187270 84516 189042
rect 87956 188796 88252 188816
rect 88012 188794 88036 188796
rect 88092 188794 88116 188796
rect 88172 188794 88196 188796
rect 88034 188742 88036 188794
rect 88098 188742 88110 188794
rect 88172 188742 88174 188794
rect 88012 188740 88036 188742
rect 88092 188740 88116 188742
rect 88172 188740 88196 188742
rect 87956 188720 88252 188740
rect 85956 188252 86252 188272
rect 86012 188250 86036 188252
rect 86092 188250 86116 188252
rect 86172 188250 86196 188252
rect 86034 188198 86036 188250
rect 86098 188198 86110 188250
rect 86172 188198 86174 188250
rect 86012 188196 86036 188198
rect 86092 188196 86116 188198
rect 86172 188196 86196 188198
rect 85956 188176 86252 188196
rect 89956 188252 90252 188272
rect 90012 188250 90036 188252
rect 90092 188250 90116 188252
rect 90172 188250 90196 188252
rect 90034 188198 90036 188250
rect 90098 188198 90110 188250
rect 90172 188198 90174 188250
rect 90012 188196 90036 188198
rect 90092 188196 90116 188198
rect 90172 188196 90196 188198
rect 89956 188176 90252 188196
rect 87956 187708 88252 187728
rect 88012 187706 88036 187708
rect 88092 187706 88116 187708
rect 88172 187706 88196 187708
rect 88034 187654 88036 187706
rect 88098 187654 88110 187706
rect 88172 187654 88174 187706
rect 88012 187652 88036 187654
rect 88092 187652 88116 187654
rect 88172 187652 88196 187654
rect 87956 187632 88252 187652
rect 84476 187264 84528 187270
rect 84476 187206 84528 187212
rect 79322 187096 79378 187105
rect 79322 187031 79378 187040
rect 79336 186862 79364 187031
rect 79324 186856 79376 186862
rect 79324 186798 79376 186804
rect 4436 186788 4488 186794
rect 4436 186730 4488 186736
rect 3956 186620 4252 186640
rect 4012 186618 4036 186620
rect 4092 186618 4116 186620
rect 4172 186618 4196 186620
rect 4034 186566 4036 186618
rect 4098 186566 4110 186618
rect 4172 186566 4174 186618
rect 4012 186564 4036 186566
rect 4092 186564 4116 186566
rect 4172 186564 4196 186566
rect 3956 186544 4252 186564
rect 1956 186076 2252 186096
rect 2012 186074 2036 186076
rect 2092 186074 2116 186076
rect 2172 186074 2196 186076
rect 2034 186022 2036 186074
rect 2098 186022 2110 186074
rect 2172 186022 2174 186074
rect 2012 186020 2036 186022
rect 2092 186020 2116 186022
rect 2172 186020 2196 186022
rect 1956 186000 2252 186020
rect 3956 185532 4252 185552
rect 4012 185530 4036 185532
rect 4092 185530 4116 185532
rect 4172 185530 4196 185532
rect 4034 185478 4036 185530
rect 4098 185478 4110 185530
rect 4172 185478 4174 185530
rect 4012 185476 4036 185478
rect 4092 185476 4116 185478
rect 4172 185476 4196 185478
rect 3956 185456 4252 185476
rect 1956 184988 2252 185008
rect 2012 184986 2036 184988
rect 2092 184986 2116 184988
rect 2172 184986 2196 184988
rect 2034 184934 2036 184986
rect 2098 184934 2110 184986
rect 2172 184934 2174 184986
rect 2012 184932 2036 184934
rect 2092 184932 2116 184934
rect 2172 184932 2196 184934
rect 1956 184912 2252 184932
rect 3956 184444 4252 184464
rect 4012 184442 4036 184444
rect 4092 184442 4116 184444
rect 4172 184442 4196 184444
rect 4034 184390 4036 184442
rect 4098 184390 4110 184442
rect 4172 184390 4174 184442
rect 4012 184388 4036 184390
rect 4092 184388 4116 184390
rect 4172 184388 4196 184390
rect 3956 184368 4252 184388
rect 1956 183900 2252 183920
rect 2012 183898 2036 183900
rect 2092 183898 2116 183900
rect 2172 183898 2196 183900
rect 2034 183846 2036 183898
rect 2098 183846 2110 183898
rect 2172 183846 2174 183898
rect 2012 183844 2036 183846
rect 2092 183844 2116 183846
rect 2172 183844 2196 183846
rect 1956 183824 2252 183844
rect 3956 183356 4252 183376
rect 4012 183354 4036 183356
rect 4092 183354 4116 183356
rect 4172 183354 4196 183356
rect 4034 183302 4036 183354
rect 4098 183302 4110 183354
rect 4172 183302 4174 183354
rect 4012 183300 4036 183302
rect 4092 183300 4116 183302
rect 4172 183300 4196 183302
rect 3956 183280 4252 183300
rect 1956 182812 2252 182832
rect 2012 182810 2036 182812
rect 2092 182810 2116 182812
rect 2172 182810 2196 182812
rect 2034 182758 2036 182810
rect 2098 182758 2110 182810
rect 2172 182758 2174 182810
rect 2012 182756 2036 182758
rect 2092 182756 2116 182758
rect 2172 182756 2196 182758
rect 1956 182736 2252 182756
rect 3956 182268 4252 182288
rect 4012 182266 4036 182268
rect 4092 182266 4116 182268
rect 4172 182266 4196 182268
rect 4034 182214 4036 182266
rect 4098 182214 4110 182266
rect 4172 182214 4174 182266
rect 4012 182212 4036 182214
rect 4092 182212 4116 182214
rect 4172 182212 4196 182214
rect 3956 182192 4252 182212
rect 1956 181724 2252 181744
rect 2012 181722 2036 181724
rect 2092 181722 2116 181724
rect 2172 181722 2196 181724
rect 2034 181670 2036 181722
rect 2098 181670 2110 181722
rect 2172 181670 2174 181722
rect 2012 181668 2036 181670
rect 2092 181668 2116 181670
rect 2172 181668 2196 181670
rect 1956 181648 2252 181668
rect 3956 181180 4252 181200
rect 4012 181178 4036 181180
rect 4092 181178 4116 181180
rect 4172 181178 4196 181180
rect 4034 181126 4036 181178
rect 4098 181126 4110 181178
rect 4172 181126 4174 181178
rect 4012 181124 4036 181126
rect 4092 181124 4116 181126
rect 4172 181124 4196 181126
rect 3956 181104 4252 181124
rect 1956 180636 2252 180656
rect 2012 180634 2036 180636
rect 2092 180634 2116 180636
rect 2172 180634 2196 180636
rect 2034 180582 2036 180634
rect 2098 180582 2110 180634
rect 2172 180582 2174 180634
rect 2012 180580 2036 180582
rect 2092 180580 2116 180582
rect 2172 180580 2196 180582
rect 1956 180560 2252 180580
rect 3956 180092 4252 180112
rect 4012 180090 4036 180092
rect 4092 180090 4116 180092
rect 4172 180090 4196 180092
rect 4034 180038 4036 180090
rect 4098 180038 4110 180090
rect 4172 180038 4174 180090
rect 4012 180036 4036 180038
rect 4092 180036 4116 180038
rect 4172 180036 4196 180038
rect 3956 180016 4252 180036
rect 1956 179548 2252 179568
rect 2012 179546 2036 179548
rect 2092 179546 2116 179548
rect 2172 179546 2196 179548
rect 2034 179494 2036 179546
rect 2098 179494 2110 179546
rect 2172 179494 2174 179546
rect 2012 179492 2036 179494
rect 2092 179492 2116 179494
rect 2172 179492 2196 179494
rect 1956 179472 2252 179492
rect 3956 179004 4252 179024
rect 4012 179002 4036 179004
rect 4092 179002 4116 179004
rect 4172 179002 4196 179004
rect 4034 178950 4036 179002
rect 4098 178950 4110 179002
rect 4172 178950 4174 179002
rect 4012 178948 4036 178950
rect 4092 178948 4116 178950
rect 4172 178948 4196 178950
rect 3956 178928 4252 178948
rect 1956 178460 2252 178480
rect 2012 178458 2036 178460
rect 2092 178458 2116 178460
rect 2172 178458 2196 178460
rect 2034 178406 2036 178458
rect 2098 178406 2110 178458
rect 2172 178406 2174 178458
rect 2012 178404 2036 178406
rect 2092 178404 2116 178406
rect 2172 178404 2196 178406
rect 1956 178384 2252 178404
rect 3956 177916 4252 177936
rect 4012 177914 4036 177916
rect 4092 177914 4116 177916
rect 4172 177914 4196 177916
rect 4034 177862 4036 177914
rect 4098 177862 4110 177914
rect 4172 177862 4174 177914
rect 4012 177860 4036 177862
rect 4092 177860 4116 177862
rect 4172 177860 4196 177862
rect 3956 177840 4252 177860
rect 1956 177372 2252 177392
rect 2012 177370 2036 177372
rect 2092 177370 2116 177372
rect 2172 177370 2196 177372
rect 2034 177318 2036 177370
rect 2098 177318 2110 177370
rect 2172 177318 2174 177370
rect 2012 177316 2036 177318
rect 2092 177316 2116 177318
rect 2172 177316 2196 177318
rect 1956 177296 2252 177316
rect 3956 176828 4252 176848
rect 4012 176826 4036 176828
rect 4092 176826 4116 176828
rect 4172 176826 4196 176828
rect 4034 176774 4036 176826
rect 4098 176774 4110 176826
rect 4172 176774 4174 176826
rect 4012 176772 4036 176774
rect 4092 176772 4116 176774
rect 4172 176772 4196 176774
rect 3956 176752 4252 176772
rect 1956 176284 2252 176304
rect 2012 176282 2036 176284
rect 2092 176282 2116 176284
rect 2172 176282 2196 176284
rect 2034 176230 2036 176282
rect 2098 176230 2110 176282
rect 2172 176230 2174 176282
rect 2012 176228 2036 176230
rect 2092 176228 2116 176230
rect 2172 176228 2196 176230
rect 1956 176208 2252 176228
rect 3956 175740 4252 175760
rect 4012 175738 4036 175740
rect 4092 175738 4116 175740
rect 4172 175738 4196 175740
rect 4034 175686 4036 175738
rect 4098 175686 4110 175738
rect 4172 175686 4174 175738
rect 4012 175684 4036 175686
rect 4092 175684 4116 175686
rect 4172 175684 4196 175686
rect 3956 175664 4252 175684
rect 1956 175196 2252 175216
rect 2012 175194 2036 175196
rect 2092 175194 2116 175196
rect 2172 175194 2196 175196
rect 2034 175142 2036 175194
rect 2098 175142 2110 175194
rect 2172 175142 2174 175194
rect 2012 175140 2036 175142
rect 2092 175140 2116 175142
rect 2172 175140 2196 175142
rect 1956 175120 2252 175140
rect 3956 174652 4252 174672
rect 4012 174650 4036 174652
rect 4092 174650 4116 174652
rect 4172 174650 4196 174652
rect 4034 174598 4036 174650
rect 4098 174598 4110 174650
rect 4172 174598 4174 174650
rect 4012 174596 4036 174598
rect 4092 174596 4116 174598
rect 4172 174596 4196 174598
rect 3956 174576 4252 174596
rect 1956 174108 2252 174128
rect 2012 174106 2036 174108
rect 2092 174106 2116 174108
rect 2172 174106 2196 174108
rect 2034 174054 2036 174106
rect 2098 174054 2110 174106
rect 2172 174054 2174 174106
rect 2012 174052 2036 174054
rect 2092 174052 2116 174054
rect 2172 174052 2196 174054
rect 1956 174032 2252 174052
rect 3956 173564 4252 173584
rect 4012 173562 4036 173564
rect 4092 173562 4116 173564
rect 4172 173562 4196 173564
rect 4034 173510 4036 173562
rect 4098 173510 4110 173562
rect 4172 173510 4174 173562
rect 4012 173508 4036 173510
rect 4092 173508 4116 173510
rect 4172 173508 4196 173510
rect 3956 173488 4252 173508
rect 1956 173020 2252 173040
rect 2012 173018 2036 173020
rect 2092 173018 2116 173020
rect 2172 173018 2196 173020
rect 2034 172966 2036 173018
rect 2098 172966 2110 173018
rect 2172 172966 2174 173018
rect 2012 172964 2036 172966
rect 2092 172964 2116 172966
rect 2172 172964 2196 172966
rect 1956 172944 2252 172964
rect 3956 172476 4252 172496
rect 4012 172474 4036 172476
rect 4092 172474 4116 172476
rect 4172 172474 4196 172476
rect 4034 172422 4036 172474
rect 4098 172422 4110 172474
rect 4172 172422 4174 172474
rect 4012 172420 4036 172422
rect 4092 172420 4116 172422
rect 4172 172420 4196 172422
rect 3956 172400 4252 172420
rect 1956 171932 2252 171952
rect 2012 171930 2036 171932
rect 2092 171930 2116 171932
rect 2172 171930 2196 171932
rect 2034 171878 2036 171930
rect 2098 171878 2110 171930
rect 2172 171878 2174 171930
rect 2012 171876 2036 171878
rect 2092 171876 2116 171878
rect 2172 171876 2196 171878
rect 1956 171856 2252 171876
rect 3956 171388 4252 171408
rect 4012 171386 4036 171388
rect 4092 171386 4116 171388
rect 4172 171386 4196 171388
rect 4034 171334 4036 171386
rect 4098 171334 4110 171386
rect 4172 171334 4174 171386
rect 4012 171332 4036 171334
rect 4092 171332 4116 171334
rect 4172 171332 4196 171334
rect 3956 171312 4252 171332
rect 1956 170844 2252 170864
rect 2012 170842 2036 170844
rect 2092 170842 2116 170844
rect 2172 170842 2196 170844
rect 2034 170790 2036 170842
rect 2098 170790 2110 170842
rect 2172 170790 2174 170842
rect 2012 170788 2036 170790
rect 2092 170788 2116 170790
rect 2172 170788 2196 170790
rect 1956 170768 2252 170788
rect 3956 170300 4252 170320
rect 4012 170298 4036 170300
rect 4092 170298 4116 170300
rect 4172 170298 4196 170300
rect 4034 170246 4036 170298
rect 4098 170246 4110 170298
rect 4172 170246 4174 170298
rect 4012 170244 4036 170246
rect 4092 170244 4116 170246
rect 4172 170244 4196 170246
rect 3956 170224 4252 170244
rect 1956 169756 2252 169776
rect 2012 169754 2036 169756
rect 2092 169754 2116 169756
rect 2172 169754 2196 169756
rect 2034 169702 2036 169754
rect 2098 169702 2110 169754
rect 2172 169702 2174 169754
rect 2012 169700 2036 169702
rect 2092 169700 2116 169702
rect 2172 169700 2196 169702
rect 1956 169680 2252 169700
rect 3956 169212 4252 169232
rect 4012 169210 4036 169212
rect 4092 169210 4116 169212
rect 4172 169210 4196 169212
rect 4034 169158 4036 169210
rect 4098 169158 4110 169210
rect 4172 169158 4174 169210
rect 4012 169156 4036 169158
rect 4092 169156 4116 169158
rect 4172 169156 4196 169158
rect 3956 169136 4252 169156
rect 1956 168668 2252 168688
rect 2012 168666 2036 168668
rect 2092 168666 2116 168668
rect 2172 168666 2196 168668
rect 2034 168614 2036 168666
rect 2098 168614 2110 168666
rect 2172 168614 2174 168666
rect 2012 168612 2036 168614
rect 2092 168612 2116 168614
rect 2172 168612 2196 168614
rect 1956 168592 2252 168612
rect 3956 168124 4252 168144
rect 4012 168122 4036 168124
rect 4092 168122 4116 168124
rect 4172 168122 4196 168124
rect 4034 168070 4036 168122
rect 4098 168070 4110 168122
rect 4172 168070 4174 168122
rect 4012 168068 4036 168070
rect 4092 168068 4116 168070
rect 4172 168068 4196 168070
rect 3956 168048 4252 168068
rect 1956 167580 2252 167600
rect 2012 167578 2036 167580
rect 2092 167578 2116 167580
rect 2172 167578 2196 167580
rect 2034 167526 2036 167578
rect 2098 167526 2110 167578
rect 2172 167526 2174 167578
rect 2012 167524 2036 167526
rect 2092 167524 2116 167526
rect 2172 167524 2196 167526
rect 1956 167504 2252 167524
rect 3956 167036 4252 167056
rect 4012 167034 4036 167036
rect 4092 167034 4116 167036
rect 4172 167034 4196 167036
rect 4034 166982 4036 167034
rect 4098 166982 4110 167034
rect 4172 166982 4174 167034
rect 4012 166980 4036 166982
rect 4092 166980 4116 166982
rect 4172 166980 4196 166982
rect 3956 166960 4252 166980
rect 1956 166492 2252 166512
rect 2012 166490 2036 166492
rect 2092 166490 2116 166492
rect 2172 166490 2196 166492
rect 2034 166438 2036 166490
rect 2098 166438 2110 166490
rect 2172 166438 2174 166490
rect 2012 166436 2036 166438
rect 2092 166436 2116 166438
rect 2172 166436 2196 166438
rect 1956 166416 2252 166436
rect 3956 165948 4252 165968
rect 4012 165946 4036 165948
rect 4092 165946 4116 165948
rect 4172 165946 4196 165948
rect 4034 165894 4036 165946
rect 4098 165894 4110 165946
rect 4172 165894 4174 165946
rect 4012 165892 4036 165894
rect 4092 165892 4116 165894
rect 4172 165892 4196 165894
rect 3956 165872 4252 165892
rect 1956 165404 2252 165424
rect 2012 165402 2036 165404
rect 2092 165402 2116 165404
rect 2172 165402 2196 165404
rect 2034 165350 2036 165402
rect 2098 165350 2110 165402
rect 2172 165350 2174 165402
rect 2012 165348 2036 165350
rect 2092 165348 2116 165350
rect 2172 165348 2196 165350
rect 1956 165328 2252 165348
rect 3956 164860 4252 164880
rect 4012 164858 4036 164860
rect 4092 164858 4116 164860
rect 4172 164858 4196 164860
rect 4034 164806 4036 164858
rect 4098 164806 4110 164858
rect 4172 164806 4174 164858
rect 4012 164804 4036 164806
rect 4092 164804 4116 164806
rect 4172 164804 4196 164806
rect 3956 164784 4252 164804
rect 1956 164316 2252 164336
rect 2012 164314 2036 164316
rect 2092 164314 2116 164316
rect 2172 164314 2196 164316
rect 2034 164262 2036 164314
rect 2098 164262 2110 164314
rect 2172 164262 2174 164314
rect 2012 164260 2036 164262
rect 2092 164260 2116 164262
rect 2172 164260 2196 164262
rect 1956 164240 2252 164260
rect 3956 163772 4252 163792
rect 4012 163770 4036 163772
rect 4092 163770 4116 163772
rect 4172 163770 4196 163772
rect 4034 163718 4036 163770
rect 4098 163718 4110 163770
rect 4172 163718 4174 163770
rect 4012 163716 4036 163718
rect 4092 163716 4116 163718
rect 4172 163716 4196 163718
rect 3956 163696 4252 163716
rect 1956 163228 2252 163248
rect 2012 163226 2036 163228
rect 2092 163226 2116 163228
rect 2172 163226 2196 163228
rect 2034 163174 2036 163226
rect 2098 163174 2110 163226
rect 2172 163174 2174 163226
rect 2012 163172 2036 163174
rect 2092 163172 2116 163174
rect 2172 163172 2196 163174
rect 1956 163152 2252 163172
rect 3956 162684 4252 162704
rect 4012 162682 4036 162684
rect 4092 162682 4116 162684
rect 4172 162682 4196 162684
rect 4034 162630 4036 162682
rect 4098 162630 4110 162682
rect 4172 162630 4174 162682
rect 4012 162628 4036 162630
rect 4092 162628 4116 162630
rect 4172 162628 4196 162630
rect 3956 162608 4252 162628
rect 1956 162140 2252 162160
rect 2012 162138 2036 162140
rect 2092 162138 2116 162140
rect 2172 162138 2196 162140
rect 2034 162086 2036 162138
rect 2098 162086 2110 162138
rect 2172 162086 2174 162138
rect 2012 162084 2036 162086
rect 2092 162084 2116 162086
rect 2172 162084 2196 162086
rect 1956 162064 2252 162084
rect 3956 161596 4252 161616
rect 4012 161594 4036 161596
rect 4092 161594 4116 161596
rect 4172 161594 4196 161596
rect 4034 161542 4036 161594
rect 4098 161542 4110 161594
rect 4172 161542 4174 161594
rect 4012 161540 4036 161542
rect 4092 161540 4116 161542
rect 4172 161540 4196 161542
rect 3956 161520 4252 161540
rect 1956 161052 2252 161072
rect 2012 161050 2036 161052
rect 2092 161050 2116 161052
rect 2172 161050 2196 161052
rect 2034 160998 2036 161050
rect 2098 160998 2110 161050
rect 2172 160998 2174 161050
rect 2012 160996 2036 160998
rect 2092 160996 2116 160998
rect 2172 160996 2196 160998
rect 1956 160976 2252 160996
rect 3956 160508 4252 160528
rect 4012 160506 4036 160508
rect 4092 160506 4116 160508
rect 4172 160506 4196 160508
rect 4034 160454 4036 160506
rect 4098 160454 4110 160506
rect 4172 160454 4174 160506
rect 4012 160452 4036 160454
rect 4092 160452 4116 160454
rect 4172 160452 4196 160454
rect 3956 160432 4252 160452
rect 1956 159964 2252 159984
rect 2012 159962 2036 159964
rect 2092 159962 2116 159964
rect 2172 159962 2196 159964
rect 2034 159910 2036 159962
rect 2098 159910 2110 159962
rect 2172 159910 2174 159962
rect 2012 159908 2036 159910
rect 2092 159908 2116 159910
rect 2172 159908 2196 159910
rect 1956 159888 2252 159908
rect 3956 159420 4252 159440
rect 4012 159418 4036 159420
rect 4092 159418 4116 159420
rect 4172 159418 4196 159420
rect 4034 159366 4036 159418
rect 4098 159366 4110 159418
rect 4172 159366 4174 159418
rect 4012 159364 4036 159366
rect 4092 159364 4116 159366
rect 4172 159364 4196 159366
rect 3956 159344 4252 159364
rect 1956 158876 2252 158896
rect 2012 158874 2036 158876
rect 2092 158874 2116 158876
rect 2172 158874 2196 158876
rect 2034 158822 2036 158874
rect 2098 158822 2110 158874
rect 2172 158822 2174 158874
rect 2012 158820 2036 158822
rect 2092 158820 2116 158822
rect 2172 158820 2196 158822
rect 1956 158800 2252 158820
rect 3956 158332 4252 158352
rect 4012 158330 4036 158332
rect 4092 158330 4116 158332
rect 4172 158330 4196 158332
rect 4034 158278 4036 158330
rect 4098 158278 4110 158330
rect 4172 158278 4174 158330
rect 4012 158276 4036 158278
rect 4092 158276 4116 158278
rect 4172 158276 4196 158278
rect 3956 158256 4252 158276
rect 1956 157788 2252 157808
rect 2012 157786 2036 157788
rect 2092 157786 2116 157788
rect 2172 157786 2196 157788
rect 2034 157734 2036 157786
rect 2098 157734 2110 157786
rect 2172 157734 2174 157786
rect 2012 157732 2036 157734
rect 2092 157732 2116 157734
rect 2172 157732 2196 157734
rect 1956 157712 2252 157732
rect 3956 157244 4252 157264
rect 4012 157242 4036 157244
rect 4092 157242 4116 157244
rect 4172 157242 4196 157244
rect 4034 157190 4036 157242
rect 4098 157190 4110 157242
rect 4172 157190 4174 157242
rect 4012 157188 4036 157190
rect 4092 157188 4116 157190
rect 4172 157188 4196 157190
rect 3956 157168 4252 157188
rect 1956 156700 2252 156720
rect 2012 156698 2036 156700
rect 2092 156698 2116 156700
rect 2172 156698 2196 156700
rect 2034 156646 2036 156698
rect 2098 156646 2110 156698
rect 2172 156646 2174 156698
rect 2012 156644 2036 156646
rect 2092 156644 2116 156646
rect 2172 156644 2196 156646
rect 1956 156624 2252 156644
rect 3956 156156 4252 156176
rect 4012 156154 4036 156156
rect 4092 156154 4116 156156
rect 4172 156154 4196 156156
rect 4034 156102 4036 156154
rect 4098 156102 4110 156154
rect 4172 156102 4174 156154
rect 4012 156100 4036 156102
rect 4092 156100 4116 156102
rect 4172 156100 4196 156102
rect 3956 156080 4252 156100
rect 1956 155612 2252 155632
rect 2012 155610 2036 155612
rect 2092 155610 2116 155612
rect 2172 155610 2196 155612
rect 2034 155558 2036 155610
rect 2098 155558 2110 155610
rect 2172 155558 2174 155610
rect 2012 155556 2036 155558
rect 2092 155556 2116 155558
rect 2172 155556 2196 155558
rect 1956 155536 2252 155556
rect 3956 155068 4252 155088
rect 4012 155066 4036 155068
rect 4092 155066 4116 155068
rect 4172 155066 4196 155068
rect 4034 155014 4036 155066
rect 4098 155014 4110 155066
rect 4172 155014 4174 155066
rect 4012 155012 4036 155014
rect 4092 155012 4116 155014
rect 4172 155012 4196 155014
rect 3956 154992 4252 155012
rect 1956 154524 2252 154544
rect 2012 154522 2036 154524
rect 2092 154522 2116 154524
rect 2172 154522 2196 154524
rect 2034 154470 2036 154522
rect 2098 154470 2110 154522
rect 2172 154470 2174 154522
rect 2012 154468 2036 154470
rect 2092 154468 2116 154470
rect 2172 154468 2196 154470
rect 1956 154448 2252 154468
rect 3956 153980 4252 154000
rect 4012 153978 4036 153980
rect 4092 153978 4116 153980
rect 4172 153978 4196 153980
rect 4034 153926 4036 153978
rect 4098 153926 4110 153978
rect 4172 153926 4174 153978
rect 4012 153924 4036 153926
rect 4092 153924 4116 153926
rect 4172 153924 4196 153926
rect 3956 153904 4252 153924
rect 1956 153436 2252 153456
rect 2012 153434 2036 153436
rect 2092 153434 2116 153436
rect 2172 153434 2196 153436
rect 2034 153382 2036 153434
rect 2098 153382 2110 153434
rect 2172 153382 2174 153434
rect 2012 153380 2036 153382
rect 2092 153380 2116 153382
rect 2172 153380 2196 153382
rect 1956 153360 2252 153380
rect 3956 152892 4252 152912
rect 4012 152890 4036 152892
rect 4092 152890 4116 152892
rect 4172 152890 4196 152892
rect 4034 152838 4036 152890
rect 4098 152838 4110 152890
rect 4172 152838 4174 152890
rect 4012 152836 4036 152838
rect 4092 152836 4116 152838
rect 4172 152836 4196 152838
rect 3956 152816 4252 152836
rect 1956 152348 2252 152368
rect 2012 152346 2036 152348
rect 2092 152346 2116 152348
rect 2172 152346 2196 152348
rect 2034 152294 2036 152346
rect 2098 152294 2110 152346
rect 2172 152294 2174 152346
rect 2012 152292 2036 152294
rect 2092 152292 2116 152294
rect 2172 152292 2196 152294
rect 1956 152272 2252 152292
rect 3956 151804 4252 151824
rect 4012 151802 4036 151804
rect 4092 151802 4116 151804
rect 4172 151802 4196 151804
rect 4034 151750 4036 151802
rect 4098 151750 4110 151802
rect 4172 151750 4174 151802
rect 4012 151748 4036 151750
rect 4092 151748 4116 151750
rect 4172 151748 4196 151750
rect 3956 151728 4252 151748
rect 1956 151260 2252 151280
rect 2012 151258 2036 151260
rect 2092 151258 2116 151260
rect 2172 151258 2196 151260
rect 2034 151206 2036 151258
rect 2098 151206 2110 151258
rect 2172 151206 2174 151258
rect 2012 151204 2036 151206
rect 2092 151204 2116 151206
rect 2172 151204 2196 151206
rect 1956 151184 2252 151204
rect 3956 150716 4252 150736
rect 4012 150714 4036 150716
rect 4092 150714 4116 150716
rect 4172 150714 4196 150716
rect 4034 150662 4036 150714
rect 4098 150662 4110 150714
rect 4172 150662 4174 150714
rect 4012 150660 4036 150662
rect 4092 150660 4116 150662
rect 4172 150660 4196 150662
rect 3956 150640 4252 150660
rect 1956 150172 2252 150192
rect 2012 150170 2036 150172
rect 2092 150170 2116 150172
rect 2172 150170 2196 150172
rect 2034 150118 2036 150170
rect 2098 150118 2110 150170
rect 2172 150118 2174 150170
rect 2012 150116 2036 150118
rect 2092 150116 2116 150118
rect 2172 150116 2196 150118
rect 1956 150096 2252 150116
rect 3956 149628 4252 149648
rect 4012 149626 4036 149628
rect 4092 149626 4116 149628
rect 4172 149626 4196 149628
rect 4034 149574 4036 149626
rect 4098 149574 4110 149626
rect 4172 149574 4174 149626
rect 4012 149572 4036 149574
rect 4092 149572 4116 149574
rect 4172 149572 4196 149574
rect 3956 149552 4252 149572
rect 1956 149084 2252 149104
rect 2012 149082 2036 149084
rect 2092 149082 2116 149084
rect 2172 149082 2196 149084
rect 2034 149030 2036 149082
rect 2098 149030 2110 149082
rect 2172 149030 2174 149082
rect 2012 149028 2036 149030
rect 2092 149028 2116 149030
rect 2172 149028 2196 149030
rect 1956 149008 2252 149028
rect 3956 148540 4252 148560
rect 4012 148538 4036 148540
rect 4092 148538 4116 148540
rect 4172 148538 4196 148540
rect 4034 148486 4036 148538
rect 4098 148486 4110 148538
rect 4172 148486 4174 148538
rect 4012 148484 4036 148486
rect 4092 148484 4116 148486
rect 4172 148484 4196 148486
rect 3956 148464 4252 148484
rect 1956 147996 2252 148016
rect 2012 147994 2036 147996
rect 2092 147994 2116 147996
rect 2172 147994 2196 147996
rect 2034 147942 2036 147994
rect 2098 147942 2110 147994
rect 2172 147942 2174 147994
rect 2012 147940 2036 147942
rect 2092 147940 2116 147942
rect 2172 147940 2196 147942
rect 1956 147920 2252 147940
rect 3956 147452 4252 147472
rect 4012 147450 4036 147452
rect 4092 147450 4116 147452
rect 4172 147450 4196 147452
rect 4034 147398 4036 147450
rect 4098 147398 4110 147450
rect 4172 147398 4174 147450
rect 4012 147396 4036 147398
rect 4092 147396 4116 147398
rect 4172 147396 4196 147398
rect 3956 147376 4252 147396
rect 1956 146908 2252 146928
rect 2012 146906 2036 146908
rect 2092 146906 2116 146908
rect 2172 146906 2196 146908
rect 2034 146854 2036 146906
rect 2098 146854 2110 146906
rect 2172 146854 2174 146906
rect 2012 146852 2036 146854
rect 2092 146852 2116 146854
rect 2172 146852 2196 146854
rect 1956 146832 2252 146852
rect 3956 146364 4252 146384
rect 4012 146362 4036 146364
rect 4092 146362 4116 146364
rect 4172 146362 4196 146364
rect 4034 146310 4036 146362
rect 4098 146310 4110 146362
rect 4172 146310 4174 146362
rect 4012 146308 4036 146310
rect 4092 146308 4116 146310
rect 4172 146308 4196 146310
rect 3956 146288 4252 146308
rect 1956 145820 2252 145840
rect 2012 145818 2036 145820
rect 2092 145818 2116 145820
rect 2172 145818 2196 145820
rect 2034 145766 2036 145818
rect 2098 145766 2110 145818
rect 2172 145766 2174 145818
rect 2012 145764 2036 145766
rect 2092 145764 2116 145766
rect 2172 145764 2196 145766
rect 1956 145744 2252 145764
rect 3956 145276 4252 145296
rect 4012 145274 4036 145276
rect 4092 145274 4116 145276
rect 4172 145274 4196 145276
rect 4034 145222 4036 145274
rect 4098 145222 4110 145274
rect 4172 145222 4174 145274
rect 4012 145220 4036 145222
rect 4092 145220 4116 145222
rect 4172 145220 4196 145222
rect 3956 145200 4252 145220
rect 1956 144732 2252 144752
rect 2012 144730 2036 144732
rect 2092 144730 2116 144732
rect 2172 144730 2196 144732
rect 2034 144678 2036 144730
rect 2098 144678 2110 144730
rect 2172 144678 2174 144730
rect 2012 144676 2036 144678
rect 2092 144676 2116 144678
rect 2172 144676 2196 144678
rect 1956 144656 2252 144676
rect 3956 144188 4252 144208
rect 4012 144186 4036 144188
rect 4092 144186 4116 144188
rect 4172 144186 4196 144188
rect 4034 144134 4036 144186
rect 4098 144134 4110 144186
rect 4172 144134 4174 144186
rect 4012 144132 4036 144134
rect 4092 144132 4116 144134
rect 4172 144132 4196 144134
rect 3956 144112 4252 144132
rect 1956 143644 2252 143664
rect 2012 143642 2036 143644
rect 2092 143642 2116 143644
rect 2172 143642 2196 143644
rect 2034 143590 2036 143642
rect 2098 143590 2110 143642
rect 2172 143590 2174 143642
rect 2012 143588 2036 143590
rect 2092 143588 2116 143590
rect 2172 143588 2196 143590
rect 1956 143568 2252 143588
rect 3956 143100 4252 143120
rect 4012 143098 4036 143100
rect 4092 143098 4116 143100
rect 4172 143098 4196 143100
rect 4034 143046 4036 143098
rect 4098 143046 4110 143098
rect 4172 143046 4174 143098
rect 4012 143044 4036 143046
rect 4092 143044 4116 143046
rect 4172 143044 4196 143046
rect 3956 143024 4252 143044
rect 1956 142556 2252 142576
rect 2012 142554 2036 142556
rect 2092 142554 2116 142556
rect 2172 142554 2196 142556
rect 2034 142502 2036 142554
rect 2098 142502 2110 142554
rect 2172 142502 2174 142554
rect 2012 142500 2036 142502
rect 2092 142500 2116 142502
rect 2172 142500 2196 142502
rect 1956 142480 2252 142500
rect 3956 142012 4252 142032
rect 4012 142010 4036 142012
rect 4092 142010 4116 142012
rect 4172 142010 4196 142012
rect 4034 141958 4036 142010
rect 4098 141958 4110 142010
rect 4172 141958 4174 142010
rect 4012 141956 4036 141958
rect 4092 141956 4116 141958
rect 4172 141956 4196 141958
rect 3956 141936 4252 141956
rect 1956 141468 2252 141488
rect 2012 141466 2036 141468
rect 2092 141466 2116 141468
rect 2172 141466 2196 141468
rect 2034 141414 2036 141466
rect 2098 141414 2110 141466
rect 2172 141414 2174 141466
rect 2012 141412 2036 141414
rect 2092 141412 2116 141414
rect 2172 141412 2196 141414
rect 1956 141392 2252 141412
rect 3956 140924 4252 140944
rect 4012 140922 4036 140924
rect 4092 140922 4116 140924
rect 4172 140922 4196 140924
rect 4034 140870 4036 140922
rect 4098 140870 4110 140922
rect 4172 140870 4174 140922
rect 4012 140868 4036 140870
rect 4092 140868 4116 140870
rect 4172 140868 4196 140870
rect 3956 140848 4252 140868
rect 1956 140380 2252 140400
rect 2012 140378 2036 140380
rect 2092 140378 2116 140380
rect 2172 140378 2196 140380
rect 2034 140326 2036 140378
rect 2098 140326 2110 140378
rect 2172 140326 2174 140378
rect 2012 140324 2036 140326
rect 2092 140324 2116 140326
rect 2172 140324 2196 140326
rect 1956 140304 2252 140324
rect 3956 139836 4252 139856
rect 4012 139834 4036 139836
rect 4092 139834 4116 139836
rect 4172 139834 4196 139836
rect 4034 139782 4036 139834
rect 4098 139782 4110 139834
rect 4172 139782 4174 139834
rect 4012 139780 4036 139782
rect 4092 139780 4116 139782
rect 4172 139780 4196 139782
rect 3956 139760 4252 139780
rect 1956 139292 2252 139312
rect 2012 139290 2036 139292
rect 2092 139290 2116 139292
rect 2172 139290 2196 139292
rect 2034 139238 2036 139290
rect 2098 139238 2110 139290
rect 2172 139238 2174 139290
rect 2012 139236 2036 139238
rect 2092 139236 2116 139238
rect 2172 139236 2196 139238
rect 1956 139216 2252 139236
rect 3956 138748 4252 138768
rect 4012 138746 4036 138748
rect 4092 138746 4116 138748
rect 4172 138746 4196 138748
rect 4034 138694 4036 138746
rect 4098 138694 4110 138746
rect 4172 138694 4174 138746
rect 4012 138692 4036 138694
rect 4092 138692 4116 138694
rect 4172 138692 4196 138694
rect 3956 138672 4252 138692
rect 1956 138204 2252 138224
rect 2012 138202 2036 138204
rect 2092 138202 2116 138204
rect 2172 138202 2196 138204
rect 2034 138150 2036 138202
rect 2098 138150 2110 138202
rect 2172 138150 2174 138202
rect 2012 138148 2036 138150
rect 2092 138148 2116 138150
rect 2172 138148 2196 138150
rect 1956 138128 2252 138148
rect 3956 137660 4252 137680
rect 4012 137658 4036 137660
rect 4092 137658 4116 137660
rect 4172 137658 4196 137660
rect 4034 137606 4036 137658
rect 4098 137606 4110 137658
rect 4172 137606 4174 137658
rect 4012 137604 4036 137606
rect 4092 137604 4116 137606
rect 4172 137604 4196 137606
rect 3956 137584 4252 137604
rect 1956 137116 2252 137136
rect 2012 137114 2036 137116
rect 2092 137114 2116 137116
rect 2172 137114 2196 137116
rect 2034 137062 2036 137114
rect 2098 137062 2110 137114
rect 2172 137062 2174 137114
rect 2012 137060 2036 137062
rect 2092 137060 2116 137062
rect 2172 137060 2196 137062
rect 1956 137040 2252 137060
rect 3956 136572 4252 136592
rect 4012 136570 4036 136572
rect 4092 136570 4116 136572
rect 4172 136570 4196 136572
rect 4034 136518 4036 136570
rect 4098 136518 4110 136570
rect 4172 136518 4174 136570
rect 4012 136516 4036 136518
rect 4092 136516 4116 136518
rect 4172 136516 4196 136518
rect 3956 136496 4252 136516
rect 1956 136028 2252 136048
rect 2012 136026 2036 136028
rect 2092 136026 2116 136028
rect 2172 136026 2196 136028
rect 2034 135974 2036 136026
rect 2098 135974 2110 136026
rect 2172 135974 2174 136026
rect 2012 135972 2036 135974
rect 2092 135972 2116 135974
rect 2172 135972 2196 135974
rect 1956 135952 2252 135972
rect 3956 135484 4252 135504
rect 4012 135482 4036 135484
rect 4092 135482 4116 135484
rect 4172 135482 4196 135484
rect 4034 135430 4036 135482
rect 4098 135430 4110 135482
rect 4172 135430 4174 135482
rect 4012 135428 4036 135430
rect 4092 135428 4116 135430
rect 4172 135428 4196 135430
rect 3956 135408 4252 135428
rect 1956 134940 2252 134960
rect 2012 134938 2036 134940
rect 2092 134938 2116 134940
rect 2172 134938 2196 134940
rect 2034 134886 2036 134938
rect 2098 134886 2110 134938
rect 2172 134886 2174 134938
rect 2012 134884 2036 134886
rect 2092 134884 2116 134886
rect 2172 134884 2196 134886
rect 1956 134864 2252 134884
rect 3956 134396 4252 134416
rect 4012 134394 4036 134396
rect 4092 134394 4116 134396
rect 4172 134394 4196 134396
rect 4034 134342 4036 134394
rect 4098 134342 4110 134394
rect 4172 134342 4174 134394
rect 4012 134340 4036 134342
rect 4092 134340 4116 134342
rect 4172 134340 4196 134342
rect 3956 134320 4252 134340
rect 1956 133852 2252 133872
rect 2012 133850 2036 133852
rect 2092 133850 2116 133852
rect 2172 133850 2196 133852
rect 2034 133798 2036 133850
rect 2098 133798 2110 133850
rect 2172 133798 2174 133850
rect 2012 133796 2036 133798
rect 2092 133796 2116 133798
rect 2172 133796 2196 133798
rect 1956 133776 2252 133796
rect 3956 133308 4252 133328
rect 4012 133306 4036 133308
rect 4092 133306 4116 133308
rect 4172 133306 4196 133308
rect 4034 133254 4036 133306
rect 4098 133254 4110 133306
rect 4172 133254 4174 133306
rect 4012 133252 4036 133254
rect 4092 133252 4116 133254
rect 4172 133252 4196 133254
rect 3956 133232 4252 133252
rect 1956 132764 2252 132784
rect 2012 132762 2036 132764
rect 2092 132762 2116 132764
rect 2172 132762 2196 132764
rect 2034 132710 2036 132762
rect 2098 132710 2110 132762
rect 2172 132710 2174 132762
rect 2012 132708 2036 132710
rect 2092 132708 2116 132710
rect 2172 132708 2196 132710
rect 1956 132688 2252 132708
rect 3956 132220 4252 132240
rect 4012 132218 4036 132220
rect 4092 132218 4116 132220
rect 4172 132218 4196 132220
rect 4034 132166 4036 132218
rect 4098 132166 4110 132218
rect 4172 132166 4174 132218
rect 4012 132164 4036 132166
rect 4092 132164 4116 132166
rect 4172 132164 4196 132166
rect 3956 132144 4252 132164
rect 1956 131676 2252 131696
rect 2012 131674 2036 131676
rect 2092 131674 2116 131676
rect 2172 131674 2196 131676
rect 2034 131622 2036 131674
rect 2098 131622 2110 131674
rect 2172 131622 2174 131674
rect 2012 131620 2036 131622
rect 2092 131620 2116 131622
rect 2172 131620 2196 131622
rect 1956 131600 2252 131620
rect 3956 131132 4252 131152
rect 4012 131130 4036 131132
rect 4092 131130 4116 131132
rect 4172 131130 4196 131132
rect 4034 131078 4036 131130
rect 4098 131078 4110 131130
rect 4172 131078 4174 131130
rect 4012 131076 4036 131078
rect 4092 131076 4116 131078
rect 4172 131076 4196 131078
rect 3956 131056 4252 131076
rect 1956 130588 2252 130608
rect 2012 130586 2036 130588
rect 2092 130586 2116 130588
rect 2172 130586 2196 130588
rect 2034 130534 2036 130586
rect 2098 130534 2110 130586
rect 2172 130534 2174 130586
rect 2012 130532 2036 130534
rect 2092 130532 2116 130534
rect 2172 130532 2196 130534
rect 1956 130512 2252 130532
rect 3956 130044 4252 130064
rect 4012 130042 4036 130044
rect 4092 130042 4116 130044
rect 4172 130042 4196 130044
rect 4034 129990 4036 130042
rect 4098 129990 4110 130042
rect 4172 129990 4174 130042
rect 4012 129988 4036 129990
rect 4092 129988 4116 129990
rect 4172 129988 4196 129990
rect 3956 129968 4252 129988
rect 1956 129500 2252 129520
rect 2012 129498 2036 129500
rect 2092 129498 2116 129500
rect 2172 129498 2196 129500
rect 2034 129446 2036 129498
rect 2098 129446 2110 129498
rect 2172 129446 2174 129498
rect 2012 129444 2036 129446
rect 2092 129444 2116 129446
rect 2172 129444 2196 129446
rect 1956 129424 2252 129444
rect 3956 128956 4252 128976
rect 4012 128954 4036 128956
rect 4092 128954 4116 128956
rect 4172 128954 4196 128956
rect 4034 128902 4036 128954
rect 4098 128902 4110 128954
rect 4172 128902 4174 128954
rect 4012 128900 4036 128902
rect 4092 128900 4116 128902
rect 4172 128900 4196 128902
rect 3956 128880 4252 128900
rect 1956 128412 2252 128432
rect 2012 128410 2036 128412
rect 2092 128410 2116 128412
rect 2172 128410 2196 128412
rect 2034 128358 2036 128410
rect 2098 128358 2110 128410
rect 2172 128358 2174 128410
rect 2012 128356 2036 128358
rect 2092 128356 2116 128358
rect 2172 128356 2196 128358
rect 1956 128336 2252 128356
rect 3956 127868 4252 127888
rect 4012 127866 4036 127868
rect 4092 127866 4116 127868
rect 4172 127866 4196 127868
rect 4034 127814 4036 127866
rect 4098 127814 4110 127866
rect 4172 127814 4174 127866
rect 4012 127812 4036 127814
rect 4092 127812 4116 127814
rect 4172 127812 4196 127814
rect 3956 127792 4252 127812
rect 1956 127324 2252 127344
rect 2012 127322 2036 127324
rect 2092 127322 2116 127324
rect 2172 127322 2196 127324
rect 2034 127270 2036 127322
rect 2098 127270 2110 127322
rect 2172 127270 2174 127322
rect 2012 127268 2036 127270
rect 2092 127268 2116 127270
rect 2172 127268 2196 127270
rect 1956 127248 2252 127268
rect 3956 126780 4252 126800
rect 4012 126778 4036 126780
rect 4092 126778 4116 126780
rect 4172 126778 4196 126780
rect 4034 126726 4036 126778
rect 4098 126726 4110 126778
rect 4172 126726 4174 126778
rect 4012 126724 4036 126726
rect 4092 126724 4116 126726
rect 4172 126724 4196 126726
rect 3956 126704 4252 126724
rect 1956 126236 2252 126256
rect 2012 126234 2036 126236
rect 2092 126234 2116 126236
rect 2172 126234 2196 126236
rect 2034 126182 2036 126234
rect 2098 126182 2110 126234
rect 2172 126182 2174 126234
rect 2012 126180 2036 126182
rect 2092 126180 2116 126182
rect 2172 126180 2196 126182
rect 1956 126160 2252 126180
rect 3956 125692 4252 125712
rect 4012 125690 4036 125692
rect 4092 125690 4116 125692
rect 4172 125690 4196 125692
rect 4034 125638 4036 125690
rect 4098 125638 4110 125690
rect 4172 125638 4174 125690
rect 4012 125636 4036 125638
rect 4092 125636 4116 125638
rect 4172 125636 4196 125638
rect 3956 125616 4252 125636
rect 1956 125148 2252 125168
rect 2012 125146 2036 125148
rect 2092 125146 2116 125148
rect 2172 125146 2196 125148
rect 2034 125094 2036 125146
rect 2098 125094 2110 125146
rect 2172 125094 2174 125146
rect 2012 125092 2036 125094
rect 2092 125092 2116 125094
rect 2172 125092 2196 125094
rect 1956 125072 2252 125092
rect 3956 124604 4252 124624
rect 4012 124602 4036 124604
rect 4092 124602 4116 124604
rect 4172 124602 4196 124604
rect 4034 124550 4036 124602
rect 4098 124550 4110 124602
rect 4172 124550 4174 124602
rect 4012 124548 4036 124550
rect 4092 124548 4116 124550
rect 4172 124548 4196 124550
rect 3956 124528 4252 124548
rect 1956 124060 2252 124080
rect 2012 124058 2036 124060
rect 2092 124058 2116 124060
rect 2172 124058 2196 124060
rect 2034 124006 2036 124058
rect 2098 124006 2110 124058
rect 2172 124006 2174 124058
rect 2012 124004 2036 124006
rect 2092 124004 2116 124006
rect 2172 124004 2196 124006
rect 1956 123984 2252 124004
rect 3956 123516 4252 123536
rect 4012 123514 4036 123516
rect 4092 123514 4116 123516
rect 4172 123514 4196 123516
rect 4034 123462 4036 123514
rect 4098 123462 4110 123514
rect 4172 123462 4174 123514
rect 4012 123460 4036 123462
rect 4092 123460 4116 123462
rect 4172 123460 4196 123462
rect 3956 123440 4252 123460
rect 1956 122972 2252 122992
rect 2012 122970 2036 122972
rect 2092 122970 2116 122972
rect 2172 122970 2196 122972
rect 2034 122918 2036 122970
rect 2098 122918 2110 122970
rect 2172 122918 2174 122970
rect 2012 122916 2036 122918
rect 2092 122916 2116 122918
rect 2172 122916 2196 122918
rect 1956 122896 2252 122916
rect 3956 122428 4252 122448
rect 4012 122426 4036 122428
rect 4092 122426 4116 122428
rect 4172 122426 4196 122428
rect 4034 122374 4036 122426
rect 4098 122374 4110 122426
rect 4172 122374 4174 122426
rect 4012 122372 4036 122374
rect 4092 122372 4116 122374
rect 4172 122372 4196 122374
rect 3956 122352 4252 122372
rect 1956 121884 2252 121904
rect 2012 121882 2036 121884
rect 2092 121882 2116 121884
rect 2172 121882 2196 121884
rect 2034 121830 2036 121882
rect 2098 121830 2110 121882
rect 2172 121830 2174 121882
rect 2012 121828 2036 121830
rect 2092 121828 2116 121830
rect 2172 121828 2196 121830
rect 1956 121808 2252 121828
rect 3956 121340 4252 121360
rect 4012 121338 4036 121340
rect 4092 121338 4116 121340
rect 4172 121338 4196 121340
rect 4034 121286 4036 121338
rect 4098 121286 4110 121338
rect 4172 121286 4174 121338
rect 4012 121284 4036 121286
rect 4092 121284 4116 121286
rect 4172 121284 4196 121286
rect 3956 121264 4252 121284
rect 1956 120796 2252 120816
rect 2012 120794 2036 120796
rect 2092 120794 2116 120796
rect 2172 120794 2196 120796
rect 2034 120742 2036 120794
rect 2098 120742 2110 120794
rect 2172 120742 2174 120794
rect 2012 120740 2036 120742
rect 2092 120740 2116 120742
rect 2172 120740 2196 120742
rect 1956 120720 2252 120740
rect 3956 120252 4252 120272
rect 4012 120250 4036 120252
rect 4092 120250 4116 120252
rect 4172 120250 4196 120252
rect 4034 120198 4036 120250
rect 4098 120198 4110 120250
rect 4172 120198 4174 120250
rect 4012 120196 4036 120198
rect 4092 120196 4116 120198
rect 4172 120196 4196 120198
rect 3956 120176 4252 120196
rect 1956 119708 2252 119728
rect 2012 119706 2036 119708
rect 2092 119706 2116 119708
rect 2172 119706 2196 119708
rect 2034 119654 2036 119706
rect 2098 119654 2110 119706
rect 2172 119654 2174 119706
rect 2012 119652 2036 119654
rect 2092 119652 2116 119654
rect 2172 119652 2196 119654
rect 1956 119632 2252 119652
rect 3956 119164 4252 119184
rect 4012 119162 4036 119164
rect 4092 119162 4116 119164
rect 4172 119162 4196 119164
rect 4034 119110 4036 119162
rect 4098 119110 4110 119162
rect 4172 119110 4174 119162
rect 4012 119108 4036 119110
rect 4092 119108 4116 119110
rect 4172 119108 4196 119110
rect 3956 119088 4252 119108
rect 1956 118620 2252 118640
rect 2012 118618 2036 118620
rect 2092 118618 2116 118620
rect 2172 118618 2196 118620
rect 2034 118566 2036 118618
rect 2098 118566 2110 118618
rect 2172 118566 2174 118618
rect 2012 118564 2036 118566
rect 2092 118564 2116 118566
rect 2172 118564 2196 118566
rect 1956 118544 2252 118564
rect 3956 118076 4252 118096
rect 4012 118074 4036 118076
rect 4092 118074 4116 118076
rect 4172 118074 4196 118076
rect 4034 118022 4036 118074
rect 4098 118022 4110 118074
rect 4172 118022 4174 118074
rect 4012 118020 4036 118022
rect 4092 118020 4116 118022
rect 4172 118020 4196 118022
rect 3956 118000 4252 118020
rect 1956 117532 2252 117552
rect 2012 117530 2036 117532
rect 2092 117530 2116 117532
rect 2172 117530 2196 117532
rect 2034 117478 2036 117530
rect 2098 117478 2110 117530
rect 2172 117478 2174 117530
rect 2012 117476 2036 117478
rect 2092 117476 2116 117478
rect 2172 117476 2196 117478
rect 1956 117456 2252 117476
rect 3956 116988 4252 117008
rect 4012 116986 4036 116988
rect 4092 116986 4116 116988
rect 4172 116986 4196 116988
rect 4034 116934 4036 116986
rect 4098 116934 4110 116986
rect 4172 116934 4174 116986
rect 4012 116932 4036 116934
rect 4092 116932 4116 116934
rect 4172 116932 4196 116934
rect 3956 116912 4252 116932
rect 1956 116444 2252 116464
rect 2012 116442 2036 116444
rect 2092 116442 2116 116444
rect 2172 116442 2196 116444
rect 2034 116390 2036 116442
rect 2098 116390 2110 116442
rect 2172 116390 2174 116442
rect 2012 116388 2036 116390
rect 2092 116388 2116 116390
rect 2172 116388 2196 116390
rect 1956 116368 2252 116388
rect 3956 115900 4252 115920
rect 4012 115898 4036 115900
rect 4092 115898 4116 115900
rect 4172 115898 4196 115900
rect 4034 115846 4036 115898
rect 4098 115846 4110 115898
rect 4172 115846 4174 115898
rect 4012 115844 4036 115846
rect 4092 115844 4116 115846
rect 4172 115844 4196 115846
rect 3956 115824 4252 115844
rect 1956 115356 2252 115376
rect 2012 115354 2036 115356
rect 2092 115354 2116 115356
rect 2172 115354 2196 115356
rect 2034 115302 2036 115354
rect 2098 115302 2110 115354
rect 2172 115302 2174 115354
rect 2012 115300 2036 115302
rect 2092 115300 2116 115302
rect 2172 115300 2196 115302
rect 1956 115280 2252 115300
rect 3956 114812 4252 114832
rect 4012 114810 4036 114812
rect 4092 114810 4116 114812
rect 4172 114810 4196 114812
rect 4034 114758 4036 114810
rect 4098 114758 4110 114810
rect 4172 114758 4174 114810
rect 4012 114756 4036 114758
rect 4092 114756 4116 114758
rect 4172 114756 4196 114758
rect 3956 114736 4252 114756
rect 1956 114268 2252 114288
rect 2012 114266 2036 114268
rect 2092 114266 2116 114268
rect 2172 114266 2196 114268
rect 2034 114214 2036 114266
rect 2098 114214 2110 114266
rect 2172 114214 2174 114266
rect 2012 114212 2036 114214
rect 2092 114212 2116 114214
rect 2172 114212 2196 114214
rect 1956 114192 2252 114212
rect 3956 113724 4252 113744
rect 4012 113722 4036 113724
rect 4092 113722 4116 113724
rect 4172 113722 4196 113724
rect 4034 113670 4036 113722
rect 4098 113670 4110 113722
rect 4172 113670 4174 113722
rect 4012 113668 4036 113670
rect 4092 113668 4116 113670
rect 4172 113668 4196 113670
rect 3956 113648 4252 113668
rect 1956 113180 2252 113200
rect 2012 113178 2036 113180
rect 2092 113178 2116 113180
rect 2172 113178 2196 113180
rect 2034 113126 2036 113178
rect 2098 113126 2110 113178
rect 2172 113126 2174 113178
rect 2012 113124 2036 113126
rect 2092 113124 2116 113126
rect 2172 113124 2196 113126
rect 1956 113104 2252 113124
rect 3956 112636 4252 112656
rect 4012 112634 4036 112636
rect 4092 112634 4116 112636
rect 4172 112634 4196 112636
rect 4034 112582 4036 112634
rect 4098 112582 4110 112634
rect 4172 112582 4174 112634
rect 4012 112580 4036 112582
rect 4092 112580 4116 112582
rect 4172 112580 4196 112582
rect 3956 112560 4252 112580
rect 1956 112092 2252 112112
rect 2012 112090 2036 112092
rect 2092 112090 2116 112092
rect 2172 112090 2196 112092
rect 2034 112038 2036 112090
rect 2098 112038 2110 112090
rect 2172 112038 2174 112090
rect 2012 112036 2036 112038
rect 2092 112036 2116 112038
rect 2172 112036 2196 112038
rect 1956 112016 2252 112036
rect 3956 111548 4252 111568
rect 4012 111546 4036 111548
rect 4092 111546 4116 111548
rect 4172 111546 4196 111548
rect 4034 111494 4036 111546
rect 4098 111494 4110 111546
rect 4172 111494 4174 111546
rect 4012 111492 4036 111494
rect 4092 111492 4116 111494
rect 4172 111492 4196 111494
rect 3956 111472 4252 111492
rect 1956 111004 2252 111024
rect 2012 111002 2036 111004
rect 2092 111002 2116 111004
rect 2172 111002 2196 111004
rect 2034 110950 2036 111002
rect 2098 110950 2110 111002
rect 2172 110950 2174 111002
rect 2012 110948 2036 110950
rect 2092 110948 2116 110950
rect 2172 110948 2196 110950
rect 1956 110928 2252 110948
rect 3956 110460 4252 110480
rect 4012 110458 4036 110460
rect 4092 110458 4116 110460
rect 4172 110458 4196 110460
rect 4034 110406 4036 110458
rect 4098 110406 4110 110458
rect 4172 110406 4174 110458
rect 4012 110404 4036 110406
rect 4092 110404 4116 110406
rect 4172 110404 4196 110406
rect 3956 110384 4252 110404
rect 1956 109916 2252 109936
rect 2012 109914 2036 109916
rect 2092 109914 2116 109916
rect 2172 109914 2196 109916
rect 2034 109862 2036 109914
rect 2098 109862 2110 109914
rect 2172 109862 2174 109914
rect 2012 109860 2036 109862
rect 2092 109860 2116 109862
rect 2172 109860 2196 109862
rect 1956 109840 2252 109860
rect 3956 109372 4252 109392
rect 4012 109370 4036 109372
rect 4092 109370 4116 109372
rect 4172 109370 4196 109372
rect 4034 109318 4036 109370
rect 4098 109318 4110 109370
rect 4172 109318 4174 109370
rect 4012 109316 4036 109318
rect 4092 109316 4116 109318
rect 4172 109316 4196 109318
rect 3956 109296 4252 109316
rect 1956 108828 2252 108848
rect 2012 108826 2036 108828
rect 2092 108826 2116 108828
rect 2172 108826 2196 108828
rect 2034 108774 2036 108826
rect 2098 108774 2110 108826
rect 2172 108774 2174 108826
rect 2012 108772 2036 108774
rect 2092 108772 2116 108774
rect 2172 108772 2196 108774
rect 1956 108752 2252 108772
rect 3956 108284 4252 108304
rect 4012 108282 4036 108284
rect 4092 108282 4116 108284
rect 4172 108282 4196 108284
rect 4034 108230 4036 108282
rect 4098 108230 4110 108282
rect 4172 108230 4174 108282
rect 4012 108228 4036 108230
rect 4092 108228 4116 108230
rect 4172 108228 4196 108230
rect 3956 108208 4252 108228
rect 1956 107740 2252 107760
rect 2012 107738 2036 107740
rect 2092 107738 2116 107740
rect 2172 107738 2196 107740
rect 2034 107686 2036 107738
rect 2098 107686 2110 107738
rect 2172 107686 2174 107738
rect 2012 107684 2036 107686
rect 2092 107684 2116 107686
rect 2172 107684 2196 107686
rect 1956 107664 2252 107684
rect 3956 107196 4252 107216
rect 4012 107194 4036 107196
rect 4092 107194 4116 107196
rect 4172 107194 4196 107196
rect 4034 107142 4036 107194
rect 4098 107142 4110 107194
rect 4172 107142 4174 107194
rect 4012 107140 4036 107142
rect 4092 107140 4116 107142
rect 4172 107140 4196 107142
rect 3956 107120 4252 107140
rect 1956 106652 2252 106672
rect 2012 106650 2036 106652
rect 2092 106650 2116 106652
rect 2172 106650 2196 106652
rect 2034 106598 2036 106650
rect 2098 106598 2110 106650
rect 2172 106598 2174 106650
rect 2012 106596 2036 106598
rect 2092 106596 2116 106598
rect 2172 106596 2196 106598
rect 1956 106576 2252 106596
rect 3956 106108 4252 106128
rect 4012 106106 4036 106108
rect 4092 106106 4116 106108
rect 4172 106106 4196 106108
rect 4034 106054 4036 106106
rect 4098 106054 4110 106106
rect 4172 106054 4174 106106
rect 4012 106052 4036 106054
rect 4092 106052 4116 106054
rect 4172 106052 4196 106054
rect 3956 106032 4252 106052
rect 4448 105874 4476 186730
rect 84384 186380 84436 186386
rect 84384 186322 84436 186328
rect 84396 186289 84424 186322
rect 84382 186280 84438 186289
rect 84382 186215 84438 186224
rect 4802 183016 4858 183025
rect 4802 182951 4804 182960
rect 4856 182951 4858 182960
rect 5170 183016 5226 183025
rect 5170 182951 5226 182960
rect 4804 182922 4856 182928
rect 4802 181928 4858 181937
rect 4802 181863 4804 181872
rect 4856 181863 4858 181872
rect 4804 181834 4856 181840
rect 4816 180794 4844 181834
rect 4816 180766 4936 180794
rect 4620 180192 4672 180198
rect 4618 180160 4620 180169
rect 4672 180160 4674 180169
rect 4618 180095 4674 180104
rect 4528 179104 4580 179110
rect 4526 179072 4528 179081
rect 4580 179072 4582 179081
rect 4526 179007 4582 179016
rect 4540 174418 4568 179007
rect 4528 174412 4580 174418
rect 4528 174354 4580 174360
rect 4632 174350 4660 180095
rect 4710 177032 4766 177041
rect 4710 176967 4766 176976
rect 4724 176934 4752 176967
rect 4712 176928 4764 176934
rect 4712 176870 4764 176876
rect 4620 174344 4672 174350
rect 4620 174286 4672 174292
rect 4436 105868 4488 105874
rect 4436 105810 4488 105816
rect 1956 105564 2252 105584
rect 2012 105562 2036 105564
rect 2092 105562 2116 105564
rect 2172 105562 2196 105564
rect 2034 105510 2036 105562
rect 2098 105510 2110 105562
rect 2172 105510 2174 105562
rect 2012 105508 2036 105510
rect 2092 105508 2116 105510
rect 2172 105508 2196 105510
rect 1956 105488 2252 105508
rect 3956 105020 4252 105040
rect 4012 105018 4036 105020
rect 4092 105018 4116 105020
rect 4172 105018 4196 105020
rect 4034 104966 4036 105018
rect 4098 104966 4110 105018
rect 4172 104966 4174 105018
rect 4012 104964 4036 104966
rect 4092 104964 4116 104966
rect 4172 104964 4196 104966
rect 3956 104944 4252 104964
rect 1956 104476 2252 104496
rect 2012 104474 2036 104476
rect 2092 104474 2116 104476
rect 2172 104474 2196 104476
rect 2034 104422 2036 104474
rect 2098 104422 2110 104474
rect 2172 104422 2174 104474
rect 2012 104420 2036 104422
rect 2092 104420 2116 104422
rect 2172 104420 2196 104422
rect 1956 104400 2252 104420
rect 3956 103932 4252 103952
rect 4012 103930 4036 103932
rect 4092 103930 4116 103932
rect 4172 103930 4196 103932
rect 4034 103878 4036 103930
rect 4098 103878 4110 103930
rect 4172 103878 4174 103930
rect 4012 103876 4036 103878
rect 4092 103876 4116 103878
rect 4172 103876 4196 103878
rect 3956 103856 4252 103876
rect 1956 103388 2252 103408
rect 2012 103386 2036 103388
rect 2092 103386 2116 103388
rect 2172 103386 2196 103388
rect 2034 103334 2036 103386
rect 2098 103334 2110 103386
rect 2172 103334 2174 103386
rect 2012 103332 2036 103334
rect 2092 103332 2116 103334
rect 2172 103332 2196 103334
rect 1956 103312 2252 103332
rect 3956 102844 4252 102864
rect 4012 102842 4036 102844
rect 4092 102842 4116 102844
rect 4172 102842 4196 102844
rect 4034 102790 4036 102842
rect 4098 102790 4110 102842
rect 4172 102790 4174 102842
rect 4012 102788 4036 102790
rect 4092 102788 4116 102790
rect 4172 102788 4196 102790
rect 3956 102768 4252 102788
rect 1956 102300 2252 102320
rect 2012 102298 2036 102300
rect 2092 102298 2116 102300
rect 2172 102298 2196 102300
rect 2034 102246 2036 102298
rect 2098 102246 2110 102298
rect 2172 102246 2174 102298
rect 2012 102244 2036 102246
rect 2092 102244 2116 102246
rect 2172 102244 2196 102246
rect 1956 102224 2252 102244
rect 3956 101756 4252 101776
rect 4012 101754 4036 101756
rect 4092 101754 4116 101756
rect 4172 101754 4196 101756
rect 4034 101702 4036 101754
rect 4098 101702 4110 101754
rect 4172 101702 4174 101754
rect 4012 101700 4036 101702
rect 4092 101700 4116 101702
rect 4172 101700 4196 101702
rect 3956 101680 4252 101700
rect 1956 101212 2252 101232
rect 2012 101210 2036 101212
rect 2092 101210 2116 101212
rect 2172 101210 2196 101212
rect 2034 101158 2036 101210
rect 2098 101158 2110 101210
rect 2172 101158 2174 101210
rect 2012 101156 2036 101158
rect 2092 101156 2116 101158
rect 2172 101156 2196 101158
rect 1956 101136 2252 101156
rect 3956 100668 4252 100688
rect 4012 100666 4036 100668
rect 4092 100666 4116 100668
rect 4172 100666 4196 100668
rect 4034 100614 4036 100666
rect 4098 100614 4110 100666
rect 4172 100614 4174 100666
rect 4012 100612 4036 100614
rect 4092 100612 4116 100614
rect 4172 100612 4196 100614
rect 3956 100592 4252 100612
rect 1956 100124 2252 100144
rect 2012 100122 2036 100124
rect 2092 100122 2116 100124
rect 2172 100122 2196 100124
rect 2034 100070 2036 100122
rect 2098 100070 2110 100122
rect 2172 100070 2174 100122
rect 2012 100068 2036 100070
rect 2092 100068 2116 100070
rect 2172 100068 2196 100070
rect 1956 100048 2252 100068
rect 3956 99580 4252 99600
rect 4012 99578 4036 99580
rect 4092 99578 4116 99580
rect 4172 99578 4196 99580
rect 4034 99526 4036 99578
rect 4098 99526 4110 99578
rect 4172 99526 4174 99578
rect 4012 99524 4036 99526
rect 4092 99524 4116 99526
rect 4172 99524 4196 99526
rect 3956 99504 4252 99524
rect 1956 99036 2252 99056
rect 2012 99034 2036 99036
rect 2092 99034 2116 99036
rect 2172 99034 2196 99036
rect 2034 98982 2036 99034
rect 2098 98982 2110 99034
rect 2172 98982 2174 99034
rect 2012 98980 2036 98982
rect 2092 98980 2116 98982
rect 2172 98980 2196 98982
rect 1956 98960 2252 98980
rect 4344 98592 4396 98598
rect 4344 98534 4396 98540
rect 3956 98492 4252 98512
rect 4012 98490 4036 98492
rect 4092 98490 4116 98492
rect 4172 98490 4196 98492
rect 4034 98438 4036 98490
rect 4098 98438 4110 98490
rect 4172 98438 4174 98490
rect 4012 98436 4036 98438
rect 4092 98436 4116 98438
rect 4172 98436 4196 98438
rect 3956 98416 4252 98436
rect 1956 97948 2252 97968
rect 2012 97946 2036 97948
rect 2092 97946 2116 97948
rect 2172 97946 2196 97948
rect 2034 97894 2036 97946
rect 2098 97894 2110 97946
rect 2172 97894 2174 97946
rect 2012 97892 2036 97894
rect 2092 97892 2116 97894
rect 2172 97892 2196 97894
rect 1956 97872 2252 97892
rect 2596 97844 2648 97850
rect 2596 97786 2648 97792
rect 2608 97306 2636 97786
rect 3332 97504 3384 97510
rect 3332 97446 3384 97452
rect 2596 97300 2648 97306
rect 2596 97242 2648 97248
rect 1956 96860 2252 96880
rect 2012 96858 2036 96860
rect 2092 96858 2116 96860
rect 2172 96858 2196 96860
rect 2034 96806 2036 96858
rect 2098 96806 2110 96858
rect 2172 96806 2174 96858
rect 2012 96804 2036 96806
rect 2092 96804 2116 96806
rect 2172 96804 2196 96806
rect 1956 96784 2252 96804
rect 1956 95772 2252 95792
rect 2012 95770 2036 95772
rect 2092 95770 2116 95772
rect 2172 95770 2196 95772
rect 2034 95718 2036 95770
rect 2098 95718 2110 95770
rect 2172 95718 2174 95770
rect 2012 95716 2036 95718
rect 2092 95716 2116 95718
rect 2172 95716 2196 95718
rect 1956 95696 2252 95716
rect 1956 94684 2252 94704
rect 2012 94682 2036 94684
rect 2092 94682 2116 94684
rect 2172 94682 2196 94684
rect 2034 94630 2036 94682
rect 2098 94630 2110 94682
rect 2172 94630 2174 94682
rect 2012 94628 2036 94630
rect 2092 94628 2116 94630
rect 2172 94628 2196 94630
rect 1956 94608 2252 94628
rect 1956 93596 2252 93616
rect 2012 93594 2036 93596
rect 2092 93594 2116 93596
rect 2172 93594 2196 93596
rect 2034 93542 2036 93594
rect 2098 93542 2110 93594
rect 2172 93542 2174 93594
rect 2012 93540 2036 93542
rect 2092 93540 2116 93542
rect 2172 93540 2196 93542
rect 1956 93520 2252 93540
rect 1956 92508 2252 92528
rect 2012 92506 2036 92508
rect 2092 92506 2116 92508
rect 2172 92506 2196 92508
rect 2034 92454 2036 92506
rect 2098 92454 2110 92506
rect 2172 92454 2174 92506
rect 2012 92452 2036 92454
rect 2092 92452 2116 92454
rect 2172 92452 2196 92454
rect 1956 92432 2252 92452
rect 1956 91420 2252 91440
rect 2012 91418 2036 91420
rect 2092 91418 2116 91420
rect 2172 91418 2196 91420
rect 2034 91366 2036 91418
rect 2098 91366 2110 91418
rect 2172 91366 2174 91418
rect 2012 91364 2036 91366
rect 2092 91364 2116 91366
rect 2172 91364 2196 91366
rect 1956 91344 2252 91364
rect 1956 90332 2252 90352
rect 2012 90330 2036 90332
rect 2092 90330 2116 90332
rect 2172 90330 2196 90332
rect 2034 90278 2036 90330
rect 2098 90278 2110 90330
rect 2172 90278 2174 90330
rect 2012 90276 2036 90278
rect 2092 90276 2116 90278
rect 2172 90276 2196 90278
rect 1956 90256 2252 90276
rect 1956 89244 2252 89264
rect 2012 89242 2036 89244
rect 2092 89242 2116 89244
rect 2172 89242 2196 89244
rect 2034 89190 2036 89242
rect 2098 89190 2110 89242
rect 2172 89190 2174 89242
rect 2012 89188 2036 89190
rect 2092 89188 2116 89190
rect 2172 89188 2196 89190
rect 1956 89168 2252 89188
rect 1956 88156 2252 88176
rect 2012 88154 2036 88156
rect 2092 88154 2116 88156
rect 2172 88154 2196 88156
rect 2034 88102 2036 88154
rect 2098 88102 2110 88154
rect 2172 88102 2174 88154
rect 2012 88100 2036 88102
rect 2092 88100 2116 88102
rect 2172 88100 2196 88102
rect 1956 88080 2252 88100
rect 1956 87068 2252 87088
rect 2012 87066 2036 87068
rect 2092 87066 2116 87068
rect 2172 87066 2196 87068
rect 2034 87014 2036 87066
rect 2098 87014 2110 87066
rect 2172 87014 2174 87066
rect 2012 87012 2036 87014
rect 2092 87012 2116 87014
rect 2172 87012 2196 87014
rect 1956 86992 2252 87012
rect 1956 85980 2252 86000
rect 2012 85978 2036 85980
rect 2092 85978 2116 85980
rect 2172 85978 2196 85980
rect 2034 85926 2036 85978
rect 2098 85926 2110 85978
rect 2172 85926 2174 85978
rect 2012 85924 2036 85926
rect 2092 85924 2116 85926
rect 2172 85924 2196 85926
rect 1956 85904 2252 85924
rect 1956 84892 2252 84912
rect 2012 84890 2036 84892
rect 2092 84890 2116 84892
rect 2172 84890 2196 84892
rect 2034 84838 2036 84890
rect 2098 84838 2110 84890
rect 2172 84838 2174 84890
rect 2012 84836 2036 84838
rect 2092 84836 2116 84838
rect 2172 84836 2196 84838
rect 1956 84816 2252 84836
rect 2608 84194 2636 97242
rect 2964 96960 3016 96966
rect 2964 96902 3016 96908
rect 2976 96694 3004 96902
rect 3344 96762 3372 97446
rect 3956 97404 4252 97424
rect 4012 97402 4036 97404
rect 4092 97402 4116 97404
rect 4172 97402 4196 97404
rect 4034 97350 4036 97402
rect 4098 97350 4110 97402
rect 4172 97350 4174 97402
rect 4012 97348 4036 97350
rect 4092 97348 4116 97350
rect 4172 97348 4196 97350
rect 3956 97328 4252 97348
rect 3608 97232 3660 97238
rect 3608 97174 3660 97180
rect 3332 96756 3384 96762
rect 3332 96698 3384 96704
rect 2964 96688 3016 96694
rect 2964 96630 3016 96636
rect 3344 96506 3372 96698
rect 3424 96688 3476 96694
rect 3424 96630 3476 96636
rect 2516 84166 2636 84194
rect 3252 96478 3372 96506
rect 1956 83804 2252 83824
rect 2012 83802 2036 83804
rect 2092 83802 2116 83804
rect 2172 83802 2196 83804
rect 2034 83750 2036 83802
rect 2098 83750 2110 83802
rect 2172 83750 2174 83802
rect 2012 83748 2036 83750
rect 2092 83748 2116 83750
rect 2172 83748 2196 83750
rect 1956 83728 2252 83748
rect 1956 82716 2252 82736
rect 2012 82714 2036 82716
rect 2092 82714 2116 82716
rect 2172 82714 2196 82716
rect 2034 82662 2036 82714
rect 2098 82662 2110 82714
rect 2172 82662 2174 82714
rect 2012 82660 2036 82662
rect 2092 82660 2116 82662
rect 2172 82660 2196 82662
rect 1956 82640 2252 82660
rect 1956 81628 2252 81648
rect 2012 81626 2036 81628
rect 2092 81626 2116 81628
rect 2172 81626 2196 81628
rect 2034 81574 2036 81626
rect 2098 81574 2110 81626
rect 2172 81574 2174 81626
rect 2012 81572 2036 81574
rect 2092 81572 2116 81574
rect 2172 81572 2196 81574
rect 1956 81552 2252 81572
rect 1956 80540 2252 80560
rect 2012 80538 2036 80540
rect 2092 80538 2116 80540
rect 2172 80538 2196 80540
rect 2034 80486 2036 80538
rect 2098 80486 2110 80538
rect 2172 80486 2174 80538
rect 2012 80484 2036 80486
rect 2092 80484 2116 80486
rect 2172 80484 2196 80486
rect 1956 80464 2252 80484
rect 1956 79452 2252 79472
rect 2012 79450 2036 79452
rect 2092 79450 2116 79452
rect 2172 79450 2196 79452
rect 2034 79398 2036 79450
rect 2098 79398 2110 79450
rect 2172 79398 2174 79450
rect 2012 79396 2036 79398
rect 2092 79396 2116 79398
rect 2172 79396 2196 79398
rect 1956 79376 2252 79396
rect 1956 78364 2252 78384
rect 2012 78362 2036 78364
rect 2092 78362 2116 78364
rect 2172 78362 2196 78364
rect 2034 78310 2036 78362
rect 2098 78310 2110 78362
rect 2172 78310 2174 78362
rect 2012 78308 2036 78310
rect 2092 78308 2116 78310
rect 2172 78308 2196 78310
rect 1956 78288 2252 78308
rect 1956 77276 2252 77296
rect 2012 77274 2036 77276
rect 2092 77274 2116 77276
rect 2172 77274 2196 77276
rect 2034 77222 2036 77274
rect 2098 77222 2110 77274
rect 2172 77222 2174 77274
rect 2012 77220 2036 77222
rect 2092 77220 2116 77222
rect 2172 77220 2196 77222
rect 1956 77200 2252 77220
rect 1956 76188 2252 76208
rect 2012 76186 2036 76188
rect 2092 76186 2116 76188
rect 2172 76186 2196 76188
rect 2034 76134 2036 76186
rect 2098 76134 2110 76186
rect 2172 76134 2174 76186
rect 2012 76132 2036 76134
rect 2092 76132 2116 76134
rect 2172 76132 2196 76134
rect 1956 76112 2252 76132
rect 1956 75100 2252 75120
rect 2012 75098 2036 75100
rect 2092 75098 2116 75100
rect 2172 75098 2196 75100
rect 2034 75046 2036 75098
rect 2098 75046 2110 75098
rect 2172 75046 2174 75098
rect 2012 75044 2036 75046
rect 2092 75044 2116 75046
rect 2172 75044 2196 75046
rect 1956 75024 2252 75044
rect 1956 74012 2252 74032
rect 2012 74010 2036 74012
rect 2092 74010 2116 74012
rect 2172 74010 2196 74012
rect 2034 73958 2036 74010
rect 2098 73958 2110 74010
rect 2172 73958 2174 74010
rect 2012 73956 2036 73958
rect 2092 73956 2116 73958
rect 2172 73956 2196 73958
rect 1956 73936 2252 73956
rect 1956 72924 2252 72944
rect 2012 72922 2036 72924
rect 2092 72922 2116 72924
rect 2172 72922 2196 72924
rect 2034 72870 2036 72922
rect 2098 72870 2110 72922
rect 2172 72870 2174 72922
rect 2012 72868 2036 72870
rect 2092 72868 2116 72870
rect 2172 72868 2196 72870
rect 1956 72848 2252 72868
rect 1956 71836 2252 71856
rect 2012 71834 2036 71836
rect 2092 71834 2116 71836
rect 2172 71834 2196 71836
rect 2034 71782 2036 71834
rect 2098 71782 2110 71834
rect 2172 71782 2174 71834
rect 2012 71780 2036 71782
rect 2092 71780 2116 71782
rect 2172 71780 2196 71782
rect 1956 71760 2252 71780
rect 1956 70748 2252 70768
rect 2012 70746 2036 70748
rect 2092 70746 2116 70748
rect 2172 70746 2196 70748
rect 2034 70694 2036 70746
rect 2098 70694 2110 70746
rect 2172 70694 2174 70746
rect 2012 70692 2036 70694
rect 2092 70692 2116 70694
rect 2172 70692 2196 70694
rect 1956 70672 2252 70692
rect 1956 69660 2252 69680
rect 2012 69658 2036 69660
rect 2092 69658 2116 69660
rect 2172 69658 2196 69660
rect 2034 69606 2036 69658
rect 2098 69606 2110 69658
rect 2172 69606 2174 69658
rect 2012 69604 2036 69606
rect 2092 69604 2116 69606
rect 2172 69604 2196 69606
rect 1956 69584 2252 69604
rect 1956 68572 2252 68592
rect 2012 68570 2036 68572
rect 2092 68570 2116 68572
rect 2172 68570 2196 68572
rect 2034 68518 2036 68570
rect 2098 68518 2110 68570
rect 2172 68518 2174 68570
rect 2012 68516 2036 68518
rect 2092 68516 2116 68518
rect 2172 68516 2196 68518
rect 1956 68496 2252 68516
rect 1956 67484 2252 67504
rect 2012 67482 2036 67484
rect 2092 67482 2116 67484
rect 2172 67482 2196 67484
rect 2034 67430 2036 67482
rect 2098 67430 2110 67482
rect 2172 67430 2174 67482
rect 2012 67428 2036 67430
rect 2092 67428 2116 67430
rect 2172 67428 2196 67430
rect 1956 67408 2252 67428
rect 1956 66396 2252 66416
rect 2012 66394 2036 66396
rect 2092 66394 2116 66396
rect 2172 66394 2196 66396
rect 2034 66342 2036 66394
rect 2098 66342 2110 66394
rect 2172 66342 2174 66394
rect 2012 66340 2036 66342
rect 2092 66340 2116 66342
rect 2172 66340 2196 66342
rect 1956 66320 2252 66340
rect 1956 65308 2252 65328
rect 2012 65306 2036 65308
rect 2092 65306 2116 65308
rect 2172 65306 2196 65308
rect 2034 65254 2036 65306
rect 2098 65254 2110 65306
rect 2172 65254 2174 65306
rect 2012 65252 2036 65254
rect 2092 65252 2116 65254
rect 2172 65252 2196 65254
rect 1956 65232 2252 65252
rect 1956 64220 2252 64240
rect 2012 64218 2036 64220
rect 2092 64218 2116 64220
rect 2172 64218 2196 64220
rect 2034 64166 2036 64218
rect 2098 64166 2110 64218
rect 2172 64166 2174 64218
rect 2012 64164 2036 64166
rect 2092 64164 2116 64166
rect 2172 64164 2196 64166
rect 1956 64144 2252 64164
rect 1956 63132 2252 63152
rect 2012 63130 2036 63132
rect 2092 63130 2116 63132
rect 2172 63130 2196 63132
rect 2034 63078 2036 63130
rect 2098 63078 2110 63130
rect 2172 63078 2174 63130
rect 2012 63076 2036 63078
rect 2092 63076 2116 63078
rect 2172 63076 2196 63078
rect 1956 63056 2252 63076
rect 1956 62044 2252 62064
rect 2012 62042 2036 62044
rect 2092 62042 2116 62044
rect 2172 62042 2196 62044
rect 2034 61990 2036 62042
rect 2098 61990 2110 62042
rect 2172 61990 2174 62042
rect 2012 61988 2036 61990
rect 2092 61988 2116 61990
rect 2172 61988 2196 61990
rect 1956 61968 2252 61988
rect 1956 60956 2252 60976
rect 2012 60954 2036 60956
rect 2092 60954 2116 60956
rect 2172 60954 2196 60956
rect 2034 60902 2036 60954
rect 2098 60902 2110 60954
rect 2172 60902 2174 60954
rect 2012 60900 2036 60902
rect 2092 60900 2116 60902
rect 2172 60900 2196 60902
rect 1956 60880 2252 60900
rect 1956 59868 2252 59888
rect 2012 59866 2036 59868
rect 2092 59866 2116 59868
rect 2172 59866 2196 59868
rect 2034 59814 2036 59866
rect 2098 59814 2110 59866
rect 2172 59814 2174 59866
rect 2012 59812 2036 59814
rect 2092 59812 2116 59814
rect 2172 59812 2196 59814
rect 1956 59792 2252 59812
rect 1956 58780 2252 58800
rect 2012 58778 2036 58780
rect 2092 58778 2116 58780
rect 2172 58778 2196 58780
rect 2034 58726 2036 58778
rect 2098 58726 2110 58778
rect 2172 58726 2174 58778
rect 2012 58724 2036 58726
rect 2092 58724 2116 58726
rect 2172 58724 2196 58726
rect 1956 58704 2252 58724
rect 1956 57692 2252 57712
rect 2012 57690 2036 57692
rect 2092 57690 2116 57692
rect 2172 57690 2196 57692
rect 2034 57638 2036 57690
rect 2098 57638 2110 57690
rect 2172 57638 2174 57690
rect 2012 57636 2036 57638
rect 2092 57636 2116 57638
rect 2172 57636 2196 57638
rect 1956 57616 2252 57636
rect 1956 56604 2252 56624
rect 2012 56602 2036 56604
rect 2092 56602 2116 56604
rect 2172 56602 2196 56604
rect 2034 56550 2036 56602
rect 2098 56550 2110 56602
rect 2172 56550 2174 56602
rect 2012 56548 2036 56550
rect 2092 56548 2116 56550
rect 2172 56548 2196 56550
rect 1956 56528 2252 56548
rect 1956 55516 2252 55536
rect 2012 55514 2036 55516
rect 2092 55514 2116 55516
rect 2172 55514 2196 55516
rect 2034 55462 2036 55514
rect 2098 55462 2110 55514
rect 2172 55462 2174 55514
rect 2012 55460 2036 55462
rect 2092 55460 2116 55462
rect 2172 55460 2196 55462
rect 1956 55440 2252 55460
rect 1956 54428 2252 54448
rect 2012 54426 2036 54428
rect 2092 54426 2116 54428
rect 2172 54426 2196 54428
rect 2034 54374 2036 54426
rect 2098 54374 2110 54426
rect 2172 54374 2174 54426
rect 2012 54372 2036 54374
rect 2092 54372 2116 54374
rect 2172 54372 2196 54374
rect 1956 54352 2252 54372
rect 1956 53340 2252 53360
rect 2012 53338 2036 53340
rect 2092 53338 2116 53340
rect 2172 53338 2196 53340
rect 2034 53286 2036 53338
rect 2098 53286 2110 53338
rect 2172 53286 2174 53338
rect 2012 53284 2036 53286
rect 2092 53284 2116 53286
rect 2172 53284 2196 53286
rect 1956 53264 2252 53284
rect 1956 52252 2252 52272
rect 2012 52250 2036 52252
rect 2092 52250 2116 52252
rect 2172 52250 2196 52252
rect 2034 52198 2036 52250
rect 2098 52198 2110 52250
rect 2172 52198 2174 52250
rect 2012 52196 2036 52198
rect 2092 52196 2116 52198
rect 2172 52196 2196 52198
rect 1956 52176 2252 52196
rect 1956 51164 2252 51184
rect 2012 51162 2036 51164
rect 2092 51162 2116 51164
rect 2172 51162 2196 51164
rect 2034 51110 2036 51162
rect 2098 51110 2110 51162
rect 2172 51110 2174 51162
rect 2012 51108 2036 51110
rect 2092 51108 2116 51110
rect 2172 51108 2196 51110
rect 1956 51088 2252 51108
rect 1956 50076 2252 50096
rect 2012 50074 2036 50076
rect 2092 50074 2116 50076
rect 2172 50074 2196 50076
rect 2034 50022 2036 50074
rect 2098 50022 2110 50074
rect 2172 50022 2174 50074
rect 2012 50020 2036 50022
rect 2092 50020 2116 50022
rect 2172 50020 2196 50022
rect 1956 50000 2252 50020
rect 1956 48988 2252 49008
rect 2012 48986 2036 48988
rect 2092 48986 2116 48988
rect 2172 48986 2196 48988
rect 2034 48934 2036 48986
rect 2098 48934 2110 48986
rect 2172 48934 2174 48986
rect 2012 48932 2036 48934
rect 2092 48932 2116 48934
rect 2172 48932 2196 48934
rect 1956 48912 2252 48932
rect 1956 47900 2252 47920
rect 2012 47898 2036 47900
rect 2092 47898 2116 47900
rect 2172 47898 2196 47900
rect 2034 47846 2036 47898
rect 2098 47846 2110 47898
rect 2172 47846 2174 47898
rect 2012 47844 2036 47846
rect 2092 47844 2116 47846
rect 2172 47844 2196 47846
rect 1956 47824 2252 47844
rect 1956 46812 2252 46832
rect 2012 46810 2036 46812
rect 2092 46810 2116 46812
rect 2172 46810 2196 46812
rect 2034 46758 2036 46810
rect 2098 46758 2110 46810
rect 2172 46758 2174 46810
rect 2012 46756 2036 46758
rect 2092 46756 2116 46758
rect 2172 46756 2196 46758
rect 1956 46736 2252 46756
rect 1956 45724 2252 45744
rect 2012 45722 2036 45724
rect 2092 45722 2116 45724
rect 2172 45722 2196 45724
rect 2034 45670 2036 45722
rect 2098 45670 2110 45722
rect 2172 45670 2174 45722
rect 2012 45668 2036 45670
rect 2092 45668 2116 45670
rect 2172 45668 2196 45670
rect 1956 45648 2252 45668
rect 1956 44636 2252 44656
rect 2012 44634 2036 44636
rect 2092 44634 2116 44636
rect 2172 44634 2196 44636
rect 2034 44582 2036 44634
rect 2098 44582 2110 44634
rect 2172 44582 2174 44634
rect 2012 44580 2036 44582
rect 2092 44580 2116 44582
rect 2172 44580 2196 44582
rect 1956 44560 2252 44580
rect 1956 43548 2252 43568
rect 2012 43546 2036 43548
rect 2092 43546 2116 43548
rect 2172 43546 2196 43548
rect 2034 43494 2036 43546
rect 2098 43494 2110 43546
rect 2172 43494 2174 43546
rect 2012 43492 2036 43494
rect 2092 43492 2116 43494
rect 2172 43492 2196 43494
rect 1956 43472 2252 43492
rect 1956 42460 2252 42480
rect 2012 42458 2036 42460
rect 2092 42458 2116 42460
rect 2172 42458 2196 42460
rect 2034 42406 2036 42458
rect 2098 42406 2110 42458
rect 2172 42406 2174 42458
rect 2012 42404 2036 42406
rect 2092 42404 2116 42406
rect 2172 42404 2196 42406
rect 1956 42384 2252 42404
rect 1956 41372 2252 41392
rect 2012 41370 2036 41372
rect 2092 41370 2116 41372
rect 2172 41370 2196 41372
rect 2034 41318 2036 41370
rect 2098 41318 2110 41370
rect 2172 41318 2174 41370
rect 2012 41316 2036 41318
rect 2092 41316 2116 41318
rect 2172 41316 2196 41318
rect 1956 41296 2252 41316
rect 1956 40284 2252 40304
rect 2012 40282 2036 40284
rect 2092 40282 2116 40284
rect 2172 40282 2196 40284
rect 2034 40230 2036 40282
rect 2098 40230 2110 40282
rect 2172 40230 2174 40282
rect 2012 40228 2036 40230
rect 2092 40228 2116 40230
rect 2172 40228 2196 40230
rect 1956 40208 2252 40228
rect 1956 39196 2252 39216
rect 2012 39194 2036 39196
rect 2092 39194 2116 39196
rect 2172 39194 2196 39196
rect 2034 39142 2036 39194
rect 2098 39142 2110 39194
rect 2172 39142 2174 39194
rect 2012 39140 2036 39142
rect 2092 39140 2116 39142
rect 2172 39140 2196 39142
rect 1956 39120 2252 39140
rect 1956 38108 2252 38128
rect 2012 38106 2036 38108
rect 2092 38106 2116 38108
rect 2172 38106 2196 38108
rect 2034 38054 2036 38106
rect 2098 38054 2110 38106
rect 2172 38054 2174 38106
rect 2012 38052 2036 38054
rect 2092 38052 2116 38054
rect 2172 38052 2196 38054
rect 1956 38032 2252 38052
rect 1956 37020 2252 37040
rect 2012 37018 2036 37020
rect 2092 37018 2116 37020
rect 2172 37018 2196 37020
rect 2034 36966 2036 37018
rect 2098 36966 2110 37018
rect 2172 36966 2174 37018
rect 2012 36964 2036 36966
rect 2092 36964 2116 36966
rect 2172 36964 2196 36966
rect 1956 36944 2252 36964
rect 1956 35932 2252 35952
rect 2012 35930 2036 35932
rect 2092 35930 2116 35932
rect 2172 35930 2196 35932
rect 2034 35878 2036 35930
rect 2098 35878 2110 35930
rect 2172 35878 2174 35930
rect 2012 35876 2036 35878
rect 2092 35876 2116 35878
rect 2172 35876 2196 35878
rect 1956 35856 2252 35876
rect 1956 34844 2252 34864
rect 2012 34842 2036 34844
rect 2092 34842 2116 34844
rect 2172 34842 2196 34844
rect 2034 34790 2036 34842
rect 2098 34790 2110 34842
rect 2172 34790 2174 34842
rect 2012 34788 2036 34790
rect 2092 34788 2116 34790
rect 2172 34788 2196 34790
rect 1956 34768 2252 34788
rect 1956 33756 2252 33776
rect 2012 33754 2036 33756
rect 2092 33754 2116 33756
rect 2172 33754 2196 33756
rect 2034 33702 2036 33754
rect 2098 33702 2110 33754
rect 2172 33702 2174 33754
rect 2012 33700 2036 33702
rect 2092 33700 2116 33702
rect 2172 33700 2196 33702
rect 1956 33680 2252 33700
rect 1956 32668 2252 32688
rect 2012 32666 2036 32668
rect 2092 32666 2116 32668
rect 2172 32666 2196 32668
rect 2034 32614 2036 32666
rect 2098 32614 2110 32666
rect 2172 32614 2174 32666
rect 2012 32612 2036 32614
rect 2092 32612 2116 32614
rect 2172 32612 2196 32614
rect 1956 32592 2252 32612
rect 1956 31580 2252 31600
rect 2012 31578 2036 31580
rect 2092 31578 2116 31580
rect 2172 31578 2196 31580
rect 2034 31526 2036 31578
rect 2098 31526 2110 31578
rect 2172 31526 2174 31578
rect 2012 31524 2036 31526
rect 2092 31524 2116 31526
rect 2172 31524 2196 31526
rect 1956 31504 2252 31524
rect 1956 30492 2252 30512
rect 2012 30490 2036 30492
rect 2092 30490 2116 30492
rect 2172 30490 2196 30492
rect 2034 30438 2036 30490
rect 2098 30438 2110 30490
rect 2172 30438 2174 30490
rect 2012 30436 2036 30438
rect 2092 30436 2116 30438
rect 2172 30436 2196 30438
rect 1956 30416 2252 30436
rect 1956 29404 2252 29424
rect 2012 29402 2036 29404
rect 2092 29402 2116 29404
rect 2172 29402 2196 29404
rect 2034 29350 2036 29402
rect 2098 29350 2110 29402
rect 2172 29350 2174 29402
rect 2012 29348 2036 29350
rect 2092 29348 2116 29350
rect 2172 29348 2196 29350
rect 1956 29328 2252 29348
rect 1956 28316 2252 28336
rect 2012 28314 2036 28316
rect 2092 28314 2116 28316
rect 2172 28314 2196 28316
rect 2034 28262 2036 28314
rect 2098 28262 2110 28314
rect 2172 28262 2174 28314
rect 2012 28260 2036 28262
rect 2092 28260 2116 28262
rect 2172 28260 2196 28262
rect 1956 28240 2252 28260
rect 1956 27228 2252 27248
rect 2012 27226 2036 27228
rect 2092 27226 2116 27228
rect 2172 27226 2196 27228
rect 2034 27174 2036 27226
rect 2098 27174 2110 27226
rect 2172 27174 2174 27226
rect 2012 27172 2036 27174
rect 2092 27172 2116 27174
rect 2172 27172 2196 27174
rect 1956 27152 2252 27172
rect 1956 26140 2252 26160
rect 2012 26138 2036 26140
rect 2092 26138 2116 26140
rect 2172 26138 2196 26140
rect 2034 26086 2036 26138
rect 2098 26086 2110 26138
rect 2172 26086 2174 26138
rect 2012 26084 2036 26086
rect 2092 26084 2116 26086
rect 2172 26084 2196 26086
rect 1956 26064 2252 26084
rect 1956 25052 2252 25072
rect 2012 25050 2036 25052
rect 2092 25050 2116 25052
rect 2172 25050 2196 25052
rect 2034 24998 2036 25050
rect 2098 24998 2110 25050
rect 2172 24998 2174 25050
rect 2012 24996 2036 24998
rect 2092 24996 2116 24998
rect 2172 24996 2196 24998
rect 1956 24976 2252 24996
rect 1956 23964 2252 23984
rect 2012 23962 2036 23964
rect 2092 23962 2116 23964
rect 2172 23962 2196 23964
rect 2034 23910 2036 23962
rect 2098 23910 2110 23962
rect 2172 23910 2174 23962
rect 2012 23908 2036 23910
rect 2092 23908 2116 23910
rect 2172 23908 2196 23910
rect 1956 23888 2252 23908
rect 1956 22876 2252 22896
rect 2012 22874 2036 22876
rect 2092 22874 2116 22876
rect 2172 22874 2196 22876
rect 2034 22822 2036 22874
rect 2098 22822 2110 22874
rect 2172 22822 2174 22874
rect 2012 22820 2036 22822
rect 2092 22820 2116 22822
rect 2172 22820 2196 22822
rect 1956 22800 2252 22820
rect 1956 21788 2252 21808
rect 2012 21786 2036 21788
rect 2092 21786 2116 21788
rect 2172 21786 2196 21788
rect 2034 21734 2036 21786
rect 2098 21734 2110 21786
rect 2172 21734 2174 21786
rect 2012 21732 2036 21734
rect 2092 21732 2116 21734
rect 2172 21732 2196 21734
rect 1956 21712 2252 21732
rect 1956 20700 2252 20720
rect 2012 20698 2036 20700
rect 2092 20698 2116 20700
rect 2172 20698 2196 20700
rect 2034 20646 2036 20698
rect 2098 20646 2110 20698
rect 2172 20646 2174 20698
rect 2012 20644 2036 20646
rect 2092 20644 2116 20646
rect 2172 20644 2196 20646
rect 1956 20624 2252 20644
rect 1956 19612 2252 19632
rect 2012 19610 2036 19612
rect 2092 19610 2116 19612
rect 2172 19610 2196 19612
rect 2034 19558 2036 19610
rect 2098 19558 2110 19610
rect 2172 19558 2174 19610
rect 2012 19556 2036 19558
rect 2092 19556 2116 19558
rect 2172 19556 2196 19558
rect 1956 19536 2252 19556
rect 1956 18524 2252 18544
rect 2012 18522 2036 18524
rect 2092 18522 2116 18524
rect 2172 18522 2196 18524
rect 2034 18470 2036 18522
rect 2098 18470 2110 18522
rect 2172 18470 2174 18522
rect 2012 18468 2036 18470
rect 2092 18468 2116 18470
rect 2172 18468 2196 18470
rect 1956 18448 2252 18468
rect 1956 17436 2252 17456
rect 2012 17434 2036 17436
rect 2092 17434 2116 17436
rect 2172 17434 2196 17436
rect 2034 17382 2036 17434
rect 2098 17382 2110 17434
rect 2172 17382 2174 17434
rect 2012 17380 2036 17382
rect 2092 17380 2116 17382
rect 2172 17380 2196 17382
rect 1956 17360 2252 17380
rect 1956 16348 2252 16368
rect 2012 16346 2036 16348
rect 2092 16346 2116 16348
rect 2172 16346 2196 16348
rect 2034 16294 2036 16346
rect 2098 16294 2110 16346
rect 2172 16294 2174 16346
rect 2012 16292 2036 16294
rect 2092 16292 2116 16294
rect 2172 16292 2196 16294
rect 1956 16272 2252 16292
rect 1956 15260 2252 15280
rect 2012 15258 2036 15260
rect 2092 15258 2116 15260
rect 2172 15258 2196 15260
rect 2034 15206 2036 15258
rect 2098 15206 2110 15258
rect 2172 15206 2174 15258
rect 2012 15204 2036 15206
rect 2092 15204 2116 15206
rect 2172 15204 2196 15206
rect 1956 15184 2252 15204
rect 1956 14172 2252 14192
rect 2012 14170 2036 14172
rect 2092 14170 2116 14172
rect 2172 14170 2196 14172
rect 2034 14118 2036 14170
rect 2098 14118 2110 14170
rect 2172 14118 2174 14170
rect 2012 14116 2036 14118
rect 2092 14116 2116 14118
rect 2172 14116 2196 14118
rect 1956 14096 2252 14116
rect 1956 13084 2252 13104
rect 2012 13082 2036 13084
rect 2092 13082 2116 13084
rect 2172 13082 2196 13084
rect 2034 13030 2036 13082
rect 2098 13030 2110 13082
rect 2172 13030 2174 13082
rect 2012 13028 2036 13030
rect 2092 13028 2116 13030
rect 2172 13028 2196 13030
rect 1956 13008 2252 13028
rect 1956 11996 2252 12016
rect 2012 11994 2036 11996
rect 2092 11994 2116 11996
rect 2172 11994 2196 11996
rect 2034 11942 2036 11994
rect 2098 11942 2110 11994
rect 2172 11942 2174 11994
rect 2012 11940 2036 11942
rect 2092 11940 2116 11942
rect 2172 11940 2196 11942
rect 1956 11920 2252 11940
rect 1956 10908 2252 10928
rect 2012 10906 2036 10908
rect 2092 10906 2116 10908
rect 2172 10906 2196 10908
rect 2034 10854 2036 10906
rect 2098 10854 2110 10906
rect 2172 10854 2174 10906
rect 2012 10852 2036 10854
rect 2092 10852 2116 10854
rect 2172 10852 2196 10854
rect 1956 10832 2252 10852
rect 1956 9820 2252 9840
rect 2012 9818 2036 9820
rect 2092 9818 2116 9820
rect 2172 9818 2196 9820
rect 2034 9766 2036 9818
rect 2098 9766 2110 9818
rect 2172 9766 2174 9818
rect 2012 9764 2036 9766
rect 2092 9764 2116 9766
rect 2172 9764 2196 9766
rect 1956 9744 2252 9764
rect 1956 8732 2252 8752
rect 2012 8730 2036 8732
rect 2092 8730 2116 8732
rect 2172 8730 2196 8732
rect 2034 8678 2036 8730
rect 2098 8678 2110 8730
rect 2172 8678 2174 8730
rect 2012 8676 2036 8678
rect 2092 8676 2116 8678
rect 2172 8676 2196 8678
rect 1956 8656 2252 8676
rect 1956 7644 2252 7664
rect 2012 7642 2036 7644
rect 2092 7642 2116 7644
rect 2172 7642 2196 7644
rect 2034 7590 2036 7642
rect 2098 7590 2110 7642
rect 2172 7590 2174 7642
rect 2012 7588 2036 7590
rect 2092 7588 2116 7590
rect 2172 7588 2196 7590
rect 1956 7568 2252 7588
rect 1956 6556 2252 6576
rect 2012 6554 2036 6556
rect 2092 6554 2116 6556
rect 2172 6554 2196 6556
rect 2034 6502 2036 6554
rect 2098 6502 2110 6554
rect 2172 6502 2174 6554
rect 2012 6500 2036 6502
rect 2092 6500 2116 6502
rect 2172 6500 2196 6502
rect 1956 6480 2252 6500
rect 1956 5468 2252 5488
rect 2012 5466 2036 5468
rect 2092 5466 2116 5468
rect 2172 5466 2196 5468
rect 2034 5414 2036 5466
rect 2098 5414 2110 5466
rect 2172 5414 2174 5466
rect 2012 5412 2036 5414
rect 2092 5412 2116 5414
rect 2172 5412 2196 5414
rect 1956 5392 2252 5412
rect 1956 4380 2252 4400
rect 2012 4378 2036 4380
rect 2092 4378 2116 4380
rect 2172 4378 2196 4380
rect 2034 4326 2036 4378
rect 2098 4326 2110 4378
rect 2172 4326 2174 4378
rect 2012 4324 2036 4326
rect 2092 4324 2116 4326
rect 2172 4324 2196 4326
rect 1956 4304 2252 4324
rect 1956 3292 2252 3312
rect 2012 3290 2036 3292
rect 2092 3290 2116 3292
rect 2172 3290 2196 3292
rect 2034 3238 2036 3290
rect 2098 3238 2110 3290
rect 2172 3238 2174 3290
rect 2012 3236 2036 3238
rect 2092 3236 2116 3238
rect 2172 3236 2196 3238
rect 1956 3216 2252 3236
rect 2516 3126 2544 84166
rect 2504 3120 2556 3126
rect 2504 3062 2556 3068
rect 3252 2582 3280 96478
rect 3332 96416 3384 96422
rect 3332 96358 3384 96364
rect 3344 96150 3372 96358
rect 3332 96144 3384 96150
rect 3332 96086 3384 96092
rect 3436 84194 3464 96630
rect 3344 84166 3464 84194
rect 3344 3738 3372 84166
rect 3620 16574 3648 97174
rect 3700 96416 3752 96422
rect 3700 96358 3752 96364
rect 3712 95402 3740 96358
rect 3956 96316 4252 96336
rect 4012 96314 4036 96316
rect 4092 96314 4116 96316
rect 4172 96314 4196 96316
rect 4034 96262 4036 96314
rect 4098 96262 4110 96314
rect 4172 96262 4174 96314
rect 4012 96260 4036 96262
rect 4092 96260 4116 96262
rect 4172 96260 4196 96262
rect 3956 96240 4252 96260
rect 3700 95396 3752 95402
rect 3700 95338 3752 95344
rect 3884 95396 3936 95402
rect 3884 95338 3936 95344
rect 3620 16546 3740 16574
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 3608 3392 3660 3398
rect 3514 3360 3570 3369
rect 3608 3334 3660 3340
rect 3514 3295 3570 3304
rect 3528 3194 3556 3295
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 3620 2961 3648 3334
rect 3712 3194 3740 16546
rect 3896 4146 3924 95338
rect 3956 95228 4252 95248
rect 4012 95226 4036 95228
rect 4092 95226 4116 95228
rect 4172 95226 4196 95228
rect 4034 95174 4036 95226
rect 4098 95174 4110 95226
rect 4172 95174 4174 95226
rect 4012 95172 4036 95174
rect 4092 95172 4116 95174
rect 4172 95172 4196 95174
rect 3956 95152 4252 95172
rect 4356 94994 4384 98534
rect 4436 98048 4488 98054
rect 4436 97990 4488 97996
rect 4528 98048 4580 98054
rect 4528 97990 4580 97996
rect 4344 94988 4396 94994
rect 4344 94930 4396 94936
rect 3956 94140 4252 94160
rect 4012 94138 4036 94140
rect 4092 94138 4116 94140
rect 4172 94138 4196 94140
rect 4034 94086 4036 94138
rect 4098 94086 4110 94138
rect 4172 94086 4174 94138
rect 4012 94084 4036 94086
rect 4092 94084 4116 94086
rect 4172 94084 4196 94086
rect 3956 94064 4252 94084
rect 3956 93052 4252 93072
rect 4012 93050 4036 93052
rect 4092 93050 4116 93052
rect 4172 93050 4196 93052
rect 4034 92998 4036 93050
rect 4098 92998 4110 93050
rect 4172 92998 4174 93050
rect 4012 92996 4036 92998
rect 4092 92996 4116 92998
rect 4172 92996 4196 92998
rect 3956 92976 4252 92996
rect 3956 91964 4252 91984
rect 4012 91962 4036 91964
rect 4092 91962 4116 91964
rect 4172 91962 4196 91964
rect 4034 91910 4036 91962
rect 4098 91910 4110 91962
rect 4172 91910 4174 91962
rect 4012 91908 4036 91910
rect 4092 91908 4116 91910
rect 4172 91908 4196 91910
rect 3956 91888 4252 91908
rect 3956 90876 4252 90896
rect 4012 90874 4036 90876
rect 4092 90874 4116 90876
rect 4172 90874 4196 90876
rect 4034 90822 4036 90874
rect 4098 90822 4110 90874
rect 4172 90822 4174 90874
rect 4012 90820 4036 90822
rect 4092 90820 4116 90822
rect 4172 90820 4196 90822
rect 3956 90800 4252 90820
rect 4356 90574 4384 94930
rect 4448 94790 4476 97990
rect 4436 94784 4488 94790
rect 4436 94726 4488 94732
rect 4448 94246 4476 94726
rect 4540 94586 4568 97990
rect 4620 96552 4672 96558
rect 4620 96494 4672 96500
rect 4528 94580 4580 94586
rect 4528 94522 4580 94528
rect 4436 94240 4488 94246
rect 4436 94182 4488 94188
rect 4540 93906 4568 94522
rect 4528 93900 4580 93906
rect 4528 93842 4580 93848
rect 4528 93696 4580 93702
rect 4528 93638 4580 93644
rect 4434 93528 4490 93537
rect 4434 93463 4490 93472
rect 4344 90568 4396 90574
rect 4344 90510 4396 90516
rect 4344 90432 4396 90438
rect 4344 90374 4396 90380
rect 3956 89788 4252 89808
rect 4012 89786 4036 89788
rect 4092 89786 4116 89788
rect 4172 89786 4196 89788
rect 4034 89734 4036 89786
rect 4098 89734 4110 89786
rect 4172 89734 4174 89786
rect 4012 89732 4036 89734
rect 4092 89732 4116 89734
rect 4172 89732 4196 89734
rect 3956 89712 4252 89732
rect 4356 89010 4384 90374
rect 4344 89004 4396 89010
rect 4344 88946 4396 88952
rect 4344 88868 4396 88874
rect 4344 88810 4396 88816
rect 3956 88700 4252 88720
rect 4012 88698 4036 88700
rect 4092 88698 4116 88700
rect 4172 88698 4196 88700
rect 4034 88646 4036 88698
rect 4098 88646 4110 88698
rect 4172 88646 4174 88698
rect 4012 88644 4036 88646
rect 4092 88644 4116 88646
rect 4172 88644 4196 88646
rect 3956 88624 4252 88644
rect 3956 87612 4252 87632
rect 4012 87610 4036 87612
rect 4092 87610 4116 87612
rect 4172 87610 4196 87612
rect 4034 87558 4036 87610
rect 4098 87558 4110 87610
rect 4172 87558 4174 87610
rect 4012 87556 4036 87558
rect 4092 87556 4116 87558
rect 4172 87556 4196 87558
rect 3956 87536 4252 87556
rect 3956 86524 4252 86544
rect 4012 86522 4036 86524
rect 4092 86522 4116 86524
rect 4172 86522 4196 86524
rect 4034 86470 4036 86522
rect 4098 86470 4110 86522
rect 4172 86470 4174 86522
rect 4012 86468 4036 86470
rect 4092 86468 4116 86470
rect 4172 86468 4196 86470
rect 3956 86448 4252 86468
rect 3956 85436 4252 85456
rect 4012 85434 4036 85436
rect 4092 85434 4116 85436
rect 4172 85434 4196 85436
rect 4034 85382 4036 85434
rect 4098 85382 4110 85434
rect 4172 85382 4174 85434
rect 4012 85380 4036 85382
rect 4092 85380 4116 85382
rect 4172 85380 4196 85382
rect 3956 85360 4252 85380
rect 3956 84348 4252 84368
rect 4012 84346 4036 84348
rect 4092 84346 4116 84348
rect 4172 84346 4196 84348
rect 4034 84294 4036 84346
rect 4098 84294 4110 84346
rect 4172 84294 4174 84346
rect 4012 84292 4036 84294
rect 4092 84292 4116 84294
rect 4172 84292 4196 84294
rect 3956 84272 4252 84292
rect 3956 83260 4252 83280
rect 4012 83258 4036 83260
rect 4092 83258 4116 83260
rect 4172 83258 4196 83260
rect 4034 83206 4036 83258
rect 4098 83206 4110 83258
rect 4172 83206 4174 83258
rect 4012 83204 4036 83206
rect 4092 83204 4116 83206
rect 4172 83204 4196 83206
rect 3956 83184 4252 83204
rect 3956 82172 4252 82192
rect 4012 82170 4036 82172
rect 4092 82170 4116 82172
rect 4172 82170 4196 82172
rect 4034 82118 4036 82170
rect 4098 82118 4110 82170
rect 4172 82118 4174 82170
rect 4012 82116 4036 82118
rect 4092 82116 4116 82118
rect 4172 82116 4196 82118
rect 3956 82096 4252 82116
rect 3956 81084 4252 81104
rect 4012 81082 4036 81084
rect 4092 81082 4116 81084
rect 4172 81082 4196 81084
rect 4034 81030 4036 81082
rect 4098 81030 4110 81082
rect 4172 81030 4174 81082
rect 4012 81028 4036 81030
rect 4092 81028 4116 81030
rect 4172 81028 4196 81030
rect 3956 81008 4252 81028
rect 3956 79996 4252 80016
rect 4012 79994 4036 79996
rect 4092 79994 4116 79996
rect 4172 79994 4196 79996
rect 4034 79942 4036 79994
rect 4098 79942 4110 79994
rect 4172 79942 4174 79994
rect 4012 79940 4036 79942
rect 4092 79940 4116 79942
rect 4172 79940 4196 79942
rect 3956 79920 4252 79940
rect 3956 78908 4252 78928
rect 4012 78906 4036 78908
rect 4092 78906 4116 78908
rect 4172 78906 4196 78908
rect 4034 78854 4036 78906
rect 4098 78854 4110 78906
rect 4172 78854 4174 78906
rect 4012 78852 4036 78854
rect 4092 78852 4116 78854
rect 4172 78852 4196 78854
rect 3956 78832 4252 78852
rect 3956 77820 4252 77840
rect 4012 77818 4036 77820
rect 4092 77818 4116 77820
rect 4172 77818 4196 77820
rect 4034 77766 4036 77818
rect 4098 77766 4110 77818
rect 4172 77766 4174 77818
rect 4012 77764 4036 77766
rect 4092 77764 4116 77766
rect 4172 77764 4196 77766
rect 3956 77744 4252 77764
rect 3956 76732 4252 76752
rect 4012 76730 4036 76732
rect 4092 76730 4116 76732
rect 4172 76730 4196 76732
rect 4034 76678 4036 76730
rect 4098 76678 4110 76730
rect 4172 76678 4174 76730
rect 4012 76676 4036 76678
rect 4092 76676 4116 76678
rect 4172 76676 4196 76678
rect 3956 76656 4252 76676
rect 3956 75644 4252 75664
rect 4012 75642 4036 75644
rect 4092 75642 4116 75644
rect 4172 75642 4196 75644
rect 4034 75590 4036 75642
rect 4098 75590 4110 75642
rect 4172 75590 4174 75642
rect 4012 75588 4036 75590
rect 4092 75588 4116 75590
rect 4172 75588 4196 75590
rect 3956 75568 4252 75588
rect 3956 74556 4252 74576
rect 4012 74554 4036 74556
rect 4092 74554 4116 74556
rect 4172 74554 4196 74556
rect 4034 74502 4036 74554
rect 4098 74502 4110 74554
rect 4172 74502 4174 74554
rect 4012 74500 4036 74502
rect 4092 74500 4116 74502
rect 4172 74500 4196 74502
rect 3956 74480 4252 74500
rect 3956 73468 4252 73488
rect 4012 73466 4036 73468
rect 4092 73466 4116 73468
rect 4172 73466 4196 73468
rect 4034 73414 4036 73466
rect 4098 73414 4110 73466
rect 4172 73414 4174 73466
rect 4012 73412 4036 73414
rect 4092 73412 4116 73414
rect 4172 73412 4196 73414
rect 3956 73392 4252 73412
rect 3956 72380 4252 72400
rect 4012 72378 4036 72380
rect 4092 72378 4116 72380
rect 4172 72378 4196 72380
rect 4034 72326 4036 72378
rect 4098 72326 4110 72378
rect 4172 72326 4174 72378
rect 4012 72324 4036 72326
rect 4092 72324 4116 72326
rect 4172 72324 4196 72326
rect 3956 72304 4252 72324
rect 3956 71292 4252 71312
rect 4012 71290 4036 71292
rect 4092 71290 4116 71292
rect 4172 71290 4196 71292
rect 4034 71238 4036 71290
rect 4098 71238 4110 71290
rect 4172 71238 4174 71290
rect 4012 71236 4036 71238
rect 4092 71236 4116 71238
rect 4172 71236 4196 71238
rect 3956 71216 4252 71236
rect 3956 70204 4252 70224
rect 4012 70202 4036 70204
rect 4092 70202 4116 70204
rect 4172 70202 4196 70204
rect 4034 70150 4036 70202
rect 4098 70150 4110 70202
rect 4172 70150 4174 70202
rect 4012 70148 4036 70150
rect 4092 70148 4116 70150
rect 4172 70148 4196 70150
rect 3956 70128 4252 70148
rect 3956 69116 4252 69136
rect 4012 69114 4036 69116
rect 4092 69114 4116 69116
rect 4172 69114 4196 69116
rect 4034 69062 4036 69114
rect 4098 69062 4110 69114
rect 4172 69062 4174 69114
rect 4012 69060 4036 69062
rect 4092 69060 4116 69062
rect 4172 69060 4196 69062
rect 3956 69040 4252 69060
rect 3956 68028 4252 68048
rect 4012 68026 4036 68028
rect 4092 68026 4116 68028
rect 4172 68026 4196 68028
rect 4034 67974 4036 68026
rect 4098 67974 4110 68026
rect 4172 67974 4174 68026
rect 4012 67972 4036 67974
rect 4092 67972 4116 67974
rect 4172 67972 4196 67974
rect 3956 67952 4252 67972
rect 3956 66940 4252 66960
rect 4012 66938 4036 66940
rect 4092 66938 4116 66940
rect 4172 66938 4196 66940
rect 4034 66886 4036 66938
rect 4098 66886 4110 66938
rect 4172 66886 4174 66938
rect 4012 66884 4036 66886
rect 4092 66884 4116 66886
rect 4172 66884 4196 66886
rect 3956 66864 4252 66884
rect 3956 65852 4252 65872
rect 4012 65850 4036 65852
rect 4092 65850 4116 65852
rect 4172 65850 4196 65852
rect 4034 65798 4036 65850
rect 4098 65798 4110 65850
rect 4172 65798 4174 65850
rect 4012 65796 4036 65798
rect 4092 65796 4116 65798
rect 4172 65796 4196 65798
rect 3956 65776 4252 65796
rect 3956 64764 4252 64784
rect 4012 64762 4036 64764
rect 4092 64762 4116 64764
rect 4172 64762 4196 64764
rect 4034 64710 4036 64762
rect 4098 64710 4110 64762
rect 4172 64710 4174 64762
rect 4012 64708 4036 64710
rect 4092 64708 4116 64710
rect 4172 64708 4196 64710
rect 3956 64688 4252 64708
rect 3956 63676 4252 63696
rect 4012 63674 4036 63676
rect 4092 63674 4116 63676
rect 4172 63674 4196 63676
rect 4034 63622 4036 63674
rect 4098 63622 4110 63674
rect 4172 63622 4174 63674
rect 4012 63620 4036 63622
rect 4092 63620 4116 63622
rect 4172 63620 4196 63622
rect 3956 63600 4252 63620
rect 3956 62588 4252 62608
rect 4012 62586 4036 62588
rect 4092 62586 4116 62588
rect 4172 62586 4196 62588
rect 4034 62534 4036 62586
rect 4098 62534 4110 62586
rect 4172 62534 4174 62586
rect 4012 62532 4036 62534
rect 4092 62532 4116 62534
rect 4172 62532 4196 62534
rect 3956 62512 4252 62532
rect 3956 61500 4252 61520
rect 4012 61498 4036 61500
rect 4092 61498 4116 61500
rect 4172 61498 4196 61500
rect 4034 61446 4036 61498
rect 4098 61446 4110 61498
rect 4172 61446 4174 61498
rect 4012 61444 4036 61446
rect 4092 61444 4116 61446
rect 4172 61444 4196 61446
rect 3956 61424 4252 61444
rect 3956 60412 4252 60432
rect 4012 60410 4036 60412
rect 4092 60410 4116 60412
rect 4172 60410 4196 60412
rect 4034 60358 4036 60410
rect 4098 60358 4110 60410
rect 4172 60358 4174 60410
rect 4012 60356 4036 60358
rect 4092 60356 4116 60358
rect 4172 60356 4196 60358
rect 3956 60336 4252 60356
rect 3956 59324 4252 59344
rect 4012 59322 4036 59324
rect 4092 59322 4116 59324
rect 4172 59322 4196 59324
rect 4034 59270 4036 59322
rect 4098 59270 4110 59322
rect 4172 59270 4174 59322
rect 4012 59268 4036 59270
rect 4092 59268 4116 59270
rect 4172 59268 4196 59270
rect 3956 59248 4252 59268
rect 3956 58236 4252 58256
rect 4012 58234 4036 58236
rect 4092 58234 4116 58236
rect 4172 58234 4196 58236
rect 4034 58182 4036 58234
rect 4098 58182 4110 58234
rect 4172 58182 4174 58234
rect 4012 58180 4036 58182
rect 4092 58180 4116 58182
rect 4172 58180 4196 58182
rect 3956 58160 4252 58180
rect 3956 57148 4252 57168
rect 4012 57146 4036 57148
rect 4092 57146 4116 57148
rect 4172 57146 4196 57148
rect 4034 57094 4036 57146
rect 4098 57094 4110 57146
rect 4172 57094 4174 57146
rect 4012 57092 4036 57094
rect 4092 57092 4116 57094
rect 4172 57092 4196 57094
rect 3956 57072 4252 57092
rect 3956 56060 4252 56080
rect 4012 56058 4036 56060
rect 4092 56058 4116 56060
rect 4172 56058 4196 56060
rect 4034 56006 4036 56058
rect 4098 56006 4110 56058
rect 4172 56006 4174 56058
rect 4012 56004 4036 56006
rect 4092 56004 4116 56006
rect 4172 56004 4196 56006
rect 3956 55984 4252 56004
rect 3956 54972 4252 54992
rect 4012 54970 4036 54972
rect 4092 54970 4116 54972
rect 4172 54970 4196 54972
rect 4034 54918 4036 54970
rect 4098 54918 4110 54970
rect 4172 54918 4174 54970
rect 4012 54916 4036 54918
rect 4092 54916 4116 54918
rect 4172 54916 4196 54918
rect 3956 54896 4252 54916
rect 3956 53884 4252 53904
rect 4012 53882 4036 53884
rect 4092 53882 4116 53884
rect 4172 53882 4196 53884
rect 4034 53830 4036 53882
rect 4098 53830 4110 53882
rect 4172 53830 4174 53882
rect 4012 53828 4036 53830
rect 4092 53828 4116 53830
rect 4172 53828 4196 53830
rect 3956 53808 4252 53828
rect 3956 52796 4252 52816
rect 4012 52794 4036 52796
rect 4092 52794 4116 52796
rect 4172 52794 4196 52796
rect 4034 52742 4036 52794
rect 4098 52742 4110 52794
rect 4172 52742 4174 52794
rect 4012 52740 4036 52742
rect 4092 52740 4116 52742
rect 4172 52740 4196 52742
rect 3956 52720 4252 52740
rect 3956 51708 4252 51728
rect 4012 51706 4036 51708
rect 4092 51706 4116 51708
rect 4172 51706 4196 51708
rect 4034 51654 4036 51706
rect 4098 51654 4110 51706
rect 4172 51654 4174 51706
rect 4012 51652 4036 51654
rect 4092 51652 4116 51654
rect 4172 51652 4196 51654
rect 3956 51632 4252 51652
rect 3956 50620 4252 50640
rect 4012 50618 4036 50620
rect 4092 50618 4116 50620
rect 4172 50618 4196 50620
rect 4034 50566 4036 50618
rect 4098 50566 4110 50618
rect 4172 50566 4174 50618
rect 4012 50564 4036 50566
rect 4092 50564 4116 50566
rect 4172 50564 4196 50566
rect 3956 50544 4252 50564
rect 3956 49532 4252 49552
rect 4012 49530 4036 49532
rect 4092 49530 4116 49532
rect 4172 49530 4196 49532
rect 4034 49478 4036 49530
rect 4098 49478 4110 49530
rect 4172 49478 4174 49530
rect 4012 49476 4036 49478
rect 4092 49476 4116 49478
rect 4172 49476 4196 49478
rect 3956 49456 4252 49476
rect 3956 48444 4252 48464
rect 4012 48442 4036 48444
rect 4092 48442 4116 48444
rect 4172 48442 4196 48444
rect 4034 48390 4036 48442
rect 4098 48390 4110 48442
rect 4172 48390 4174 48442
rect 4012 48388 4036 48390
rect 4092 48388 4116 48390
rect 4172 48388 4196 48390
rect 3956 48368 4252 48388
rect 3956 47356 4252 47376
rect 4012 47354 4036 47356
rect 4092 47354 4116 47356
rect 4172 47354 4196 47356
rect 4034 47302 4036 47354
rect 4098 47302 4110 47354
rect 4172 47302 4174 47354
rect 4012 47300 4036 47302
rect 4092 47300 4116 47302
rect 4172 47300 4196 47302
rect 3956 47280 4252 47300
rect 3956 46268 4252 46288
rect 4012 46266 4036 46268
rect 4092 46266 4116 46268
rect 4172 46266 4196 46268
rect 4034 46214 4036 46266
rect 4098 46214 4110 46266
rect 4172 46214 4174 46266
rect 4012 46212 4036 46214
rect 4092 46212 4116 46214
rect 4172 46212 4196 46214
rect 3956 46192 4252 46212
rect 3956 45180 4252 45200
rect 4012 45178 4036 45180
rect 4092 45178 4116 45180
rect 4172 45178 4196 45180
rect 4034 45126 4036 45178
rect 4098 45126 4110 45178
rect 4172 45126 4174 45178
rect 4012 45124 4036 45126
rect 4092 45124 4116 45126
rect 4172 45124 4196 45126
rect 3956 45104 4252 45124
rect 3956 44092 4252 44112
rect 4012 44090 4036 44092
rect 4092 44090 4116 44092
rect 4172 44090 4196 44092
rect 4034 44038 4036 44090
rect 4098 44038 4110 44090
rect 4172 44038 4174 44090
rect 4012 44036 4036 44038
rect 4092 44036 4116 44038
rect 4172 44036 4196 44038
rect 3956 44016 4252 44036
rect 3956 43004 4252 43024
rect 4012 43002 4036 43004
rect 4092 43002 4116 43004
rect 4172 43002 4196 43004
rect 4034 42950 4036 43002
rect 4098 42950 4110 43002
rect 4172 42950 4174 43002
rect 4012 42948 4036 42950
rect 4092 42948 4116 42950
rect 4172 42948 4196 42950
rect 3956 42928 4252 42948
rect 3956 41916 4252 41936
rect 4012 41914 4036 41916
rect 4092 41914 4116 41916
rect 4172 41914 4196 41916
rect 4034 41862 4036 41914
rect 4098 41862 4110 41914
rect 4172 41862 4174 41914
rect 4012 41860 4036 41862
rect 4092 41860 4116 41862
rect 4172 41860 4196 41862
rect 3956 41840 4252 41860
rect 3956 40828 4252 40848
rect 4012 40826 4036 40828
rect 4092 40826 4116 40828
rect 4172 40826 4196 40828
rect 4034 40774 4036 40826
rect 4098 40774 4110 40826
rect 4172 40774 4174 40826
rect 4012 40772 4036 40774
rect 4092 40772 4116 40774
rect 4172 40772 4196 40774
rect 3956 40752 4252 40772
rect 3956 39740 4252 39760
rect 4012 39738 4036 39740
rect 4092 39738 4116 39740
rect 4172 39738 4196 39740
rect 4034 39686 4036 39738
rect 4098 39686 4110 39738
rect 4172 39686 4174 39738
rect 4012 39684 4036 39686
rect 4092 39684 4116 39686
rect 4172 39684 4196 39686
rect 3956 39664 4252 39684
rect 3956 38652 4252 38672
rect 4012 38650 4036 38652
rect 4092 38650 4116 38652
rect 4172 38650 4196 38652
rect 4034 38598 4036 38650
rect 4098 38598 4110 38650
rect 4172 38598 4174 38650
rect 4012 38596 4036 38598
rect 4092 38596 4116 38598
rect 4172 38596 4196 38598
rect 3956 38576 4252 38596
rect 3956 37564 4252 37584
rect 4012 37562 4036 37564
rect 4092 37562 4116 37564
rect 4172 37562 4196 37564
rect 4034 37510 4036 37562
rect 4098 37510 4110 37562
rect 4172 37510 4174 37562
rect 4012 37508 4036 37510
rect 4092 37508 4116 37510
rect 4172 37508 4196 37510
rect 3956 37488 4252 37508
rect 3956 36476 4252 36496
rect 4012 36474 4036 36476
rect 4092 36474 4116 36476
rect 4172 36474 4196 36476
rect 4034 36422 4036 36474
rect 4098 36422 4110 36474
rect 4172 36422 4174 36474
rect 4012 36420 4036 36422
rect 4092 36420 4116 36422
rect 4172 36420 4196 36422
rect 3956 36400 4252 36420
rect 3956 35388 4252 35408
rect 4012 35386 4036 35388
rect 4092 35386 4116 35388
rect 4172 35386 4196 35388
rect 4034 35334 4036 35386
rect 4098 35334 4110 35386
rect 4172 35334 4174 35386
rect 4012 35332 4036 35334
rect 4092 35332 4116 35334
rect 4172 35332 4196 35334
rect 3956 35312 4252 35332
rect 3956 34300 4252 34320
rect 4012 34298 4036 34300
rect 4092 34298 4116 34300
rect 4172 34298 4196 34300
rect 4034 34246 4036 34298
rect 4098 34246 4110 34298
rect 4172 34246 4174 34298
rect 4012 34244 4036 34246
rect 4092 34244 4116 34246
rect 4172 34244 4196 34246
rect 3956 34224 4252 34244
rect 3956 33212 4252 33232
rect 4012 33210 4036 33212
rect 4092 33210 4116 33212
rect 4172 33210 4196 33212
rect 4034 33158 4036 33210
rect 4098 33158 4110 33210
rect 4172 33158 4174 33210
rect 4012 33156 4036 33158
rect 4092 33156 4116 33158
rect 4172 33156 4196 33158
rect 3956 33136 4252 33156
rect 3956 32124 4252 32144
rect 4012 32122 4036 32124
rect 4092 32122 4116 32124
rect 4172 32122 4196 32124
rect 4034 32070 4036 32122
rect 4098 32070 4110 32122
rect 4172 32070 4174 32122
rect 4012 32068 4036 32070
rect 4092 32068 4116 32070
rect 4172 32068 4196 32070
rect 3956 32048 4252 32068
rect 3956 31036 4252 31056
rect 4012 31034 4036 31036
rect 4092 31034 4116 31036
rect 4172 31034 4196 31036
rect 4034 30982 4036 31034
rect 4098 30982 4110 31034
rect 4172 30982 4174 31034
rect 4012 30980 4036 30982
rect 4092 30980 4116 30982
rect 4172 30980 4196 30982
rect 3956 30960 4252 30980
rect 3956 29948 4252 29968
rect 4012 29946 4036 29948
rect 4092 29946 4116 29948
rect 4172 29946 4196 29948
rect 4034 29894 4036 29946
rect 4098 29894 4110 29946
rect 4172 29894 4174 29946
rect 4012 29892 4036 29894
rect 4092 29892 4116 29894
rect 4172 29892 4196 29894
rect 3956 29872 4252 29892
rect 3956 28860 4252 28880
rect 4012 28858 4036 28860
rect 4092 28858 4116 28860
rect 4172 28858 4196 28860
rect 4034 28806 4036 28858
rect 4098 28806 4110 28858
rect 4172 28806 4174 28858
rect 4012 28804 4036 28806
rect 4092 28804 4116 28806
rect 4172 28804 4196 28806
rect 3956 28784 4252 28804
rect 3956 27772 4252 27792
rect 4012 27770 4036 27772
rect 4092 27770 4116 27772
rect 4172 27770 4196 27772
rect 4034 27718 4036 27770
rect 4098 27718 4110 27770
rect 4172 27718 4174 27770
rect 4012 27716 4036 27718
rect 4092 27716 4116 27718
rect 4172 27716 4196 27718
rect 3956 27696 4252 27716
rect 3956 26684 4252 26704
rect 4012 26682 4036 26684
rect 4092 26682 4116 26684
rect 4172 26682 4196 26684
rect 4034 26630 4036 26682
rect 4098 26630 4110 26682
rect 4172 26630 4174 26682
rect 4012 26628 4036 26630
rect 4092 26628 4116 26630
rect 4172 26628 4196 26630
rect 3956 26608 4252 26628
rect 3956 25596 4252 25616
rect 4012 25594 4036 25596
rect 4092 25594 4116 25596
rect 4172 25594 4196 25596
rect 4034 25542 4036 25594
rect 4098 25542 4110 25594
rect 4172 25542 4174 25594
rect 4012 25540 4036 25542
rect 4092 25540 4116 25542
rect 4172 25540 4196 25542
rect 3956 25520 4252 25540
rect 3956 24508 4252 24528
rect 4012 24506 4036 24508
rect 4092 24506 4116 24508
rect 4172 24506 4196 24508
rect 4034 24454 4036 24506
rect 4098 24454 4110 24506
rect 4172 24454 4174 24506
rect 4012 24452 4036 24454
rect 4092 24452 4116 24454
rect 4172 24452 4196 24454
rect 3956 24432 4252 24452
rect 3956 23420 4252 23440
rect 4012 23418 4036 23420
rect 4092 23418 4116 23420
rect 4172 23418 4196 23420
rect 4034 23366 4036 23418
rect 4098 23366 4110 23418
rect 4172 23366 4174 23418
rect 4012 23364 4036 23366
rect 4092 23364 4116 23366
rect 4172 23364 4196 23366
rect 3956 23344 4252 23364
rect 3956 22332 4252 22352
rect 4012 22330 4036 22332
rect 4092 22330 4116 22332
rect 4172 22330 4196 22332
rect 4034 22278 4036 22330
rect 4098 22278 4110 22330
rect 4172 22278 4174 22330
rect 4012 22276 4036 22278
rect 4092 22276 4116 22278
rect 4172 22276 4196 22278
rect 3956 22256 4252 22276
rect 3956 21244 4252 21264
rect 4012 21242 4036 21244
rect 4092 21242 4116 21244
rect 4172 21242 4196 21244
rect 4034 21190 4036 21242
rect 4098 21190 4110 21242
rect 4172 21190 4174 21242
rect 4012 21188 4036 21190
rect 4092 21188 4116 21190
rect 4172 21188 4196 21190
rect 3956 21168 4252 21188
rect 3956 20156 4252 20176
rect 4012 20154 4036 20156
rect 4092 20154 4116 20156
rect 4172 20154 4196 20156
rect 4034 20102 4036 20154
rect 4098 20102 4110 20154
rect 4172 20102 4174 20154
rect 4012 20100 4036 20102
rect 4092 20100 4116 20102
rect 4172 20100 4196 20102
rect 3956 20080 4252 20100
rect 3956 19068 4252 19088
rect 4012 19066 4036 19068
rect 4092 19066 4116 19068
rect 4172 19066 4196 19068
rect 4034 19014 4036 19066
rect 4098 19014 4110 19066
rect 4172 19014 4174 19066
rect 4012 19012 4036 19014
rect 4092 19012 4116 19014
rect 4172 19012 4196 19014
rect 3956 18992 4252 19012
rect 3956 17980 4252 18000
rect 4012 17978 4036 17980
rect 4092 17978 4116 17980
rect 4172 17978 4196 17980
rect 4034 17926 4036 17978
rect 4098 17926 4110 17978
rect 4172 17926 4174 17978
rect 4012 17924 4036 17926
rect 4092 17924 4116 17926
rect 4172 17924 4196 17926
rect 3956 17904 4252 17924
rect 3956 16892 4252 16912
rect 4012 16890 4036 16892
rect 4092 16890 4116 16892
rect 4172 16890 4196 16892
rect 4034 16838 4036 16890
rect 4098 16838 4110 16890
rect 4172 16838 4174 16890
rect 4012 16836 4036 16838
rect 4092 16836 4116 16838
rect 4172 16836 4196 16838
rect 3956 16816 4252 16836
rect 3956 15804 4252 15824
rect 4012 15802 4036 15804
rect 4092 15802 4116 15804
rect 4172 15802 4196 15804
rect 4034 15750 4036 15802
rect 4098 15750 4110 15802
rect 4172 15750 4174 15802
rect 4012 15748 4036 15750
rect 4092 15748 4116 15750
rect 4172 15748 4196 15750
rect 3956 15728 4252 15748
rect 3956 14716 4252 14736
rect 4012 14714 4036 14716
rect 4092 14714 4116 14716
rect 4172 14714 4196 14716
rect 4034 14662 4036 14714
rect 4098 14662 4110 14714
rect 4172 14662 4174 14714
rect 4012 14660 4036 14662
rect 4092 14660 4116 14662
rect 4172 14660 4196 14662
rect 3956 14640 4252 14660
rect 3956 13628 4252 13648
rect 4012 13626 4036 13628
rect 4092 13626 4116 13628
rect 4172 13626 4196 13628
rect 4034 13574 4036 13626
rect 4098 13574 4110 13626
rect 4172 13574 4174 13626
rect 4012 13572 4036 13574
rect 4092 13572 4116 13574
rect 4172 13572 4196 13574
rect 3956 13552 4252 13572
rect 3956 12540 4252 12560
rect 4012 12538 4036 12540
rect 4092 12538 4116 12540
rect 4172 12538 4196 12540
rect 4034 12486 4036 12538
rect 4098 12486 4110 12538
rect 4172 12486 4174 12538
rect 4012 12484 4036 12486
rect 4092 12484 4116 12486
rect 4172 12484 4196 12486
rect 3956 12464 4252 12484
rect 3956 11452 4252 11472
rect 4012 11450 4036 11452
rect 4092 11450 4116 11452
rect 4172 11450 4196 11452
rect 4034 11398 4036 11450
rect 4098 11398 4110 11450
rect 4172 11398 4174 11450
rect 4012 11396 4036 11398
rect 4092 11396 4116 11398
rect 4172 11396 4196 11398
rect 3956 11376 4252 11396
rect 3956 10364 4252 10384
rect 4012 10362 4036 10364
rect 4092 10362 4116 10364
rect 4172 10362 4196 10364
rect 4034 10310 4036 10362
rect 4098 10310 4110 10362
rect 4172 10310 4174 10362
rect 4012 10308 4036 10310
rect 4092 10308 4116 10310
rect 4172 10308 4196 10310
rect 3956 10288 4252 10308
rect 3956 9276 4252 9296
rect 4012 9274 4036 9276
rect 4092 9274 4116 9276
rect 4172 9274 4196 9276
rect 4034 9222 4036 9274
rect 4098 9222 4110 9274
rect 4172 9222 4174 9274
rect 4012 9220 4036 9222
rect 4092 9220 4116 9222
rect 4172 9220 4196 9222
rect 3956 9200 4252 9220
rect 3956 8188 4252 8208
rect 4012 8186 4036 8188
rect 4092 8186 4116 8188
rect 4172 8186 4196 8188
rect 4034 8134 4036 8186
rect 4098 8134 4110 8186
rect 4172 8134 4174 8186
rect 4012 8132 4036 8134
rect 4092 8132 4116 8134
rect 4172 8132 4196 8134
rect 3956 8112 4252 8132
rect 3956 7100 4252 7120
rect 4012 7098 4036 7100
rect 4092 7098 4116 7100
rect 4172 7098 4196 7100
rect 4034 7046 4036 7098
rect 4098 7046 4110 7098
rect 4172 7046 4174 7098
rect 4012 7044 4036 7046
rect 4092 7044 4116 7046
rect 4172 7044 4196 7046
rect 3956 7024 4252 7044
rect 3956 6012 4252 6032
rect 4012 6010 4036 6012
rect 4092 6010 4116 6012
rect 4172 6010 4196 6012
rect 4034 5958 4036 6010
rect 4098 5958 4110 6010
rect 4172 5958 4174 6010
rect 4012 5956 4036 5958
rect 4092 5956 4116 5958
rect 4172 5956 4196 5958
rect 3956 5936 4252 5956
rect 3956 4924 4252 4944
rect 4012 4922 4036 4924
rect 4092 4922 4116 4924
rect 4172 4922 4196 4924
rect 4034 4870 4036 4922
rect 4098 4870 4110 4922
rect 4172 4870 4174 4922
rect 4012 4868 4036 4870
rect 4092 4868 4116 4870
rect 4172 4868 4196 4870
rect 3956 4848 4252 4868
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3804 3398 3832 3878
rect 3792 3392 3844 3398
rect 3792 3334 3844 3340
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 3606 2952 3662 2961
rect 3606 2887 3662 2896
rect 3240 2576 3292 2582
rect 3240 2518 3292 2524
rect 1956 2204 2252 2224
rect 2012 2202 2036 2204
rect 2092 2202 2116 2204
rect 2172 2202 2196 2204
rect 2034 2150 2036 2202
rect 2098 2150 2110 2202
rect 2172 2150 2174 2202
rect 2012 2148 2036 2150
rect 2092 2148 2116 2150
rect 2172 2148 2196 2150
rect 1956 2128 2252 2148
rect 3712 746 3740 3130
rect 3790 3088 3846 3097
rect 3790 3023 3846 3032
rect 3804 2990 3832 3023
rect 3896 2990 3924 4082
rect 3956 3836 4252 3856
rect 4012 3834 4036 3836
rect 4092 3834 4116 3836
rect 4172 3834 4196 3836
rect 4034 3782 4036 3834
rect 4098 3782 4110 3834
rect 4172 3782 4174 3834
rect 4012 3780 4036 3782
rect 4092 3780 4116 3782
rect 4172 3780 4196 3782
rect 3956 3760 4252 3780
rect 4356 3346 4384 88810
rect 4448 49978 4476 93463
rect 4540 57934 4568 93638
rect 4528 57928 4580 57934
rect 4528 57870 4580 57876
rect 4436 49972 4488 49978
rect 4436 49914 4488 49920
rect 4434 10160 4490 10169
rect 4434 10095 4436 10104
rect 4488 10095 4490 10104
rect 4436 10066 4488 10072
rect 4528 4140 4580 4146
rect 4528 4082 4580 4088
rect 4436 3664 4488 3670
rect 4436 3606 4488 3612
rect 4264 3318 4384 3346
rect 3792 2984 3844 2990
rect 3792 2926 3844 2932
rect 3884 2984 3936 2990
rect 3884 2926 3936 2932
rect 4264 2836 4292 3318
rect 4342 3224 4398 3233
rect 4342 3159 4398 3168
rect 4356 2854 4384 3159
rect 3896 2808 4292 2836
rect 4344 2848 4396 2854
rect 3896 2650 3924 2808
rect 4344 2790 4396 2796
rect 3956 2748 4252 2768
rect 4012 2746 4036 2748
rect 4092 2746 4116 2748
rect 4172 2746 4196 2748
rect 4034 2694 4036 2746
rect 4098 2694 4110 2746
rect 4172 2694 4174 2746
rect 4012 2692 4036 2694
rect 4092 2692 4116 2694
rect 4172 2692 4196 2694
rect 3956 2672 4252 2692
rect 3884 2644 3936 2650
rect 3884 2586 3936 2592
rect 3896 950 3924 2586
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 4172 1970 4200 2382
rect 4160 1964 4212 1970
rect 4160 1906 4212 1912
rect 4448 1086 4476 3606
rect 4540 3126 4568 4082
rect 4632 3233 4660 96494
rect 4724 92449 4752 176870
rect 4802 176216 4858 176225
rect 4802 176151 4804 176160
rect 4856 176151 4858 176160
rect 4804 176122 4856 176128
rect 4802 174584 4858 174593
rect 4802 174519 4804 174528
rect 4856 174519 4858 174528
rect 4804 174490 4856 174496
rect 4804 174412 4856 174418
rect 4804 174354 4856 174360
rect 4710 92440 4766 92449
rect 4710 92375 4766 92384
rect 4710 91080 4766 91089
rect 4710 91015 4766 91024
rect 4724 89321 4752 91015
rect 4710 89312 4766 89321
rect 4710 89247 4766 89256
rect 4816 89162 4844 174354
rect 4908 95946 4936 180766
rect 5184 175930 5212 182951
rect 83740 180872 83792 180878
rect 83740 180814 83792 180820
rect 5262 176216 5318 176225
rect 5262 176151 5318 176160
rect 5092 175902 5212 175930
rect 4988 174344 5040 174350
rect 4988 174286 5040 174292
rect 4896 95940 4948 95946
rect 4896 95882 4948 95888
rect 5000 95554 5028 174286
rect 5092 97170 5120 175902
rect 5276 174706 5304 176151
rect 5184 174678 5304 174706
rect 5080 97164 5132 97170
rect 5080 97106 5132 97112
rect 4908 95526 5028 95554
rect 4908 94518 4936 95526
rect 5092 95418 5120 97106
rect 5000 95390 5120 95418
rect 4896 94512 4948 94518
rect 4896 94454 4948 94460
rect 4908 90794 4936 94454
rect 5000 90930 5028 95390
rect 5184 94738 5212 174678
rect 5262 174584 5318 174593
rect 5262 174519 5318 174528
rect 5092 94710 5212 94738
rect 5092 91089 5120 94710
rect 5276 94602 5304 174519
rect 83556 167136 83608 167142
rect 83556 167078 83608 167084
rect 82452 162920 82504 162926
rect 82452 162862 82504 162868
rect 5446 121544 5502 121553
rect 5446 121479 5502 121488
rect 5354 116648 5410 116657
rect 5354 116583 5356 116592
rect 5408 116583 5410 116592
rect 5356 116554 5408 116560
rect 5460 116498 5488 121479
rect 5368 116470 5488 116498
rect 5368 98054 5396 116470
rect 5446 115016 5502 115025
rect 5446 114951 5448 114960
rect 5500 114951 5502 114960
rect 5448 114922 5500 114928
rect 5356 98048 5408 98054
rect 5356 97990 5408 97996
rect 5460 96626 5488 114922
rect 6736 98592 6788 98598
rect 6736 98534 6788 98540
rect 5816 97776 5868 97782
rect 5816 97718 5868 97724
rect 5724 97708 5776 97714
rect 5724 97650 5776 97656
rect 5632 97504 5684 97510
rect 5632 97446 5684 97452
rect 5540 97096 5592 97102
rect 5540 97038 5592 97044
rect 5448 96620 5500 96626
rect 5448 96562 5500 96568
rect 5448 95940 5500 95946
rect 5448 95882 5500 95888
rect 5356 95328 5408 95334
rect 5356 95270 5408 95276
rect 5184 94574 5304 94602
rect 5078 91080 5134 91089
rect 5078 91015 5134 91024
rect 5000 90902 5120 90930
rect 4908 90766 5028 90794
rect 4896 90704 4948 90710
rect 4896 90646 4948 90652
rect 4724 89134 4844 89162
rect 4908 89162 4936 90646
rect 5000 89298 5028 90766
rect 5092 89418 5120 90902
rect 5184 89457 5212 94574
rect 5264 94240 5316 94246
rect 5264 94182 5316 94188
rect 5170 89448 5226 89457
rect 5080 89412 5132 89418
rect 5170 89383 5226 89392
rect 5080 89354 5132 89360
rect 5000 89270 5212 89298
rect 5078 89176 5134 89185
rect 4908 89134 5028 89162
rect 4724 86737 4752 89134
rect 4804 89072 4856 89078
rect 4802 89040 4804 89049
rect 4856 89040 4858 89049
rect 4802 88975 4858 88984
rect 4896 89004 4948 89010
rect 4896 88946 4948 88952
rect 4802 88904 4858 88913
rect 4802 88839 4858 88848
rect 4710 86728 4766 86737
rect 4710 86663 4766 86672
rect 4724 85338 4752 86663
rect 4712 85332 4764 85338
rect 4712 85274 4764 85280
rect 4724 85241 4752 85274
rect 4710 85232 4766 85241
rect 4710 85167 4766 85176
rect 4816 83366 4844 88839
rect 4804 83360 4856 83366
rect 4802 83328 4804 83337
rect 4856 83328 4858 83337
rect 4802 83263 4858 83272
rect 4804 82272 4856 82278
rect 4802 82240 4804 82249
rect 4856 82240 4858 82249
rect 4802 82175 4858 82184
rect 4802 80472 4858 80481
rect 4802 80407 4804 80416
rect 4856 80407 4858 80416
rect 4804 80378 4856 80384
rect 4712 22432 4764 22438
rect 4710 22400 4712 22409
rect 4764 22400 4766 22409
rect 4710 22335 4766 22344
rect 4618 3224 4674 3233
rect 4618 3159 4674 3168
rect 4528 3120 4580 3126
rect 4528 3062 4580 3068
rect 4436 1080 4488 1086
rect 4436 1022 4488 1028
rect 4540 1018 4568 3062
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 4632 1358 4660 2790
rect 4724 2650 4752 22335
rect 4802 20904 4858 20913
rect 4802 20839 4804 20848
rect 4856 20839 4858 20848
rect 4804 20810 4856 20816
rect 4908 12434 4936 88946
rect 5000 88058 5028 89134
rect 5078 89111 5134 89120
rect 4988 88052 5040 88058
rect 4988 87994 5040 88000
rect 5000 87825 5028 87994
rect 4986 87816 5042 87825
rect 4986 87751 5042 87760
rect 5092 84194 5120 89111
rect 5184 86426 5212 89270
rect 5276 88874 5304 94182
rect 5264 88868 5316 88874
rect 5264 88810 5316 88816
rect 5262 88768 5318 88777
rect 5262 88703 5318 88712
rect 5172 86420 5224 86426
rect 5172 86362 5224 86368
rect 5184 86329 5212 86362
rect 5170 86320 5226 86329
rect 5170 86255 5226 86264
rect 5092 84166 5212 84194
rect 5184 82249 5212 84166
rect 5170 82240 5226 82249
rect 5170 82175 5226 82184
rect 5276 80481 5304 88703
rect 5262 80472 5318 80481
rect 5262 80407 5318 80416
rect 4988 20868 5040 20874
rect 4988 20810 5040 20816
rect 4816 12406 4936 12434
rect 4816 3942 4844 12406
rect 4804 3936 4856 3942
rect 4802 3904 4804 3913
rect 4856 3904 4858 3913
rect 4802 3839 4858 3848
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4620 1352 4672 1358
rect 4620 1294 4672 1300
rect 4816 1290 4844 3674
rect 4894 3088 4950 3097
rect 4894 3023 4950 3032
rect 4908 2854 4936 3023
rect 4896 2848 4948 2854
rect 4896 2790 4948 2796
rect 5000 2446 5028 20810
rect 5368 7818 5396 95270
rect 5460 90710 5488 95882
rect 5448 90704 5500 90710
rect 5448 90646 5500 90652
rect 5448 90568 5500 90574
rect 5448 90510 5500 90516
rect 5356 7812 5408 7818
rect 5356 7754 5408 7760
rect 5460 7698 5488 90510
rect 5276 7670 5488 7698
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 4804 1284 4856 1290
rect 4804 1226 4856 1232
rect 4528 1012 4580 1018
rect 4528 954 4580 960
rect 3884 944 3936 950
rect 3884 886 3936 892
rect 3700 740 3752 746
rect 3700 682 3752 688
rect 5092 678 5120 4762
rect 5172 4752 5224 4758
rect 5172 4694 5224 4700
rect 5184 814 5212 4694
rect 5276 1970 5304 7670
rect 5356 7608 5408 7614
rect 5356 7550 5408 7556
rect 5368 2825 5396 7550
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5354 2816 5410 2825
rect 5354 2751 5410 2760
rect 5264 1964 5316 1970
rect 5264 1906 5316 1912
rect 5460 1426 5488 4966
rect 5552 3194 5580 97038
rect 5644 96898 5672 97446
rect 5736 96937 5764 97650
rect 5722 96928 5778 96937
rect 5632 96892 5684 96898
rect 5722 96863 5778 96872
rect 5632 96834 5684 96840
rect 5644 3738 5672 96834
rect 5828 96665 5856 97718
rect 6748 97374 6776 98534
rect 6828 98116 6880 98122
rect 6828 98058 6880 98064
rect 6736 97368 6788 97374
rect 6736 97310 6788 97316
rect 5908 97300 5960 97306
rect 5908 97242 5960 97248
rect 5920 96801 5948 97242
rect 6460 96960 6512 96966
rect 6182 96928 6238 96937
rect 6460 96902 6512 96908
rect 6182 96863 6238 96872
rect 5906 96792 5962 96801
rect 5906 96727 5962 96736
rect 5814 96656 5870 96665
rect 5736 96614 5814 96642
rect 5736 4826 5764 96614
rect 5814 96591 5870 96600
rect 5908 96416 5960 96422
rect 5908 96358 5960 96364
rect 5816 95872 5868 95878
rect 5816 95814 5868 95820
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5552 2774 5580 3130
rect 5644 2961 5672 3470
rect 5736 3097 5764 4014
rect 5828 3670 5856 95814
rect 5920 4146 5948 96358
rect 6092 96144 6144 96150
rect 6092 96086 6144 96092
rect 6104 84194 6132 96086
rect 6012 84166 6132 84194
rect 6012 4758 6040 84166
rect 6000 4752 6052 4758
rect 6000 4694 6052 4700
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 5816 3664 5868 3670
rect 5816 3606 5868 3612
rect 5906 3360 5962 3369
rect 5906 3295 5962 3304
rect 5722 3088 5778 3097
rect 5920 3058 5948 3295
rect 5722 3023 5778 3032
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 5630 2952 5686 2961
rect 5630 2887 5686 2896
rect 5552 2746 5672 2774
rect 5448 1420 5500 1426
rect 5448 1362 5500 1368
rect 5644 882 5672 2746
rect 6196 2514 6224 96863
rect 6276 96824 6328 96830
rect 6276 96766 6328 96772
rect 6366 96792 6422 96801
rect 6184 2508 6236 2514
rect 6184 2450 6236 2456
rect 6196 2174 6224 2450
rect 6288 2310 6316 96766
rect 6366 96727 6422 96736
rect 6380 4078 6408 96727
rect 6472 94654 6500 96902
rect 6552 95532 6604 95538
rect 6552 95474 6604 95480
rect 6460 94648 6512 94654
rect 6460 94590 6512 94596
rect 6368 4072 6420 4078
rect 6368 4014 6420 4020
rect 6276 2304 6328 2310
rect 6276 2246 6328 2252
rect 6184 2168 6236 2174
rect 6184 2110 6236 2116
rect 6288 2038 6316 2246
rect 6276 2032 6328 2038
rect 6276 1974 6328 1980
rect 6472 1358 6500 94590
rect 6564 2961 6592 95474
rect 6748 89714 6776 97310
rect 6840 95606 6868 98058
rect 22928 97300 22980 97306
rect 22928 97242 22980 97248
rect 21916 97232 21968 97238
rect 21914 97200 21916 97209
rect 21968 97200 21970 97209
rect 21914 97135 21970 97144
rect 22650 97200 22706 97209
rect 22650 97135 22706 97144
rect 18052 97096 18104 97102
rect 14646 97064 14702 97073
rect 14646 96999 14648 97008
rect 14700 96999 14702 97008
rect 17130 97064 17186 97073
rect 17130 96999 17132 97008
rect 14648 96970 14700 96976
rect 17184 96999 17186 97008
rect 18050 97064 18052 97073
rect 18104 97064 18106 97073
rect 22664 97034 22692 97135
rect 18050 96999 18106 97008
rect 22652 97028 22704 97034
rect 17132 96970 17184 96976
rect 22652 96970 22704 96976
rect 22940 96694 22968 97242
rect 78954 97200 79010 97209
rect 78692 97158 78954 97186
rect 78692 97073 78720 97158
rect 80150 97200 80206 97209
rect 78954 97135 79010 97144
rect 80072 97158 80150 97186
rect 24306 97064 24362 97073
rect 24306 96999 24362 97008
rect 25410 97064 25466 97073
rect 25410 96999 25466 97008
rect 30102 97064 30158 97073
rect 30102 96999 30158 97008
rect 32034 97064 32090 97073
rect 32034 96999 32090 97008
rect 33138 97064 33194 97073
rect 33138 96999 33194 97008
rect 77390 97064 77446 97073
rect 77390 96999 77446 97008
rect 78678 97064 78734 97073
rect 78678 96999 78734 97008
rect 24320 96762 24348 96999
rect 24308 96756 24360 96762
rect 24308 96698 24360 96704
rect 25424 96694 25452 96999
rect 30116 96898 30144 96999
rect 30104 96892 30156 96898
rect 30104 96834 30156 96840
rect 32048 96830 32076 96999
rect 33152 96966 33180 96999
rect 33140 96960 33192 96966
rect 33140 96902 33192 96908
rect 54850 96928 54906 96937
rect 54850 96863 54906 96872
rect 60462 96928 60518 96937
rect 60462 96863 60518 96872
rect 60646 96928 60702 96937
rect 77114 96928 77170 96937
rect 60646 96863 60702 96872
rect 61764 96886 62068 96914
rect 32036 96824 32088 96830
rect 32036 96766 32088 96772
rect 22100 96688 22152 96694
rect 22100 96630 22152 96636
rect 22928 96688 22980 96694
rect 22928 96630 22980 96636
rect 25412 96688 25464 96694
rect 25412 96630 25464 96636
rect 53746 96656 53802 96665
rect 16486 96520 16542 96529
rect 16486 96455 16488 96464
rect 16540 96455 16542 96464
rect 16488 96426 16540 96432
rect 15750 96384 15806 96393
rect 15750 96319 15752 96328
rect 15804 96319 15806 96328
rect 15752 96290 15804 96296
rect 9586 96248 9642 96257
rect 9586 96183 9588 96192
rect 9640 96183 9642 96192
rect 9588 96154 9640 96160
rect 6920 96008 6972 96014
rect 6920 95950 6972 95956
rect 6828 95600 6880 95606
rect 6828 95542 6880 95548
rect 6748 89686 6868 89714
rect 6840 12434 6868 89686
rect 6748 12406 6868 12434
rect 6748 3262 6776 12406
rect 6736 3256 6788 3262
rect 6736 3198 6788 3204
rect 6550 2952 6606 2961
rect 6550 2887 6606 2896
rect 6932 2854 6960 95950
rect 9600 93906 9628 96154
rect 15764 95810 15792 96290
rect 15752 95804 15804 95810
rect 15752 95746 15804 95752
rect 16500 95606 16528 96426
rect 22112 96257 22140 96630
rect 53746 96591 53802 96600
rect 39580 96552 39632 96558
rect 39580 96494 39632 96500
rect 29184 96416 29236 96422
rect 29184 96358 29236 96364
rect 29196 96257 29224 96358
rect 37832 96280 37884 96286
rect 22098 96248 22154 96257
rect 22098 96183 22154 96192
rect 27986 96248 28042 96257
rect 27986 96183 28042 96192
rect 29182 96248 29238 96257
rect 37832 96222 37884 96228
rect 29182 96183 29238 96192
rect 28000 96150 28028 96183
rect 27988 96144 28040 96150
rect 20994 96112 21050 96121
rect 20994 96047 21050 96056
rect 26790 96112 26846 96121
rect 27988 96086 28040 96092
rect 28908 96144 28960 96150
rect 28908 96086 28960 96092
rect 26790 96047 26846 96056
rect 16488 95600 16540 95606
rect 16488 95542 16540 95548
rect 21008 95402 21036 96047
rect 24584 95804 24636 95810
rect 24584 95746 24636 95752
rect 20996 95396 21048 95402
rect 20996 95338 21048 95344
rect 24596 95305 24624 95746
rect 26804 95334 26832 96047
rect 27528 95600 27580 95606
rect 27528 95542 27580 95548
rect 27540 95334 27568 95542
rect 28920 95470 28948 96086
rect 28908 95464 28960 95470
rect 28908 95406 28960 95412
rect 26792 95328 26844 95334
rect 24582 95296 24638 95305
rect 26792 95270 26844 95276
rect 27528 95328 27580 95334
rect 27528 95270 27580 95276
rect 24582 95231 24638 95240
rect 24768 95192 24820 95198
rect 12806 95160 12862 95169
rect 12806 95095 12862 95104
rect 19338 95160 19394 95169
rect 19338 95095 19340 95104
rect 12820 94654 12848 95095
rect 19392 95095 19394 95104
rect 24766 95160 24768 95169
rect 24820 95160 24822 95169
rect 24766 95095 24822 95104
rect 25962 95160 26018 95169
rect 25962 95095 26018 95104
rect 19340 95066 19392 95072
rect 19352 94790 19380 95066
rect 25976 95062 26004 95095
rect 25964 95056 26016 95062
rect 23386 95024 23442 95033
rect 25964 94998 26016 95004
rect 29196 94994 29224 96183
rect 31482 96112 31538 96121
rect 31482 96047 31538 96056
rect 34978 96112 35034 96121
rect 34978 96047 35034 96056
rect 31496 95674 31524 96047
rect 34992 95742 35020 96047
rect 34980 95736 35032 95742
rect 34980 95678 35032 95684
rect 31484 95668 31536 95674
rect 31484 95610 31536 95616
rect 37844 95305 37872 96222
rect 39592 95985 39620 96494
rect 46846 96384 46902 96393
rect 46846 96319 46902 96328
rect 50342 96384 50398 96393
rect 50342 96319 50398 96328
rect 51170 96384 51226 96393
rect 51170 96319 51226 96328
rect 41144 96280 41196 96286
rect 41144 96222 41196 96228
rect 41970 96248 42026 96257
rect 39578 95976 39634 95985
rect 39578 95911 39634 95920
rect 38474 95840 38530 95849
rect 38474 95775 38530 95784
rect 38488 95538 38516 95775
rect 38476 95532 38528 95538
rect 38476 95474 38528 95480
rect 41156 95305 41184 96222
rect 41970 96183 42026 96192
rect 44178 96248 44234 96257
rect 44178 96183 44234 96192
rect 41984 96014 42012 96183
rect 41972 96008 42024 96014
rect 41972 95950 42024 95956
rect 37830 95296 37886 95305
rect 37830 95231 37886 95240
rect 41142 95296 41198 95305
rect 41142 95231 41198 95240
rect 38566 95160 38622 95169
rect 38566 95095 38622 95104
rect 44086 95160 44142 95169
rect 44086 95095 44142 95104
rect 30286 95024 30342 95033
rect 23386 94959 23442 94968
rect 29184 94988 29236 94994
rect 20626 94888 20682 94897
rect 20626 94823 20628 94832
rect 20680 94823 20682 94832
rect 20628 94794 20680 94800
rect 19340 94784 19392 94790
rect 19340 94726 19392 94732
rect 23400 94654 23428 94959
rect 30286 94959 30288 94968
rect 29184 94930 29236 94936
rect 30340 94959 30342 94968
rect 31666 95024 31722 95033
rect 31666 94959 31722 94968
rect 30288 94930 30340 94936
rect 31680 94926 31708 94959
rect 31668 94920 31720 94926
rect 31668 94862 31720 94868
rect 38580 94722 38608 95095
rect 38568 94716 38620 94722
rect 38568 94658 38620 94664
rect 12808 94648 12860 94654
rect 12808 94590 12860 94596
rect 13728 94648 13780 94654
rect 13728 94590 13780 94596
rect 23388 94648 23440 94654
rect 23388 94590 23440 94596
rect 37278 94616 37334 94625
rect 13740 93974 13768 94590
rect 37278 94551 37280 94560
rect 37332 94551 37334 94560
rect 37280 94522 37332 94528
rect 42706 94480 42762 94489
rect 42706 94415 42762 94424
rect 42720 94178 42748 94415
rect 44100 94246 44128 95095
rect 44192 94858 44220 96183
rect 45374 95296 45430 95305
rect 45374 95231 45376 95240
rect 45428 95231 45430 95240
rect 45376 95202 45428 95208
rect 45190 95160 45246 95169
rect 45190 95095 45246 95104
rect 45558 95160 45614 95169
rect 45558 95095 45614 95104
rect 46662 95160 46718 95169
rect 46662 95095 46718 95104
rect 45204 94858 45232 95095
rect 44180 94852 44232 94858
rect 44180 94794 44232 94800
rect 45192 94852 45244 94858
rect 45192 94794 45244 94800
rect 45572 94790 45600 95095
rect 45560 94784 45612 94790
rect 45560 94726 45612 94732
rect 46676 94586 46704 95095
rect 46860 94722 46888 96319
rect 50356 96218 50384 96319
rect 51184 96218 51212 96319
rect 50344 96212 50396 96218
rect 50344 96154 50396 96160
rect 51172 96212 51224 96218
rect 51172 96154 51224 96160
rect 52184 95872 52236 95878
rect 52184 95814 52236 95820
rect 47950 95296 48006 95305
rect 47950 95231 48006 95240
rect 48226 95296 48282 95305
rect 48226 95231 48282 95240
rect 49516 95260 49568 95266
rect 47964 94722 47992 95231
rect 48134 95160 48190 95169
rect 48134 95095 48190 95104
rect 46848 94716 46900 94722
rect 46848 94658 46900 94664
rect 47952 94716 48004 94722
rect 47952 94658 48004 94664
rect 46664 94580 46716 94586
rect 46664 94522 46716 94528
rect 45098 94480 45154 94489
rect 45098 94415 45154 94424
rect 45112 94314 45140 94415
rect 45100 94308 45152 94314
rect 45100 94250 45152 94256
rect 44088 94240 44140 94246
rect 44088 94182 44140 94188
rect 48148 94178 48176 95095
rect 48240 94654 48268 95231
rect 49516 95202 49568 95208
rect 49608 95260 49660 95266
rect 49608 95202 49660 95208
rect 48228 94648 48280 94654
rect 48228 94590 48280 94596
rect 42708 94172 42760 94178
rect 42708 94114 42760 94120
rect 48136 94172 48188 94178
rect 48136 94114 48188 94120
rect 49056 94036 49108 94042
rect 49056 93978 49108 93984
rect 13728 93968 13780 93974
rect 13728 93910 13780 93916
rect 9588 93900 9640 93906
rect 9588 93842 9640 93848
rect 49068 93673 49096 93978
rect 49528 93770 49556 95202
rect 49516 93764 49568 93770
rect 49516 93706 49568 93712
rect 49620 93673 49648 95202
rect 50802 95160 50858 95169
rect 50802 95095 50858 95104
rect 50816 94654 50844 95095
rect 49884 94648 49936 94654
rect 49884 94590 49936 94596
rect 50804 94648 50856 94654
rect 50804 94590 50856 94596
rect 49896 94489 49924 94590
rect 49882 94480 49938 94489
rect 50158 94480 50214 94489
rect 49882 94415 49938 94424
rect 49976 94444 50028 94450
rect 50158 94415 50214 94424
rect 49976 94386 50028 94392
rect 49988 93673 50016 94386
rect 50172 94217 50200 94415
rect 51448 94376 51500 94382
rect 51448 94318 51500 94324
rect 50158 94208 50214 94217
rect 50158 94143 50214 94152
rect 50988 94172 51040 94178
rect 50988 94114 51040 94120
rect 51000 94081 51028 94114
rect 50986 94072 51042 94081
rect 50986 94007 51042 94016
rect 50620 93832 50672 93838
rect 50620 93774 50672 93780
rect 50632 93673 50660 93774
rect 51460 93673 51488 94318
rect 52196 93673 52224 95814
rect 52552 94648 52604 94654
rect 52552 94590 52604 94596
rect 52564 93673 52592 94590
rect 53760 94314 53788 96591
rect 54576 96008 54628 96014
rect 54576 95950 54628 95956
rect 53748 94308 53800 94314
rect 53748 94250 53800 94256
rect 54024 94308 54076 94314
rect 54024 94250 54076 94256
rect 53288 94172 53340 94178
rect 53288 94114 53340 94120
rect 53300 93673 53328 94114
rect 54036 93673 54064 94250
rect 54588 93673 54616 95950
rect 54864 94246 54892 96863
rect 60476 96665 60504 96863
rect 57610 96656 57666 96665
rect 57610 96591 57666 96600
rect 57886 96656 57942 96665
rect 57886 96591 57942 96600
rect 58070 96656 58126 96665
rect 58070 96591 58126 96600
rect 59542 96656 59598 96665
rect 59542 96591 59598 96600
rect 59726 96656 59782 96665
rect 59726 96591 59782 96600
rect 59910 96656 59966 96665
rect 59910 96591 59966 96600
rect 60462 96656 60518 96665
rect 60462 96591 60518 96600
rect 57624 96218 57652 96591
rect 57612 96212 57664 96218
rect 57612 96154 57664 96160
rect 57900 96082 57928 96591
rect 57888 96076 57940 96082
rect 57888 96018 57940 96024
rect 58084 95538 58112 96591
rect 59360 96280 59412 96286
rect 59360 96222 59412 96228
rect 58072 95532 58124 95538
rect 58072 95474 58124 95480
rect 54852 94240 54904 94246
rect 54852 94182 54904 94188
rect 54944 94240 54996 94246
rect 54944 94182 54996 94188
rect 54956 93673 54984 94182
rect 40866 93664 40922 93673
rect 40866 93599 40922 93608
rect 42614 93664 42670 93673
rect 42614 93599 42670 93608
rect 44086 93664 44142 93673
rect 44086 93599 44142 93608
rect 46662 93664 46718 93673
rect 46662 93599 46718 93608
rect 47950 93664 48006 93673
rect 47950 93599 48006 93608
rect 48778 93664 48834 93673
rect 48778 93599 48780 93608
rect 40880 93401 40908 93599
rect 40866 93392 40922 93401
rect 40866 93327 40922 93336
rect 40590 93256 40646 93265
rect 40590 93191 40646 93200
rect 39948 93084 40000 93090
rect 39948 93026 40000 93032
rect 38384 93016 38436 93022
rect 38384 92958 38436 92964
rect 35256 92948 35308 92954
rect 35256 92890 35308 92896
rect 35268 92857 35296 92890
rect 36728 92880 36780 92886
rect 32862 92848 32918 92857
rect 32862 92783 32864 92792
rect 32916 92783 32918 92792
rect 34150 92848 34206 92857
rect 34150 92783 34152 92792
rect 32864 92754 32916 92760
rect 34204 92783 34206 92792
rect 35254 92848 35310 92857
rect 35254 92783 35310 92792
rect 36726 92848 36728 92857
rect 38396 92857 38424 92958
rect 39960 92857 39988 93026
rect 40604 92857 40632 93191
rect 42628 93158 42656 93599
rect 44100 93226 44128 93599
rect 46676 93294 46704 93599
rect 47964 93362 47992 93599
rect 48832 93599 48834 93608
rect 49054 93664 49110 93673
rect 49054 93599 49110 93608
rect 49606 93664 49662 93673
rect 49606 93599 49662 93608
rect 49974 93664 50030 93673
rect 49974 93599 50030 93608
rect 50618 93664 50674 93673
rect 50618 93599 50674 93608
rect 51262 93664 51318 93673
rect 51262 93599 51318 93608
rect 51446 93664 51502 93673
rect 51446 93599 51502 93608
rect 52182 93664 52238 93673
rect 52182 93599 52238 93608
rect 52550 93664 52606 93673
rect 52550 93599 52606 93608
rect 53286 93664 53342 93673
rect 53286 93599 53342 93608
rect 53746 93664 53802 93673
rect 53746 93599 53802 93608
rect 54022 93664 54078 93673
rect 54022 93599 54078 93608
rect 54206 93664 54262 93673
rect 54206 93599 54208 93608
rect 48780 93570 48832 93576
rect 51276 93498 51304 93599
rect 51264 93492 51316 93498
rect 51264 93434 51316 93440
rect 53760 93430 53788 93599
rect 54260 93599 54262 93608
rect 54574 93664 54630 93673
rect 54574 93599 54630 93608
rect 54942 93664 54998 93673
rect 54942 93599 54998 93608
rect 54208 93570 54260 93576
rect 59372 93566 59400 96222
rect 59556 96218 59584 96591
rect 59544 96212 59596 96218
rect 59544 96154 59596 96160
rect 59740 96150 59768 96591
rect 59728 96144 59780 96150
rect 59728 96086 59780 96092
rect 59924 94178 59952 96591
rect 60660 96286 60688 96863
rect 61764 96801 61792 96886
rect 61566 96792 61622 96801
rect 61566 96727 61622 96736
rect 61750 96792 61806 96801
rect 61750 96727 61806 96736
rect 61934 96792 61990 96801
rect 62040 96778 62068 96886
rect 77114 96863 77170 96872
rect 62040 96750 62160 96778
rect 61934 96727 61990 96736
rect 61580 96286 61608 96727
rect 60648 96280 60700 96286
rect 60648 96222 60700 96228
rect 61568 96280 61620 96286
rect 61568 96222 61620 96228
rect 59912 94172 59964 94178
rect 59912 94114 59964 94120
rect 61948 94110 61976 96727
rect 62132 95810 62160 96750
rect 76932 96756 76984 96762
rect 76932 96698 76984 96704
rect 76944 96665 76972 96698
rect 77128 96665 77156 96863
rect 76930 96656 76986 96665
rect 76930 96591 76986 96600
rect 77114 96656 77170 96665
rect 77114 96591 77170 96600
rect 62304 96552 62356 96558
rect 77404 96506 77432 96999
rect 79506 96792 79562 96801
rect 79244 96750 79506 96778
rect 79244 96665 79272 96750
rect 80072 96762 80100 97158
rect 80150 97135 80206 97144
rect 79506 96727 79562 96736
rect 80060 96756 80112 96762
rect 80060 96698 80112 96704
rect 79230 96656 79286 96665
rect 79230 96591 79286 96600
rect 82174 96656 82230 96665
rect 82174 96591 82230 96600
rect 62304 96494 62356 96500
rect 62028 95804 62080 95810
rect 62028 95746 62080 95752
rect 62120 95804 62172 95810
rect 62120 95746 62172 95752
rect 62040 94178 62068 95746
rect 62028 94172 62080 94178
rect 62028 94114 62080 94120
rect 62316 94110 62344 96494
rect 76668 96490 77432 96506
rect 82188 96490 82216 96591
rect 76656 96484 77432 96490
rect 76708 96478 77432 96484
rect 82176 96484 82228 96490
rect 76656 96426 76708 96432
rect 82176 96426 82228 96432
rect 80150 96384 80206 96393
rect 80206 96342 80468 96370
rect 80150 96319 80206 96328
rect 75184 96212 75236 96218
rect 75184 96154 75236 96160
rect 74632 96144 74684 96150
rect 74632 96086 74684 96092
rect 74644 95985 74672 96086
rect 74630 95976 74686 95985
rect 74630 95911 74686 95920
rect 74814 95976 74870 95985
rect 74814 95911 74870 95920
rect 74828 95713 74856 95911
rect 74814 95704 74870 95713
rect 74814 95639 74870 95648
rect 75196 95577 75224 96154
rect 80152 96144 80204 96150
rect 79506 96112 79562 96121
rect 79506 96047 79562 96056
rect 79690 96112 79746 96121
rect 80152 96086 80204 96092
rect 79690 96047 79746 96056
rect 76840 96008 76892 96014
rect 76838 95976 76840 95985
rect 76892 95976 76894 95985
rect 76838 95911 76894 95920
rect 77022 95976 77078 95985
rect 77022 95911 77078 95920
rect 75182 95568 75238 95577
rect 75182 95503 75238 95512
rect 76102 95568 76158 95577
rect 76102 95503 76158 95512
rect 64144 95328 64196 95334
rect 63958 95296 64014 95305
rect 63958 95231 64014 95240
rect 64142 95296 64144 95305
rect 64196 95296 64198 95305
rect 64326 95296 64382 95305
rect 64142 95231 64198 95240
rect 64248 95254 64326 95282
rect 63972 95146 64000 95231
rect 64248 95146 64276 95254
rect 64326 95231 64382 95240
rect 64788 95260 64840 95266
rect 64788 95202 64840 95208
rect 63972 95118 64276 95146
rect 61936 94104 61988 94110
rect 61936 94046 61988 94052
rect 62304 94104 62356 94110
rect 62304 94046 62356 94052
rect 64800 93634 64828 95202
rect 74540 94920 74592 94926
rect 74540 94862 74592 94868
rect 74552 94738 74580 94862
rect 76116 94790 76144 95503
rect 76104 94784 76156 94790
rect 74552 94710 74672 94738
rect 76104 94726 76156 94732
rect 74644 94586 74672 94710
rect 74540 94580 74592 94586
rect 74540 94522 74592 94528
rect 74632 94580 74684 94586
rect 74632 94522 74684 94528
rect 74552 94466 74580 94522
rect 74552 94450 74856 94466
rect 74552 94444 74868 94450
rect 74552 94438 74816 94444
rect 74816 94386 74868 94392
rect 77036 93673 77064 95911
rect 79520 95441 79548 96047
rect 79704 96014 79732 96047
rect 79692 96008 79744 96014
rect 79692 95950 79744 95956
rect 79784 96008 79836 96014
rect 79784 95950 79836 95956
rect 79506 95432 79562 95441
rect 79506 95367 79562 95376
rect 79796 95146 79824 95950
rect 80164 95860 80192 96086
rect 80336 96008 80388 96014
rect 80242 95976 80298 95985
rect 80298 95956 80336 95962
rect 80440 95985 80468 96342
rect 80518 96248 80574 96257
rect 80518 96183 80574 96192
rect 82188 96206 82400 96234
rect 80298 95950 80388 95956
rect 80426 95976 80482 95985
rect 80298 95934 80376 95950
rect 80242 95911 80298 95920
rect 80426 95911 80482 95920
rect 80532 95860 80560 96183
rect 80164 95832 80560 95860
rect 80152 95464 80204 95470
rect 79888 95424 80152 95452
rect 79888 95266 79916 95424
rect 80152 95406 80204 95412
rect 79876 95260 79928 95266
rect 79876 95202 79928 95208
rect 79428 95118 79824 95146
rect 80152 95192 80204 95198
rect 80204 95152 80652 95180
rect 80152 95134 80204 95140
rect 79428 94874 79456 95118
rect 79506 95024 79562 95033
rect 79506 94959 79562 94968
rect 80058 95024 80114 95033
rect 80518 95024 80574 95033
rect 80114 94994 80192 95010
rect 80114 94988 80204 94994
rect 80114 94982 80152 94988
rect 80058 94959 80114 94968
rect 78232 94858 79456 94874
rect 78220 94852 79456 94858
rect 78272 94846 79456 94852
rect 78220 94794 78272 94800
rect 79232 94172 79284 94178
rect 79232 94114 79284 94120
rect 79244 94081 79272 94114
rect 79230 94072 79286 94081
rect 79230 94007 79286 94016
rect 79520 93945 79548 94959
rect 80152 94930 80204 94936
rect 80428 94988 80480 94994
rect 80518 94959 80574 94968
rect 80428 94930 80480 94936
rect 80244 94920 80296 94926
rect 80244 94862 80296 94868
rect 80256 94722 80284 94862
rect 80244 94716 80296 94722
rect 80244 94658 80296 94664
rect 80440 94586 80468 94930
rect 80532 94722 80560 94959
rect 80624 94790 80652 95152
rect 81438 95024 81494 95033
rect 81438 94959 81494 94968
rect 80612 94784 80664 94790
rect 80612 94726 80664 94732
rect 80520 94716 80572 94722
rect 80520 94658 80572 94664
rect 80428 94580 80480 94586
rect 80428 94522 80480 94528
rect 81452 94178 81480 94959
rect 82188 94625 82216 96206
rect 82372 96150 82400 96206
rect 82360 96144 82412 96150
rect 82360 96086 82412 96092
rect 82464 95713 82492 162862
rect 82542 154048 82598 154057
rect 82542 153983 82598 153992
rect 82556 132297 82584 153983
rect 82542 132288 82598 132297
rect 82542 132223 82598 132232
rect 83372 127016 83424 127022
rect 83372 126958 83424 126964
rect 83280 125860 83332 125866
rect 83280 125802 83332 125808
rect 83188 122868 83240 122874
rect 83188 122810 83240 122816
rect 83096 121508 83148 121514
rect 83096 121450 83148 121456
rect 83004 120148 83056 120154
rect 83004 120090 83056 120096
rect 82912 118720 82964 118726
rect 82912 118662 82964 118668
rect 82634 114336 82690 114345
rect 82634 114271 82690 114280
rect 82544 110356 82596 110362
rect 82544 110298 82596 110304
rect 82450 95704 82506 95713
rect 82450 95639 82506 95648
rect 82556 95062 82584 110298
rect 82648 96801 82676 114271
rect 82728 99340 82780 99346
rect 82728 99282 82780 99288
rect 82740 98326 82768 99282
rect 82728 98320 82780 98326
rect 82728 98262 82780 98268
rect 82728 98184 82780 98190
rect 82728 98126 82780 98132
rect 82634 96792 82690 96801
rect 82634 96727 82690 96736
rect 82740 96354 82768 98126
rect 82818 97608 82874 97617
rect 82818 97543 82874 97552
rect 82832 96490 82860 97543
rect 82924 96898 82952 118662
rect 82912 96892 82964 96898
rect 82912 96834 82964 96840
rect 82910 96792 82966 96801
rect 82910 96727 82966 96736
rect 82820 96484 82872 96490
rect 82820 96426 82872 96432
rect 82728 96348 82780 96354
rect 82728 96290 82780 96296
rect 82728 95872 82780 95878
rect 82728 95814 82780 95820
rect 82544 95056 82596 95062
rect 82544 94998 82596 95004
rect 82360 94784 82412 94790
rect 82360 94726 82412 94732
rect 82372 94625 82400 94726
rect 82174 94616 82230 94625
rect 82174 94551 82230 94560
rect 82358 94616 82414 94625
rect 82358 94551 82414 94560
rect 81440 94172 81492 94178
rect 81440 94114 81492 94120
rect 79506 93936 79562 93945
rect 79506 93871 79562 93880
rect 82634 93800 82690 93809
rect 82096 93758 82634 93786
rect 79416 93696 79468 93702
rect 77022 93664 77078 93673
rect 64788 93628 64840 93634
rect 77022 93599 77078 93608
rect 77298 93664 77354 93673
rect 77298 93599 77354 93608
rect 79046 93664 79102 93673
rect 79102 93644 79416 93650
rect 79102 93638 79468 93644
rect 79102 93622 79456 93638
rect 79046 93599 79102 93608
rect 64788 93570 64840 93576
rect 59360 93560 59412 93566
rect 59360 93502 59412 93508
rect 77312 93430 77340 93599
rect 53748 93424 53800 93430
rect 53748 93366 53800 93372
rect 77300 93424 77352 93430
rect 77300 93366 77352 93372
rect 79506 93392 79562 93401
rect 47952 93356 48004 93362
rect 79506 93327 79562 93336
rect 47952 93298 48004 93304
rect 79520 93294 79548 93327
rect 46664 93288 46716 93294
rect 46664 93230 46716 93236
rect 77484 93288 77536 93294
rect 77484 93230 77536 93236
rect 79508 93288 79560 93294
rect 79508 93230 79560 93236
rect 44088 93220 44140 93226
rect 44088 93162 44140 93168
rect 42616 93152 42668 93158
rect 77496 93129 77524 93230
rect 42616 93094 42668 93100
rect 77482 93120 77538 93129
rect 77482 93055 77538 93064
rect 77666 93120 77722 93129
rect 77666 93055 77722 93064
rect 77680 92857 77708 93055
rect 82096 92857 82124 93758
rect 82634 93735 82690 93744
rect 82452 93356 82504 93362
rect 82452 93298 82504 93304
rect 36780 92848 36782 92857
rect 36726 92783 36782 92792
rect 38382 92848 38438 92857
rect 38382 92783 38438 92792
rect 39946 92848 40002 92857
rect 39946 92783 40002 92792
rect 40590 92848 40646 92857
rect 40590 92783 40646 92792
rect 77666 92848 77722 92857
rect 77666 92783 77722 92792
rect 82082 92848 82138 92857
rect 82082 92783 82138 92792
rect 34152 92754 34204 92760
rect 82464 74458 82492 93298
rect 82740 93106 82768 95814
rect 82924 95033 82952 96727
rect 83016 95674 83044 120090
rect 83108 96830 83136 121450
rect 83200 96966 83228 122810
rect 83292 97073 83320 125802
rect 83278 97064 83334 97073
rect 83278 96999 83334 97008
rect 83188 96960 83240 96966
rect 83188 96902 83240 96908
rect 83096 96824 83148 96830
rect 83096 96766 83148 96772
rect 83280 96824 83332 96830
rect 83280 96766 83332 96772
rect 83004 95668 83056 95674
rect 83004 95610 83056 95616
rect 83188 95600 83240 95606
rect 83188 95542 83240 95548
rect 83292 95554 83320 96766
rect 83384 95849 83412 126958
rect 83464 98116 83516 98122
rect 83464 98058 83516 98064
rect 83476 97374 83504 98058
rect 83464 97368 83516 97374
rect 83464 97310 83516 97316
rect 83464 96960 83516 96966
rect 83464 96902 83516 96908
rect 83476 95996 83504 96902
rect 83568 96121 83596 167078
rect 83648 107364 83700 107370
rect 83648 107306 83700 107312
rect 83660 97102 83688 107306
rect 83648 97096 83700 97102
rect 83648 97038 83700 97044
rect 83648 96892 83700 96898
rect 83648 96834 83700 96840
rect 83554 96112 83610 96121
rect 83554 96047 83610 96056
rect 83476 95968 83596 95996
rect 83370 95840 83426 95849
rect 83370 95775 83426 95784
rect 83004 95396 83056 95402
rect 83004 95338 83056 95344
rect 82910 95024 82966 95033
rect 82910 94959 82966 94968
rect 82820 94920 82872 94926
rect 82820 94862 82872 94868
rect 82832 93362 82860 94862
rect 82912 93696 82964 93702
rect 82912 93638 82964 93644
rect 82820 93356 82872 93362
rect 82820 93298 82872 93304
rect 82740 93078 82860 93106
rect 82726 92984 82782 92993
rect 82726 92919 82782 92928
rect 82452 74452 82504 74458
rect 82452 74394 82504 74400
rect 82450 55312 82506 55321
rect 82450 55247 82506 55256
rect 82464 45529 82492 55247
rect 82740 49706 82768 92919
rect 82832 92274 82860 93078
rect 82820 92268 82872 92274
rect 82820 92210 82872 92216
rect 82820 92132 82872 92138
rect 82820 92074 82872 92080
rect 82728 49700 82780 49706
rect 82728 49642 82780 49648
rect 82450 45520 82506 45529
rect 82450 45455 82506 45464
rect 82450 16688 82506 16697
rect 82450 16623 82506 16632
rect 15292 3256 15344 3262
rect 15292 3198 15344 3204
rect 25044 3256 25096 3262
rect 52552 3256 52604 3262
rect 25044 3198 25096 3204
rect 47766 3224 47822 3233
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 13924 2854 13952 2994
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 8116 2848 8168 2854
rect 8116 2790 8168 2796
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 8128 2689 8156 2790
rect 8114 2680 8170 2689
rect 8114 2615 8170 2624
rect 9772 2372 9824 2378
rect 9772 2314 9824 2320
rect 9784 2281 9812 2314
rect 13924 2281 13952 2790
rect 15304 2689 15332 3198
rect 22100 3188 22152 3194
rect 22100 3130 22152 3136
rect 16304 3120 16356 3126
rect 16304 3062 16356 3068
rect 15290 2680 15346 2689
rect 15290 2615 15346 2624
rect 16316 2281 16344 3062
rect 20720 2984 20772 2990
rect 20720 2926 20772 2932
rect 20732 2689 20760 2926
rect 20718 2680 20774 2689
rect 20718 2615 20774 2624
rect 22112 2281 22140 3130
rect 24124 2916 24176 2922
rect 24124 2858 24176 2864
rect 22650 2544 22706 2553
rect 22650 2479 22652 2488
rect 22704 2479 22706 2488
rect 22652 2450 22704 2456
rect 24136 2281 24164 2858
rect 25056 2689 25084 3198
rect 47766 3159 47822 3168
rect 48686 3224 48742 3233
rect 52552 3198 52604 3204
rect 48686 3159 48742 3168
rect 49976 3188 50028 3194
rect 47780 2922 47808 3159
rect 48700 2961 48728 3159
rect 49976 3130 50028 3136
rect 49988 2961 50016 3130
rect 48686 2952 48742 2961
rect 47768 2916 47820 2922
rect 48686 2887 48742 2896
rect 49974 2952 50030 2961
rect 49974 2887 50030 2896
rect 47768 2858 47820 2864
rect 25042 2680 25098 2689
rect 25042 2615 25098 2624
rect 50344 2576 50396 2582
rect 50344 2518 50396 2524
rect 45928 2508 45980 2514
rect 45928 2450 45980 2456
rect 41420 2440 41472 2446
rect 41420 2382 41472 2388
rect 9770 2272 9826 2281
rect 9770 2207 9826 2216
rect 13910 2272 13966 2281
rect 13910 2207 13966 2216
rect 16302 2272 16358 2281
rect 16302 2207 16358 2216
rect 22098 2272 22154 2281
rect 22098 2207 22154 2216
rect 24122 2272 24178 2281
rect 24122 2207 24178 2216
rect 32678 2272 32734 2281
rect 32678 2207 32734 2216
rect 36174 2272 36230 2281
rect 36174 2207 36230 2216
rect 37462 2272 37518 2281
rect 37462 2207 37464 2216
rect 9784 1465 9812 2207
rect 32692 2038 32720 2207
rect 36188 2174 36216 2207
rect 37516 2207 37518 2216
rect 37464 2178 37516 2184
rect 36176 2168 36228 2174
rect 32770 2136 32826 2145
rect 32770 2071 32826 2080
rect 33966 2136 34022 2145
rect 36268 2168 36320 2174
rect 36176 2110 36228 2116
rect 36266 2136 36268 2145
rect 36320 2136 36322 2145
rect 33966 2071 33968 2080
rect 32784 2038 32812 2071
rect 34020 2071 34022 2080
rect 36266 2071 36322 2080
rect 33968 2042 34020 2048
rect 32680 2032 32732 2038
rect 29090 2000 29146 2009
rect 29090 1935 29092 1944
rect 29144 1935 29146 1944
rect 30470 2000 30526 2009
rect 30470 1935 30472 1944
rect 29092 1906 29144 1912
rect 30524 1935 30526 1944
rect 31666 2000 31722 2009
rect 32680 1974 32732 1980
rect 32772 2032 32824 2038
rect 32772 1974 32824 1980
rect 31666 1935 31722 1944
rect 30472 1906 30524 1912
rect 31680 1902 31708 1935
rect 31668 1896 31720 1902
rect 17498 1864 17554 1873
rect 17498 1799 17554 1808
rect 21086 1864 21142 1873
rect 21086 1799 21142 1808
rect 22282 1864 22338 1873
rect 22282 1799 22338 1808
rect 25778 1864 25834 1873
rect 25778 1799 25780 1808
rect 9770 1456 9826 1465
rect 17512 1426 17540 1799
rect 21100 1630 21128 1799
rect 21088 1624 21140 1630
rect 21088 1566 21140 1572
rect 22296 1562 22324 1799
rect 25832 1799 25834 1808
rect 26974 1864 27030 1873
rect 26974 1799 27030 1808
rect 28170 1864 28226 1873
rect 31668 1838 31720 1844
rect 28170 1799 28226 1808
rect 25780 1770 25832 1776
rect 26988 1698 27016 1799
rect 28184 1766 28212 1799
rect 28172 1760 28224 1766
rect 28172 1702 28224 1708
rect 26976 1692 27028 1698
rect 26976 1634 27028 1640
rect 22284 1556 22336 1562
rect 22284 1498 22336 1504
rect 19248 1488 19300 1494
rect 19248 1430 19300 1436
rect 9770 1391 9826 1400
rect 17500 1420 17552 1426
rect 17500 1362 17552 1368
rect 6460 1352 6512 1358
rect 12440 1352 12492 1358
rect 6460 1294 6512 1300
rect 12438 1320 12440 1329
rect 19260 1329 19288 1430
rect 35532 1352 35584 1358
rect 12492 1320 12494 1329
rect 12438 1255 12494 1264
rect 19246 1320 19302 1329
rect 30286 1320 30342 1329
rect 19246 1255 19302 1264
rect 29000 1284 29052 1290
rect 30286 1255 30342 1264
rect 35530 1320 35532 1329
rect 35584 1320 35586 1329
rect 35530 1255 35586 1264
rect 39854 1320 39910 1329
rect 39854 1255 39910 1264
rect 29000 1226 29052 1232
rect 29012 1193 29040 1226
rect 30300 1222 30328 1255
rect 30288 1216 30340 1222
rect 17958 1184 18014 1193
rect 17958 1119 18014 1128
rect 19338 1184 19394 1193
rect 19338 1119 19394 1128
rect 28998 1184 29054 1193
rect 30288 1158 30340 1164
rect 34518 1184 34574 1193
rect 28998 1119 29054 1128
rect 34518 1119 34574 1128
rect 17972 882 18000 1119
rect 19352 950 19380 1119
rect 34532 1086 34560 1119
rect 39868 1086 39896 1255
rect 39946 1184 40002 1193
rect 39946 1119 39948 1128
rect 40000 1119 40002 1128
rect 39948 1090 40000 1096
rect 34520 1080 34572 1086
rect 24766 1048 24822 1057
rect 24766 983 24822 992
rect 30378 1048 30434 1057
rect 34520 1022 34572 1028
rect 39856 1080 39908 1086
rect 39856 1022 39908 1028
rect 41326 1048 41382 1057
rect 30378 983 30380 992
rect 24780 950 24808 983
rect 30432 983 30434 992
rect 41326 983 41328 992
rect 30380 954 30432 960
rect 41380 983 41382 992
rect 41328 954 41380 960
rect 41432 950 41460 2382
rect 45940 1358 45968 2450
rect 45928 1352 45980 1358
rect 44914 1320 44970 1329
rect 48228 1352 48280 1358
rect 45928 1294 45980 1300
rect 48226 1320 48228 1329
rect 48280 1320 48282 1329
rect 44914 1255 44916 1264
rect 44968 1255 44970 1264
rect 50356 1290 50384 2518
rect 51356 2304 51408 2310
rect 51354 2272 51356 2281
rect 52564 2281 52592 3198
rect 53472 3052 53524 3058
rect 53472 2994 53524 3000
rect 53484 2961 53512 2994
rect 53470 2952 53526 2961
rect 82464 2922 82492 16623
rect 82832 4146 82860 92074
rect 82924 84590 82952 93638
rect 83016 86358 83044 95338
rect 83096 95260 83148 95266
rect 83096 95202 83148 95208
rect 83004 86352 83056 86358
rect 83004 86294 83056 86300
rect 82912 84584 82964 84590
rect 82912 84526 82964 84532
rect 83108 84182 83136 95202
rect 83096 84176 83148 84182
rect 83096 84118 83148 84124
rect 83200 82006 83228 95542
rect 83292 95526 83504 95554
rect 83280 95328 83332 95334
rect 83280 95270 83332 95276
rect 83188 82000 83240 82006
rect 83188 81942 83240 81948
rect 83292 80918 83320 95270
rect 83372 95192 83424 95198
rect 83372 95134 83424 95140
rect 83384 94314 83412 95134
rect 83476 94874 83504 95526
rect 83568 95198 83596 95968
rect 83556 95192 83608 95198
rect 83556 95134 83608 95140
rect 83660 94926 83688 96834
rect 83752 95169 83780 180814
rect 83924 173936 83976 173942
rect 83924 173878 83976 173884
rect 83832 164416 83884 164422
rect 83832 164358 83884 164364
rect 83844 95554 83872 164358
rect 83936 95690 83964 173878
rect 84106 169960 84162 169969
rect 84106 169895 84162 169904
rect 84016 168428 84068 168434
rect 84016 168370 84068 168376
rect 84028 161474 84056 168370
rect 84120 164121 84148 169895
rect 84106 164112 84162 164121
rect 84106 164047 84162 164056
rect 84028 161446 84148 161474
rect 84016 128512 84068 128518
rect 84016 128454 84068 128460
rect 84028 96257 84056 128454
rect 84014 96248 84070 96257
rect 84014 96183 84070 96192
rect 83936 95662 84056 95690
rect 83844 95526 83964 95554
rect 83832 95464 83884 95470
rect 83832 95406 83884 95412
rect 83738 95160 83794 95169
rect 83738 95095 83794 95104
rect 83648 94920 83700 94926
rect 83476 94846 83596 94874
rect 83648 94862 83700 94868
rect 83568 94738 83596 94846
rect 83568 94722 83688 94738
rect 83556 94716 83688 94722
rect 83608 94710 83688 94716
rect 83556 94658 83608 94664
rect 83568 94627 83596 94658
rect 83372 94308 83424 94314
rect 83372 94250 83424 94256
rect 83464 94308 83516 94314
rect 83464 94250 83516 94256
rect 83280 80912 83332 80918
rect 83280 80854 83332 80860
rect 83384 80054 83412 94250
rect 83476 94178 83504 94250
rect 83464 94172 83516 94178
rect 83464 94114 83516 94120
rect 83476 93922 83504 94114
rect 83476 93894 83596 93922
rect 83464 93628 83516 93634
rect 83464 93570 83516 93576
rect 82924 80026 83412 80054
rect 82924 16574 82952 80026
rect 83372 23588 83424 23594
rect 83372 23530 83424 23536
rect 83280 20800 83332 20806
rect 83280 20742 83332 20748
rect 82924 16546 83044 16574
rect 82912 11076 82964 11082
rect 82912 11018 82964 11024
rect 82820 4140 82872 4146
rect 82820 4082 82872 4088
rect 82728 4072 82780 4078
rect 82728 4014 82780 4020
rect 82636 4004 82688 4010
rect 82636 3946 82688 3952
rect 82544 3460 82596 3466
rect 82544 3402 82596 3408
rect 53470 2887 53526 2896
rect 82452 2916 82504 2922
rect 82452 2858 82504 2864
rect 81440 2848 81492 2854
rect 81440 2790 81492 2796
rect 81348 2712 81400 2718
rect 81348 2654 81400 2660
rect 53840 2644 53892 2650
rect 53840 2586 53892 2592
rect 51408 2272 51410 2281
rect 51354 2207 51410 2216
rect 52550 2272 52606 2281
rect 52550 2207 52606 2216
rect 53852 1358 53880 2586
rect 53840 1352 53892 1358
rect 53840 1294 53892 1300
rect 48226 1255 48282 1264
rect 50344 1284 50396 1290
rect 44916 1226 44968 1232
rect 50344 1226 50396 1232
rect 52366 1184 52422 1193
rect 52366 1119 52422 1128
rect 42706 1048 42762 1057
rect 42706 983 42762 992
rect 46754 1048 46810 1057
rect 46754 983 46810 992
rect 49606 1048 49662 1057
rect 49606 983 49662 992
rect 42720 950 42748 983
rect 19340 944 19392 950
rect 19340 886 19392 892
rect 24768 944 24820 950
rect 41420 944 41472 950
rect 24768 886 24820 892
rect 27618 912 27674 921
rect 5632 876 5684 882
rect 5632 818 5684 824
rect 17960 876 18012 882
rect 41420 886 41472 892
rect 42708 944 42760 950
rect 42708 886 42760 892
rect 42798 912 42854 921
rect 27618 847 27674 856
rect 42798 847 42854 856
rect 44086 912 44142 921
rect 44086 847 44088 856
rect 17960 818 18012 824
rect 27632 814 27660 847
rect 5172 808 5224 814
rect 27620 808 27672 814
rect 5172 750 5224 756
rect 24766 776 24822 785
rect 27620 750 27672 756
rect 33138 776 33194 785
rect 24766 711 24822 720
rect 33138 711 33140 720
rect 5080 672 5132 678
rect 5080 614 5132 620
rect 20626 232 20682 241
rect 20626 167 20628 176
rect 20680 167 20682 176
rect 20628 138 20680 144
rect 24780 134 24808 711
rect 33192 711 33194 720
rect 33140 682 33192 688
rect 42812 678 42840 847
rect 44140 847 44142 856
rect 44088 818 44140 824
rect 46768 746 46796 983
rect 46846 912 46902 921
rect 46846 847 46902 856
rect 46860 814 46888 847
rect 46848 808 46900 814
rect 46848 750 46900 756
rect 46756 740 46808 746
rect 46756 682 46808 688
rect 49620 678 49648 983
rect 50986 776 51042 785
rect 50986 711 51042 720
rect 42800 672 42852 678
rect 42800 614 42852 620
rect 49608 672 49660 678
rect 49608 614 49660 620
rect 51000 610 51028 711
rect 50988 604 51040 610
rect 50988 546 51040 552
rect 52380 542 52408 1119
rect 54666 1048 54722 1057
rect 54666 983 54722 992
rect 52368 536 52420 542
rect 52368 478 52420 484
rect 53746 504 53802 513
rect 53746 439 53748 448
rect 53800 439 53802 448
rect 53748 410 53800 416
rect 54680 338 54708 983
rect 55034 776 55090 785
rect 55034 711 55090 720
rect 54668 332 54720 338
rect 54668 274 54720 280
rect 55048 270 55076 711
rect 55126 504 55182 513
rect 55126 439 55182 448
rect 55140 406 55168 439
rect 55128 400 55180 406
rect 55128 342 55180 348
rect 81360 270 81388 2654
rect 81452 338 81480 2790
rect 82452 2780 82504 2786
rect 82556 2774 82584 3402
rect 82504 2746 82584 2774
rect 82452 2722 82504 2728
rect 82648 610 82676 3946
rect 82636 604 82688 610
rect 82636 546 82688 552
rect 82740 542 82768 4014
rect 82832 3262 82860 4082
rect 82820 3256 82872 3262
rect 82820 3198 82872 3204
rect 82924 2825 82952 11018
rect 83016 2961 83044 16546
rect 83096 8356 83148 8362
rect 83096 8298 83148 8304
rect 83002 2952 83058 2961
rect 83002 2887 83004 2896
rect 83056 2887 83058 2896
rect 83004 2858 83056 2864
rect 83016 2827 83044 2858
rect 82910 2816 82966 2825
rect 82910 2751 82966 2760
rect 83108 1494 83136 8298
rect 83188 4412 83240 4418
rect 83188 4354 83240 4360
rect 83200 3233 83228 4354
rect 83186 3224 83242 3233
rect 83186 3159 83242 3168
rect 83200 3058 83228 3159
rect 83188 3052 83240 3058
rect 83188 2994 83240 3000
rect 83186 2816 83242 2825
rect 83186 2751 83242 2760
rect 83200 1630 83228 2751
rect 83292 1970 83320 20742
rect 83384 2038 83412 23530
rect 83476 4418 83504 93570
rect 83464 4412 83516 4418
rect 83464 4354 83516 4360
rect 83464 3732 83516 3738
rect 83464 3674 83516 3680
rect 83476 3097 83504 3674
rect 83568 3262 83596 93894
rect 83660 4350 83688 94710
rect 83740 93220 83792 93226
rect 83740 93162 83792 93168
rect 83752 63510 83780 93162
rect 83844 85270 83872 95406
rect 83936 94654 83964 95526
rect 83924 94648 83976 94654
rect 83924 94590 83976 94596
rect 84028 94489 84056 95662
rect 84120 94761 84148 161446
rect 84396 153882 84424 186215
rect 84488 167482 84516 187206
rect 85956 187164 86252 187184
rect 86012 187162 86036 187164
rect 86092 187162 86116 187164
rect 86172 187162 86196 187164
rect 86034 187110 86036 187162
rect 86098 187110 86110 187162
rect 86172 187110 86174 187162
rect 86012 187108 86036 187110
rect 86092 187108 86116 187110
rect 86172 187108 86196 187110
rect 85956 187088 86252 187108
rect 89956 187164 90252 187184
rect 90012 187162 90036 187164
rect 90092 187162 90116 187164
rect 90172 187162 90196 187164
rect 90034 187110 90036 187162
rect 90098 187110 90110 187162
rect 90172 187110 90174 187162
rect 90012 187108 90036 187110
rect 90092 187108 90116 187110
rect 90172 187108 90196 187110
rect 89956 187088 90252 187108
rect 87956 186620 88252 186640
rect 88012 186618 88036 186620
rect 88092 186618 88116 186620
rect 88172 186618 88196 186620
rect 88034 186566 88036 186618
rect 88098 186566 88110 186618
rect 88172 186566 88174 186618
rect 88012 186564 88036 186566
rect 88092 186564 88116 186566
rect 88172 186564 88196 186566
rect 87956 186544 88252 186564
rect 85956 186076 86252 186096
rect 86012 186074 86036 186076
rect 86092 186074 86116 186076
rect 86172 186074 86196 186076
rect 86034 186022 86036 186074
rect 86098 186022 86110 186074
rect 86172 186022 86174 186074
rect 86012 186020 86036 186022
rect 86092 186020 86116 186022
rect 86172 186020 86196 186022
rect 85956 186000 86252 186020
rect 89956 186076 90252 186096
rect 90012 186074 90036 186076
rect 90092 186074 90116 186076
rect 90172 186074 90196 186076
rect 90034 186022 90036 186074
rect 90098 186022 90110 186074
rect 90172 186022 90174 186074
rect 90012 186020 90036 186022
rect 90092 186020 90116 186022
rect 90172 186020 90196 186022
rect 89956 186000 90252 186020
rect 87956 185532 88252 185552
rect 88012 185530 88036 185532
rect 88092 185530 88116 185532
rect 88172 185530 88196 185532
rect 88034 185478 88036 185530
rect 88098 185478 88110 185530
rect 88172 185478 88174 185530
rect 88012 185476 88036 185478
rect 88092 185476 88116 185478
rect 88172 185476 88196 185478
rect 87956 185456 88252 185476
rect 85956 184988 86252 185008
rect 86012 184986 86036 184988
rect 86092 184986 86116 184988
rect 86172 184986 86196 184988
rect 86034 184934 86036 184986
rect 86098 184934 86110 184986
rect 86172 184934 86174 184986
rect 86012 184932 86036 184934
rect 86092 184932 86116 184934
rect 86172 184932 86196 184934
rect 85956 184912 86252 184932
rect 89956 184988 90252 185008
rect 90012 184986 90036 184988
rect 90092 184986 90116 184988
rect 90172 184986 90196 184988
rect 90034 184934 90036 184986
rect 90098 184934 90110 184986
rect 90172 184934 90174 184986
rect 90012 184932 90036 184934
rect 90092 184932 90116 184934
rect 90172 184932 90196 184934
rect 89956 184912 90252 184932
rect 87956 184444 88252 184464
rect 88012 184442 88036 184444
rect 88092 184442 88116 184444
rect 88172 184442 88196 184444
rect 88034 184390 88036 184442
rect 88098 184390 88110 184442
rect 88172 184390 88174 184442
rect 88012 184388 88036 184390
rect 88092 184388 88116 184390
rect 88172 184388 88196 184390
rect 87956 184368 88252 184388
rect 85956 183900 86252 183920
rect 86012 183898 86036 183900
rect 86092 183898 86116 183900
rect 86172 183898 86196 183900
rect 86034 183846 86036 183898
rect 86098 183846 86110 183898
rect 86172 183846 86174 183898
rect 86012 183844 86036 183846
rect 86092 183844 86116 183846
rect 86172 183844 86196 183846
rect 85956 183824 86252 183844
rect 89956 183900 90252 183920
rect 90012 183898 90036 183900
rect 90092 183898 90116 183900
rect 90172 183898 90196 183900
rect 90034 183846 90036 183898
rect 90098 183846 90110 183898
rect 90172 183846 90174 183898
rect 90012 183844 90036 183846
rect 90092 183844 90116 183846
rect 90172 183844 90196 183846
rect 89956 183824 90252 183844
rect 87956 183356 88252 183376
rect 88012 183354 88036 183356
rect 88092 183354 88116 183356
rect 88172 183354 88196 183356
rect 88034 183302 88036 183354
rect 88098 183302 88110 183354
rect 88172 183302 88174 183354
rect 88012 183300 88036 183302
rect 88092 183300 88116 183302
rect 88172 183300 88196 183302
rect 87956 183280 88252 183300
rect 85956 182812 86252 182832
rect 86012 182810 86036 182812
rect 86092 182810 86116 182812
rect 86172 182810 86196 182812
rect 86034 182758 86036 182810
rect 86098 182758 86110 182810
rect 86172 182758 86174 182810
rect 86012 182756 86036 182758
rect 86092 182756 86116 182758
rect 86172 182756 86196 182758
rect 85956 182736 86252 182756
rect 89956 182812 90252 182832
rect 90012 182810 90036 182812
rect 90092 182810 90116 182812
rect 90172 182810 90196 182812
rect 90034 182758 90036 182810
rect 90098 182758 90110 182810
rect 90172 182758 90174 182810
rect 90012 182756 90036 182758
rect 90092 182756 90116 182758
rect 90172 182756 90196 182758
rect 89956 182736 90252 182756
rect 87956 182268 88252 182288
rect 88012 182266 88036 182268
rect 88092 182266 88116 182268
rect 88172 182266 88196 182268
rect 88034 182214 88036 182266
rect 88098 182214 88110 182266
rect 88172 182214 88174 182266
rect 88012 182212 88036 182214
rect 88092 182212 88116 182214
rect 88172 182212 88196 182214
rect 87956 182192 88252 182212
rect 85956 181724 86252 181744
rect 86012 181722 86036 181724
rect 86092 181722 86116 181724
rect 86172 181722 86196 181724
rect 86034 181670 86036 181722
rect 86098 181670 86110 181722
rect 86172 181670 86174 181722
rect 86012 181668 86036 181670
rect 86092 181668 86116 181670
rect 86172 181668 86196 181670
rect 85956 181648 86252 181668
rect 89956 181724 90252 181744
rect 90012 181722 90036 181724
rect 90092 181722 90116 181724
rect 90172 181722 90196 181724
rect 90034 181670 90036 181722
rect 90098 181670 90110 181722
rect 90172 181670 90174 181722
rect 90012 181668 90036 181670
rect 90092 181668 90116 181670
rect 90172 181668 90196 181670
rect 89956 181648 90252 181668
rect 87694 181520 87750 181529
rect 87694 181455 87750 181464
rect 87708 180878 87736 181455
rect 87956 181180 88252 181200
rect 88012 181178 88036 181180
rect 88092 181178 88116 181180
rect 88172 181178 88196 181180
rect 88034 181126 88036 181178
rect 88098 181126 88110 181178
rect 88172 181126 88174 181178
rect 88012 181124 88036 181126
rect 88092 181124 88116 181126
rect 88172 181124 88196 181126
rect 87956 181104 88252 181124
rect 87696 180872 87748 180878
rect 87696 180814 87748 180820
rect 85956 180636 86252 180656
rect 86012 180634 86036 180636
rect 86092 180634 86116 180636
rect 86172 180634 86196 180636
rect 86034 180582 86036 180634
rect 86098 180582 86110 180634
rect 86172 180582 86174 180634
rect 86012 180580 86036 180582
rect 86092 180580 86116 180582
rect 86172 180580 86196 180582
rect 85956 180560 86252 180580
rect 89956 180636 90252 180656
rect 90012 180634 90036 180636
rect 90092 180634 90116 180636
rect 90172 180634 90196 180636
rect 90034 180582 90036 180634
rect 90098 180582 90110 180634
rect 90172 180582 90174 180634
rect 90012 180580 90036 180582
rect 90092 180580 90116 180582
rect 90172 180580 90196 180582
rect 89956 180560 90252 180580
rect 87956 180092 88252 180112
rect 88012 180090 88036 180092
rect 88092 180090 88116 180092
rect 88172 180090 88196 180092
rect 88034 180038 88036 180090
rect 88098 180038 88110 180090
rect 88172 180038 88174 180090
rect 88012 180036 88036 180038
rect 88092 180036 88116 180038
rect 88172 180036 88196 180038
rect 87956 180016 88252 180036
rect 84568 179648 84620 179654
rect 84568 179590 84620 179596
rect 84476 167476 84528 167482
rect 84476 167418 84528 167424
rect 84476 160132 84528 160138
rect 84476 160074 84528 160080
rect 84384 153876 84436 153882
rect 84384 153818 84436 153824
rect 84200 141228 84252 141234
rect 84200 141170 84252 141176
rect 84212 99521 84240 141170
rect 84488 132494 84516 160074
rect 84396 132466 84516 132494
rect 84396 123418 84424 132466
rect 84580 125882 84608 179590
rect 85956 179548 86252 179568
rect 86012 179546 86036 179548
rect 86092 179546 86116 179548
rect 86172 179546 86196 179548
rect 86034 179494 86036 179546
rect 86098 179494 86110 179546
rect 86172 179494 86174 179546
rect 86012 179492 86036 179494
rect 86092 179492 86116 179494
rect 86172 179492 86196 179494
rect 85956 179472 86252 179492
rect 89956 179548 90252 179568
rect 90012 179546 90036 179548
rect 90092 179546 90116 179548
rect 90172 179546 90196 179548
rect 90034 179494 90036 179546
rect 90098 179494 90110 179546
rect 90172 179494 90174 179546
rect 90012 179492 90036 179494
rect 90092 179492 90116 179494
rect 90172 179492 90196 179494
rect 89956 179472 90252 179492
rect 87956 179004 88252 179024
rect 88012 179002 88036 179004
rect 88092 179002 88116 179004
rect 88172 179002 88196 179004
rect 88034 178950 88036 179002
rect 88098 178950 88110 179002
rect 88172 178950 88174 179002
rect 88012 178948 88036 178950
rect 88092 178948 88116 178950
rect 88172 178948 88196 178950
rect 87956 178928 88252 178948
rect 85956 178460 86252 178480
rect 86012 178458 86036 178460
rect 86092 178458 86116 178460
rect 86172 178458 86196 178460
rect 86034 178406 86036 178458
rect 86098 178406 86110 178458
rect 86172 178406 86174 178458
rect 86012 178404 86036 178406
rect 86092 178404 86116 178406
rect 86172 178404 86196 178406
rect 85956 178384 86252 178404
rect 89956 178460 90252 178480
rect 90012 178458 90036 178460
rect 90092 178458 90116 178460
rect 90172 178458 90196 178460
rect 90034 178406 90036 178458
rect 90098 178406 90110 178458
rect 90172 178406 90174 178458
rect 90012 178404 90036 178406
rect 90092 178404 90116 178406
rect 90172 178404 90196 178406
rect 89956 178384 90252 178404
rect 87956 177916 88252 177936
rect 88012 177914 88036 177916
rect 88092 177914 88116 177916
rect 88172 177914 88196 177916
rect 88034 177862 88036 177914
rect 88098 177862 88110 177914
rect 88172 177862 88174 177914
rect 88012 177860 88036 177862
rect 88092 177860 88116 177862
rect 88172 177860 88196 177862
rect 87956 177840 88252 177860
rect 87786 177712 87842 177721
rect 87786 177647 87842 177656
rect 85956 177372 86252 177392
rect 86012 177370 86036 177372
rect 86092 177370 86116 177372
rect 86172 177370 86196 177372
rect 86034 177318 86036 177370
rect 86098 177318 86110 177370
rect 86172 177318 86174 177370
rect 86012 177316 86036 177318
rect 86092 177316 86116 177318
rect 86172 177316 86196 177318
rect 85956 177296 86252 177316
rect 85956 176284 86252 176304
rect 86012 176282 86036 176284
rect 86092 176282 86116 176284
rect 86172 176282 86196 176284
rect 86034 176230 86036 176282
rect 86098 176230 86110 176282
rect 86172 176230 86174 176282
rect 86012 176228 86036 176230
rect 86092 176228 86116 176230
rect 86172 176228 86196 176230
rect 85956 176208 86252 176228
rect 85956 175196 86252 175216
rect 86012 175194 86036 175196
rect 86092 175194 86116 175196
rect 86172 175194 86196 175196
rect 86034 175142 86036 175194
rect 86098 175142 86110 175194
rect 86172 175142 86174 175194
rect 86012 175140 86036 175142
rect 86092 175140 86116 175142
rect 86172 175140 86196 175142
rect 85956 175120 86252 175140
rect 87418 174312 87474 174321
rect 87418 174247 87474 174256
rect 85956 174108 86252 174128
rect 86012 174106 86036 174108
rect 86092 174106 86116 174108
rect 86172 174106 86196 174108
rect 86034 174054 86036 174106
rect 86098 174054 86110 174106
rect 86172 174054 86174 174106
rect 86012 174052 86036 174054
rect 86092 174052 86116 174054
rect 86172 174052 86196 174054
rect 85956 174032 86252 174052
rect 87432 173942 87460 174247
rect 87420 173936 87472 173942
rect 87420 173878 87472 173884
rect 87602 173224 87658 173233
rect 87602 173159 87658 173168
rect 85956 173020 86252 173040
rect 86012 173018 86036 173020
rect 86092 173018 86116 173020
rect 86172 173018 86196 173020
rect 86034 172966 86036 173018
rect 86098 172966 86110 173018
rect 86172 172966 86174 173018
rect 86012 172964 86036 172966
rect 86092 172964 86116 172966
rect 86172 172964 86196 172966
rect 85956 172944 86252 172964
rect 85956 171932 86252 171952
rect 86012 171930 86036 171932
rect 86092 171930 86116 171932
rect 86172 171930 86196 171932
rect 86034 171878 86036 171930
rect 86098 171878 86110 171930
rect 86172 171878 86174 171930
rect 86012 171876 86036 171878
rect 86092 171876 86116 171878
rect 86172 171876 86196 171878
rect 85956 171856 86252 171876
rect 85956 170844 86252 170864
rect 86012 170842 86036 170844
rect 86092 170842 86116 170844
rect 86172 170842 86196 170844
rect 86034 170790 86036 170842
rect 86098 170790 86110 170842
rect 86172 170790 86174 170842
rect 86012 170788 86036 170790
rect 86092 170788 86116 170790
rect 86172 170788 86196 170790
rect 85956 170768 86252 170788
rect 85956 169756 86252 169776
rect 86012 169754 86036 169756
rect 86092 169754 86116 169756
rect 86172 169754 86196 169756
rect 86034 169702 86036 169754
rect 86098 169702 86110 169754
rect 86172 169702 86174 169754
rect 86012 169700 86036 169702
rect 86092 169700 86116 169702
rect 86172 169700 86196 169702
rect 85956 169680 86252 169700
rect 85956 168668 86252 168688
rect 86012 168666 86036 168668
rect 86092 168666 86116 168668
rect 86172 168666 86196 168668
rect 86034 168614 86036 168666
rect 86098 168614 86110 168666
rect 86172 168614 86174 168666
rect 86012 168612 86036 168614
rect 86092 168612 86116 168614
rect 86172 168612 86196 168614
rect 85956 168592 86252 168612
rect 87050 168328 87106 168337
rect 87050 168263 87106 168272
rect 85956 167580 86252 167600
rect 86012 167578 86036 167580
rect 86092 167578 86116 167580
rect 86172 167578 86196 167580
rect 86034 167526 86036 167578
rect 86098 167526 86110 167578
rect 86172 167526 86174 167578
rect 86012 167524 86036 167526
rect 86092 167524 86116 167526
rect 86172 167524 86196 167526
rect 85956 167504 86252 167524
rect 87064 167142 87092 168263
rect 87052 167136 87104 167142
rect 87052 167078 87104 167084
rect 85956 166492 86252 166512
rect 86012 166490 86036 166492
rect 86092 166490 86116 166492
rect 86172 166490 86196 166492
rect 86034 166438 86036 166490
rect 86098 166438 86110 166490
rect 86172 166438 86174 166490
rect 86012 166436 86036 166438
rect 86092 166436 86116 166438
rect 86172 166436 86196 166438
rect 85956 166416 86252 166436
rect 87510 165744 87566 165753
rect 87510 165679 87566 165688
rect 85956 165404 86252 165424
rect 86012 165402 86036 165404
rect 86092 165402 86116 165404
rect 86172 165402 86196 165404
rect 86034 165350 86036 165402
rect 86098 165350 86110 165402
rect 86172 165350 86174 165402
rect 86012 165348 86036 165350
rect 86092 165348 86116 165350
rect 86172 165348 86196 165350
rect 85956 165328 86252 165348
rect 85956 164316 86252 164336
rect 86012 164314 86036 164316
rect 86092 164314 86116 164316
rect 86172 164314 86196 164316
rect 86034 164262 86036 164314
rect 86098 164262 86110 164314
rect 86172 164262 86174 164314
rect 86012 164260 86036 164262
rect 86092 164260 86116 164262
rect 86172 164260 86196 164262
rect 85956 164240 86252 164260
rect 85956 163228 86252 163248
rect 86012 163226 86036 163228
rect 86092 163226 86116 163228
rect 86172 163226 86196 163228
rect 86034 163174 86036 163226
rect 86098 163174 86110 163226
rect 86172 163174 86174 163226
rect 86012 163172 86036 163174
rect 86092 163172 86116 163174
rect 86172 163172 86196 163174
rect 85956 163152 86252 163172
rect 84660 162444 84712 162450
rect 84660 162386 84712 162392
rect 84672 162042 84700 162386
rect 85120 162376 85172 162382
rect 85120 162318 85172 162324
rect 84660 162036 84712 162042
rect 84660 161978 84712 161984
rect 84672 141098 84700 161978
rect 85132 161809 85160 162318
rect 85956 162140 86252 162160
rect 86012 162138 86036 162140
rect 86092 162138 86116 162140
rect 86172 162138 86196 162140
rect 86034 162086 86036 162138
rect 86098 162086 86110 162138
rect 86172 162086 86174 162138
rect 86012 162084 86036 162086
rect 86092 162084 86116 162086
rect 86172 162084 86196 162086
rect 85956 162064 86252 162084
rect 85118 161800 85174 161809
rect 85118 161735 85174 161744
rect 85956 161052 86252 161072
rect 86012 161050 86036 161052
rect 86092 161050 86116 161052
rect 86172 161050 86196 161052
rect 86034 160998 86036 161050
rect 86098 160998 86110 161050
rect 86172 160998 86174 161050
rect 86012 160996 86036 160998
rect 86092 160996 86116 160998
rect 86172 160996 86196 160998
rect 85956 160976 86252 160996
rect 85956 159964 86252 159984
rect 86012 159962 86036 159964
rect 86092 159962 86116 159964
rect 86172 159962 86196 159964
rect 86034 159910 86036 159962
rect 86098 159910 86110 159962
rect 86172 159910 86174 159962
rect 86012 159908 86036 159910
rect 86092 159908 86116 159910
rect 86172 159908 86196 159910
rect 85956 159888 86252 159908
rect 87418 159760 87474 159769
rect 87418 159695 87474 159704
rect 85956 158876 86252 158896
rect 86012 158874 86036 158876
rect 86092 158874 86116 158876
rect 86172 158874 86196 158876
rect 86034 158822 86036 158874
rect 86098 158822 86110 158874
rect 86172 158822 86174 158874
rect 86012 158820 86036 158822
rect 86092 158820 86116 158822
rect 86172 158820 86196 158822
rect 85956 158800 86252 158820
rect 86590 158536 86646 158545
rect 86590 158471 86646 158480
rect 85956 157788 86252 157808
rect 86012 157786 86036 157788
rect 86092 157786 86116 157788
rect 86172 157786 86196 157788
rect 86034 157734 86036 157786
rect 86098 157734 86110 157786
rect 86172 157734 86174 157786
rect 86012 157732 86036 157734
rect 86092 157732 86116 157734
rect 86172 157732 86196 157734
rect 85956 157712 86252 157732
rect 85956 156700 86252 156720
rect 86012 156698 86036 156700
rect 86092 156698 86116 156700
rect 86172 156698 86196 156700
rect 86034 156646 86036 156698
rect 86098 156646 86110 156698
rect 86172 156646 86174 156698
rect 86012 156644 86036 156646
rect 86092 156644 86116 156646
rect 86172 156644 86196 156646
rect 85956 156624 86252 156644
rect 85956 155612 86252 155632
rect 86012 155610 86036 155612
rect 86092 155610 86116 155612
rect 86172 155610 86196 155612
rect 86034 155558 86036 155610
rect 86098 155558 86110 155610
rect 86172 155558 86174 155610
rect 86012 155556 86036 155558
rect 86092 155556 86116 155558
rect 86172 155556 86196 155558
rect 85956 155536 86252 155556
rect 85956 154524 86252 154544
rect 86012 154522 86036 154524
rect 86092 154522 86116 154524
rect 86172 154522 86196 154524
rect 86034 154470 86036 154522
rect 86098 154470 86110 154522
rect 86172 154470 86174 154522
rect 86012 154468 86036 154470
rect 86092 154468 86116 154470
rect 86172 154468 86196 154470
rect 85956 154448 86252 154468
rect 85956 153436 86252 153456
rect 86012 153434 86036 153436
rect 86092 153434 86116 153436
rect 86172 153434 86196 153436
rect 86034 153382 86036 153434
rect 86098 153382 86110 153434
rect 86172 153382 86174 153434
rect 86012 153380 86036 153382
rect 86092 153380 86116 153382
rect 86172 153380 86196 153382
rect 85956 153360 86252 153380
rect 85956 152348 86252 152368
rect 86012 152346 86036 152348
rect 86092 152346 86116 152348
rect 86172 152346 86196 152348
rect 86034 152294 86036 152346
rect 86098 152294 86110 152346
rect 86172 152294 86174 152346
rect 86012 152292 86036 152294
rect 86092 152292 86116 152294
rect 86172 152292 86196 152294
rect 85956 152272 86252 152292
rect 85956 151260 86252 151280
rect 86012 151258 86036 151260
rect 86092 151258 86116 151260
rect 86172 151258 86196 151260
rect 86034 151206 86036 151258
rect 86098 151206 86110 151258
rect 86172 151206 86174 151258
rect 86012 151204 86036 151206
rect 86092 151204 86116 151206
rect 86172 151204 86196 151206
rect 85956 151184 86252 151204
rect 85956 150172 86252 150192
rect 86012 150170 86036 150172
rect 86092 150170 86116 150172
rect 86172 150170 86196 150172
rect 86034 150118 86036 150170
rect 86098 150118 86110 150170
rect 86172 150118 86174 150170
rect 86012 150116 86036 150118
rect 86092 150116 86116 150118
rect 86172 150116 86196 150118
rect 85956 150096 86252 150116
rect 85956 149084 86252 149104
rect 86012 149082 86036 149084
rect 86092 149082 86116 149084
rect 86172 149082 86196 149084
rect 86034 149030 86036 149082
rect 86098 149030 86110 149082
rect 86172 149030 86174 149082
rect 86012 149028 86036 149030
rect 86092 149028 86116 149030
rect 86172 149028 86196 149030
rect 85956 149008 86252 149028
rect 85956 147996 86252 148016
rect 86012 147994 86036 147996
rect 86092 147994 86116 147996
rect 86172 147994 86196 147996
rect 86034 147942 86036 147994
rect 86098 147942 86110 147994
rect 86172 147942 86174 147994
rect 86012 147940 86036 147942
rect 86092 147940 86116 147942
rect 86172 147940 86196 147942
rect 85956 147920 86252 147940
rect 85956 146908 86252 146928
rect 86012 146906 86036 146908
rect 86092 146906 86116 146908
rect 86172 146906 86196 146908
rect 86034 146854 86036 146906
rect 86098 146854 86110 146906
rect 86172 146854 86174 146906
rect 86012 146852 86036 146854
rect 86092 146852 86116 146854
rect 86172 146852 86196 146854
rect 85956 146832 86252 146852
rect 85956 145820 86252 145840
rect 86012 145818 86036 145820
rect 86092 145818 86116 145820
rect 86172 145818 86196 145820
rect 86034 145766 86036 145818
rect 86098 145766 86110 145818
rect 86172 145766 86174 145818
rect 86012 145764 86036 145766
rect 86092 145764 86116 145766
rect 86172 145764 86196 145766
rect 85956 145744 86252 145764
rect 84752 144968 84804 144974
rect 84752 144910 84804 144916
rect 84660 141092 84712 141098
rect 84660 141034 84712 141040
rect 84488 125854 84608 125882
rect 84488 124506 84516 125854
rect 84568 125792 84620 125798
rect 84566 125760 84568 125769
rect 84620 125760 84622 125769
rect 84566 125695 84622 125704
rect 84476 124500 84528 124506
rect 84476 124442 84528 124448
rect 84488 124137 84516 124442
rect 84474 124128 84530 124137
rect 84474 124063 84530 124072
rect 84384 123412 84436 123418
rect 84384 123354 84436 123360
rect 84396 123049 84424 123354
rect 84382 123040 84438 123049
rect 84382 122975 84438 122984
rect 84474 121000 84530 121009
rect 84474 120935 84530 120944
rect 84488 120902 84516 120935
rect 84476 120896 84528 120902
rect 84476 120838 84528 120844
rect 84382 118280 84438 118289
rect 84382 118215 84438 118224
rect 84396 118182 84424 118215
rect 84384 118176 84436 118182
rect 84384 118118 84436 118124
rect 84292 108996 84344 109002
rect 84292 108938 84344 108944
rect 84198 99512 84254 99521
rect 84198 99447 84254 99456
rect 84304 97510 84332 108938
rect 84292 97504 84344 97510
rect 84292 97446 84344 97452
rect 84304 96966 84332 97446
rect 84292 96960 84344 96966
rect 84292 96902 84344 96908
rect 84106 94752 84162 94761
rect 84106 94687 84162 94696
rect 84014 94480 84070 94489
rect 84014 94415 84070 94424
rect 84016 93560 84068 93566
rect 84016 93502 84068 93508
rect 83924 93016 83976 93022
rect 83924 92958 83976 92964
rect 83832 85264 83884 85270
rect 83832 85206 83884 85212
rect 83936 84946 83964 92958
rect 83844 84918 83964 84946
rect 83844 66230 83872 84918
rect 84028 84810 84056 93502
rect 84108 93288 84160 93294
rect 84108 93230 84160 93236
rect 83936 84782 84056 84810
rect 83936 69018 83964 84782
rect 84120 84674 84148 93230
rect 84200 93152 84252 93158
rect 84200 93094 84252 93100
rect 84028 84646 84148 84674
rect 84028 70378 84056 84646
rect 84108 84584 84160 84590
rect 84108 84526 84160 84532
rect 84120 77178 84148 84526
rect 84108 77172 84160 77178
rect 84108 77114 84160 77120
rect 84016 70372 84068 70378
rect 84016 70314 84068 70320
rect 83924 69012 83976 69018
rect 83924 68954 83976 68960
rect 83832 66224 83884 66230
rect 83832 66166 83884 66172
rect 84212 66162 84240 93094
rect 84292 92948 84344 92954
rect 84292 92890 84344 92896
rect 84200 66156 84252 66162
rect 84200 66098 84252 66104
rect 83740 63504 83792 63510
rect 83740 63446 83792 63452
rect 84304 61946 84332 92890
rect 84292 61940 84344 61946
rect 84292 61882 84344 61888
rect 83740 45620 83792 45626
rect 83740 45562 83792 45568
rect 83648 4344 83700 4350
rect 83648 4286 83700 4292
rect 83648 4208 83700 4214
rect 83648 4150 83700 4156
rect 83660 3330 83688 4150
rect 83648 3324 83700 3330
rect 83648 3266 83700 3272
rect 83556 3256 83608 3262
rect 83556 3198 83608 3204
rect 83462 3088 83518 3097
rect 83462 3023 83518 3032
rect 83556 2780 83608 2786
rect 83556 2722 83608 2728
rect 83568 2310 83596 2722
rect 83556 2304 83608 2310
rect 83556 2246 83608 2252
rect 83372 2032 83424 2038
rect 83372 1974 83424 1980
rect 83280 1964 83332 1970
rect 83280 1906 83332 1912
rect 83188 1624 83240 1630
rect 83568 1601 83596 2246
rect 83188 1566 83240 1572
rect 83554 1592 83610 1601
rect 83554 1527 83610 1536
rect 83096 1488 83148 1494
rect 83096 1430 83148 1436
rect 82728 536 82780 542
rect 82728 478 82780 484
rect 83752 406 83780 45562
rect 83832 44192 83884 44198
rect 83832 44134 83884 44140
rect 83844 474 83872 44134
rect 84396 39098 84424 118118
rect 84384 39092 84436 39098
rect 84384 39034 84436 39040
rect 83924 27668 83976 27674
rect 83924 27610 83976 27616
rect 83936 2242 83964 27610
rect 84016 26308 84068 26314
rect 84016 26250 84068 26256
rect 83924 2236 83976 2242
rect 83924 2178 83976 2184
rect 84028 2174 84056 26250
rect 84290 24440 84346 24449
rect 84290 24375 84292 24384
rect 84344 24375 84346 24384
rect 84292 24346 84344 24352
rect 84108 23520 84160 23526
rect 84108 23462 84160 23468
rect 84016 2168 84068 2174
rect 84016 2110 84068 2116
rect 84120 2106 84148 23462
rect 84290 23352 84346 23361
rect 84290 23287 84292 23296
rect 84344 23287 84346 23296
rect 84292 23258 84344 23264
rect 84488 17746 84516 120838
rect 84566 120184 84622 120193
rect 84566 120119 84622 120128
rect 84580 120086 84608 120119
rect 84568 120080 84620 120086
rect 84568 120022 84620 120028
rect 84566 117328 84622 117337
rect 84566 117263 84622 117272
rect 84580 117094 84608 117263
rect 84568 117088 84620 117094
rect 84568 117030 84620 117036
rect 84580 93430 84608 117030
rect 84568 93424 84620 93430
rect 84568 93366 84620 93372
rect 84566 93256 84622 93265
rect 84566 93191 84622 93200
rect 84580 84998 84608 93191
rect 84568 84992 84620 84998
rect 84568 84934 84620 84940
rect 84568 29300 84620 29306
rect 84568 29242 84620 29248
rect 84580 28937 84608 29242
rect 84566 28928 84622 28937
rect 84566 28863 84622 28872
rect 84568 27600 84620 27606
rect 84566 27568 84568 27577
rect 84620 27568 84622 27577
rect 84566 27503 84622 27512
rect 84568 26580 84620 26586
rect 84568 26522 84620 26528
rect 84580 26217 84608 26522
rect 84566 26208 84622 26217
rect 84566 26143 84622 26152
rect 84568 22228 84620 22234
rect 84568 22170 84620 22176
rect 84476 17740 84528 17746
rect 84476 17682 84528 17688
rect 84476 15360 84528 15366
rect 84476 15302 84528 15308
rect 84108 2100 84160 2106
rect 84108 2042 84160 2048
rect 84488 1834 84516 15302
rect 84580 1902 84608 22170
rect 84672 14618 84700 141034
rect 84764 97481 84792 144910
rect 85956 144732 86252 144752
rect 86012 144730 86036 144732
rect 86092 144730 86116 144732
rect 86172 144730 86196 144732
rect 86034 144678 86036 144730
rect 86098 144678 86110 144730
rect 86172 144678 86174 144730
rect 86012 144676 86036 144678
rect 86092 144676 86116 144678
rect 86172 144676 86196 144678
rect 85956 144656 86252 144676
rect 85764 143744 85816 143750
rect 85764 143686 85816 143692
rect 85212 141024 85264 141030
rect 85212 140966 85264 140972
rect 85120 140004 85172 140010
rect 85120 139946 85172 139952
rect 84844 138916 84896 138922
rect 84844 138858 84896 138864
rect 84856 97850 84884 138858
rect 84936 131232 84988 131238
rect 84936 131174 84988 131180
rect 84948 98054 84976 131174
rect 85028 99680 85080 99686
rect 85028 99622 85080 99628
rect 84936 98048 84988 98054
rect 84936 97990 84988 97996
rect 84844 97844 84896 97850
rect 84844 97786 84896 97792
rect 85040 97730 85068 99622
rect 85132 99521 85160 139946
rect 85224 109614 85252 140966
rect 85580 131300 85632 131306
rect 85580 131242 85632 131248
rect 85486 118416 85542 118425
rect 85486 118351 85542 118360
rect 85396 113892 85448 113898
rect 85396 113834 85448 113840
rect 85304 111852 85356 111858
rect 85304 111794 85356 111800
rect 85212 109608 85264 109614
rect 85212 109550 85264 109556
rect 85212 108656 85264 108662
rect 85212 108598 85264 108604
rect 85118 99512 85174 99521
rect 85118 99447 85174 99456
rect 85118 99376 85174 99385
rect 85118 99311 85174 99320
rect 84948 97702 85068 97730
rect 84844 97504 84896 97510
rect 84750 97472 84806 97481
rect 84844 97446 84896 97452
rect 84750 97407 84806 97416
rect 84752 97300 84804 97306
rect 84752 97242 84804 97248
rect 84764 96218 84792 97242
rect 84856 96422 84884 97446
rect 84948 96966 84976 97702
rect 85026 97472 85082 97481
rect 85026 97407 85082 97416
rect 84936 96960 84988 96966
rect 84936 96902 84988 96908
rect 84844 96416 84896 96422
rect 84844 96358 84896 96364
rect 84752 96212 84804 96218
rect 84752 96154 84804 96160
rect 84764 93430 84792 96154
rect 84856 94314 84884 96358
rect 84948 94489 84976 96902
rect 85040 95878 85068 97407
rect 85132 96422 85160 99311
rect 85120 96416 85172 96422
rect 85120 96358 85172 96364
rect 85028 95872 85080 95878
rect 85028 95814 85080 95820
rect 85224 95130 85252 108598
rect 85316 97034 85344 111794
rect 85408 99686 85436 113834
rect 85500 110362 85528 118351
rect 85488 110356 85540 110362
rect 85488 110298 85540 110304
rect 85488 104576 85540 104582
rect 85488 104518 85540 104524
rect 85500 99686 85528 104518
rect 85396 99680 85448 99686
rect 85396 99622 85448 99628
rect 85488 99680 85540 99686
rect 85488 99622 85540 99628
rect 85592 99498 85620 131242
rect 85672 114572 85724 114578
rect 85672 114514 85724 114520
rect 85684 104310 85712 114514
rect 85672 104304 85724 104310
rect 85672 104246 85724 104252
rect 85670 104136 85726 104145
rect 85670 104071 85726 104080
rect 85684 99770 85712 104071
rect 85776 100026 85804 143686
rect 85956 143644 86252 143664
rect 86012 143642 86036 143644
rect 86092 143642 86116 143644
rect 86172 143642 86196 143644
rect 86034 143590 86036 143642
rect 86098 143590 86110 143642
rect 86172 143590 86174 143642
rect 86012 143588 86036 143590
rect 86092 143588 86116 143590
rect 86172 143588 86196 143590
rect 85956 143568 86252 143588
rect 85956 142556 86252 142576
rect 86012 142554 86036 142556
rect 86092 142554 86116 142556
rect 86172 142554 86196 142556
rect 86034 142502 86036 142554
rect 86098 142502 86110 142554
rect 86172 142502 86174 142554
rect 86012 142500 86036 142502
rect 86092 142500 86116 142502
rect 86172 142500 86196 142502
rect 85956 142480 86252 142500
rect 85856 142452 85908 142458
rect 85856 142394 85908 142400
rect 85868 131238 85896 142394
rect 85956 141468 86252 141488
rect 86012 141466 86036 141468
rect 86092 141466 86116 141468
rect 86172 141466 86196 141468
rect 86034 141414 86036 141466
rect 86098 141414 86110 141466
rect 86172 141414 86174 141466
rect 86012 141412 86036 141414
rect 86092 141412 86116 141414
rect 86172 141412 86196 141414
rect 85956 141392 86252 141412
rect 85956 140380 86252 140400
rect 86012 140378 86036 140380
rect 86092 140378 86116 140380
rect 86172 140378 86196 140380
rect 86034 140326 86036 140378
rect 86098 140326 86110 140378
rect 86172 140326 86174 140378
rect 86012 140324 86036 140326
rect 86092 140324 86116 140326
rect 86172 140324 86196 140326
rect 85956 140304 86252 140324
rect 85956 139292 86252 139312
rect 86012 139290 86036 139292
rect 86092 139290 86116 139292
rect 86172 139290 86196 139292
rect 86034 139238 86036 139290
rect 86098 139238 86110 139290
rect 86172 139238 86174 139290
rect 86012 139236 86036 139238
rect 86092 139236 86116 139238
rect 86172 139236 86196 139238
rect 85956 139216 86252 139236
rect 85956 138204 86252 138224
rect 86012 138202 86036 138204
rect 86092 138202 86116 138204
rect 86172 138202 86196 138204
rect 86034 138150 86036 138202
rect 86098 138150 86110 138202
rect 86172 138150 86174 138202
rect 86012 138148 86036 138150
rect 86092 138148 86116 138150
rect 86172 138148 86196 138150
rect 85956 138128 86252 138148
rect 86498 137864 86554 137873
rect 86498 137799 86554 137808
rect 85956 137116 86252 137136
rect 86012 137114 86036 137116
rect 86092 137114 86116 137116
rect 86172 137114 86196 137116
rect 86034 137062 86036 137114
rect 86098 137062 86110 137114
rect 86172 137062 86174 137114
rect 86012 137060 86036 137062
rect 86092 137060 86116 137062
rect 86172 137060 86196 137062
rect 85956 137040 86252 137060
rect 86314 136368 86370 136377
rect 86314 136303 86370 136312
rect 85956 136028 86252 136048
rect 86012 136026 86036 136028
rect 86092 136026 86116 136028
rect 86172 136026 86196 136028
rect 86034 135974 86036 136026
rect 86098 135974 86110 136026
rect 86172 135974 86174 136026
rect 86012 135972 86036 135974
rect 86092 135972 86116 135974
rect 86172 135972 86196 135974
rect 85956 135952 86252 135972
rect 85956 134940 86252 134960
rect 86012 134938 86036 134940
rect 86092 134938 86116 134940
rect 86172 134938 86196 134940
rect 86034 134886 86036 134938
rect 86098 134886 86110 134938
rect 86172 134886 86174 134938
rect 86012 134884 86036 134886
rect 86092 134884 86116 134886
rect 86172 134884 86196 134886
rect 85956 134864 86252 134884
rect 85956 133852 86252 133872
rect 86012 133850 86036 133852
rect 86092 133850 86116 133852
rect 86172 133850 86196 133852
rect 86034 133798 86036 133850
rect 86098 133798 86110 133850
rect 86172 133798 86174 133850
rect 86012 133796 86036 133798
rect 86092 133796 86116 133798
rect 86172 133796 86196 133798
rect 85956 133776 86252 133796
rect 85956 132764 86252 132784
rect 86012 132762 86036 132764
rect 86092 132762 86116 132764
rect 86172 132762 86196 132764
rect 86034 132710 86036 132762
rect 86098 132710 86110 132762
rect 86172 132710 86174 132762
rect 86012 132708 86036 132710
rect 86092 132708 86116 132710
rect 86172 132708 86196 132710
rect 85956 132688 86252 132708
rect 85956 131676 86252 131696
rect 86012 131674 86036 131676
rect 86092 131674 86116 131676
rect 86172 131674 86196 131676
rect 86034 131622 86036 131674
rect 86098 131622 86110 131674
rect 86172 131622 86174 131674
rect 86012 131620 86036 131622
rect 86092 131620 86116 131622
rect 86172 131620 86196 131622
rect 85956 131600 86252 131620
rect 85856 131232 85908 131238
rect 85856 131174 85908 131180
rect 85956 130588 86252 130608
rect 86012 130586 86036 130588
rect 86092 130586 86116 130588
rect 86172 130586 86196 130588
rect 86034 130534 86036 130586
rect 86098 130534 86110 130586
rect 86172 130534 86174 130586
rect 86012 130532 86036 130534
rect 86092 130532 86116 130534
rect 86172 130532 86196 130534
rect 85956 130512 86252 130532
rect 85956 129500 86252 129520
rect 86012 129498 86036 129500
rect 86092 129498 86116 129500
rect 86172 129498 86196 129500
rect 86034 129446 86036 129498
rect 86098 129446 86110 129498
rect 86172 129446 86174 129498
rect 86012 129444 86036 129446
rect 86092 129444 86116 129446
rect 86172 129444 86196 129446
rect 85956 129424 86252 129444
rect 85956 128412 86252 128432
rect 86012 128410 86036 128412
rect 86092 128410 86116 128412
rect 86172 128410 86196 128412
rect 86034 128358 86036 128410
rect 86098 128358 86110 128410
rect 86172 128358 86174 128410
rect 86012 128356 86036 128358
rect 86092 128356 86116 128358
rect 86172 128356 86196 128358
rect 85956 128336 86252 128356
rect 85956 127324 86252 127344
rect 86012 127322 86036 127324
rect 86092 127322 86116 127324
rect 86172 127322 86196 127324
rect 86034 127270 86036 127322
rect 86098 127270 86110 127322
rect 86172 127270 86174 127322
rect 86012 127268 86036 127270
rect 86092 127268 86116 127270
rect 86172 127268 86196 127270
rect 85956 127248 86252 127268
rect 85956 126236 86252 126256
rect 86012 126234 86036 126236
rect 86092 126234 86116 126236
rect 86172 126234 86196 126236
rect 86034 126182 86036 126234
rect 86098 126182 86110 126234
rect 86172 126182 86174 126234
rect 86012 126180 86036 126182
rect 86092 126180 86116 126182
rect 86172 126180 86196 126182
rect 85956 126160 86252 126180
rect 85956 125148 86252 125168
rect 86012 125146 86036 125148
rect 86092 125146 86116 125148
rect 86172 125146 86196 125148
rect 86034 125094 86036 125146
rect 86098 125094 86110 125146
rect 86172 125094 86174 125146
rect 86012 125092 86036 125094
rect 86092 125092 86116 125094
rect 86172 125092 86196 125094
rect 85956 125072 86252 125092
rect 85956 124060 86252 124080
rect 86012 124058 86036 124060
rect 86092 124058 86116 124060
rect 86172 124058 86196 124060
rect 86034 124006 86036 124058
rect 86098 124006 86110 124058
rect 86172 124006 86174 124058
rect 86012 124004 86036 124006
rect 86092 124004 86116 124006
rect 86172 124004 86196 124006
rect 85956 123984 86252 124004
rect 85956 122972 86252 122992
rect 86012 122970 86036 122972
rect 86092 122970 86116 122972
rect 86172 122970 86196 122972
rect 86034 122918 86036 122970
rect 86098 122918 86110 122970
rect 86172 122918 86174 122970
rect 86012 122916 86036 122918
rect 86092 122916 86116 122918
rect 86172 122916 86196 122918
rect 85956 122896 86252 122916
rect 86328 122834 86356 136303
rect 86406 135280 86462 135289
rect 86406 135215 86462 135224
rect 85868 122806 86356 122834
rect 85868 109698 85896 122806
rect 85956 121884 86252 121904
rect 86012 121882 86036 121884
rect 86092 121882 86116 121884
rect 86172 121882 86196 121884
rect 86034 121830 86036 121882
rect 86098 121830 86110 121882
rect 86172 121830 86174 121882
rect 86012 121828 86036 121830
rect 86092 121828 86116 121830
rect 86172 121828 86196 121830
rect 85956 121808 86252 121828
rect 85956 120796 86252 120816
rect 86012 120794 86036 120796
rect 86092 120794 86116 120796
rect 86172 120794 86196 120796
rect 86034 120742 86036 120794
rect 86098 120742 86110 120794
rect 86172 120742 86174 120794
rect 86012 120740 86036 120742
rect 86092 120740 86116 120742
rect 86172 120740 86196 120742
rect 85956 120720 86252 120740
rect 85956 119708 86252 119728
rect 86012 119706 86036 119708
rect 86092 119706 86116 119708
rect 86172 119706 86196 119708
rect 86034 119654 86036 119706
rect 86098 119654 86110 119706
rect 86172 119654 86174 119706
rect 86012 119652 86036 119654
rect 86092 119652 86116 119654
rect 86172 119652 86196 119654
rect 85956 119632 86252 119652
rect 85956 118620 86252 118640
rect 86012 118618 86036 118620
rect 86092 118618 86116 118620
rect 86172 118618 86196 118620
rect 86034 118566 86036 118618
rect 86098 118566 86110 118618
rect 86172 118566 86174 118618
rect 86012 118564 86036 118566
rect 86092 118564 86116 118566
rect 86172 118564 86196 118566
rect 85956 118544 86252 118564
rect 85956 117532 86252 117552
rect 86012 117530 86036 117532
rect 86092 117530 86116 117532
rect 86172 117530 86196 117532
rect 86034 117478 86036 117530
rect 86098 117478 86110 117530
rect 86172 117478 86174 117530
rect 86012 117476 86036 117478
rect 86092 117476 86116 117478
rect 86172 117476 86196 117478
rect 85956 117456 86252 117476
rect 85956 116444 86252 116464
rect 86012 116442 86036 116444
rect 86092 116442 86116 116444
rect 86172 116442 86196 116444
rect 86034 116390 86036 116442
rect 86098 116390 86110 116442
rect 86172 116390 86174 116442
rect 86012 116388 86036 116390
rect 86092 116388 86116 116390
rect 86172 116388 86196 116390
rect 85956 116368 86252 116388
rect 86314 116104 86370 116113
rect 86314 116039 86370 116048
rect 85956 115356 86252 115376
rect 86012 115354 86036 115356
rect 86092 115354 86116 115356
rect 86172 115354 86196 115356
rect 86034 115302 86036 115354
rect 86098 115302 86110 115354
rect 86172 115302 86174 115354
rect 86012 115300 86036 115302
rect 86092 115300 86116 115302
rect 86172 115300 86196 115302
rect 85956 115280 86252 115300
rect 85956 114268 86252 114288
rect 86012 114266 86036 114268
rect 86092 114266 86116 114268
rect 86172 114266 86196 114268
rect 86034 114214 86036 114266
rect 86098 114214 86110 114266
rect 86172 114214 86174 114266
rect 86012 114212 86036 114214
rect 86092 114212 86116 114214
rect 86172 114212 86196 114214
rect 85956 114192 86252 114212
rect 85956 113180 86252 113200
rect 86012 113178 86036 113180
rect 86092 113178 86116 113180
rect 86172 113178 86196 113180
rect 86034 113126 86036 113178
rect 86098 113126 86110 113178
rect 86172 113126 86174 113178
rect 86012 113124 86036 113126
rect 86092 113124 86116 113126
rect 86172 113124 86196 113126
rect 85956 113104 86252 113124
rect 85956 112092 86252 112112
rect 86012 112090 86036 112092
rect 86092 112090 86116 112092
rect 86172 112090 86196 112092
rect 86034 112038 86036 112090
rect 86098 112038 86110 112090
rect 86172 112038 86174 112090
rect 86012 112036 86036 112038
rect 86092 112036 86116 112038
rect 86172 112036 86196 112038
rect 85956 112016 86252 112036
rect 85956 111004 86252 111024
rect 86012 111002 86036 111004
rect 86092 111002 86116 111004
rect 86172 111002 86196 111004
rect 86034 110950 86036 111002
rect 86098 110950 86110 111002
rect 86172 110950 86174 111002
rect 86012 110948 86036 110950
rect 86092 110948 86116 110950
rect 86172 110948 86196 110950
rect 85956 110928 86252 110948
rect 85956 109916 86252 109936
rect 86012 109914 86036 109916
rect 86092 109914 86116 109916
rect 86172 109914 86196 109916
rect 86034 109862 86036 109914
rect 86098 109862 86110 109914
rect 86172 109862 86174 109914
rect 86012 109860 86036 109862
rect 86092 109860 86116 109862
rect 86172 109860 86196 109862
rect 85956 109840 86252 109860
rect 85868 109670 85988 109698
rect 85856 109608 85908 109614
rect 85856 109550 85908 109556
rect 85764 100020 85816 100026
rect 85764 99962 85816 99968
rect 85868 99890 85896 109550
rect 85960 109002 85988 109670
rect 85948 108996 86000 109002
rect 85948 108938 86000 108944
rect 85956 108828 86252 108848
rect 86012 108826 86036 108828
rect 86092 108826 86116 108828
rect 86172 108826 86196 108828
rect 86034 108774 86036 108826
rect 86098 108774 86110 108826
rect 86172 108774 86174 108826
rect 86012 108772 86036 108774
rect 86092 108772 86116 108774
rect 86172 108772 86196 108774
rect 85956 108752 86252 108772
rect 85956 107740 86252 107760
rect 86012 107738 86036 107740
rect 86092 107738 86116 107740
rect 86172 107738 86196 107740
rect 86034 107686 86036 107738
rect 86098 107686 86110 107738
rect 86172 107686 86174 107738
rect 86012 107684 86036 107686
rect 86092 107684 86116 107686
rect 86172 107684 86196 107686
rect 85956 107664 86252 107684
rect 85956 106652 86252 106672
rect 86012 106650 86036 106652
rect 86092 106650 86116 106652
rect 86172 106650 86196 106652
rect 86034 106598 86036 106650
rect 86098 106598 86110 106650
rect 86172 106598 86174 106650
rect 86012 106596 86036 106598
rect 86092 106596 86116 106598
rect 86172 106596 86196 106598
rect 85956 106576 86252 106596
rect 86328 106554 86356 116039
rect 86316 106548 86368 106554
rect 86316 106490 86368 106496
rect 86420 106434 86448 135215
rect 86512 113898 86540 137799
rect 86500 113892 86552 113898
rect 86500 113834 86552 113840
rect 86498 113520 86554 113529
rect 86498 113455 86554 113464
rect 86236 106406 86448 106434
rect 86236 105738 86264 106406
rect 86316 106344 86368 106350
rect 86316 106286 86368 106292
rect 86406 106312 86462 106321
rect 86224 105732 86276 105738
rect 86224 105674 86276 105680
rect 85956 105564 86252 105584
rect 86012 105562 86036 105564
rect 86092 105562 86116 105564
rect 86172 105562 86196 105564
rect 86034 105510 86036 105562
rect 86098 105510 86110 105562
rect 86172 105510 86174 105562
rect 86012 105508 86036 105510
rect 86092 105508 86116 105510
rect 86172 105508 86196 105510
rect 85956 105488 86252 105508
rect 85956 104476 86252 104496
rect 86012 104474 86036 104476
rect 86092 104474 86116 104476
rect 86172 104474 86196 104476
rect 86034 104422 86036 104474
rect 86098 104422 86110 104474
rect 86172 104422 86174 104474
rect 86012 104420 86036 104422
rect 86092 104420 86116 104422
rect 86172 104420 86196 104422
rect 85956 104400 86252 104420
rect 86328 104394 86356 106286
rect 86406 106247 86462 106256
rect 86420 104582 86448 106247
rect 86512 104582 86540 113455
rect 86408 104576 86460 104582
rect 86408 104518 86460 104524
rect 86500 104576 86552 104582
rect 86500 104518 86552 104524
rect 86328 104366 86540 104394
rect 85956 103388 86252 103408
rect 86012 103386 86036 103388
rect 86092 103386 86116 103388
rect 86172 103386 86196 103388
rect 86034 103334 86036 103386
rect 86098 103334 86110 103386
rect 86172 103334 86174 103386
rect 86012 103332 86036 103334
rect 86092 103332 86116 103334
rect 86172 103332 86196 103334
rect 85956 103312 86252 103332
rect 85956 102300 86252 102320
rect 86012 102298 86036 102300
rect 86092 102298 86116 102300
rect 86172 102298 86196 102300
rect 86034 102246 86036 102298
rect 86098 102246 86110 102298
rect 86172 102246 86174 102298
rect 86012 102244 86036 102246
rect 86092 102244 86116 102246
rect 86172 102244 86196 102246
rect 85956 102224 86252 102244
rect 85956 101212 86252 101232
rect 86012 101210 86036 101212
rect 86092 101210 86116 101212
rect 86172 101210 86196 101212
rect 86034 101158 86036 101210
rect 86098 101158 86110 101210
rect 86172 101158 86174 101210
rect 86012 101156 86036 101158
rect 86092 101156 86116 101158
rect 86172 101156 86196 101158
rect 85956 101136 86252 101156
rect 85956 100124 86252 100144
rect 86012 100122 86036 100124
rect 86092 100122 86116 100124
rect 86172 100122 86196 100124
rect 86034 100070 86036 100122
rect 86098 100070 86110 100122
rect 86172 100070 86174 100122
rect 86012 100068 86036 100070
rect 86092 100068 86116 100070
rect 86172 100068 86196 100070
rect 85956 100048 86252 100068
rect 86408 100020 86460 100026
rect 86408 99962 86460 99968
rect 86132 99952 86184 99958
rect 86132 99894 86184 99900
rect 85856 99884 85908 99890
rect 85856 99826 85908 99832
rect 85684 99742 85804 99770
rect 85672 99680 85724 99686
rect 85672 99622 85724 99628
rect 85396 99476 85448 99482
rect 85396 99418 85448 99424
rect 85500 99470 85620 99498
rect 85408 99278 85436 99418
rect 85396 99272 85448 99278
rect 85396 99214 85448 99220
rect 85394 99104 85450 99113
rect 85394 99039 85450 99048
rect 85408 97850 85436 99039
rect 85396 97844 85448 97850
rect 85396 97786 85448 97792
rect 85304 97028 85356 97034
rect 85304 96970 85356 96976
rect 85408 96506 85436 97786
rect 85316 96478 85436 96506
rect 85500 96506 85528 99470
rect 85580 99408 85632 99414
rect 85580 99350 85632 99356
rect 85592 96694 85620 99350
rect 85580 96688 85632 96694
rect 85580 96630 85632 96636
rect 85500 96478 85620 96506
rect 85212 95124 85264 95130
rect 85212 95066 85264 95072
rect 84934 94480 84990 94489
rect 84934 94415 84990 94424
rect 85316 94382 85344 96478
rect 85396 96416 85448 96422
rect 85396 96358 85448 96364
rect 85408 94450 85436 96358
rect 85488 95872 85540 95878
rect 85488 95814 85540 95820
rect 85500 94586 85528 95814
rect 85592 95441 85620 96478
rect 85578 95432 85634 95441
rect 85578 95367 85634 95376
rect 85488 94580 85540 94586
rect 85488 94522 85540 94528
rect 85396 94444 85448 94450
rect 85396 94386 85448 94392
rect 85304 94376 85356 94382
rect 85304 94318 85356 94324
rect 84844 94308 84896 94314
rect 84844 94250 84896 94256
rect 85316 94058 85344 94318
rect 85224 94030 85344 94058
rect 84936 93968 84988 93974
rect 84936 93910 84988 93916
rect 84752 93424 84804 93430
rect 84752 93366 84804 93372
rect 84752 92880 84804 92886
rect 84752 92822 84804 92828
rect 84764 57934 84792 92822
rect 84844 92744 84896 92750
rect 84844 92686 84896 92692
rect 84856 85134 84884 92686
rect 84948 88330 84976 93910
rect 85118 93664 85174 93673
rect 85118 93599 85174 93608
rect 85026 93528 85082 93537
rect 85026 93463 85082 93472
rect 84936 88324 84988 88330
rect 84936 88266 84988 88272
rect 85040 85377 85068 93463
rect 85132 93430 85160 93599
rect 85120 93424 85172 93430
rect 85120 93366 85172 93372
rect 85224 92834 85252 94030
rect 85304 93900 85356 93906
rect 85304 93842 85356 93848
rect 85132 92806 85252 92834
rect 85026 85368 85082 85377
rect 85026 85303 85082 85312
rect 84844 85128 84896 85134
rect 85132 85082 85160 92806
rect 85212 92744 85264 92750
rect 85212 92686 85264 92692
rect 84844 85070 84896 85076
rect 84948 85054 85160 85082
rect 84844 84992 84896 84998
rect 84844 84934 84896 84940
rect 84752 57928 84804 57934
rect 84752 57870 84804 57876
rect 84856 53786 84884 84934
rect 84844 53780 84896 53786
rect 84844 53722 84896 53728
rect 84844 40112 84896 40118
rect 84844 40054 84896 40060
rect 84750 32056 84806 32065
rect 84750 31991 84752 32000
rect 84804 31991 84806 32000
rect 84752 31962 84804 31968
rect 84752 30320 84804 30326
rect 84750 30288 84752 30297
rect 84804 30288 84806 30297
rect 84750 30223 84806 30232
rect 84752 29028 84804 29034
rect 84752 28970 84804 28976
rect 84660 14612 84712 14618
rect 84660 14554 84712 14560
rect 84672 13870 84700 14554
rect 84660 13864 84712 13870
rect 84660 13806 84712 13812
rect 84568 1896 84620 1902
rect 84568 1838 84620 1844
rect 84476 1828 84528 1834
rect 84476 1770 84528 1776
rect 84764 1086 84792 28970
rect 84752 1080 84804 1086
rect 84752 1022 84804 1028
rect 84856 678 84884 40054
rect 84948 3738 84976 85054
rect 85026 84960 85082 84969
rect 85224 84946 85252 92686
rect 85026 84895 85082 84904
rect 85132 84918 85252 84946
rect 85040 84794 85068 84895
rect 85028 84788 85080 84794
rect 85028 84730 85080 84736
rect 85026 84688 85082 84697
rect 85026 84623 85082 84632
rect 84936 3732 84988 3738
rect 84936 3674 84988 3680
rect 84948 3194 84976 3674
rect 84936 3188 84988 3194
rect 84936 3130 84988 3136
rect 85040 2378 85068 84623
rect 85132 56438 85160 84918
rect 85212 84788 85264 84794
rect 85212 84730 85264 84736
rect 85120 56432 85172 56438
rect 85120 56374 85172 56380
rect 85224 54670 85252 84730
rect 85212 54664 85264 54670
rect 85212 54606 85264 54612
rect 85120 36372 85172 36378
rect 85120 36314 85172 36320
rect 85028 2372 85080 2378
rect 85028 2314 85080 2320
rect 85132 746 85160 36314
rect 85212 34536 85264 34542
rect 85212 34478 85264 34484
rect 85224 882 85252 34478
rect 85316 13938 85344 93842
rect 85408 85105 85436 94386
rect 85394 85096 85450 85105
rect 85394 85031 85450 85040
rect 85500 84946 85528 94522
rect 85580 92064 85632 92070
rect 85578 92032 85580 92041
rect 85632 92032 85634 92041
rect 85578 91967 85634 91976
rect 85580 85128 85632 85134
rect 85580 85070 85632 85076
rect 85408 84918 85528 84946
rect 85304 13932 85356 13938
rect 85304 13874 85356 13880
rect 85304 12640 85356 12646
rect 85304 12582 85356 12588
rect 85316 1562 85344 12582
rect 85408 3738 85436 84918
rect 85592 84810 85620 85070
rect 85500 84782 85620 84810
rect 85500 56506 85528 84782
rect 85488 56500 85540 56506
rect 85488 56442 85540 56448
rect 85488 31816 85540 31822
rect 85488 31758 85540 31764
rect 85396 3732 85448 3738
rect 85396 3674 85448 3680
rect 85304 1556 85356 1562
rect 85304 1498 85356 1504
rect 85500 1018 85528 31758
rect 85684 23322 85712 99622
rect 85776 96558 85804 99742
rect 86144 99414 86172 99894
rect 86224 99884 86276 99890
rect 86224 99826 86276 99832
rect 86132 99408 86184 99414
rect 86132 99350 86184 99356
rect 86236 99328 86264 99826
rect 86236 99300 86356 99328
rect 85856 99272 85908 99278
rect 85856 99214 85908 99220
rect 85764 96552 85816 96558
rect 85764 96494 85816 96500
rect 85868 96082 85896 99214
rect 85956 99036 86252 99056
rect 86012 99034 86036 99036
rect 86092 99034 86116 99036
rect 86172 99034 86196 99036
rect 86034 98982 86036 99034
rect 86098 98982 86110 99034
rect 86172 98982 86174 99034
rect 86012 98980 86036 98982
rect 86092 98980 86116 98982
rect 86172 98980 86196 98982
rect 85956 98960 86252 98980
rect 85956 97948 86252 97968
rect 86012 97946 86036 97948
rect 86092 97946 86116 97948
rect 86172 97946 86196 97948
rect 86034 97894 86036 97946
rect 86098 97894 86110 97946
rect 86172 97894 86174 97946
rect 86012 97892 86036 97894
rect 86092 97892 86116 97894
rect 86172 97892 86196 97894
rect 85956 97872 86252 97892
rect 85956 96860 86252 96880
rect 86012 96858 86036 96860
rect 86092 96858 86116 96860
rect 86172 96858 86196 96860
rect 86034 96806 86036 96858
rect 86098 96806 86110 96858
rect 86172 96806 86174 96858
rect 86012 96804 86036 96806
rect 86092 96804 86116 96806
rect 86172 96804 86196 96806
rect 85956 96784 86252 96804
rect 85948 96688 86000 96694
rect 85948 96630 86000 96636
rect 85856 96076 85908 96082
rect 85856 96018 85908 96024
rect 85960 95860 85988 96630
rect 85776 95832 85988 95860
rect 85776 94790 85804 95832
rect 85956 95772 86252 95792
rect 86012 95770 86036 95772
rect 86092 95770 86116 95772
rect 86172 95770 86196 95772
rect 86034 95718 86036 95770
rect 86098 95718 86110 95770
rect 86172 95718 86174 95770
rect 86012 95716 86036 95718
rect 86092 95716 86116 95718
rect 86172 95716 86196 95718
rect 85956 95696 86252 95716
rect 85856 94988 85908 94994
rect 85856 94930 85908 94936
rect 85764 94784 85816 94790
rect 85764 94726 85816 94732
rect 85672 23316 85724 23322
rect 85672 23258 85724 23264
rect 85776 3534 85804 94726
rect 85868 24410 85896 94930
rect 86328 94858 86356 99300
rect 86420 97102 86448 99962
rect 86512 99482 86540 104366
rect 86604 104242 86632 158471
rect 87326 157040 87382 157049
rect 87326 156975 87382 156984
rect 87142 154864 87198 154873
rect 87142 154799 87198 154808
rect 86774 152552 86830 152561
rect 86774 152487 86830 152496
rect 86682 151056 86738 151065
rect 86682 150991 86738 151000
rect 86696 104689 86724 150991
rect 86682 104680 86738 104689
rect 86682 104615 86738 104624
rect 86684 104576 86736 104582
rect 86684 104518 86736 104524
rect 86592 104236 86644 104242
rect 86592 104178 86644 104184
rect 86590 101416 86646 101425
rect 86590 101351 86646 101360
rect 86500 99476 86552 99482
rect 86500 99418 86552 99424
rect 86498 99376 86554 99385
rect 86498 99311 86554 99320
rect 86408 97096 86460 97102
rect 86408 97038 86460 97044
rect 86420 96694 86448 97038
rect 86408 96688 86460 96694
rect 86408 96630 86460 96636
rect 86316 94852 86368 94858
rect 86316 94794 86368 94800
rect 86512 94738 86540 99311
rect 86328 94710 86540 94738
rect 85956 94684 86252 94704
rect 86012 94682 86036 94684
rect 86092 94682 86116 94684
rect 86172 94682 86196 94684
rect 86034 94630 86036 94682
rect 86098 94630 86110 94682
rect 86172 94630 86174 94682
rect 86012 94628 86036 94630
rect 86092 94628 86116 94630
rect 86172 94628 86196 94630
rect 85956 94608 86252 94628
rect 85956 93596 86252 93616
rect 86012 93594 86036 93596
rect 86092 93594 86116 93596
rect 86172 93594 86196 93596
rect 86034 93542 86036 93594
rect 86098 93542 86110 93594
rect 86172 93542 86174 93594
rect 86012 93540 86036 93542
rect 86092 93540 86116 93542
rect 86172 93540 86196 93542
rect 85956 93520 86252 93540
rect 85956 92508 86252 92528
rect 86012 92506 86036 92508
rect 86092 92506 86116 92508
rect 86172 92506 86196 92508
rect 86034 92454 86036 92506
rect 86098 92454 86110 92506
rect 86172 92454 86174 92506
rect 86012 92452 86036 92454
rect 86092 92452 86116 92454
rect 86172 92452 86196 92454
rect 85956 92432 86252 92452
rect 85956 91420 86252 91440
rect 86012 91418 86036 91420
rect 86092 91418 86116 91420
rect 86172 91418 86196 91420
rect 86034 91366 86036 91418
rect 86098 91366 86110 91418
rect 86172 91366 86174 91418
rect 86012 91364 86036 91366
rect 86092 91364 86116 91366
rect 86172 91364 86196 91366
rect 85956 91344 86252 91364
rect 85956 90332 86252 90352
rect 86012 90330 86036 90332
rect 86092 90330 86116 90332
rect 86172 90330 86196 90332
rect 86034 90278 86036 90330
rect 86098 90278 86110 90330
rect 86172 90278 86174 90330
rect 86012 90276 86036 90278
rect 86092 90276 86116 90278
rect 86172 90276 86196 90278
rect 85956 90256 86252 90276
rect 85956 89244 86252 89264
rect 86012 89242 86036 89244
rect 86092 89242 86116 89244
rect 86172 89242 86196 89244
rect 86034 89190 86036 89242
rect 86098 89190 86110 89242
rect 86172 89190 86174 89242
rect 86012 89188 86036 89190
rect 86092 89188 86116 89190
rect 86172 89188 86196 89190
rect 85956 89168 86252 89188
rect 85956 88156 86252 88176
rect 86012 88154 86036 88156
rect 86092 88154 86116 88156
rect 86172 88154 86196 88156
rect 86034 88102 86036 88154
rect 86098 88102 86110 88154
rect 86172 88102 86174 88154
rect 86012 88100 86036 88102
rect 86092 88100 86116 88102
rect 86172 88100 86196 88102
rect 85956 88080 86252 88100
rect 85956 87068 86252 87088
rect 86012 87066 86036 87068
rect 86092 87066 86116 87068
rect 86172 87066 86196 87068
rect 86034 87014 86036 87066
rect 86098 87014 86110 87066
rect 86172 87014 86174 87066
rect 86012 87012 86036 87014
rect 86092 87012 86116 87014
rect 86172 87012 86196 87014
rect 85956 86992 86252 87012
rect 85956 85980 86252 86000
rect 86012 85978 86036 85980
rect 86092 85978 86116 85980
rect 86172 85978 86196 85980
rect 86034 85926 86036 85978
rect 86098 85926 86110 85978
rect 86172 85926 86174 85978
rect 86012 85924 86036 85926
rect 86092 85924 86116 85926
rect 86172 85924 86196 85926
rect 85956 85904 86252 85924
rect 85956 84892 86252 84912
rect 86012 84890 86036 84892
rect 86092 84890 86116 84892
rect 86172 84890 86196 84892
rect 86034 84838 86036 84890
rect 86098 84838 86110 84890
rect 86172 84838 86174 84890
rect 86012 84836 86036 84838
rect 86092 84836 86116 84838
rect 86172 84836 86196 84838
rect 85956 84816 86252 84836
rect 85956 83804 86252 83824
rect 86012 83802 86036 83804
rect 86092 83802 86116 83804
rect 86172 83802 86196 83804
rect 86034 83750 86036 83802
rect 86098 83750 86110 83802
rect 86172 83750 86174 83802
rect 86012 83748 86036 83750
rect 86092 83748 86116 83750
rect 86172 83748 86196 83750
rect 85956 83728 86252 83748
rect 85956 82716 86252 82736
rect 86012 82714 86036 82716
rect 86092 82714 86116 82716
rect 86172 82714 86196 82716
rect 86034 82662 86036 82714
rect 86098 82662 86110 82714
rect 86172 82662 86174 82714
rect 86012 82660 86036 82662
rect 86092 82660 86116 82662
rect 86172 82660 86196 82662
rect 85956 82640 86252 82660
rect 85956 81628 86252 81648
rect 86012 81626 86036 81628
rect 86092 81626 86116 81628
rect 86172 81626 86196 81628
rect 86034 81574 86036 81626
rect 86098 81574 86110 81626
rect 86172 81574 86174 81626
rect 86012 81572 86036 81574
rect 86092 81572 86116 81574
rect 86172 81572 86196 81574
rect 85956 81552 86252 81572
rect 85956 80540 86252 80560
rect 86012 80538 86036 80540
rect 86092 80538 86116 80540
rect 86172 80538 86196 80540
rect 86034 80486 86036 80538
rect 86098 80486 86110 80538
rect 86172 80486 86174 80538
rect 86012 80484 86036 80486
rect 86092 80484 86116 80486
rect 86172 80484 86196 80486
rect 85956 80464 86252 80484
rect 85956 79452 86252 79472
rect 86012 79450 86036 79452
rect 86092 79450 86116 79452
rect 86172 79450 86196 79452
rect 86034 79398 86036 79450
rect 86098 79398 86110 79450
rect 86172 79398 86174 79450
rect 86012 79396 86036 79398
rect 86092 79396 86116 79398
rect 86172 79396 86196 79398
rect 85956 79376 86252 79396
rect 85956 78364 86252 78384
rect 86012 78362 86036 78364
rect 86092 78362 86116 78364
rect 86172 78362 86196 78364
rect 86034 78310 86036 78362
rect 86098 78310 86110 78362
rect 86172 78310 86174 78362
rect 86012 78308 86036 78310
rect 86092 78308 86116 78310
rect 86172 78308 86196 78310
rect 85956 78288 86252 78308
rect 85956 77276 86252 77296
rect 86012 77274 86036 77276
rect 86092 77274 86116 77276
rect 86172 77274 86196 77276
rect 86034 77222 86036 77274
rect 86098 77222 86110 77274
rect 86172 77222 86174 77274
rect 86012 77220 86036 77222
rect 86092 77220 86116 77222
rect 86172 77220 86196 77222
rect 85956 77200 86252 77220
rect 85956 76188 86252 76208
rect 86012 76186 86036 76188
rect 86092 76186 86116 76188
rect 86172 76186 86196 76188
rect 86034 76134 86036 76186
rect 86098 76134 86110 76186
rect 86172 76134 86174 76186
rect 86012 76132 86036 76134
rect 86092 76132 86116 76134
rect 86172 76132 86196 76134
rect 85956 76112 86252 76132
rect 85956 75100 86252 75120
rect 86012 75098 86036 75100
rect 86092 75098 86116 75100
rect 86172 75098 86196 75100
rect 86034 75046 86036 75098
rect 86098 75046 86110 75098
rect 86172 75046 86174 75098
rect 86012 75044 86036 75046
rect 86092 75044 86116 75046
rect 86172 75044 86196 75046
rect 85956 75024 86252 75044
rect 85956 74012 86252 74032
rect 86012 74010 86036 74012
rect 86092 74010 86116 74012
rect 86172 74010 86196 74012
rect 86034 73958 86036 74010
rect 86098 73958 86110 74010
rect 86172 73958 86174 74010
rect 86012 73956 86036 73958
rect 86092 73956 86116 73958
rect 86172 73956 86196 73958
rect 85956 73936 86252 73956
rect 85956 72924 86252 72944
rect 86012 72922 86036 72924
rect 86092 72922 86116 72924
rect 86172 72922 86196 72924
rect 86034 72870 86036 72922
rect 86098 72870 86110 72922
rect 86172 72870 86174 72922
rect 86012 72868 86036 72870
rect 86092 72868 86116 72870
rect 86172 72868 86196 72870
rect 85956 72848 86252 72868
rect 85956 71836 86252 71856
rect 86012 71834 86036 71836
rect 86092 71834 86116 71836
rect 86172 71834 86196 71836
rect 86034 71782 86036 71834
rect 86098 71782 86110 71834
rect 86172 71782 86174 71834
rect 86012 71780 86036 71782
rect 86092 71780 86116 71782
rect 86172 71780 86196 71782
rect 85956 71760 86252 71780
rect 85956 70748 86252 70768
rect 86012 70746 86036 70748
rect 86092 70746 86116 70748
rect 86172 70746 86196 70748
rect 86034 70694 86036 70746
rect 86098 70694 86110 70746
rect 86172 70694 86174 70746
rect 86012 70692 86036 70694
rect 86092 70692 86116 70694
rect 86172 70692 86196 70694
rect 85956 70672 86252 70692
rect 85956 69660 86252 69680
rect 86012 69658 86036 69660
rect 86092 69658 86116 69660
rect 86172 69658 86196 69660
rect 86034 69606 86036 69658
rect 86098 69606 86110 69658
rect 86172 69606 86174 69658
rect 86012 69604 86036 69606
rect 86092 69604 86116 69606
rect 86172 69604 86196 69606
rect 85956 69584 86252 69604
rect 85956 68572 86252 68592
rect 86012 68570 86036 68572
rect 86092 68570 86116 68572
rect 86172 68570 86196 68572
rect 86034 68518 86036 68570
rect 86098 68518 86110 68570
rect 86172 68518 86174 68570
rect 86012 68516 86036 68518
rect 86092 68516 86116 68518
rect 86172 68516 86196 68518
rect 85956 68496 86252 68516
rect 85956 67484 86252 67504
rect 86012 67482 86036 67484
rect 86092 67482 86116 67484
rect 86172 67482 86196 67484
rect 86034 67430 86036 67482
rect 86098 67430 86110 67482
rect 86172 67430 86174 67482
rect 86012 67428 86036 67430
rect 86092 67428 86116 67430
rect 86172 67428 86196 67430
rect 85956 67408 86252 67428
rect 85956 66396 86252 66416
rect 86012 66394 86036 66396
rect 86092 66394 86116 66396
rect 86172 66394 86196 66396
rect 86034 66342 86036 66394
rect 86098 66342 86110 66394
rect 86172 66342 86174 66394
rect 86012 66340 86036 66342
rect 86092 66340 86116 66342
rect 86172 66340 86196 66342
rect 85956 66320 86252 66340
rect 85956 65308 86252 65328
rect 86012 65306 86036 65308
rect 86092 65306 86116 65308
rect 86172 65306 86196 65308
rect 86034 65254 86036 65306
rect 86098 65254 86110 65306
rect 86172 65254 86174 65306
rect 86012 65252 86036 65254
rect 86092 65252 86116 65254
rect 86172 65252 86196 65254
rect 85956 65232 86252 65252
rect 85956 64220 86252 64240
rect 86012 64218 86036 64220
rect 86092 64218 86116 64220
rect 86172 64218 86196 64220
rect 86034 64166 86036 64218
rect 86098 64166 86110 64218
rect 86172 64166 86174 64218
rect 86012 64164 86036 64166
rect 86092 64164 86116 64166
rect 86172 64164 86196 64166
rect 85956 64144 86252 64164
rect 85956 63132 86252 63152
rect 86012 63130 86036 63132
rect 86092 63130 86116 63132
rect 86172 63130 86196 63132
rect 86034 63078 86036 63130
rect 86098 63078 86110 63130
rect 86172 63078 86174 63130
rect 86012 63076 86036 63078
rect 86092 63076 86116 63078
rect 86172 63076 86196 63078
rect 85956 63056 86252 63076
rect 85956 62044 86252 62064
rect 86012 62042 86036 62044
rect 86092 62042 86116 62044
rect 86172 62042 86196 62044
rect 86034 61990 86036 62042
rect 86098 61990 86110 62042
rect 86172 61990 86174 62042
rect 86012 61988 86036 61990
rect 86092 61988 86116 61990
rect 86172 61988 86196 61990
rect 85956 61968 86252 61988
rect 85956 60956 86252 60976
rect 86012 60954 86036 60956
rect 86092 60954 86116 60956
rect 86172 60954 86196 60956
rect 86034 60902 86036 60954
rect 86098 60902 86110 60954
rect 86172 60902 86174 60954
rect 86012 60900 86036 60902
rect 86092 60900 86116 60902
rect 86172 60900 86196 60902
rect 85956 60880 86252 60900
rect 85956 59868 86252 59888
rect 86012 59866 86036 59868
rect 86092 59866 86116 59868
rect 86172 59866 86196 59868
rect 86034 59814 86036 59866
rect 86098 59814 86110 59866
rect 86172 59814 86174 59866
rect 86012 59812 86036 59814
rect 86092 59812 86116 59814
rect 86172 59812 86196 59814
rect 85956 59792 86252 59812
rect 85956 58780 86252 58800
rect 86012 58778 86036 58780
rect 86092 58778 86116 58780
rect 86172 58778 86196 58780
rect 86034 58726 86036 58778
rect 86098 58726 86110 58778
rect 86172 58726 86174 58778
rect 86012 58724 86036 58726
rect 86092 58724 86116 58726
rect 86172 58724 86196 58726
rect 85956 58704 86252 58724
rect 85956 57692 86252 57712
rect 86012 57690 86036 57692
rect 86092 57690 86116 57692
rect 86172 57690 86196 57692
rect 86034 57638 86036 57690
rect 86098 57638 86110 57690
rect 86172 57638 86174 57690
rect 86012 57636 86036 57638
rect 86092 57636 86116 57638
rect 86172 57636 86196 57638
rect 85956 57616 86252 57636
rect 85956 56604 86252 56624
rect 86012 56602 86036 56604
rect 86092 56602 86116 56604
rect 86172 56602 86196 56604
rect 86034 56550 86036 56602
rect 86098 56550 86110 56602
rect 86172 56550 86174 56602
rect 86012 56548 86036 56550
rect 86092 56548 86116 56550
rect 86172 56548 86196 56550
rect 85956 56528 86252 56548
rect 85956 55516 86252 55536
rect 86012 55514 86036 55516
rect 86092 55514 86116 55516
rect 86172 55514 86196 55516
rect 86034 55462 86036 55514
rect 86098 55462 86110 55514
rect 86172 55462 86174 55514
rect 86012 55460 86036 55462
rect 86092 55460 86116 55462
rect 86172 55460 86196 55462
rect 85956 55440 86252 55460
rect 85956 54428 86252 54448
rect 86012 54426 86036 54428
rect 86092 54426 86116 54428
rect 86172 54426 86196 54428
rect 86034 54374 86036 54426
rect 86098 54374 86110 54426
rect 86172 54374 86174 54426
rect 86012 54372 86036 54374
rect 86092 54372 86116 54374
rect 86172 54372 86196 54374
rect 85956 54352 86252 54372
rect 85956 53340 86252 53360
rect 86012 53338 86036 53340
rect 86092 53338 86116 53340
rect 86172 53338 86196 53340
rect 86034 53286 86036 53338
rect 86098 53286 86110 53338
rect 86172 53286 86174 53338
rect 86012 53284 86036 53286
rect 86092 53284 86116 53286
rect 86172 53284 86196 53286
rect 85956 53264 86252 53284
rect 85956 52252 86252 52272
rect 86012 52250 86036 52252
rect 86092 52250 86116 52252
rect 86172 52250 86196 52252
rect 86034 52198 86036 52250
rect 86098 52198 86110 52250
rect 86172 52198 86174 52250
rect 86012 52196 86036 52198
rect 86092 52196 86116 52198
rect 86172 52196 86196 52198
rect 85956 52176 86252 52196
rect 85956 51164 86252 51184
rect 86012 51162 86036 51164
rect 86092 51162 86116 51164
rect 86172 51162 86196 51164
rect 86034 51110 86036 51162
rect 86098 51110 86110 51162
rect 86172 51110 86174 51162
rect 86012 51108 86036 51110
rect 86092 51108 86116 51110
rect 86172 51108 86196 51110
rect 85956 51088 86252 51108
rect 85956 50076 86252 50096
rect 86012 50074 86036 50076
rect 86092 50074 86116 50076
rect 86172 50074 86196 50076
rect 86034 50022 86036 50074
rect 86098 50022 86110 50074
rect 86172 50022 86174 50074
rect 86012 50020 86036 50022
rect 86092 50020 86116 50022
rect 86172 50020 86196 50022
rect 85956 50000 86252 50020
rect 85956 48988 86252 49008
rect 86012 48986 86036 48988
rect 86092 48986 86116 48988
rect 86172 48986 86196 48988
rect 86034 48934 86036 48986
rect 86098 48934 86110 48986
rect 86172 48934 86174 48986
rect 86012 48932 86036 48934
rect 86092 48932 86116 48934
rect 86172 48932 86196 48934
rect 85956 48912 86252 48932
rect 85956 47900 86252 47920
rect 86012 47898 86036 47900
rect 86092 47898 86116 47900
rect 86172 47898 86196 47900
rect 86034 47846 86036 47898
rect 86098 47846 86110 47898
rect 86172 47846 86174 47898
rect 86012 47844 86036 47846
rect 86092 47844 86116 47846
rect 86172 47844 86196 47846
rect 85956 47824 86252 47844
rect 85956 46812 86252 46832
rect 86012 46810 86036 46812
rect 86092 46810 86116 46812
rect 86172 46810 86196 46812
rect 86034 46758 86036 46810
rect 86098 46758 86110 46810
rect 86172 46758 86174 46810
rect 86012 46756 86036 46758
rect 86092 46756 86116 46758
rect 86172 46756 86196 46758
rect 85956 46736 86252 46756
rect 85956 45724 86252 45744
rect 86012 45722 86036 45724
rect 86092 45722 86116 45724
rect 86172 45722 86196 45724
rect 86034 45670 86036 45722
rect 86098 45670 86110 45722
rect 86172 45670 86174 45722
rect 86012 45668 86036 45670
rect 86092 45668 86116 45670
rect 86172 45668 86196 45670
rect 85956 45648 86252 45668
rect 85956 44636 86252 44656
rect 86012 44634 86036 44636
rect 86092 44634 86116 44636
rect 86172 44634 86196 44636
rect 86034 44582 86036 44634
rect 86098 44582 86110 44634
rect 86172 44582 86174 44634
rect 86012 44580 86036 44582
rect 86092 44580 86116 44582
rect 86172 44580 86196 44582
rect 85956 44560 86252 44580
rect 85956 43548 86252 43568
rect 86012 43546 86036 43548
rect 86092 43546 86116 43548
rect 86172 43546 86196 43548
rect 86034 43494 86036 43546
rect 86098 43494 86110 43546
rect 86172 43494 86174 43546
rect 86012 43492 86036 43494
rect 86092 43492 86116 43494
rect 86172 43492 86196 43494
rect 85956 43472 86252 43492
rect 85956 42460 86252 42480
rect 86012 42458 86036 42460
rect 86092 42458 86116 42460
rect 86172 42458 86196 42460
rect 86034 42406 86036 42458
rect 86098 42406 86110 42458
rect 86172 42406 86174 42458
rect 86012 42404 86036 42406
rect 86092 42404 86116 42406
rect 86172 42404 86196 42406
rect 85956 42384 86252 42404
rect 85956 41372 86252 41392
rect 86012 41370 86036 41372
rect 86092 41370 86116 41372
rect 86172 41370 86196 41372
rect 86034 41318 86036 41370
rect 86098 41318 86110 41370
rect 86172 41318 86174 41370
rect 86012 41316 86036 41318
rect 86092 41316 86116 41318
rect 86172 41316 86196 41318
rect 85956 41296 86252 41316
rect 85956 40284 86252 40304
rect 86012 40282 86036 40284
rect 86092 40282 86116 40284
rect 86172 40282 86196 40284
rect 86034 40230 86036 40282
rect 86098 40230 86110 40282
rect 86172 40230 86174 40282
rect 86012 40228 86036 40230
rect 86092 40228 86116 40230
rect 86172 40228 86196 40230
rect 85956 40208 86252 40228
rect 85956 39196 86252 39216
rect 86012 39194 86036 39196
rect 86092 39194 86116 39196
rect 86172 39194 86196 39196
rect 86034 39142 86036 39194
rect 86098 39142 86110 39194
rect 86172 39142 86174 39194
rect 86012 39140 86036 39142
rect 86092 39140 86116 39142
rect 86172 39140 86196 39142
rect 85956 39120 86252 39140
rect 85956 38108 86252 38128
rect 86012 38106 86036 38108
rect 86092 38106 86116 38108
rect 86172 38106 86196 38108
rect 86034 38054 86036 38106
rect 86098 38054 86110 38106
rect 86172 38054 86174 38106
rect 86012 38052 86036 38054
rect 86092 38052 86116 38054
rect 86172 38052 86196 38054
rect 85956 38032 86252 38052
rect 85956 37020 86252 37040
rect 86012 37018 86036 37020
rect 86092 37018 86116 37020
rect 86172 37018 86196 37020
rect 86034 36966 86036 37018
rect 86098 36966 86110 37018
rect 86172 36966 86174 37018
rect 86012 36964 86036 36966
rect 86092 36964 86116 36966
rect 86172 36964 86196 36966
rect 85956 36944 86252 36964
rect 85956 35932 86252 35952
rect 86012 35930 86036 35932
rect 86092 35930 86116 35932
rect 86172 35930 86196 35932
rect 86034 35878 86036 35930
rect 86098 35878 86110 35930
rect 86172 35878 86174 35930
rect 86012 35876 86036 35878
rect 86092 35876 86116 35878
rect 86172 35876 86196 35878
rect 85956 35856 86252 35876
rect 85956 34844 86252 34864
rect 86012 34842 86036 34844
rect 86092 34842 86116 34844
rect 86172 34842 86196 34844
rect 86034 34790 86036 34842
rect 86098 34790 86110 34842
rect 86172 34790 86174 34842
rect 86012 34788 86036 34790
rect 86092 34788 86116 34790
rect 86172 34788 86196 34790
rect 85956 34768 86252 34788
rect 85956 33756 86252 33776
rect 86012 33754 86036 33756
rect 86092 33754 86116 33756
rect 86172 33754 86196 33756
rect 86034 33702 86036 33754
rect 86098 33702 86110 33754
rect 86172 33702 86174 33754
rect 86012 33700 86036 33702
rect 86092 33700 86116 33702
rect 86172 33700 86196 33702
rect 85956 33680 86252 33700
rect 85956 32668 86252 32688
rect 86012 32666 86036 32668
rect 86092 32666 86116 32668
rect 86172 32666 86196 32668
rect 86034 32614 86036 32666
rect 86098 32614 86110 32666
rect 86172 32614 86174 32666
rect 86012 32612 86036 32614
rect 86092 32612 86116 32614
rect 86172 32612 86196 32614
rect 85956 32592 86252 32612
rect 85956 31580 86252 31600
rect 86012 31578 86036 31580
rect 86092 31578 86116 31580
rect 86172 31578 86196 31580
rect 86034 31526 86036 31578
rect 86098 31526 86110 31578
rect 86172 31526 86174 31578
rect 86012 31524 86036 31526
rect 86092 31524 86116 31526
rect 86172 31524 86196 31526
rect 85956 31504 86252 31524
rect 85956 30492 86252 30512
rect 86012 30490 86036 30492
rect 86092 30490 86116 30492
rect 86172 30490 86196 30492
rect 86034 30438 86036 30490
rect 86098 30438 86110 30490
rect 86172 30438 86174 30490
rect 86012 30436 86036 30438
rect 86092 30436 86116 30438
rect 86172 30436 86196 30438
rect 85956 30416 86252 30436
rect 85956 29404 86252 29424
rect 86012 29402 86036 29404
rect 86092 29402 86116 29404
rect 86172 29402 86196 29404
rect 86034 29350 86036 29402
rect 86098 29350 86110 29402
rect 86172 29350 86174 29402
rect 86012 29348 86036 29350
rect 86092 29348 86116 29350
rect 86172 29348 86196 29350
rect 85956 29328 86252 29348
rect 85956 28316 86252 28336
rect 86012 28314 86036 28316
rect 86092 28314 86116 28316
rect 86172 28314 86196 28316
rect 86034 28262 86036 28314
rect 86098 28262 86110 28314
rect 86172 28262 86174 28314
rect 86012 28260 86036 28262
rect 86092 28260 86116 28262
rect 86172 28260 86196 28262
rect 85956 28240 86252 28260
rect 85956 27228 86252 27248
rect 86012 27226 86036 27228
rect 86092 27226 86116 27228
rect 86172 27226 86196 27228
rect 86034 27174 86036 27226
rect 86098 27174 86110 27226
rect 86172 27174 86174 27226
rect 86012 27172 86036 27174
rect 86092 27172 86116 27174
rect 86172 27172 86196 27174
rect 85956 27152 86252 27172
rect 86328 26586 86356 94710
rect 86604 94058 86632 101351
rect 86696 99958 86724 104518
rect 86684 99952 86736 99958
rect 86684 99894 86736 99900
rect 86682 99512 86738 99521
rect 86682 99447 86738 99456
rect 86512 94030 86632 94058
rect 86408 90772 86460 90778
rect 86408 90714 86460 90720
rect 86420 27606 86448 90714
rect 86512 29306 86540 94030
rect 86592 93968 86644 93974
rect 86592 93910 86644 93916
rect 86604 32026 86632 93910
rect 86696 90778 86724 99447
rect 86788 97238 86816 152487
rect 86958 148880 87014 148889
rect 86958 148815 87014 148824
rect 86866 134192 86922 134201
rect 86866 134127 86922 134136
rect 86880 104378 86908 134127
rect 86868 104372 86920 104378
rect 86868 104314 86920 104320
rect 86868 104236 86920 104242
rect 86868 104178 86920 104184
rect 86880 99793 86908 104178
rect 86866 99784 86922 99793
rect 86866 99719 86922 99728
rect 86868 99680 86920 99686
rect 86868 99622 86920 99628
rect 86776 97232 86828 97238
rect 86776 97174 86828 97180
rect 86776 97096 86828 97102
rect 86776 97038 86828 97044
rect 86788 95577 86816 97038
rect 86774 95568 86830 95577
rect 86774 95503 86830 95512
rect 86880 94994 86908 99622
rect 86972 98122 87000 148815
rect 87050 146568 87106 146577
rect 87050 146503 87106 146512
rect 86960 98116 87012 98122
rect 86960 98058 87012 98064
rect 86958 97744 87014 97753
rect 86958 97679 87014 97688
rect 86972 97306 87000 97679
rect 86960 97300 87012 97306
rect 86960 97242 87012 97248
rect 86960 97164 87012 97170
rect 86960 97106 87012 97112
rect 86972 96665 87000 97106
rect 86958 96656 87014 96665
rect 87064 96626 87092 146503
rect 87156 104281 87184 154799
rect 87234 149968 87290 149977
rect 87234 149903 87290 149912
rect 87248 122369 87276 149903
rect 87234 122360 87290 122369
rect 87234 122295 87290 122304
rect 87236 122188 87288 122194
rect 87236 122130 87288 122136
rect 87248 118697 87276 122130
rect 87234 118688 87290 118697
rect 87234 118623 87290 118632
rect 87234 118552 87290 118561
rect 87234 118487 87290 118496
rect 87248 109177 87276 118487
rect 87234 109168 87290 109177
rect 87234 109103 87290 109112
rect 87340 109034 87368 156975
rect 87248 109006 87368 109034
rect 87248 108633 87276 109006
rect 87326 108760 87382 108769
rect 87326 108695 87382 108704
rect 87234 108624 87290 108633
rect 87234 108559 87290 108568
rect 87236 108520 87288 108526
rect 87236 108462 87288 108468
rect 87142 104272 87198 104281
rect 87142 104207 87198 104216
rect 87144 104168 87196 104174
rect 87144 104110 87196 104116
rect 87156 99498 87184 104110
rect 87248 99958 87276 108462
rect 87340 104378 87368 108695
rect 87328 104372 87380 104378
rect 87328 104314 87380 104320
rect 87326 104272 87382 104281
rect 87326 104207 87382 104216
rect 87236 99952 87288 99958
rect 87236 99894 87288 99900
rect 87156 99470 87276 99498
rect 87142 99388 87198 99397
rect 87142 99323 87198 99332
rect 87156 97102 87184 99323
rect 87248 98190 87276 99470
rect 87236 98184 87288 98190
rect 87236 98126 87288 98132
rect 87234 97880 87290 97889
rect 87234 97815 87290 97824
rect 87144 97096 87196 97102
rect 87144 97038 87196 97044
rect 86958 96591 87014 96600
rect 87052 96620 87104 96626
rect 87052 96562 87104 96568
rect 87248 96014 87276 97815
rect 87340 96393 87368 104207
rect 87432 99346 87460 159695
rect 87420 99340 87472 99346
rect 87420 99282 87472 99288
rect 87524 99278 87552 165679
rect 87616 108594 87644 173159
rect 87694 171728 87750 171737
rect 87694 171663 87750 171672
rect 87604 108588 87656 108594
rect 87604 108530 87656 108536
rect 87604 108452 87656 108458
rect 87604 108394 87656 108400
rect 87616 99890 87644 108394
rect 87604 99884 87656 99890
rect 87604 99826 87656 99832
rect 87604 99748 87656 99754
rect 87604 99690 87656 99696
rect 87512 99272 87564 99278
rect 87512 99214 87564 99220
rect 87420 99204 87472 99210
rect 87420 99146 87472 99152
rect 87326 96384 87382 96393
rect 87326 96319 87382 96328
rect 87236 96008 87288 96014
rect 87236 95950 87288 95956
rect 86960 95940 87012 95946
rect 86960 95882 87012 95888
rect 86972 95441 87000 95882
rect 86958 95432 87014 95441
rect 86958 95367 87014 95376
rect 87432 95334 87460 99146
rect 87512 99136 87564 99142
rect 87512 99078 87564 99084
rect 87524 95674 87552 99078
rect 87616 98938 87644 99690
rect 87708 98938 87736 171663
rect 87800 104378 87828 177647
rect 89956 177372 90252 177392
rect 90012 177370 90036 177372
rect 90092 177370 90116 177372
rect 90172 177370 90196 177372
rect 90034 177318 90036 177370
rect 90098 177318 90110 177370
rect 90172 177318 90174 177370
rect 90012 177316 90036 177318
rect 90092 177316 90116 177318
rect 90172 177316 90196 177318
rect 89956 177296 90252 177316
rect 87956 176828 88252 176848
rect 88012 176826 88036 176828
rect 88092 176826 88116 176828
rect 88172 176826 88196 176828
rect 88034 176774 88036 176826
rect 88098 176774 88110 176826
rect 88172 176774 88174 176826
rect 88012 176772 88036 176774
rect 88092 176772 88116 176774
rect 88172 176772 88196 176774
rect 87956 176752 88252 176772
rect 89956 176284 90252 176304
rect 90012 176282 90036 176284
rect 90092 176282 90116 176284
rect 90172 176282 90196 176284
rect 90034 176230 90036 176282
rect 90098 176230 90110 176282
rect 90172 176230 90174 176282
rect 90012 176228 90036 176230
rect 90092 176228 90116 176230
rect 90172 176228 90196 176230
rect 89956 176208 90252 176228
rect 87956 175740 88252 175760
rect 88012 175738 88036 175740
rect 88092 175738 88116 175740
rect 88172 175738 88196 175740
rect 88034 175686 88036 175738
rect 88098 175686 88110 175738
rect 88172 175686 88174 175738
rect 88012 175684 88036 175686
rect 88092 175684 88116 175686
rect 88172 175684 88196 175686
rect 87956 175664 88252 175684
rect 89956 175196 90252 175216
rect 90012 175194 90036 175196
rect 90092 175194 90116 175196
rect 90172 175194 90196 175196
rect 90034 175142 90036 175194
rect 90098 175142 90110 175194
rect 90172 175142 90174 175194
rect 90012 175140 90036 175142
rect 90092 175140 90116 175142
rect 90172 175140 90196 175142
rect 89956 175120 90252 175140
rect 87956 174652 88252 174672
rect 88012 174650 88036 174652
rect 88092 174650 88116 174652
rect 88172 174650 88196 174652
rect 88034 174598 88036 174650
rect 88098 174598 88110 174650
rect 88172 174598 88174 174650
rect 88012 174596 88036 174598
rect 88092 174596 88116 174598
rect 88172 174596 88196 174598
rect 87956 174576 88252 174596
rect 89956 174108 90252 174128
rect 90012 174106 90036 174108
rect 90092 174106 90116 174108
rect 90172 174106 90196 174108
rect 90034 174054 90036 174106
rect 90098 174054 90110 174106
rect 90172 174054 90174 174106
rect 90012 174052 90036 174054
rect 90092 174052 90116 174054
rect 90172 174052 90196 174054
rect 89956 174032 90252 174052
rect 87956 173564 88252 173584
rect 88012 173562 88036 173564
rect 88092 173562 88116 173564
rect 88172 173562 88196 173564
rect 88034 173510 88036 173562
rect 88098 173510 88110 173562
rect 88172 173510 88174 173562
rect 88012 173508 88036 173510
rect 88092 173508 88116 173510
rect 88172 173508 88196 173510
rect 87956 173488 88252 173508
rect 89956 173020 90252 173040
rect 90012 173018 90036 173020
rect 90092 173018 90116 173020
rect 90172 173018 90196 173020
rect 90034 172966 90036 173018
rect 90098 172966 90110 173018
rect 90172 172966 90174 173018
rect 90012 172964 90036 172966
rect 90092 172964 90116 172966
rect 90172 172964 90196 172966
rect 89956 172944 90252 172964
rect 87956 172476 88252 172496
rect 88012 172474 88036 172476
rect 88092 172474 88116 172476
rect 88172 172474 88196 172476
rect 88034 172422 88036 172474
rect 88098 172422 88110 172474
rect 88172 172422 88174 172474
rect 88012 172420 88036 172422
rect 88092 172420 88116 172422
rect 88172 172420 88196 172422
rect 87956 172400 88252 172420
rect 89956 171932 90252 171952
rect 90012 171930 90036 171932
rect 90092 171930 90116 171932
rect 90172 171930 90196 171932
rect 90034 171878 90036 171930
rect 90098 171878 90110 171930
rect 90172 171878 90174 171930
rect 90012 171876 90036 171878
rect 90092 171876 90116 171878
rect 90172 171876 90196 171878
rect 89956 171856 90252 171876
rect 87956 171388 88252 171408
rect 88012 171386 88036 171388
rect 88092 171386 88116 171388
rect 88172 171386 88196 171388
rect 88034 171334 88036 171386
rect 88098 171334 88110 171386
rect 88172 171334 88174 171386
rect 88012 171332 88036 171334
rect 88092 171332 88116 171334
rect 88172 171332 88196 171334
rect 87956 171312 88252 171332
rect 89956 170844 90252 170864
rect 90012 170842 90036 170844
rect 90092 170842 90116 170844
rect 90172 170842 90196 170844
rect 90034 170790 90036 170842
rect 90098 170790 90110 170842
rect 90172 170790 90174 170842
rect 90012 170788 90036 170790
rect 90092 170788 90116 170790
rect 90172 170788 90196 170790
rect 89956 170768 90252 170788
rect 87956 170300 88252 170320
rect 88012 170298 88036 170300
rect 88092 170298 88116 170300
rect 88172 170298 88196 170300
rect 88034 170246 88036 170298
rect 88098 170246 88110 170298
rect 88172 170246 88174 170298
rect 88012 170244 88036 170246
rect 88092 170244 88116 170246
rect 88172 170244 88196 170246
rect 87956 170224 88252 170244
rect 89956 169756 90252 169776
rect 90012 169754 90036 169756
rect 90092 169754 90116 169756
rect 90172 169754 90196 169756
rect 90034 169702 90036 169754
rect 90098 169702 90110 169754
rect 90172 169702 90174 169754
rect 90012 169700 90036 169702
rect 90092 169700 90116 169702
rect 90172 169700 90196 169702
rect 89956 169680 90252 169700
rect 87878 169552 87934 169561
rect 87878 169487 87934 169496
rect 87892 168434 87920 169487
rect 87956 169212 88252 169232
rect 88012 169210 88036 169212
rect 88092 169210 88116 169212
rect 88172 169210 88196 169212
rect 88034 169158 88036 169210
rect 88098 169158 88110 169210
rect 88172 169158 88174 169210
rect 88012 169156 88036 169158
rect 88092 169156 88116 169158
rect 88172 169156 88196 169158
rect 87956 169136 88252 169156
rect 89956 168668 90252 168688
rect 90012 168666 90036 168668
rect 90092 168666 90116 168668
rect 90172 168666 90196 168668
rect 90034 168614 90036 168666
rect 90098 168614 90110 168666
rect 90172 168614 90174 168666
rect 90012 168612 90036 168614
rect 90092 168612 90116 168614
rect 90172 168612 90196 168614
rect 89956 168592 90252 168612
rect 87880 168428 87932 168434
rect 87880 168370 87932 168376
rect 87956 168124 88252 168144
rect 88012 168122 88036 168124
rect 88092 168122 88116 168124
rect 88172 168122 88196 168124
rect 88034 168070 88036 168122
rect 88098 168070 88110 168122
rect 88172 168070 88174 168122
rect 88012 168068 88036 168070
rect 88092 168068 88116 168070
rect 88172 168068 88196 168070
rect 87956 168048 88252 168068
rect 89956 167580 90252 167600
rect 90012 167578 90036 167580
rect 90092 167578 90116 167580
rect 90172 167578 90196 167580
rect 90034 167526 90036 167578
rect 90098 167526 90110 167578
rect 90172 167526 90174 167578
rect 90012 167524 90036 167526
rect 90092 167524 90116 167526
rect 90172 167524 90196 167526
rect 89956 167504 90252 167524
rect 87956 167036 88252 167056
rect 88012 167034 88036 167036
rect 88092 167034 88116 167036
rect 88172 167034 88196 167036
rect 88034 166982 88036 167034
rect 88098 166982 88110 167034
rect 88172 166982 88174 167034
rect 88012 166980 88036 166982
rect 88092 166980 88116 166982
rect 88172 166980 88196 166982
rect 87956 166960 88252 166980
rect 89956 166492 90252 166512
rect 90012 166490 90036 166492
rect 90092 166490 90116 166492
rect 90172 166490 90196 166492
rect 90034 166438 90036 166490
rect 90098 166438 90110 166490
rect 90172 166438 90174 166490
rect 90012 166436 90036 166438
rect 90092 166436 90116 166438
rect 90172 166436 90196 166438
rect 89956 166416 90252 166436
rect 87956 165948 88252 165968
rect 88012 165946 88036 165948
rect 88092 165946 88116 165948
rect 88172 165946 88196 165948
rect 88034 165894 88036 165946
rect 88098 165894 88110 165946
rect 88172 165894 88174 165946
rect 88012 165892 88036 165894
rect 88092 165892 88116 165894
rect 88172 165892 88196 165894
rect 87956 165872 88252 165892
rect 89956 165404 90252 165424
rect 90012 165402 90036 165404
rect 90092 165402 90116 165404
rect 90172 165402 90196 165404
rect 90034 165350 90036 165402
rect 90098 165350 90110 165402
rect 90172 165350 90174 165402
rect 90012 165348 90036 165350
rect 90092 165348 90116 165350
rect 90172 165348 90196 165350
rect 89956 165328 90252 165348
rect 87956 164860 88252 164880
rect 88012 164858 88036 164860
rect 88092 164858 88116 164860
rect 88172 164858 88196 164860
rect 88034 164806 88036 164858
rect 88098 164806 88110 164858
rect 88172 164806 88174 164858
rect 88012 164804 88036 164806
rect 88092 164804 88116 164806
rect 88172 164804 88196 164806
rect 87956 164784 88252 164804
rect 87878 164656 87934 164665
rect 87878 164591 87934 164600
rect 87892 164422 87920 164591
rect 87880 164416 87932 164422
rect 87880 164358 87932 164364
rect 89956 164316 90252 164336
rect 90012 164314 90036 164316
rect 90092 164314 90116 164316
rect 90172 164314 90196 164316
rect 90034 164262 90036 164314
rect 90098 164262 90110 164314
rect 90172 164262 90174 164314
rect 90012 164260 90036 164262
rect 90092 164260 90116 164262
rect 90172 164260 90196 164262
rect 89956 164240 90252 164260
rect 87956 163772 88252 163792
rect 88012 163770 88036 163772
rect 88092 163770 88116 163772
rect 88172 163770 88196 163772
rect 88034 163718 88036 163770
rect 88098 163718 88110 163770
rect 88172 163718 88174 163770
rect 88012 163716 88036 163718
rect 88092 163716 88116 163718
rect 88172 163716 88196 163718
rect 87956 163696 88252 163716
rect 87878 163432 87934 163441
rect 87878 163367 87934 163376
rect 87892 162926 87920 163367
rect 89956 163228 90252 163248
rect 90012 163226 90036 163228
rect 90092 163226 90116 163228
rect 90172 163226 90196 163228
rect 90034 163174 90036 163226
rect 90098 163174 90110 163226
rect 90172 163174 90174 163226
rect 90012 163172 90036 163174
rect 90092 163172 90116 163174
rect 90172 163172 90196 163174
rect 89956 163152 90252 163172
rect 87880 162920 87932 162926
rect 87880 162862 87932 162868
rect 87956 162684 88252 162704
rect 88012 162682 88036 162684
rect 88092 162682 88116 162684
rect 88172 162682 88196 162684
rect 88034 162630 88036 162682
rect 88098 162630 88110 162682
rect 88172 162630 88174 162682
rect 88012 162628 88036 162630
rect 88092 162628 88116 162630
rect 88172 162628 88196 162630
rect 87956 162608 88252 162628
rect 89956 162140 90252 162160
rect 90012 162138 90036 162140
rect 90092 162138 90116 162140
rect 90172 162138 90196 162140
rect 90034 162086 90036 162138
rect 90098 162086 90110 162138
rect 90172 162086 90174 162138
rect 90012 162084 90036 162086
rect 90092 162084 90116 162086
rect 90172 162084 90196 162086
rect 89956 162064 90252 162084
rect 87956 161596 88252 161616
rect 88012 161594 88036 161596
rect 88092 161594 88116 161596
rect 88172 161594 88196 161596
rect 88034 161542 88036 161594
rect 88098 161542 88110 161594
rect 88172 161542 88174 161594
rect 88012 161540 88036 161542
rect 88092 161540 88116 161542
rect 88172 161540 88196 161542
rect 87956 161520 88252 161540
rect 89956 161052 90252 161072
rect 90012 161050 90036 161052
rect 90092 161050 90116 161052
rect 90172 161050 90196 161052
rect 90034 160998 90036 161050
rect 90098 160998 90110 161050
rect 90172 160998 90174 161050
rect 90012 160996 90036 160998
rect 90092 160996 90116 160998
rect 90172 160996 90196 160998
rect 89956 160976 90252 160996
rect 87878 160848 87934 160857
rect 87878 160783 87934 160792
rect 87892 122194 87920 160783
rect 87956 160508 88252 160528
rect 88012 160506 88036 160508
rect 88092 160506 88116 160508
rect 88172 160506 88196 160508
rect 88034 160454 88036 160506
rect 88098 160454 88110 160506
rect 88172 160454 88174 160506
rect 88012 160452 88036 160454
rect 88092 160452 88116 160454
rect 88172 160452 88196 160454
rect 87956 160432 88252 160452
rect 89956 159964 90252 159984
rect 90012 159962 90036 159964
rect 90092 159962 90116 159964
rect 90172 159962 90196 159964
rect 90034 159910 90036 159962
rect 90098 159910 90110 159962
rect 90172 159910 90174 159962
rect 90012 159908 90036 159910
rect 90092 159908 90116 159910
rect 90172 159908 90196 159910
rect 89956 159888 90252 159908
rect 87956 159420 88252 159440
rect 88012 159418 88036 159420
rect 88092 159418 88116 159420
rect 88172 159418 88196 159420
rect 88034 159366 88036 159418
rect 88098 159366 88110 159418
rect 88172 159366 88174 159418
rect 88012 159364 88036 159366
rect 88092 159364 88116 159366
rect 88172 159364 88196 159366
rect 87956 159344 88252 159364
rect 89956 158876 90252 158896
rect 90012 158874 90036 158876
rect 90092 158874 90116 158876
rect 90172 158874 90196 158876
rect 90034 158822 90036 158874
rect 90098 158822 90110 158874
rect 90172 158822 90174 158874
rect 90012 158820 90036 158822
rect 90092 158820 90116 158822
rect 90172 158820 90196 158822
rect 89956 158800 90252 158820
rect 87956 158332 88252 158352
rect 88012 158330 88036 158332
rect 88092 158330 88116 158332
rect 88172 158330 88196 158332
rect 88034 158278 88036 158330
rect 88098 158278 88110 158330
rect 88172 158278 88174 158330
rect 88012 158276 88036 158278
rect 88092 158276 88116 158278
rect 88172 158276 88196 158278
rect 87956 158256 88252 158276
rect 89956 157788 90252 157808
rect 90012 157786 90036 157788
rect 90092 157786 90116 157788
rect 90172 157786 90196 157788
rect 90034 157734 90036 157786
rect 90098 157734 90110 157786
rect 90172 157734 90174 157786
rect 90012 157732 90036 157734
rect 90092 157732 90116 157734
rect 90172 157732 90196 157734
rect 89956 157712 90252 157732
rect 87956 157244 88252 157264
rect 88012 157242 88036 157244
rect 88092 157242 88116 157244
rect 88172 157242 88196 157244
rect 88034 157190 88036 157242
rect 88098 157190 88110 157242
rect 88172 157190 88174 157242
rect 88012 157188 88036 157190
rect 88092 157188 88116 157190
rect 88172 157188 88196 157190
rect 87956 157168 88252 157188
rect 89956 156700 90252 156720
rect 90012 156698 90036 156700
rect 90092 156698 90116 156700
rect 90172 156698 90196 156700
rect 90034 156646 90036 156698
rect 90098 156646 90110 156698
rect 90172 156646 90174 156698
rect 90012 156644 90036 156646
rect 90092 156644 90116 156646
rect 90172 156644 90196 156646
rect 89956 156624 90252 156644
rect 87956 156156 88252 156176
rect 88012 156154 88036 156156
rect 88092 156154 88116 156156
rect 88172 156154 88196 156156
rect 88034 156102 88036 156154
rect 88098 156102 88110 156154
rect 88172 156102 88174 156154
rect 88012 156100 88036 156102
rect 88092 156100 88116 156102
rect 88172 156100 88196 156102
rect 87956 156080 88252 156100
rect 89956 155612 90252 155632
rect 90012 155610 90036 155612
rect 90092 155610 90116 155612
rect 90172 155610 90196 155612
rect 90034 155558 90036 155610
rect 90098 155558 90110 155610
rect 90172 155558 90174 155610
rect 90012 155556 90036 155558
rect 90092 155556 90116 155558
rect 90172 155556 90196 155558
rect 89956 155536 90252 155556
rect 87956 155068 88252 155088
rect 88012 155066 88036 155068
rect 88092 155066 88116 155068
rect 88172 155066 88196 155068
rect 88034 155014 88036 155066
rect 88098 155014 88110 155066
rect 88172 155014 88174 155066
rect 88012 155012 88036 155014
rect 88092 155012 88116 155014
rect 88172 155012 88196 155014
rect 87956 154992 88252 155012
rect 89956 154524 90252 154544
rect 90012 154522 90036 154524
rect 90092 154522 90116 154524
rect 90172 154522 90196 154524
rect 90034 154470 90036 154522
rect 90098 154470 90110 154522
rect 90172 154470 90174 154522
rect 90012 154468 90036 154470
rect 90092 154468 90116 154470
rect 90172 154468 90196 154470
rect 89956 154448 90252 154468
rect 87956 153980 88252 154000
rect 88012 153978 88036 153980
rect 88092 153978 88116 153980
rect 88172 153978 88196 153980
rect 88034 153926 88036 153978
rect 88098 153926 88110 153978
rect 88172 153926 88174 153978
rect 88012 153924 88036 153926
rect 88092 153924 88116 153926
rect 88172 153924 88196 153926
rect 87956 153904 88252 153924
rect 89956 153436 90252 153456
rect 90012 153434 90036 153436
rect 90092 153434 90116 153436
rect 90172 153434 90196 153436
rect 90034 153382 90036 153434
rect 90098 153382 90110 153434
rect 90172 153382 90174 153434
rect 90012 153380 90036 153382
rect 90092 153380 90116 153382
rect 90172 153380 90196 153382
rect 89956 153360 90252 153380
rect 87956 152892 88252 152912
rect 88012 152890 88036 152892
rect 88092 152890 88116 152892
rect 88172 152890 88196 152892
rect 88034 152838 88036 152890
rect 88098 152838 88110 152890
rect 88172 152838 88174 152890
rect 88012 152836 88036 152838
rect 88092 152836 88116 152838
rect 88172 152836 88196 152838
rect 87956 152816 88252 152836
rect 89956 152348 90252 152368
rect 90012 152346 90036 152348
rect 90092 152346 90116 152348
rect 90172 152346 90196 152348
rect 90034 152294 90036 152346
rect 90098 152294 90110 152346
rect 90172 152294 90174 152346
rect 90012 152292 90036 152294
rect 90092 152292 90116 152294
rect 90172 152292 90196 152294
rect 89956 152272 90252 152292
rect 87956 151804 88252 151824
rect 88012 151802 88036 151804
rect 88092 151802 88116 151804
rect 88172 151802 88196 151804
rect 88034 151750 88036 151802
rect 88098 151750 88110 151802
rect 88172 151750 88174 151802
rect 88012 151748 88036 151750
rect 88092 151748 88116 151750
rect 88172 151748 88196 151750
rect 87956 151728 88252 151748
rect 89956 151260 90252 151280
rect 90012 151258 90036 151260
rect 90092 151258 90116 151260
rect 90172 151258 90196 151260
rect 90034 151206 90036 151258
rect 90098 151206 90110 151258
rect 90172 151206 90174 151258
rect 90012 151204 90036 151206
rect 90092 151204 90116 151206
rect 90172 151204 90196 151206
rect 89956 151184 90252 151204
rect 87956 150716 88252 150736
rect 88012 150714 88036 150716
rect 88092 150714 88116 150716
rect 88172 150714 88196 150716
rect 88034 150662 88036 150714
rect 88098 150662 88110 150714
rect 88172 150662 88174 150714
rect 88012 150660 88036 150662
rect 88092 150660 88116 150662
rect 88172 150660 88196 150662
rect 87956 150640 88252 150660
rect 89956 150172 90252 150192
rect 90012 150170 90036 150172
rect 90092 150170 90116 150172
rect 90172 150170 90196 150172
rect 90034 150118 90036 150170
rect 90098 150118 90110 150170
rect 90172 150118 90174 150170
rect 90012 150116 90036 150118
rect 90092 150116 90116 150118
rect 90172 150116 90196 150118
rect 89956 150096 90252 150116
rect 87956 149628 88252 149648
rect 88012 149626 88036 149628
rect 88092 149626 88116 149628
rect 88172 149626 88196 149628
rect 88034 149574 88036 149626
rect 88098 149574 88110 149626
rect 88172 149574 88174 149626
rect 88012 149572 88036 149574
rect 88092 149572 88116 149574
rect 88172 149572 88196 149574
rect 87956 149552 88252 149572
rect 89956 149084 90252 149104
rect 90012 149082 90036 149084
rect 90092 149082 90116 149084
rect 90172 149082 90196 149084
rect 90034 149030 90036 149082
rect 90098 149030 90110 149082
rect 90172 149030 90174 149082
rect 90012 149028 90036 149030
rect 90092 149028 90116 149030
rect 90172 149028 90196 149030
rect 89956 149008 90252 149028
rect 87956 148540 88252 148560
rect 88012 148538 88036 148540
rect 88092 148538 88116 148540
rect 88172 148538 88196 148540
rect 88034 148486 88036 148538
rect 88098 148486 88110 148538
rect 88172 148486 88174 148538
rect 88012 148484 88036 148486
rect 88092 148484 88116 148486
rect 88172 148484 88196 148486
rect 87956 148464 88252 148484
rect 89956 147996 90252 148016
rect 90012 147994 90036 147996
rect 90092 147994 90116 147996
rect 90172 147994 90196 147996
rect 90034 147942 90036 147994
rect 90098 147942 90110 147994
rect 90172 147942 90174 147994
rect 90012 147940 90036 147942
rect 90092 147940 90116 147942
rect 90172 147940 90196 147942
rect 89956 147920 90252 147940
rect 87956 147452 88252 147472
rect 88012 147450 88036 147452
rect 88092 147450 88116 147452
rect 88172 147450 88196 147452
rect 88034 147398 88036 147450
rect 88098 147398 88110 147450
rect 88172 147398 88174 147450
rect 88012 147396 88036 147398
rect 88092 147396 88116 147398
rect 88172 147396 88196 147398
rect 87956 147376 88252 147396
rect 89956 146908 90252 146928
rect 90012 146906 90036 146908
rect 90092 146906 90116 146908
rect 90172 146906 90196 146908
rect 90034 146854 90036 146906
rect 90098 146854 90110 146906
rect 90172 146854 90174 146906
rect 90012 146852 90036 146854
rect 90092 146852 90116 146854
rect 90172 146852 90196 146854
rect 89956 146832 90252 146852
rect 87956 146364 88252 146384
rect 88012 146362 88036 146364
rect 88092 146362 88116 146364
rect 88172 146362 88196 146364
rect 88034 146310 88036 146362
rect 88098 146310 88110 146362
rect 88172 146310 88174 146362
rect 88012 146308 88036 146310
rect 88092 146308 88116 146310
rect 88172 146308 88196 146310
rect 87956 146288 88252 146308
rect 89956 145820 90252 145840
rect 90012 145818 90036 145820
rect 90092 145818 90116 145820
rect 90172 145818 90196 145820
rect 90034 145766 90036 145818
rect 90098 145766 90110 145818
rect 90172 145766 90174 145818
rect 90012 145764 90036 145766
rect 90092 145764 90116 145766
rect 90172 145764 90196 145766
rect 89956 145744 90252 145764
rect 87956 145276 88252 145296
rect 88012 145274 88036 145276
rect 88092 145274 88116 145276
rect 88172 145274 88196 145276
rect 88034 145222 88036 145274
rect 88098 145222 88110 145274
rect 88172 145222 88174 145274
rect 88012 145220 88036 145222
rect 88092 145220 88116 145222
rect 88172 145220 88196 145222
rect 87956 145200 88252 145220
rect 87970 145072 88026 145081
rect 87970 145007 88026 145016
rect 87984 144974 88012 145007
rect 87972 144968 88024 144974
rect 87972 144910 88024 144916
rect 89956 144732 90252 144752
rect 90012 144730 90036 144732
rect 90092 144730 90116 144732
rect 90172 144730 90196 144732
rect 90034 144678 90036 144730
rect 90098 144678 90110 144730
rect 90172 144678 90174 144730
rect 90012 144676 90036 144678
rect 90092 144676 90116 144678
rect 90172 144676 90196 144678
rect 89956 144656 90252 144676
rect 87956 144188 88252 144208
rect 88012 144186 88036 144188
rect 88092 144186 88116 144188
rect 88172 144186 88196 144188
rect 88034 144134 88036 144186
rect 88098 144134 88110 144186
rect 88172 144134 88174 144186
rect 88012 144132 88036 144134
rect 88092 144132 88116 144134
rect 88172 144132 88196 144134
rect 87956 144112 88252 144132
rect 88062 143984 88118 143993
rect 88062 143919 88118 143928
rect 88076 143750 88104 143919
rect 88064 143744 88116 143750
rect 88064 143686 88116 143692
rect 89956 143644 90252 143664
rect 90012 143642 90036 143644
rect 90092 143642 90116 143644
rect 90172 143642 90196 143644
rect 90034 143590 90036 143642
rect 90098 143590 90110 143642
rect 90172 143590 90174 143642
rect 90012 143588 90036 143590
rect 90092 143588 90116 143590
rect 90172 143588 90196 143590
rect 89956 143568 90252 143588
rect 87956 143100 88252 143120
rect 88012 143098 88036 143100
rect 88092 143098 88116 143100
rect 88172 143098 88196 143100
rect 88034 143046 88036 143098
rect 88098 143046 88110 143098
rect 88172 143046 88174 143098
rect 88012 143044 88036 143046
rect 88092 143044 88116 143046
rect 88172 143044 88196 143046
rect 87956 143024 88252 143044
rect 87970 142760 88026 142769
rect 87970 142695 88026 142704
rect 87984 142458 88012 142695
rect 89956 142556 90252 142576
rect 90012 142554 90036 142556
rect 90092 142554 90116 142556
rect 90172 142554 90196 142556
rect 90034 142502 90036 142554
rect 90098 142502 90110 142554
rect 90172 142502 90174 142554
rect 90012 142500 90036 142502
rect 90092 142500 90116 142502
rect 90172 142500 90196 142502
rect 89956 142480 90252 142500
rect 87972 142452 88024 142458
rect 87972 142394 88024 142400
rect 87956 142012 88252 142032
rect 88012 142010 88036 142012
rect 88092 142010 88116 142012
rect 88172 142010 88196 142012
rect 88034 141958 88036 142010
rect 88098 141958 88110 142010
rect 88172 141958 88174 142010
rect 88012 141956 88036 141958
rect 88092 141956 88116 141958
rect 88172 141956 88196 141958
rect 87956 141936 88252 141956
rect 89956 141468 90252 141488
rect 90012 141466 90036 141468
rect 90092 141466 90116 141468
rect 90172 141466 90196 141468
rect 90034 141414 90036 141466
rect 90098 141414 90110 141466
rect 90172 141414 90174 141466
rect 90012 141412 90036 141414
rect 90092 141412 90116 141414
rect 90172 141412 90196 141414
rect 89956 141392 90252 141412
rect 87970 141264 88026 141273
rect 87970 141199 87972 141208
rect 88024 141199 88026 141208
rect 87972 141170 88024 141176
rect 87956 140924 88252 140944
rect 88012 140922 88036 140924
rect 88092 140922 88116 140924
rect 88172 140922 88196 140924
rect 88034 140870 88036 140922
rect 88098 140870 88110 140922
rect 88172 140870 88174 140922
rect 88012 140868 88036 140870
rect 88092 140868 88116 140870
rect 88172 140868 88196 140870
rect 87956 140848 88252 140868
rect 89956 140380 90252 140400
rect 90012 140378 90036 140380
rect 90092 140378 90116 140380
rect 90172 140378 90196 140380
rect 90034 140326 90036 140378
rect 90098 140326 90110 140378
rect 90172 140326 90174 140378
rect 90012 140324 90036 140326
rect 90092 140324 90116 140326
rect 90172 140324 90196 140326
rect 89956 140304 90252 140324
rect 88246 140176 88302 140185
rect 88246 140111 88302 140120
rect 88260 140010 88288 140111
rect 88248 140004 88300 140010
rect 88248 139946 88300 139952
rect 87956 139836 88252 139856
rect 88012 139834 88036 139836
rect 88092 139834 88116 139836
rect 88172 139834 88196 139836
rect 88034 139782 88036 139834
rect 88098 139782 88110 139834
rect 88172 139782 88174 139834
rect 88012 139780 88036 139782
rect 88092 139780 88116 139782
rect 88172 139780 88196 139782
rect 87956 139760 88252 139780
rect 89956 139292 90252 139312
rect 90012 139290 90036 139292
rect 90092 139290 90116 139292
rect 90172 139290 90196 139292
rect 90034 139238 90036 139290
rect 90098 139238 90110 139290
rect 90172 139238 90174 139290
rect 90012 139236 90036 139238
rect 90092 139236 90116 139238
rect 90172 139236 90196 139238
rect 89956 139216 90252 139236
rect 88062 139088 88118 139097
rect 88062 139023 88118 139032
rect 88076 138922 88104 139023
rect 88064 138916 88116 138922
rect 88064 138858 88116 138864
rect 87956 138748 88252 138768
rect 88012 138746 88036 138748
rect 88092 138746 88116 138748
rect 88172 138746 88196 138748
rect 88034 138694 88036 138746
rect 88098 138694 88110 138746
rect 88172 138694 88174 138746
rect 88012 138692 88036 138694
rect 88092 138692 88116 138694
rect 88172 138692 88196 138694
rect 87956 138672 88252 138692
rect 89956 138204 90252 138224
rect 90012 138202 90036 138204
rect 90092 138202 90116 138204
rect 90172 138202 90196 138204
rect 90034 138150 90036 138202
rect 90098 138150 90110 138202
rect 90172 138150 90174 138202
rect 90012 138148 90036 138150
rect 90092 138148 90116 138150
rect 90172 138148 90196 138150
rect 89956 138128 90252 138148
rect 87956 137660 88252 137680
rect 88012 137658 88036 137660
rect 88092 137658 88116 137660
rect 88172 137658 88196 137660
rect 88034 137606 88036 137658
rect 88098 137606 88110 137658
rect 88172 137606 88174 137658
rect 88012 137604 88036 137606
rect 88092 137604 88116 137606
rect 88172 137604 88196 137606
rect 87956 137584 88252 137604
rect 89956 137116 90252 137136
rect 90012 137114 90036 137116
rect 90092 137114 90116 137116
rect 90172 137114 90196 137116
rect 90034 137062 90036 137114
rect 90098 137062 90110 137114
rect 90172 137062 90174 137114
rect 90012 137060 90036 137062
rect 90092 137060 90116 137062
rect 90172 137060 90196 137062
rect 89956 137040 90252 137060
rect 87956 136572 88252 136592
rect 88012 136570 88036 136572
rect 88092 136570 88116 136572
rect 88172 136570 88196 136572
rect 88034 136518 88036 136570
rect 88098 136518 88110 136570
rect 88172 136518 88174 136570
rect 88012 136516 88036 136518
rect 88092 136516 88116 136518
rect 88172 136516 88196 136518
rect 87956 136496 88252 136516
rect 89956 136028 90252 136048
rect 90012 136026 90036 136028
rect 90092 136026 90116 136028
rect 90172 136026 90196 136028
rect 90034 135974 90036 136026
rect 90098 135974 90110 136026
rect 90172 135974 90174 136026
rect 90012 135972 90036 135974
rect 90092 135972 90116 135974
rect 90172 135972 90196 135974
rect 89956 135952 90252 135972
rect 87956 135484 88252 135504
rect 88012 135482 88036 135484
rect 88092 135482 88116 135484
rect 88172 135482 88196 135484
rect 88034 135430 88036 135482
rect 88098 135430 88110 135482
rect 88172 135430 88174 135482
rect 88012 135428 88036 135430
rect 88092 135428 88116 135430
rect 88172 135428 88196 135430
rect 87956 135408 88252 135428
rect 89956 134940 90252 134960
rect 90012 134938 90036 134940
rect 90092 134938 90116 134940
rect 90172 134938 90196 134940
rect 90034 134886 90036 134938
rect 90098 134886 90110 134938
rect 90172 134886 90174 134938
rect 90012 134884 90036 134886
rect 90092 134884 90116 134886
rect 90172 134884 90196 134886
rect 89956 134864 90252 134884
rect 87956 134396 88252 134416
rect 88012 134394 88036 134396
rect 88092 134394 88116 134396
rect 88172 134394 88196 134396
rect 88034 134342 88036 134394
rect 88098 134342 88110 134394
rect 88172 134342 88174 134394
rect 88012 134340 88036 134342
rect 88092 134340 88116 134342
rect 88172 134340 88196 134342
rect 87956 134320 88252 134340
rect 89956 133852 90252 133872
rect 90012 133850 90036 133852
rect 90092 133850 90116 133852
rect 90172 133850 90196 133852
rect 90034 133798 90036 133850
rect 90098 133798 90110 133850
rect 90172 133798 90174 133850
rect 90012 133796 90036 133798
rect 90092 133796 90116 133798
rect 90172 133796 90196 133798
rect 89956 133776 90252 133796
rect 87956 133308 88252 133328
rect 88012 133306 88036 133308
rect 88092 133306 88116 133308
rect 88172 133306 88196 133308
rect 88034 133254 88036 133306
rect 88098 133254 88110 133306
rect 88172 133254 88174 133306
rect 88012 133252 88036 133254
rect 88092 133252 88116 133254
rect 88172 133252 88196 133254
rect 87956 133232 88252 133252
rect 89956 132764 90252 132784
rect 90012 132762 90036 132764
rect 90092 132762 90116 132764
rect 90172 132762 90196 132764
rect 90034 132710 90036 132762
rect 90098 132710 90110 132762
rect 90172 132710 90174 132762
rect 90012 132708 90036 132710
rect 90092 132708 90116 132710
rect 90172 132708 90196 132710
rect 89956 132688 90252 132708
rect 87956 132220 88252 132240
rect 88012 132218 88036 132220
rect 88092 132218 88116 132220
rect 88172 132218 88196 132220
rect 88034 132166 88036 132218
rect 88098 132166 88110 132218
rect 88172 132166 88174 132218
rect 88012 132164 88036 132166
rect 88092 132164 88116 132166
rect 88172 132164 88196 132166
rect 87956 132144 88252 132164
rect 88246 131880 88302 131889
rect 88246 131815 88302 131824
rect 88260 131306 88288 131815
rect 89956 131676 90252 131696
rect 90012 131674 90036 131676
rect 90092 131674 90116 131676
rect 90172 131674 90196 131676
rect 90034 131622 90036 131674
rect 90098 131622 90110 131674
rect 90172 131622 90174 131674
rect 90012 131620 90036 131622
rect 90092 131620 90116 131622
rect 90172 131620 90196 131622
rect 89956 131600 90252 131620
rect 88248 131300 88300 131306
rect 88248 131242 88300 131248
rect 87956 131132 88252 131152
rect 88012 131130 88036 131132
rect 88092 131130 88116 131132
rect 88172 131130 88196 131132
rect 88034 131078 88036 131130
rect 88098 131078 88110 131130
rect 88172 131078 88174 131130
rect 88012 131076 88036 131078
rect 88092 131076 88116 131078
rect 88172 131076 88196 131078
rect 87956 131056 88252 131076
rect 89956 130588 90252 130608
rect 90012 130586 90036 130588
rect 90092 130586 90116 130588
rect 90172 130586 90196 130588
rect 90034 130534 90036 130586
rect 90098 130534 90110 130586
rect 90172 130534 90174 130586
rect 90012 130532 90036 130534
rect 90092 130532 90116 130534
rect 90172 130532 90196 130534
rect 89956 130512 90252 130532
rect 87956 130044 88252 130064
rect 88012 130042 88036 130044
rect 88092 130042 88116 130044
rect 88172 130042 88196 130044
rect 88034 129990 88036 130042
rect 88098 129990 88110 130042
rect 88172 129990 88174 130042
rect 88012 129988 88036 129990
rect 88092 129988 88116 129990
rect 88172 129988 88196 129990
rect 87956 129968 88252 129988
rect 89956 129500 90252 129520
rect 90012 129498 90036 129500
rect 90092 129498 90116 129500
rect 90172 129498 90196 129500
rect 90034 129446 90036 129498
rect 90098 129446 90110 129498
rect 90172 129446 90174 129498
rect 90012 129444 90036 129446
rect 90092 129444 90116 129446
rect 90172 129444 90196 129446
rect 89956 129424 90252 129444
rect 88246 129296 88302 129305
rect 88246 129231 88302 129240
rect 88260 129146 88288 129231
rect 88260 129118 88380 129146
rect 87956 128956 88252 128976
rect 88012 128954 88036 128956
rect 88092 128954 88116 128956
rect 88172 128954 88196 128956
rect 88034 128902 88036 128954
rect 88098 128902 88110 128954
rect 88172 128902 88174 128954
rect 88012 128900 88036 128902
rect 88092 128900 88116 128902
rect 88172 128900 88196 128902
rect 87956 128880 88252 128900
rect 88352 128738 88380 129118
rect 88260 128710 88380 128738
rect 88260 128518 88288 128710
rect 88248 128512 88300 128518
rect 88248 128454 88300 128460
rect 89956 128412 90252 128432
rect 90012 128410 90036 128412
rect 90092 128410 90116 128412
rect 90172 128410 90196 128412
rect 90034 128358 90036 128410
rect 90098 128358 90110 128410
rect 90172 128358 90174 128410
rect 90012 128356 90036 128358
rect 90092 128356 90116 128358
rect 90172 128356 90196 128358
rect 89956 128336 90252 128356
rect 88246 128208 88302 128217
rect 88246 128143 88302 128152
rect 88260 128058 88288 128143
rect 88260 128030 88380 128058
rect 87956 127868 88252 127888
rect 88012 127866 88036 127868
rect 88092 127866 88116 127868
rect 88172 127866 88196 127868
rect 88034 127814 88036 127866
rect 88098 127814 88110 127866
rect 88172 127814 88174 127866
rect 88012 127812 88036 127814
rect 88092 127812 88116 127814
rect 88172 127812 88196 127814
rect 87956 127792 88252 127812
rect 88352 127650 88380 128030
rect 88260 127622 88380 127650
rect 88260 127022 88288 127622
rect 89956 127324 90252 127344
rect 90012 127322 90036 127324
rect 90092 127322 90116 127324
rect 90172 127322 90196 127324
rect 90034 127270 90036 127322
rect 90098 127270 90110 127322
rect 90172 127270 90174 127322
rect 90012 127268 90036 127270
rect 90092 127268 90116 127270
rect 90172 127268 90196 127270
rect 89956 127248 90252 127268
rect 88248 127016 88300 127022
rect 88248 126958 88300 126964
rect 87956 126780 88252 126800
rect 88012 126778 88036 126780
rect 88092 126778 88116 126780
rect 88172 126778 88196 126780
rect 88034 126726 88036 126778
rect 88098 126726 88110 126778
rect 88172 126726 88174 126778
rect 88012 126724 88036 126726
rect 88092 126724 88116 126726
rect 88172 126724 88196 126726
rect 87956 126704 88252 126724
rect 89956 126236 90252 126256
rect 90012 126234 90036 126236
rect 90092 126234 90116 126236
rect 90172 126234 90196 126236
rect 90034 126182 90036 126234
rect 90098 126182 90110 126234
rect 90172 126182 90174 126234
rect 90012 126180 90036 126182
rect 90092 126180 90116 126182
rect 90172 126180 90196 126182
rect 89956 126160 90252 126180
rect 87970 125896 88026 125905
rect 87970 125831 87972 125840
rect 88024 125831 88026 125840
rect 87972 125802 88024 125808
rect 87956 125692 88252 125712
rect 88012 125690 88036 125692
rect 88092 125690 88116 125692
rect 88172 125690 88196 125692
rect 88034 125638 88036 125690
rect 88098 125638 88110 125690
rect 88172 125638 88174 125690
rect 88012 125636 88036 125638
rect 88092 125636 88116 125638
rect 88172 125636 88196 125638
rect 87956 125616 88252 125636
rect 89956 125148 90252 125168
rect 90012 125146 90036 125148
rect 90092 125146 90116 125148
rect 90172 125146 90196 125148
rect 90034 125094 90036 125146
rect 90098 125094 90110 125146
rect 90172 125094 90174 125146
rect 90012 125092 90036 125094
rect 90092 125092 90116 125094
rect 90172 125092 90196 125094
rect 89956 125072 90252 125092
rect 87956 124604 88252 124624
rect 88012 124602 88036 124604
rect 88092 124602 88116 124604
rect 88172 124602 88196 124604
rect 88034 124550 88036 124602
rect 88098 124550 88110 124602
rect 88172 124550 88174 124602
rect 88012 124548 88036 124550
rect 88092 124548 88116 124550
rect 88172 124548 88196 124550
rect 87956 124528 88252 124548
rect 88246 124400 88302 124409
rect 88246 124335 88302 124344
rect 88260 123706 88288 124335
rect 89956 124060 90252 124080
rect 90012 124058 90036 124060
rect 90092 124058 90116 124060
rect 90172 124058 90196 124060
rect 90034 124006 90036 124058
rect 90098 124006 90110 124058
rect 90172 124006 90174 124058
rect 90012 124004 90036 124006
rect 90092 124004 90116 124006
rect 90172 124004 90196 124006
rect 89956 123984 90252 124004
rect 88260 123678 88380 123706
rect 87956 123516 88252 123536
rect 88012 123514 88036 123516
rect 88092 123514 88116 123516
rect 88172 123514 88196 123516
rect 88034 123462 88036 123514
rect 88098 123462 88110 123514
rect 88172 123462 88174 123514
rect 88012 123460 88036 123462
rect 88092 123460 88116 123462
rect 88172 123460 88196 123462
rect 87956 123440 88252 123460
rect 87970 123312 88026 123321
rect 87970 123247 88026 123256
rect 87984 122874 88012 123247
rect 87972 122868 88024 122874
rect 87972 122810 88024 122816
rect 87956 122428 88252 122448
rect 88012 122426 88036 122428
rect 88092 122426 88116 122428
rect 88172 122426 88196 122428
rect 88034 122374 88036 122426
rect 88098 122374 88110 122426
rect 88172 122374 88174 122426
rect 88012 122372 88036 122374
rect 88092 122372 88116 122374
rect 88172 122372 88196 122374
rect 87956 122352 88252 122372
rect 88352 122210 88380 123678
rect 89956 122972 90252 122992
rect 90012 122970 90036 122972
rect 90092 122970 90116 122972
rect 90172 122970 90196 122972
rect 90034 122918 90036 122970
rect 90098 122918 90110 122970
rect 90172 122918 90174 122970
rect 90012 122916 90036 122918
rect 90092 122916 90116 122918
rect 90172 122916 90196 122918
rect 89956 122896 90252 122916
rect 87880 122188 87932 122194
rect 87880 122130 87932 122136
rect 88260 122182 88380 122210
rect 87878 122088 87934 122097
rect 87878 122023 87934 122032
rect 87892 121514 87920 122023
rect 88260 121530 88288 122182
rect 89956 121884 90252 121904
rect 90012 121882 90036 121884
rect 90092 121882 90116 121884
rect 90172 121882 90196 121884
rect 90034 121830 90036 121882
rect 90098 121830 90110 121882
rect 90172 121830 90174 121882
rect 90012 121828 90036 121830
rect 90092 121828 90116 121830
rect 90172 121828 90196 121830
rect 89956 121808 90252 121828
rect 87880 121508 87932 121514
rect 88260 121502 88380 121530
rect 87880 121450 87932 121456
rect 87956 121340 88252 121360
rect 88012 121338 88036 121340
rect 88092 121338 88116 121340
rect 88172 121338 88196 121340
rect 88034 121286 88036 121338
rect 88098 121286 88110 121338
rect 88172 121286 88174 121338
rect 88012 121284 88036 121286
rect 88092 121284 88116 121286
rect 88172 121284 88196 121286
rect 87956 121264 88252 121284
rect 88352 121122 88380 121502
rect 88260 121094 88380 121122
rect 87878 120592 87934 120601
rect 87878 120527 87934 120536
rect 87892 120154 87920 120527
rect 88260 120442 88288 121094
rect 89956 120796 90252 120816
rect 90012 120794 90036 120796
rect 90092 120794 90116 120796
rect 90172 120794 90196 120796
rect 90034 120742 90036 120794
rect 90098 120742 90110 120794
rect 90172 120742 90174 120794
rect 90012 120740 90036 120742
rect 90092 120740 90116 120742
rect 90172 120740 90196 120742
rect 89956 120720 90252 120740
rect 88260 120414 88380 120442
rect 87956 120252 88252 120272
rect 88012 120250 88036 120252
rect 88092 120250 88116 120252
rect 88172 120250 88196 120252
rect 88034 120198 88036 120250
rect 88098 120198 88110 120250
rect 88172 120198 88174 120250
rect 88012 120196 88036 120198
rect 88092 120196 88116 120198
rect 88172 120196 88196 120198
rect 87956 120176 88252 120196
rect 87880 120148 87932 120154
rect 87880 120090 87932 120096
rect 88352 120034 88380 120414
rect 88260 120006 88380 120034
rect 87878 119504 87934 119513
rect 87878 119439 87934 119448
rect 87892 118726 87920 119439
rect 88260 119354 88288 120006
rect 89956 119708 90252 119728
rect 90012 119706 90036 119708
rect 90092 119706 90116 119708
rect 90172 119706 90196 119708
rect 90034 119654 90036 119706
rect 90098 119654 90110 119706
rect 90172 119654 90174 119706
rect 90012 119652 90036 119654
rect 90092 119652 90116 119654
rect 90172 119652 90196 119654
rect 89956 119632 90252 119652
rect 88260 119326 88380 119354
rect 87956 119164 88252 119184
rect 88012 119162 88036 119164
rect 88092 119162 88116 119164
rect 88172 119162 88196 119164
rect 88034 119110 88036 119162
rect 88098 119110 88110 119162
rect 88172 119110 88174 119162
rect 88012 119108 88036 119110
rect 88092 119108 88116 119110
rect 88172 119108 88196 119110
rect 87956 119088 88252 119108
rect 88352 118946 88380 119326
rect 87984 118918 88380 118946
rect 87880 118720 87932 118726
rect 87880 118662 87932 118668
rect 87984 118266 88012 118918
rect 89956 118620 90252 118640
rect 90012 118618 90036 118620
rect 90092 118618 90116 118620
rect 90172 118618 90196 118620
rect 90034 118566 90036 118618
rect 90098 118566 90110 118618
rect 90172 118566 90174 118618
rect 90012 118564 90036 118566
rect 90092 118564 90116 118566
rect 90172 118564 90196 118566
rect 89956 118544 90252 118564
rect 88982 118416 89038 118425
rect 88982 118351 89038 118360
rect 87892 118238 88012 118266
rect 87788 104372 87840 104378
rect 87788 104314 87840 104320
rect 87892 104258 87920 118238
rect 87956 118076 88252 118096
rect 88012 118074 88036 118076
rect 88092 118074 88116 118076
rect 88172 118074 88196 118076
rect 88034 118022 88036 118074
rect 88098 118022 88110 118074
rect 88172 118022 88174 118074
rect 88012 118020 88036 118022
rect 88092 118020 88116 118022
rect 88172 118020 88196 118022
rect 87956 118000 88252 118020
rect 87956 116988 88252 117008
rect 88012 116986 88036 116988
rect 88092 116986 88116 116988
rect 88172 116986 88196 116988
rect 88034 116934 88036 116986
rect 88098 116934 88110 116986
rect 88172 116934 88174 116986
rect 88012 116932 88036 116934
rect 88092 116932 88116 116934
rect 88172 116932 88196 116934
rect 87956 116912 88252 116932
rect 88246 116784 88302 116793
rect 88246 116719 88302 116728
rect 88260 116090 88288 116719
rect 88260 116062 88380 116090
rect 88352 115934 88380 116062
rect 87956 115900 88252 115920
rect 88352 115906 88564 115934
rect 88012 115898 88036 115900
rect 88092 115898 88116 115900
rect 88172 115898 88196 115900
rect 88034 115846 88036 115898
rect 88098 115846 88110 115898
rect 88172 115846 88174 115898
rect 88012 115844 88036 115846
rect 88092 115844 88116 115846
rect 88172 115844 88196 115846
rect 87956 115824 88252 115844
rect 87956 114812 88252 114832
rect 88012 114810 88036 114812
rect 88092 114810 88116 114812
rect 88172 114810 88196 114812
rect 88034 114758 88036 114810
rect 88098 114758 88110 114810
rect 88172 114758 88174 114810
rect 88012 114756 88036 114758
rect 88092 114756 88116 114758
rect 88172 114756 88196 114758
rect 87956 114736 88252 114756
rect 87970 114608 88026 114617
rect 87970 114543 87972 114552
rect 88024 114543 88026 114552
rect 87972 114514 88024 114520
rect 87956 113724 88252 113744
rect 88012 113722 88036 113724
rect 88092 113722 88116 113724
rect 88172 113722 88196 113724
rect 88034 113670 88036 113722
rect 88098 113670 88110 113722
rect 88172 113670 88174 113722
rect 88012 113668 88036 113670
rect 88092 113668 88116 113670
rect 88172 113668 88196 113670
rect 87956 113648 88252 113668
rect 87956 112636 88252 112656
rect 88012 112634 88036 112636
rect 88092 112634 88116 112636
rect 88172 112634 88196 112636
rect 88034 112582 88036 112634
rect 88098 112582 88110 112634
rect 88172 112582 88174 112634
rect 88012 112580 88036 112582
rect 88092 112580 88116 112582
rect 88172 112580 88196 112582
rect 87956 112560 88252 112580
rect 87970 112432 88026 112441
rect 87970 112367 88026 112376
rect 87984 111858 88012 112367
rect 87972 111852 88024 111858
rect 87972 111794 88024 111800
rect 87956 111548 88252 111568
rect 88012 111546 88036 111548
rect 88092 111546 88116 111548
rect 88172 111546 88196 111548
rect 88034 111494 88036 111546
rect 88098 111494 88110 111546
rect 88172 111494 88174 111546
rect 88012 111492 88036 111494
rect 88092 111492 88116 111494
rect 88172 111492 88196 111494
rect 87956 111472 88252 111492
rect 88246 111208 88302 111217
rect 88246 111143 88302 111152
rect 88260 110650 88288 111143
rect 88260 110622 88380 110650
rect 87956 110460 88252 110480
rect 88012 110458 88036 110460
rect 88092 110458 88116 110460
rect 88172 110458 88196 110460
rect 88034 110406 88036 110458
rect 88098 110406 88110 110458
rect 88172 110406 88174 110458
rect 88012 110404 88036 110406
rect 88092 110404 88116 110406
rect 88172 110404 88196 110406
rect 87956 110384 88252 110404
rect 88352 110242 88380 110622
rect 88260 110214 88380 110242
rect 88260 109562 88288 110214
rect 88260 109534 88472 109562
rect 87956 109372 88252 109392
rect 88012 109370 88036 109372
rect 88092 109370 88116 109372
rect 88172 109370 88196 109372
rect 88034 109318 88036 109370
rect 88098 109318 88110 109370
rect 88172 109318 88174 109370
rect 88012 109316 88036 109318
rect 88092 109316 88116 109318
rect 88172 109316 88196 109318
rect 87956 109296 88252 109316
rect 88246 109168 88302 109177
rect 88246 109103 88302 109112
rect 87972 108656 88024 108662
rect 87970 108624 87972 108633
rect 88024 108624 88026 108633
rect 87970 108559 88026 108568
rect 88260 108458 88288 109103
rect 88340 108588 88392 108594
rect 88340 108530 88392 108536
rect 88248 108452 88300 108458
rect 88248 108394 88300 108400
rect 87956 108284 88252 108304
rect 88012 108282 88036 108284
rect 88092 108282 88116 108284
rect 88172 108282 88196 108284
rect 88034 108230 88036 108282
rect 88098 108230 88110 108282
rect 88172 108230 88174 108282
rect 88012 108228 88036 108230
rect 88092 108228 88116 108230
rect 88172 108228 88196 108230
rect 87956 108208 88252 108228
rect 88352 108066 88380 108530
rect 88260 108038 88380 108066
rect 87970 107536 88026 107545
rect 87970 107471 88026 107480
rect 87984 107370 88012 107471
rect 88260 107386 88288 108038
rect 87972 107364 88024 107370
rect 88260 107358 88380 107386
rect 87972 107306 88024 107312
rect 87956 107196 88252 107216
rect 88012 107194 88036 107196
rect 88092 107194 88116 107196
rect 88172 107194 88196 107196
rect 88034 107142 88036 107194
rect 88098 107142 88110 107194
rect 88172 107142 88174 107194
rect 88012 107140 88036 107142
rect 88092 107140 88116 107142
rect 88172 107140 88196 107142
rect 87956 107120 88252 107140
rect 88352 106978 88380 107358
rect 88260 106950 88380 106978
rect 88260 106298 88288 106950
rect 88260 106270 88380 106298
rect 87956 106108 88252 106128
rect 88012 106106 88036 106108
rect 88092 106106 88116 106108
rect 88172 106106 88196 106108
rect 88034 106054 88036 106106
rect 88098 106054 88110 106106
rect 88172 106054 88174 106106
rect 88012 106052 88036 106054
rect 88092 106052 88116 106054
rect 88172 106052 88196 106054
rect 87956 106032 88252 106052
rect 87956 105020 88252 105040
rect 88012 105018 88036 105020
rect 88092 105018 88116 105020
rect 88172 105018 88196 105020
rect 88034 104966 88036 105018
rect 88098 104966 88110 105018
rect 88172 104966 88174 105018
rect 88012 104964 88036 104966
rect 88092 104964 88116 104966
rect 88172 104964 88196 104966
rect 87956 104944 88252 104964
rect 87800 104230 87920 104258
rect 87604 98932 87656 98938
rect 87604 98874 87656 98880
rect 87696 98932 87748 98938
rect 87696 98874 87748 98880
rect 87602 98832 87658 98841
rect 87800 98818 87828 104230
rect 87956 103932 88252 103952
rect 88012 103930 88036 103932
rect 88092 103930 88116 103932
rect 88172 103930 88196 103932
rect 88034 103878 88036 103930
rect 88098 103878 88110 103930
rect 88172 103878 88174 103930
rect 88012 103876 88036 103878
rect 88092 103876 88116 103878
rect 88172 103876 88196 103878
rect 87956 103856 88252 103876
rect 87956 102844 88252 102864
rect 88012 102842 88036 102844
rect 88092 102842 88116 102844
rect 88172 102842 88196 102844
rect 88034 102790 88036 102842
rect 88098 102790 88110 102842
rect 88172 102790 88174 102842
rect 88012 102788 88036 102790
rect 88092 102788 88116 102790
rect 88172 102788 88196 102790
rect 87956 102768 88252 102788
rect 87956 101756 88252 101776
rect 88012 101754 88036 101756
rect 88092 101754 88116 101756
rect 88172 101754 88196 101756
rect 88034 101702 88036 101754
rect 88098 101702 88110 101754
rect 88172 101702 88174 101754
rect 88012 101700 88036 101702
rect 88092 101700 88116 101702
rect 88172 101700 88196 101702
rect 87956 101680 88252 101700
rect 87880 101108 87932 101114
rect 87880 101050 87932 101056
rect 87892 99754 87920 101050
rect 87956 100668 88252 100688
rect 88012 100666 88036 100668
rect 88092 100666 88116 100668
rect 88172 100666 88196 100668
rect 88034 100614 88036 100666
rect 88098 100614 88110 100666
rect 88172 100614 88174 100666
rect 88012 100612 88036 100614
rect 88092 100612 88116 100614
rect 88172 100612 88196 100614
rect 87956 100592 88252 100612
rect 87880 99748 87932 99754
rect 87880 99690 87932 99696
rect 87956 99580 88252 99600
rect 88012 99578 88036 99580
rect 88092 99578 88116 99580
rect 88172 99578 88196 99580
rect 88034 99526 88036 99578
rect 88098 99526 88110 99578
rect 88172 99526 88174 99578
rect 88012 99524 88036 99526
rect 88092 99524 88116 99526
rect 88172 99524 88196 99526
rect 87956 99504 88252 99524
rect 87880 98932 87932 98938
rect 87880 98874 87932 98880
rect 87602 98767 87658 98776
rect 87708 98790 87828 98818
rect 87512 95668 87564 95674
rect 87512 95610 87564 95616
rect 87420 95328 87472 95334
rect 87420 95270 87472 95276
rect 86868 94988 86920 94994
rect 86868 94930 86920 94936
rect 86868 94852 86920 94858
rect 86868 94794 86920 94800
rect 86776 92064 86828 92070
rect 86776 92006 86828 92012
rect 86684 90772 86736 90778
rect 86684 90714 86736 90720
rect 86684 90092 86736 90098
rect 86684 90034 86736 90040
rect 86696 89593 86724 90034
rect 86682 89584 86738 89593
rect 86682 89519 86738 89528
rect 86684 89480 86736 89486
rect 86684 89422 86736 89428
rect 86696 86873 86724 89422
rect 86682 86864 86738 86873
rect 86682 86799 86738 86808
rect 86788 84946 86816 92006
rect 86880 89690 86908 94794
rect 86960 94512 87012 94518
rect 86960 94454 87012 94460
rect 86972 94353 87000 94454
rect 86958 94344 87014 94353
rect 86958 94279 87014 94288
rect 87512 94240 87564 94246
rect 87512 94182 87564 94188
rect 87524 93786 87552 94182
rect 87616 93974 87644 98767
rect 87708 97578 87736 98790
rect 87788 98728 87840 98734
rect 87788 98670 87840 98676
rect 87696 97572 87748 97578
rect 87696 97514 87748 97520
rect 87800 95985 87828 98670
rect 87892 97866 87920 98874
rect 88352 98734 88380 106270
rect 88444 101114 88472 109534
rect 88536 108526 88564 115906
rect 88524 108520 88576 108526
rect 88524 108462 88576 108468
rect 88522 105088 88578 105097
rect 88522 105023 88578 105032
rect 88432 101108 88484 101114
rect 88432 101050 88484 101056
rect 88432 99884 88484 99890
rect 88432 99826 88484 99832
rect 88444 99210 88472 99826
rect 88536 99822 88564 105023
rect 88708 104372 88760 104378
rect 88708 104314 88760 104320
rect 88616 99952 88668 99958
rect 88616 99894 88668 99900
rect 88524 99816 88576 99822
rect 88524 99758 88576 99764
rect 88432 99204 88484 99210
rect 88432 99146 88484 99152
rect 88628 99142 88656 99894
rect 88616 99136 88668 99142
rect 88616 99078 88668 99084
rect 88340 98728 88392 98734
rect 88340 98670 88392 98676
rect 87956 98492 88252 98512
rect 88012 98490 88036 98492
rect 88092 98490 88116 98492
rect 88172 98490 88196 98492
rect 88034 98438 88036 98490
rect 88098 98438 88110 98490
rect 88172 98438 88174 98490
rect 88012 98436 88036 98438
rect 88092 98436 88116 98438
rect 88172 98436 88196 98438
rect 87956 98416 88252 98436
rect 87892 97838 88012 97866
rect 87880 97708 87932 97714
rect 87880 97650 87932 97656
rect 87786 95976 87842 95985
rect 87786 95911 87842 95920
rect 87788 94036 87840 94042
rect 87788 93978 87840 93984
rect 87604 93968 87656 93974
rect 87604 93910 87656 93916
rect 87696 93832 87748 93838
rect 86960 93764 87012 93770
rect 87524 93758 87644 93786
rect 87696 93774 87748 93780
rect 86960 93706 87012 93712
rect 86972 90098 87000 93706
rect 87236 93696 87288 93702
rect 87236 93638 87288 93644
rect 87052 92404 87104 92410
rect 87052 92346 87104 92352
rect 86960 90092 87012 90098
rect 86960 90034 87012 90040
rect 87064 89978 87092 92346
rect 87144 92336 87196 92342
rect 87144 92278 87196 92284
rect 86972 89950 87092 89978
rect 86868 89684 86920 89690
rect 86868 89626 86920 89632
rect 86866 89584 86922 89593
rect 86866 89519 86922 89528
rect 86696 84918 86816 84946
rect 86696 70394 86724 84918
rect 86880 80209 86908 89519
rect 86972 84946 87000 89950
rect 87156 89842 87184 92278
rect 87064 89814 87184 89842
rect 87064 89714 87092 89814
rect 87064 89686 87184 89714
rect 87050 89584 87106 89593
rect 87050 89519 87106 89528
rect 87064 85105 87092 89519
rect 87050 85096 87106 85105
rect 87050 85031 87106 85040
rect 86972 84918 87092 84946
rect 86960 84788 87012 84794
rect 86960 84730 87012 84736
rect 86866 80200 86922 80209
rect 86776 80164 86828 80170
rect 86866 80135 86922 80144
rect 86776 80106 86828 80112
rect 86788 79642 86816 80106
rect 86972 80073 87000 84730
rect 86958 80064 87014 80073
rect 86958 79999 87014 80008
rect 86788 79614 87000 79642
rect 86972 74769 87000 79614
rect 87064 78577 87092 84918
rect 87050 78568 87106 78577
rect 87050 78503 87106 78512
rect 87052 77172 87104 77178
rect 87052 77114 87104 77120
rect 87064 75993 87092 77114
rect 87156 77081 87184 89686
rect 87248 84794 87276 93638
rect 87328 93492 87380 93498
rect 87328 93434 87380 93440
rect 87340 84946 87368 93434
rect 87420 92676 87472 92682
rect 87420 92618 87472 92624
rect 87432 85105 87460 92618
rect 87512 92268 87564 92274
rect 87512 92210 87564 92216
rect 87524 89865 87552 92210
rect 87510 89856 87566 89865
rect 87510 89791 87566 89800
rect 87512 89684 87564 89690
rect 87512 89626 87564 89632
rect 87418 85096 87474 85105
rect 87418 85031 87474 85040
rect 87340 84918 87460 84946
rect 87236 84788 87288 84794
rect 87236 84730 87288 84736
rect 87234 84688 87290 84697
rect 87234 84623 87290 84632
rect 87142 77072 87198 77081
rect 87142 77007 87198 77016
rect 87050 75984 87106 75993
rect 87050 75919 87106 75928
rect 87144 75540 87196 75546
rect 87144 75482 87196 75488
rect 86958 74760 87014 74769
rect 86958 74695 87014 74704
rect 86960 74452 87012 74458
rect 86960 74394 87012 74400
rect 86972 73681 87000 74394
rect 86958 73672 87014 73681
rect 86958 73607 87014 73616
rect 87156 71097 87184 75482
rect 87248 72593 87276 84623
rect 87326 84552 87382 84561
rect 87326 84487 87382 84496
rect 87340 80170 87368 84487
rect 87328 80164 87380 80170
rect 87328 80106 87380 80112
rect 87326 80068 87382 80077
rect 87432 80054 87460 84918
rect 87524 80170 87552 89626
rect 87512 80164 87564 80170
rect 87512 80106 87564 80112
rect 87432 80026 87552 80054
rect 87326 80003 87382 80012
rect 87234 72584 87290 72593
rect 87234 72519 87290 72528
rect 87142 71088 87198 71097
rect 87142 71023 87198 71032
rect 86696 70366 86908 70394
rect 86682 38312 86738 38321
rect 86682 38247 86738 38256
rect 86592 32020 86644 32026
rect 86592 31962 86644 31968
rect 86590 30832 86646 30841
rect 86590 30767 86646 30776
rect 86500 29300 86552 29306
rect 86500 29242 86552 29248
rect 86408 27600 86460 27606
rect 86408 27542 86460 27548
rect 86316 26580 86368 26586
rect 86316 26522 86368 26528
rect 85956 26140 86252 26160
rect 86012 26138 86036 26140
rect 86092 26138 86116 26140
rect 86172 26138 86196 26140
rect 86034 26086 86036 26138
rect 86098 26086 86110 26138
rect 86172 26086 86174 26138
rect 86012 26084 86036 26086
rect 86092 26084 86116 26086
rect 86172 26084 86196 26086
rect 85956 26064 86252 26084
rect 85956 25052 86252 25072
rect 86012 25050 86036 25052
rect 86092 25050 86116 25052
rect 86172 25050 86196 25052
rect 86034 24998 86036 25050
rect 86098 24998 86110 25050
rect 86172 24998 86174 25050
rect 86012 24996 86036 24998
rect 86092 24996 86116 24998
rect 86172 24996 86196 24998
rect 85956 24976 86252 24996
rect 85856 24404 85908 24410
rect 85856 24346 85908 24352
rect 85956 23964 86252 23984
rect 86012 23962 86036 23964
rect 86092 23962 86116 23964
rect 86172 23962 86196 23964
rect 86034 23910 86036 23962
rect 86098 23910 86110 23962
rect 86172 23910 86174 23962
rect 86012 23908 86036 23910
rect 86092 23908 86116 23910
rect 86172 23908 86196 23910
rect 85956 23888 86252 23908
rect 85956 22876 86252 22896
rect 86012 22874 86036 22876
rect 86092 22874 86116 22876
rect 86172 22874 86196 22876
rect 86034 22822 86036 22874
rect 86098 22822 86110 22874
rect 86172 22822 86174 22874
rect 86012 22820 86036 22822
rect 86092 22820 86116 22822
rect 86172 22820 86196 22822
rect 85956 22800 86252 22820
rect 85956 21788 86252 21808
rect 86012 21786 86036 21788
rect 86092 21786 86116 21788
rect 86172 21786 86196 21788
rect 86034 21734 86036 21786
rect 86098 21734 86110 21786
rect 86172 21734 86174 21786
rect 86012 21732 86036 21734
rect 86092 21732 86116 21734
rect 86172 21732 86196 21734
rect 85956 21712 86252 21732
rect 85956 20700 86252 20720
rect 86012 20698 86036 20700
rect 86092 20698 86116 20700
rect 86172 20698 86196 20700
rect 86034 20646 86036 20698
rect 86098 20646 86110 20698
rect 86172 20646 86174 20698
rect 86012 20644 86036 20646
rect 86092 20644 86116 20646
rect 86172 20644 86196 20646
rect 85956 20624 86252 20644
rect 86314 19952 86370 19961
rect 86314 19887 86370 19896
rect 85956 19612 86252 19632
rect 86012 19610 86036 19612
rect 86092 19610 86116 19612
rect 86172 19610 86196 19612
rect 86034 19558 86036 19610
rect 86098 19558 86110 19610
rect 86172 19558 86174 19610
rect 86012 19556 86036 19558
rect 86092 19556 86116 19558
rect 86172 19556 86196 19558
rect 85956 19536 86252 19556
rect 85956 18524 86252 18544
rect 86012 18522 86036 18524
rect 86092 18522 86116 18524
rect 86172 18522 86196 18524
rect 86034 18470 86036 18522
rect 86098 18470 86110 18522
rect 86172 18470 86174 18522
rect 86012 18468 86036 18470
rect 86092 18468 86116 18470
rect 86172 18468 86196 18470
rect 85956 18448 86252 18468
rect 85956 17436 86252 17456
rect 86012 17434 86036 17436
rect 86092 17434 86116 17436
rect 86172 17434 86196 17436
rect 86034 17382 86036 17434
rect 86098 17382 86110 17434
rect 86172 17382 86174 17434
rect 86012 17380 86036 17382
rect 86092 17380 86116 17382
rect 86172 17380 86196 17382
rect 85956 17360 86252 17380
rect 85956 16348 86252 16368
rect 86012 16346 86036 16348
rect 86092 16346 86116 16348
rect 86172 16346 86196 16348
rect 86034 16294 86036 16346
rect 86098 16294 86110 16346
rect 86172 16294 86174 16346
rect 86012 16292 86036 16294
rect 86092 16292 86116 16294
rect 86172 16292 86196 16294
rect 85956 16272 86252 16292
rect 85956 15260 86252 15280
rect 86012 15258 86036 15260
rect 86092 15258 86116 15260
rect 86172 15258 86196 15260
rect 86034 15206 86036 15258
rect 86098 15206 86110 15258
rect 86172 15206 86174 15258
rect 86012 15204 86036 15206
rect 86092 15204 86116 15206
rect 86172 15204 86196 15206
rect 85956 15184 86252 15204
rect 85956 14172 86252 14192
rect 86012 14170 86036 14172
rect 86092 14170 86116 14172
rect 86172 14170 86196 14172
rect 86034 14118 86036 14170
rect 86098 14118 86110 14170
rect 86172 14118 86174 14170
rect 86012 14116 86036 14118
rect 86092 14116 86116 14118
rect 86172 14116 86196 14118
rect 85956 14096 86252 14116
rect 85956 13084 86252 13104
rect 86012 13082 86036 13084
rect 86092 13082 86116 13084
rect 86172 13082 86196 13084
rect 86034 13030 86036 13082
rect 86098 13030 86110 13082
rect 86172 13030 86174 13082
rect 86012 13028 86036 13030
rect 86092 13028 86116 13030
rect 86172 13028 86196 13030
rect 85956 13008 86252 13028
rect 85956 11996 86252 12016
rect 86012 11994 86036 11996
rect 86092 11994 86116 11996
rect 86172 11994 86196 11996
rect 86034 11942 86036 11994
rect 86098 11942 86110 11994
rect 86172 11942 86174 11994
rect 86012 11940 86036 11942
rect 86092 11940 86116 11942
rect 86172 11940 86196 11942
rect 85956 11920 86252 11940
rect 85956 10908 86252 10928
rect 86012 10906 86036 10908
rect 86092 10906 86116 10908
rect 86172 10906 86196 10908
rect 86034 10854 86036 10906
rect 86098 10854 86110 10906
rect 86172 10854 86174 10906
rect 86012 10852 86036 10854
rect 86092 10852 86116 10854
rect 86172 10852 86196 10854
rect 85956 10832 86252 10852
rect 85956 9820 86252 9840
rect 86012 9818 86036 9820
rect 86092 9818 86116 9820
rect 86172 9818 86196 9820
rect 86034 9766 86036 9818
rect 86098 9766 86110 9818
rect 86172 9766 86174 9818
rect 86012 9764 86036 9766
rect 86092 9764 86116 9766
rect 86172 9764 86196 9766
rect 85956 9744 86252 9764
rect 85956 8732 86252 8752
rect 86012 8730 86036 8732
rect 86092 8730 86116 8732
rect 86172 8730 86196 8732
rect 86034 8678 86036 8730
rect 86098 8678 86110 8730
rect 86172 8678 86174 8730
rect 86012 8676 86036 8678
rect 86092 8676 86116 8678
rect 86172 8676 86196 8678
rect 85956 8656 86252 8676
rect 85956 7644 86252 7664
rect 86012 7642 86036 7644
rect 86092 7642 86116 7644
rect 86172 7642 86196 7644
rect 86034 7590 86036 7642
rect 86098 7590 86110 7642
rect 86172 7590 86174 7642
rect 86012 7588 86036 7590
rect 86092 7588 86116 7590
rect 86172 7588 86196 7590
rect 85956 7568 86252 7588
rect 85956 6556 86252 6576
rect 86012 6554 86036 6556
rect 86092 6554 86116 6556
rect 86172 6554 86196 6556
rect 86034 6502 86036 6554
rect 86098 6502 86110 6554
rect 86172 6502 86174 6554
rect 86012 6500 86036 6502
rect 86092 6500 86116 6502
rect 86172 6500 86196 6502
rect 85956 6480 86252 6500
rect 85956 5468 86252 5488
rect 86012 5466 86036 5468
rect 86092 5466 86116 5468
rect 86172 5466 86196 5468
rect 86034 5414 86036 5466
rect 86098 5414 86110 5466
rect 86172 5414 86174 5466
rect 86012 5412 86036 5414
rect 86092 5412 86116 5414
rect 86172 5412 86196 5414
rect 85956 5392 86252 5412
rect 85856 5364 85908 5370
rect 85856 5306 85908 5312
rect 85868 3602 85896 5306
rect 85956 4380 86252 4400
rect 86012 4378 86036 4380
rect 86092 4378 86116 4380
rect 86172 4378 86196 4380
rect 86034 4326 86036 4378
rect 86098 4326 86110 4378
rect 86172 4326 86174 4378
rect 86012 4324 86036 4326
rect 86092 4324 86116 4326
rect 86172 4324 86196 4326
rect 85956 4304 86252 4324
rect 85856 3596 85908 3602
rect 85856 3538 85908 3544
rect 85764 3528 85816 3534
rect 85764 3470 85816 3476
rect 85776 3194 85804 3470
rect 85956 3292 86252 3312
rect 86012 3290 86036 3292
rect 86092 3290 86116 3292
rect 86172 3290 86196 3292
rect 86034 3238 86036 3290
rect 86098 3238 86110 3290
rect 86172 3238 86174 3290
rect 86012 3236 86036 3238
rect 86092 3236 86116 3238
rect 86172 3236 86196 3238
rect 85956 3216 86252 3236
rect 85764 3188 85816 3194
rect 85764 3130 85816 3136
rect 85956 2204 86252 2224
rect 86012 2202 86036 2204
rect 86092 2202 86116 2204
rect 86172 2202 86196 2204
rect 86034 2150 86036 2202
rect 86098 2150 86110 2202
rect 86172 2150 86174 2202
rect 86012 2148 86036 2150
rect 86092 2148 86116 2150
rect 86172 2148 86196 2150
rect 85956 2128 86252 2148
rect 86328 1222 86356 19887
rect 86406 13968 86462 13977
rect 86406 13903 86462 13912
rect 86316 1216 86368 1222
rect 86316 1158 86368 1164
rect 85488 1012 85540 1018
rect 85488 954 85540 960
rect 85212 876 85264 882
rect 85212 818 85264 824
rect 85120 740 85172 746
rect 85120 682 85172 688
rect 84844 672 84896 678
rect 84844 614 84896 620
rect 83832 468 83884 474
rect 83832 410 83884 416
rect 83740 400 83792 406
rect 83740 342 83792 348
rect 81440 332 81492 338
rect 81440 274 81492 280
rect 55036 264 55088 270
rect 55036 206 55088 212
rect 81348 264 81400 270
rect 81348 206 81400 212
rect 86420 134 86448 13903
rect 86498 10160 86554 10169
rect 86498 10095 86554 10104
rect 86512 202 86540 10095
rect 86604 1154 86632 30767
rect 86592 1148 86644 1154
rect 86592 1090 86644 1096
rect 86696 814 86724 38247
rect 86774 33416 86830 33425
rect 86774 33351 86830 33360
rect 86788 950 86816 33351
rect 86880 1737 86908 70366
rect 87144 69012 87196 69018
rect 87144 68954 87196 68960
rect 87156 68785 87184 68954
rect 87142 68776 87198 68785
rect 87142 68711 87198 68720
rect 87340 67289 87368 80003
rect 87418 79928 87474 79937
rect 87418 79863 87474 79872
rect 87432 75546 87460 79863
rect 87420 75540 87472 75546
rect 87420 75482 87472 75488
rect 87420 75268 87472 75274
rect 87420 75210 87472 75216
rect 87326 67280 87382 67289
rect 87326 67215 87382 67224
rect 87328 66156 87380 66162
rect 87328 66098 87380 66104
rect 87340 64977 87368 66098
rect 87326 64968 87382 64977
rect 87326 64903 87382 64912
rect 87432 58993 87460 75210
rect 87524 63889 87552 80026
rect 87510 63880 87566 63889
rect 87510 63815 87566 63824
rect 87418 58984 87474 58993
rect 87418 58919 87474 58928
rect 86960 57928 87012 57934
rect 86958 57896 86960 57905
rect 87012 57896 87014 57905
rect 86958 57831 87014 57840
rect 86960 56500 87012 56506
rect 86960 56442 87012 56448
rect 86972 55321 87000 56442
rect 87052 56432 87104 56438
rect 87050 56400 87052 56409
rect 87104 56400 87106 56409
rect 87050 56335 87106 56344
rect 86958 55312 87014 55321
rect 86958 55247 87014 55256
rect 86960 54664 87012 54670
rect 86960 54606 87012 54612
rect 86972 54097 87000 54606
rect 86958 54088 87014 54097
rect 86958 54023 87014 54032
rect 86960 53780 87012 53786
rect 86960 53722 87012 53728
rect 86972 53009 87000 53722
rect 86958 53000 87014 53009
rect 86958 52935 87014 52944
rect 87616 48113 87644 93758
rect 87708 85241 87736 93774
rect 87694 85232 87750 85241
rect 87694 85167 87750 85176
rect 87800 84946 87828 93978
rect 87708 84918 87828 84946
rect 87708 60081 87736 84918
rect 87786 84824 87842 84833
rect 87786 84759 87842 84768
rect 87800 75274 87828 84759
rect 87788 75268 87840 75274
rect 87788 75210 87840 75216
rect 87788 70372 87840 70378
rect 87788 70314 87840 70320
rect 87800 69873 87828 70314
rect 87786 69864 87842 69873
rect 87786 69799 87842 69808
rect 87788 66224 87840 66230
rect 87786 66192 87788 66201
rect 87840 66192 87842 66201
rect 87786 66127 87842 66136
rect 87788 63504 87840 63510
rect 87788 63446 87840 63452
rect 87800 62801 87828 63446
rect 87786 62792 87842 62801
rect 87786 62727 87842 62736
rect 87788 61940 87840 61946
rect 87788 61882 87840 61888
rect 87800 61305 87828 61882
rect 87786 61296 87842 61305
rect 87786 61231 87842 61240
rect 87694 60072 87750 60081
rect 87694 60007 87750 60016
rect 87696 49700 87748 49706
rect 87696 49642 87748 49648
rect 87708 49201 87736 49642
rect 87694 49192 87750 49201
rect 87694 49127 87750 49136
rect 87602 48104 87658 48113
rect 87602 48039 87658 48048
rect 87694 46608 87750 46617
rect 87694 46543 87750 46552
rect 87708 45626 87736 46543
rect 87696 45620 87748 45626
rect 87696 45562 87748 45568
rect 87602 45520 87658 45529
rect 87602 45455 87658 45464
rect 87328 40724 87380 40730
rect 87328 40666 87380 40672
rect 86958 36816 87014 36825
rect 86958 36751 87014 36760
rect 86972 36378 87000 36751
rect 86960 36372 87012 36378
rect 86960 36314 87012 36320
rect 87340 35894 87368 40666
rect 87510 39400 87566 39409
rect 87510 39335 87566 39344
rect 87248 35866 87368 35894
rect 86958 34640 87014 34649
rect 86958 34575 87014 34584
rect 86972 34542 87000 34575
rect 86960 34536 87012 34542
rect 86960 34478 87012 34484
rect 86958 31920 87014 31929
rect 86958 31855 87014 31864
rect 86972 31822 87000 31855
rect 86960 31816 87012 31822
rect 86960 31758 87012 31764
rect 87248 30326 87276 35866
rect 87326 35728 87382 35737
rect 87326 35663 87382 35672
rect 87340 31754 87368 35663
rect 87340 31726 87460 31754
rect 87236 30320 87288 30326
rect 87236 30262 87288 30268
rect 86958 29744 87014 29753
rect 86958 29679 87014 29688
rect 86972 29034 87000 29679
rect 86960 29028 87012 29034
rect 86960 28970 87012 28976
rect 86958 28520 87014 28529
rect 86958 28455 87014 28464
rect 86972 27674 87000 28455
rect 86960 27668 87012 27674
rect 86960 27610 87012 27616
rect 86958 27024 87014 27033
rect 86958 26959 87014 26968
rect 86972 26314 87000 26959
rect 86960 26308 87012 26314
rect 86960 26250 87012 26256
rect 87234 25936 87290 25945
rect 87234 25871 87290 25880
rect 86958 24848 87014 24857
rect 86958 24783 87014 24792
rect 86972 23526 87000 24783
rect 87050 23624 87106 23633
rect 87050 23559 87052 23568
rect 87104 23559 87106 23568
rect 87052 23530 87104 23536
rect 86960 23520 87012 23526
rect 86960 23462 87012 23468
rect 87142 22536 87198 22545
rect 87142 22471 87198 22480
rect 87156 22234 87184 22471
rect 87144 22228 87196 22234
rect 87144 22170 87196 22176
rect 87248 20602 87276 25871
rect 87236 20596 87288 20602
rect 87236 20538 87288 20544
rect 87142 18864 87198 18873
rect 87142 18799 87198 18808
rect 87052 16584 87104 16590
rect 87052 16526 87104 16532
rect 87064 15178 87092 16526
rect 87156 16402 87184 18799
rect 87234 17640 87290 17649
rect 87234 17575 87290 17584
rect 87248 16590 87276 17575
rect 87236 16584 87288 16590
rect 87236 16526 87288 16532
rect 87156 16374 87368 16402
rect 87142 16144 87198 16153
rect 87142 16079 87198 16088
rect 87156 15366 87184 16079
rect 87144 15360 87196 15366
rect 87144 15302 87196 15308
rect 87064 15150 87276 15178
rect 87142 15056 87198 15065
rect 87142 14991 87198 15000
rect 86958 12744 87014 12753
rect 86958 12679 87014 12688
rect 86972 12646 87000 12679
rect 86960 12640 87012 12646
rect 86960 12582 87012 12588
rect 86958 11248 87014 11257
rect 86958 11183 87014 11192
rect 86972 11082 87000 11183
rect 86960 11076 87012 11082
rect 86960 11018 87012 11024
rect 86958 9072 87014 9081
rect 86958 9007 87014 9016
rect 86972 8362 87000 9007
rect 86960 8356 87012 8362
rect 86960 8298 87012 8304
rect 87052 8288 87104 8294
rect 87052 8230 87104 8236
rect 86960 7540 87012 7546
rect 86960 7482 87012 7488
rect 86972 2666 87000 7482
rect 87064 5370 87092 8230
rect 87052 5364 87104 5370
rect 87052 5306 87104 5312
rect 87050 5264 87106 5273
rect 87050 5199 87106 5208
rect 87064 4214 87092 5199
rect 87052 4208 87104 4214
rect 87052 4150 87104 4156
rect 87052 3460 87104 3466
rect 87052 3402 87104 3408
rect 87064 2961 87092 3402
rect 87050 2952 87106 2961
rect 87050 2887 87106 2896
rect 86972 2638 87092 2666
rect 86960 2440 87012 2446
rect 86960 2382 87012 2388
rect 86866 1728 86922 1737
rect 86866 1663 86922 1672
rect 86776 944 86828 950
rect 86776 886 86828 892
rect 86684 808 86736 814
rect 86684 750 86736 756
rect 86972 649 87000 2382
rect 87064 1698 87092 2638
rect 87156 2582 87184 14991
rect 87248 7546 87276 15150
rect 87340 7546 87368 16374
rect 87236 7540 87288 7546
rect 87236 7482 87288 7488
rect 87328 7540 87380 7546
rect 87328 7482 87380 7488
rect 87236 7404 87288 7410
rect 87236 7346 87288 7352
rect 87144 2576 87196 2582
rect 87144 2518 87196 2524
rect 87248 2514 87276 7346
rect 87326 6352 87382 6361
rect 87326 6287 87382 6296
rect 87340 3126 87368 6287
rect 87328 3120 87380 3126
rect 87328 3062 87380 3068
rect 87328 2916 87380 2922
rect 87328 2858 87380 2864
rect 87340 2650 87368 2858
rect 87328 2644 87380 2650
rect 87328 2586 87380 2592
rect 87236 2508 87288 2514
rect 87236 2450 87288 2456
rect 87432 1766 87460 31726
rect 87524 2922 87552 39335
rect 87616 8294 87644 45455
rect 87694 44296 87750 44305
rect 87694 44231 87750 44240
rect 87708 44198 87736 44231
rect 87696 44192 87748 44198
rect 87696 44134 87748 44140
rect 87694 43208 87750 43217
rect 87694 43143 87750 43152
rect 87604 8288 87656 8294
rect 87604 8230 87656 8236
rect 87708 8106 87736 43143
rect 87786 41712 87842 41721
rect 87786 41647 87842 41656
rect 87616 8078 87736 8106
rect 87800 8090 87828 41647
rect 87892 40730 87920 97650
rect 87984 97646 88012 97838
rect 87972 97640 88024 97646
rect 88720 97617 88748 104314
rect 87972 97582 88024 97588
rect 88706 97608 88762 97617
rect 88706 97543 88762 97552
rect 87956 97404 88252 97424
rect 88012 97402 88036 97404
rect 88092 97402 88116 97404
rect 88172 97402 88196 97404
rect 88034 97350 88036 97402
rect 88098 97350 88110 97402
rect 88172 97350 88174 97402
rect 88012 97348 88036 97350
rect 88092 97348 88116 97350
rect 88172 97348 88196 97350
rect 87956 97328 88252 97348
rect 88996 96490 89024 118351
rect 89956 117532 90252 117552
rect 90012 117530 90036 117532
rect 90092 117530 90116 117532
rect 90172 117530 90196 117532
rect 90034 117478 90036 117530
rect 90098 117478 90110 117530
rect 90172 117478 90174 117530
rect 90012 117476 90036 117478
rect 90092 117476 90116 117478
rect 90172 117476 90196 117478
rect 89956 117456 90252 117476
rect 89956 116444 90252 116464
rect 90012 116442 90036 116444
rect 90092 116442 90116 116444
rect 90172 116442 90196 116444
rect 90034 116390 90036 116442
rect 90098 116390 90110 116442
rect 90172 116390 90174 116442
rect 90012 116388 90036 116390
rect 90092 116388 90116 116390
rect 90172 116388 90196 116390
rect 89956 116368 90252 116388
rect 89956 115356 90252 115376
rect 90012 115354 90036 115356
rect 90092 115354 90116 115356
rect 90172 115354 90196 115356
rect 90034 115302 90036 115354
rect 90098 115302 90110 115354
rect 90172 115302 90174 115354
rect 90012 115300 90036 115302
rect 90092 115300 90116 115302
rect 90172 115300 90196 115302
rect 89956 115280 90252 115300
rect 89956 114268 90252 114288
rect 90012 114266 90036 114268
rect 90092 114266 90116 114268
rect 90172 114266 90196 114268
rect 90034 114214 90036 114266
rect 90098 114214 90110 114266
rect 90172 114214 90174 114266
rect 90012 114212 90036 114214
rect 90092 114212 90116 114214
rect 90172 114212 90196 114214
rect 89956 114192 90252 114212
rect 89956 113180 90252 113200
rect 90012 113178 90036 113180
rect 90092 113178 90116 113180
rect 90172 113178 90196 113180
rect 90034 113126 90036 113178
rect 90098 113126 90110 113178
rect 90172 113126 90174 113178
rect 90012 113124 90036 113126
rect 90092 113124 90116 113126
rect 90172 113124 90196 113126
rect 89956 113104 90252 113124
rect 89956 112092 90252 112112
rect 90012 112090 90036 112092
rect 90092 112090 90116 112092
rect 90172 112090 90196 112092
rect 90034 112038 90036 112090
rect 90098 112038 90110 112090
rect 90172 112038 90174 112090
rect 90012 112036 90036 112038
rect 90092 112036 90116 112038
rect 90172 112036 90196 112038
rect 89956 112016 90252 112036
rect 89956 111004 90252 111024
rect 90012 111002 90036 111004
rect 90092 111002 90116 111004
rect 90172 111002 90196 111004
rect 90034 110950 90036 111002
rect 90098 110950 90110 111002
rect 90172 110950 90174 111002
rect 90012 110948 90036 110950
rect 90092 110948 90116 110950
rect 90172 110948 90196 110950
rect 89956 110928 90252 110948
rect 89956 109916 90252 109936
rect 90012 109914 90036 109916
rect 90092 109914 90116 109916
rect 90172 109914 90196 109916
rect 90034 109862 90036 109914
rect 90098 109862 90110 109914
rect 90172 109862 90174 109914
rect 90012 109860 90036 109862
rect 90092 109860 90116 109862
rect 90172 109860 90196 109862
rect 89956 109840 90252 109860
rect 89956 108828 90252 108848
rect 90012 108826 90036 108828
rect 90092 108826 90116 108828
rect 90172 108826 90196 108828
rect 90034 108774 90036 108826
rect 90098 108774 90110 108826
rect 90172 108774 90174 108826
rect 90012 108772 90036 108774
rect 90092 108772 90116 108774
rect 90172 108772 90196 108774
rect 89956 108752 90252 108772
rect 89956 107740 90252 107760
rect 90012 107738 90036 107740
rect 90092 107738 90116 107740
rect 90172 107738 90196 107740
rect 90034 107686 90036 107738
rect 90098 107686 90110 107738
rect 90172 107686 90174 107738
rect 90012 107684 90036 107686
rect 90092 107684 90116 107686
rect 90172 107684 90196 107686
rect 89956 107664 90252 107684
rect 89956 106652 90252 106672
rect 90012 106650 90036 106652
rect 90092 106650 90116 106652
rect 90172 106650 90196 106652
rect 90034 106598 90036 106650
rect 90098 106598 90110 106650
rect 90172 106598 90174 106650
rect 90012 106596 90036 106598
rect 90092 106596 90116 106598
rect 90172 106596 90196 106598
rect 89956 106576 90252 106596
rect 89956 105564 90252 105584
rect 90012 105562 90036 105564
rect 90092 105562 90116 105564
rect 90172 105562 90196 105564
rect 90034 105510 90036 105562
rect 90098 105510 90110 105562
rect 90172 105510 90174 105562
rect 90012 105508 90036 105510
rect 90092 105508 90116 105510
rect 90172 105508 90196 105510
rect 89956 105488 90252 105508
rect 89956 104476 90252 104496
rect 90012 104474 90036 104476
rect 90092 104474 90116 104476
rect 90172 104474 90196 104476
rect 90034 104422 90036 104474
rect 90098 104422 90110 104474
rect 90172 104422 90174 104474
rect 90012 104420 90036 104422
rect 90092 104420 90116 104422
rect 90172 104420 90196 104422
rect 89956 104400 90252 104420
rect 89956 103388 90252 103408
rect 90012 103386 90036 103388
rect 90092 103386 90116 103388
rect 90172 103386 90196 103388
rect 90034 103334 90036 103386
rect 90098 103334 90110 103386
rect 90172 103334 90174 103386
rect 90012 103332 90036 103334
rect 90092 103332 90116 103334
rect 90172 103332 90196 103334
rect 89956 103312 90252 103332
rect 89956 102300 90252 102320
rect 90012 102298 90036 102300
rect 90092 102298 90116 102300
rect 90172 102298 90196 102300
rect 90034 102246 90036 102298
rect 90098 102246 90110 102298
rect 90172 102246 90174 102298
rect 90012 102244 90036 102246
rect 90092 102244 90116 102246
rect 90172 102244 90196 102246
rect 89956 102224 90252 102244
rect 89956 101212 90252 101232
rect 90012 101210 90036 101212
rect 90092 101210 90116 101212
rect 90172 101210 90196 101212
rect 90034 101158 90036 101210
rect 90098 101158 90110 101210
rect 90172 101158 90174 101210
rect 90012 101156 90036 101158
rect 90092 101156 90116 101158
rect 90172 101156 90196 101158
rect 89956 101136 90252 101156
rect 90362 100192 90418 100201
rect 89956 100124 90252 100144
rect 90362 100127 90418 100136
rect 90012 100122 90036 100124
rect 90092 100122 90116 100124
rect 90172 100122 90196 100124
rect 90034 100070 90036 100122
rect 90098 100070 90110 100122
rect 90172 100070 90174 100122
rect 90012 100068 90036 100070
rect 90092 100068 90116 100070
rect 90172 100068 90196 100070
rect 89956 100048 90252 100068
rect 89956 99036 90252 99056
rect 90012 99034 90036 99036
rect 90092 99034 90116 99036
rect 90172 99034 90196 99036
rect 90034 98982 90036 99034
rect 90098 98982 90110 99034
rect 90172 98982 90174 99034
rect 90012 98980 90036 98982
rect 90092 98980 90116 98982
rect 90172 98980 90196 98982
rect 89956 98960 90252 98980
rect 89956 97948 90252 97968
rect 90012 97946 90036 97948
rect 90092 97946 90116 97948
rect 90172 97946 90196 97948
rect 90034 97894 90036 97946
rect 90098 97894 90110 97946
rect 90172 97894 90174 97946
rect 90012 97892 90036 97894
rect 90092 97892 90116 97894
rect 90172 97892 90196 97894
rect 89956 97872 90252 97892
rect 90376 97714 90404 100127
rect 90364 97708 90416 97714
rect 90364 97650 90416 97656
rect 89956 96860 90252 96880
rect 90012 96858 90036 96860
rect 90092 96858 90116 96860
rect 90172 96858 90196 96860
rect 90034 96806 90036 96858
rect 90098 96806 90110 96858
rect 90172 96806 90174 96858
rect 90012 96804 90036 96806
rect 90092 96804 90116 96806
rect 90172 96804 90196 96806
rect 89956 96784 90252 96804
rect 88984 96484 89036 96490
rect 88984 96426 89036 96432
rect 87956 96316 88252 96336
rect 88012 96314 88036 96316
rect 88092 96314 88116 96316
rect 88172 96314 88196 96316
rect 88034 96262 88036 96314
rect 88098 96262 88110 96314
rect 88172 96262 88174 96314
rect 88012 96260 88036 96262
rect 88092 96260 88116 96262
rect 88172 96260 88196 96262
rect 87956 96240 88252 96260
rect 89956 95772 90252 95792
rect 90012 95770 90036 95772
rect 90092 95770 90116 95772
rect 90172 95770 90196 95772
rect 90034 95718 90036 95770
rect 90098 95718 90110 95770
rect 90172 95718 90174 95770
rect 90012 95716 90036 95718
rect 90092 95716 90116 95718
rect 90172 95716 90196 95718
rect 89956 95696 90252 95716
rect 87956 95228 88252 95248
rect 88012 95226 88036 95228
rect 88092 95226 88116 95228
rect 88172 95226 88196 95228
rect 88034 95174 88036 95226
rect 88098 95174 88110 95226
rect 88172 95174 88174 95226
rect 88012 95172 88036 95174
rect 88092 95172 88116 95174
rect 88172 95172 88196 95174
rect 87956 95152 88252 95172
rect 89956 94684 90252 94704
rect 90012 94682 90036 94684
rect 90092 94682 90116 94684
rect 90172 94682 90196 94684
rect 90034 94630 90036 94682
rect 90098 94630 90110 94682
rect 90172 94630 90174 94682
rect 90012 94628 90036 94630
rect 90092 94628 90116 94630
rect 90172 94628 90196 94630
rect 89956 94608 90252 94628
rect 87956 94140 88252 94160
rect 88012 94138 88036 94140
rect 88092 94138 88116 94140
rect 88172 94138 88196 94140
rect 88034 94086 88036 94138
rect 88098 94086 88110 94138
rect 88172 94086 88174 94138
rect 88012 94084 88036 94086
rect 88092 94084 88116 94086
rect 88172 94084 88196 94086
rect 87956 94064 88252 94084
rect 89956 93596 90252 93616
rect 90012 93594 90036 93596
rect 90092 93594 90116 93596
rect 90172 93594 90196 93596
rect 90034 93542 90036 93594
rect 90098 93542 90110 93594
rect 90172 93542 90174 93594
rect 90012 93540 90036 93542
rect 90092 93540 90116 93542
rect 90172 93540 90196 93542
rect 89956 93520 90252 93540
rect 87956 93052 88252 93072
rect 88012 93050 88036 93052
rect 88092 93050 88116 93052
rect 88172 93050 88196 93052
rect 88034 92998 88036 93050
rect 88098 92998 88110 93050
rect 88172 92998 88174 93050
rect 88012 92996 88036 92998
rect 88092 92996 88116 92998
rect 88172 92996 88196 92998
rect 87956 92976 88252 92996
rect 89956 92508 90252 92528
rect 90012 92506 90036 92508
rect 90092 92506 90116 92508
rect 90172 92506 90196 92508
rect 90034 92454 90036 92506
rect 90098 92454 90110 92506
rect 90172 92454 90174 92506
rect 90012 92452 90036 92454
rect 90092 92452 90116 92454
rect 90172 92452 90196 92454
rect 89956 92432 90252 92452
rect 87956 91964 88252 91984
rect 88012 91962 88036 91964
rect 88092 91962 88116 91964
rect 88172 91962 88196 91964
rect 88034 91910 88036 91962
rect 88098 91910 88110 91962
rect 88172 91910 88174 91962
rect 88012 91908 88036 91910
rect 88092 91908 88116 91910
rect 88172 91908 88196 91910
rect 87956 91888 88252 91908
rect 88340 91792 88392 91798
rect 88340 91734 88392 91740
rect 87956 90876 88252 90896
rect 88012 90874 88036 90876
rect 88092 90874 88116 90876
rect 88172 90874 88196 90876
rect 88034 90822 88036 90874
rect 88098 90822 88110 90874
rect 88172 90822 88174 90874
rect 88012 90820 88036 90822
rect 88092 90820 88116 90822
rect 88172 90820 88196 90822
rect 87956 90800 88252 90820
rect 87956 89788 88252 89808
rect 88012 89786 88036 89788
rect 88092 89786 88116 89788
rect 88172 89786 88196 89788
rect 88034 89734 88036 89786
rect 88098 89734 88110 89786
rect 88172 89734 88174 89786
rect 88012 89732 88036 89734
rect 88092 89732 88116 89734
rect 88172 89732 88196 89734
rect 87956 89712 88252 89732
rect 88352 89690 88380 91734
rect 89956 91420 90252 91440
rect 90012 91418 90036 91420
rect 90092 91418 90116 91420
rect 90172 91418 90196 91420
rect 90034 91366 90036 91418
rect 90098 91366 90110 91418
rect 90172 91366 90174 91418
rect 90012 91364 90036 91366
rect 90092 91364 90116 91366
rect 90172 91364 90196 91366
rect 89956 91344 90252 91364
rect 89956 90332 90252 90352
rect 90012 90330 90036 90332
rect 90092 90330 90116 90332
rect 90172 90330 90196 90332
rect 90034 90278 90036 90330
rect 90098 90278 90110 90330
rect 90172 90278 90174 90330
rect 90012 90276 90036 90278
rect 90092 90276 90116 90278
rect 90172 90276 90196 90278
rect 89956 90256 90252 90276
rect 88340 89684 88392 89690
rect 88340 89626 88392 89632
rect 89956 89244 90252 89264
rect 90012 89242 90036 89244
rect 90092 89242 90116 89244
rect 90172 89242 90196 89244
rect 90034 89190 90036 89242
rect 90098 89190 90110 89242
rect 90172 89190 90174 89242
rect 90012 89188 90036 89190
rect 90092 89188 90116 89190
rect 90172 89188 90196 89190
rect 89956 89168 90252 89188
rect 87956 88700 88252 88720
rect 88012 88698 88036 88700
rect 88092 88698 88116 88700
rect 88172 88698 88196 88700
rect 88034 88646 88036 88698
rect 88098 88646 88110 88698
rect 88172 88646 88174 88698
rect 88012 88644 88036 88646
rect 88092 88644 88116 88646
rect 88172 88644 88196 88646
rect 87956 88624 88252 88644
rect 87972 88324 88024 88330
rect 87972 88266 88024 88272
rect 87984 87961 88012 88266
rect 89956 88156 90252 88176
rect 90012 88154 90036 88156
rect 90092 88154 90116 88156
rect 90172 88154 90196 88156
rect 90034 88102 90036 88154
rect 90098 88102 90110 88154
rect 90172 88102 90174 88154
rect 90012 88100 90036 88102
rect 90092 88100 90116 88102
rect 90172 88100 90196 88102
rect 89956 88080 90252 88100
rect 87970 87952 88026 87961
rect 87970 87887 88026 87896
rect 87956 87612 88252 87632
rect 88012 87610 88036 87612
rect 88092 87610 88116 87612
rect 88172 87610 88196 87612
rect 88034 87558 88036 87610
rect 88098 87558 88110 87610
rect 88172 87558 88174 87610
rect 88012 87556 88036 87558
rect 88092 87556 88116 87558
rect 88172 87556 88196 87558
rect 87956 87536 88252 87556
rect 89956 87068 90252 87088
rect 90012 87066 90036 87068
rect 90092 87066 90116 87068
rect 90172 87066 90196 87068
rect 90034 87014 90036 87066
rect 90098 87014 90110 87066
rect 90172 87014 90174 87066
rect 90012 87012 90036 87014
rect 90092 87012 90116 87014
rect 90172 87012 90196 87014
rect 89956 86992 90252 87012
rect 87956 86524 88252 86544
rect 88012 86522 88036 86524
rect 88092 86522 88116 86524
rect 88172 86522 88196 86524
rect 88034 86470 88036 86522
rect 88098 86470 88110 86522
rect 88172 86470 88174 86522
rect 88012 86468 88036 86470
rect 88092 86468 88116 86470
rect 88172 86468 88196 86470
rect 87956 86448 88252 86468
rect 87972 86352 88024 86358
rect 87972 86294 88024 86300
rect 87984 85649 88012 86294
rect 89956 85980 90252 86000
rect 90012 85978 90036 85980
rect 90092 85978 90116 85980
rect 90172 85978 90196 85980
rect 90034 85926 90036 85978
rect 90098 85926 90110 85978
rect 90172 85926 90174 85978
rect 90012 85924 90036 85926
rect 90092 85924 90116 85926
rect 90172 85924 90196 85926
rect 89956 85904 90252 85924
rect 87970 85640 88026 85649
rect 87970 85575 88026 85584
rect 87956 85436 88252 85456
rect 88012 85434 88036 85436
rect 88092 85434 88116 85436
rect 88172 85434 88196 85436
rect 88034 85382 88036 85434
rect 88098 85382 88110 85434
rect 88172 85382 88174 85434
rect 88012 85380 88036 85382
rect 88092 85380 88116 85382
rect 88172 85380 88196 85382
rect 87956 85360 88252 85380
rect 87972 85264 88024 85270
rect 87972 85206 88024 85212
rect 87984 84561 88012 85206
rect 89956 84892 90252 84912
rect 90012 84890 90036 84892
rect 90092 84890 90116 84892
rect 90172 84890 90196 84892
rect 90034 84838 90036 84890
rect 90098 84838 90110 84890
rect 90172 84838 90174 84890
rect 90012 84836 90036 84838
rect 90092 84836 90116 84838
rect 90172 84836 90196 84838
rect 89956 84816 90252 84836
rect 87970 84552 88026 84561
rect 87970 84487 88026 84496
rect 87956 84348 88252 84368
rect 88012 84346 88036 84348
rect 88092 84346 88116 84348
rect 88172 84346 88196 84348
rect 88034 84294 88036 84346
rect 88098 84294 88110 84346
rect 88172 84294 88174 84346
rect 88012 84292 88036 84294
rect 88092 84292 88116 84294
rect 88172 84292 88196 84294
rect 87956 84272 88252 84292
rect 87972 84176 88024 84182
rect 87972 84118 88024 84124
rect 87984 83473 88012 84118
rect 89956 83804 90252 83824
rect 90012 83802 90036 83804
rect 90092 83802 90116 83804
rect 90172 83802 90196 83804
rect 90034 83750 90036 83802
rect 90098 83750 90110 83802
rect 90172 83750 90174 83802
rect 90012 83748 90036 83750
rect 90092 83748 90116 83750
rect 90172 83748 90196 83750
rect 89956 83728 90252 83748
rect 87970 83464 88026 83473
rect 87970 83399 88026 83408
rect 87956 83260 88252 83280
rect 88012 83258 88036 83260
rect 88092 83258 88116 83260
rect 88172 83258 88196 83260
rect 88034 83206 88036 83258
rect 88098 83206 88110 83258
rect 88172 83206 88174 83258
rect 88012 83204 88036 83206
rect 88092 83204 88116 83206
rect 88172 83204 88196 83206
rect 87956 83184 88252 83204
rect 89956 82716 90252 82736
rect 90012 82714 90036 82716
rect 90092 82714 90116 82716
rect 90172 82714 90196 82716
rect 90034 82662 90036 82714
rect 90098 82662 90110 82714
rect 90172 82662 90174 82714
rect 90012 82660 90036 82662
rect 90092 82660 90116 82662
rect 90172 82660 90196 82662
rect 89956 82640 90252 82660
rect 87956 82172 88252 82192
rect 88012 82170 88036 82172
rect 88092 82170 88116 82172
rect 88172 82170 88196 82172
rect 88034 82118 88036 82170
rect 88098 82118 88110 82170
rect 88172 82118 88174 82170
rect 88012 82116 88036 82118
rect 88092 82116 88116 82118
rect 88172 82116 88196 82118
rect 87956 82096 88252 82116
rect 87972 82000 88024 82006
rect 87970 81968 87972 81977
rect 88024 81968 88026 81977
rect 87970 81903 88026 81912
rect 89956 81628 90252 81648
rect 90012 81626 90036 81628
rect 90092 81626 90116 81628
rect 90172 81626 90196 81628
rect 90034 81574 90036 81626
rect 90098 81574 90110 81626
rect 90172 81574 90174 81626
rect 90012 81572 90036 81574
rect 90092 81572 90116 81574
rect 90172 81572 90196 81574
rect 89956 81552 90252 81572
rect 87956 81084 88252 81104
rect 88012 81082 88036 81084
rect 88092 81082 88116 81084
rect 88172 81082 88196 81084
rect 88034 81030 88036 81082
rect 88098 81030 88110 81082
rect 88172 81030 88174 81082
rect 88012 81028 88036 81030
rect 88092 81028 88116 81030
rect 88172 81028 88196 81030
rect 87956 81008 88252 81028
rect 87972 80912 88024 80918
rect 87972 80854 88024 80860
rect 87984 80753 88012 80854
rect 87970 80744 88026 80753
rect 87970 80679 88026 80688
rect 89956 80540 90252 80560
rect 90012 80538 90036 80540
rect 90092 80538 90116 80540
rect 90172 80538 90196 80540
rect 90034 80486 90036 80538
rect 90098 80486 90110 80538
rect 90172 80486 90174 80538
rect 90012 80484 90036 80486
rect 90092 80484 90116 80486
rect 90172 80484 90196 80486
rect 89956 80464 90252 80484
rect 88340 80164 88392 80170
rect 88340 80106 88392 80112
rect 87956 79996 88252 80016
rect 88012 79994 88036 79996
rect 88092 79994 88116 79996
rect 88172 79994 88196 79996
rect 88034 79942 88036 79994
rect 88098 79942 88110 79994
rect 88172 79942 88174 79994
rect 88012 79940 88036 79942
rect 88092 79940 88116 79942
rect 88172 79940 88196 79942
rect 87956 79920 88252 79940
rect 88352 79778 88380 80106
rect 88260 79750 88380 79778
rect 88260 79665 88288 79750
rect 88246 79656 88302 79665
rect 88246 79591 88302 79600
rect 89956 79452 90252 79472
rect 90012 79450 90036 79452
rect 90092 79450 90116 79452
rect 90172 79450 90196 79452
rect 90034 79398 90036 79450
rect 90098 79398 90110 79450
rect 90172 79398 90174 79450
rect 90012 79396 90036 79398
rect 90092 79396 90116 79398
rect 90172 79396 90196 79398
rect 89956 79376 90252 79396
rect 87956 78908 88252 78928
rect 88012 78906 88036 78908
rect 88092 78906 88116 78908
rect 88172 78906 88196 78908
rect 88034 78854 88036 78906
rect 88098 78854 88110 78906
rect 88172 78854 88174 78906
rect 88012 78852 88036 78854
rect 88092 78852 88116 78854
rect 88172 78852 88196 78854
rect 87956 78832 88252 78852
rect 89956 78364 90252 78384
rect 90012 78362 90036 78364
rect 90092 78362 90116 78364
rect 90172 78362 90196 78364
rect 90034 78310 90036 78362
rect 90098 78310 90110 78362
rect 90172 78310 90174 78362
rect 90012 78308 90036 78310
rect 90092 78308 90116 78310
rect 90172 78308 90196 78310
rect 89956 78288 90252 78308
rect 87956 77820 88252 77840
rect 88012 77818 88036 77820
rect 88092 77818 88116 77820
rect 88172 77818 88196 77820
rect 88034 77766 88036 77818
rect 88098 77766 88110 77818
rect 88172 77766 88174 77818
rect 88012 77764 88036 77766
rect 88092 77764 88116 77766
rect 88172 77764 88196 77766
rect 87956 77744 88252 77764
rect 89956 77276 90252 77296
rect 90012 77274 90036 77276
rect 90092 77274 90116 77276
rect 90172 77274 90196 77276
rect 90034 77222 90036 77274
rect 90098 77222 90110 77274
rect 90172 77222 90174 77274
rect 90012 77220 90036 77222
rect 90092 77220 90116 77222
rect 90172 77220 90196 77222
rect 89956 77200 90252 77220
rect 87956 76732 88252 76752
rect 88012 76730 88036 76732
rect 88092 76730 88116 76732
rect 88172 76730 88196 76732
rect 88034 76678 88036 76730
rect 88098 76678 88110 76730
rect 88172 76678 88174 76730
rect 88012 76676 88036 76678
rect 88092 76676 88116 76678
rect 88172 76676 88196 76678
rect 87956 76656 88252 76676
rect 89956 76188 90252 76208
rect 90012 76186 90036 76188
rect 90092 76186 90116 76188
rect 90172 76186 90196 76188
rect 90034 76134 90036 76186
rect 90098 76134 90110 76186
rect 90172 76134 90174 76186
rect 90012 76132 90036 76134
rect 90092 76132 90116 76134
rect 90172 76132 90196 76134
rect 89956 76112 90252 76132
rect 87956 75644 88252 75664
rect 88012 75642 88036 75644
rect 88092 75642 88116 75644
rect 88172 75642 88196 75644
rect 88034 75590 88036 75642
rect 88098 75590 88110 75642
rect 88172 75590 88174 75642
rect 88012 75588 88036 75590
rect 88092 75588 88116 75590
rect 88172 75588 88196 75590
rect 87956 75568 88252 75588
rect 89956 75100 90252 75120
rect 90012 75098 90036 75100
rect 90092 75098 90116 75100
rect 90172 75098 90196 75100
rect 90034 75046 90036 75098
rect 90098 75046 90110 75098
rect 90172 75046 90174 75098
rect 90012 75044 90036 75046
rect 90092 75044 90116 75046
rect 90172 75044 90196 75046
rect 89956 75024 90252 75044
rect 87956 74556 88252 74576
rect 88012 74554 88036 74556
rect 88092 74554 88116 74556
rect 88172 74554 88196 74556
rect 88034 74502 88036 74554
rect 88098 74502 88110 74554
rect 88172 74502 88174 74554
rect 88012 74500 88036 74502
rect 88092 74500 88116 74502
rect 88172 74500 88196 74502
rect 87956 74480 88252 74500
rect 89956 74012 90252 74032
rect 90012 74010 90036 74012
rect 90092 74010 90116 74012
rect 90172 74010 90196 74012
rect 90034 73958 90036 74010
rect 90098 73958 90110 74010
rect 90172 73958 90174 74010
rect 90012 73956 90036 73958
rect 90092 73956 90116 73958
rect 90172 73956 90196 73958
rect 89956 73936 90252 73956
rect 87956 73468 88252 73488
rect 88012 73466 88036 73468
rect 88092 73466 88116 73468
rect 88172 73466 88196 73468
rect 88034 73414 88036 73466
rect 88098 73414 88110 73466
rect 88172 73414 88174 73466
rect 88012 73412 88036 73414
rect 88092 73412 88116 73414
rect 88172 73412 88196 73414
rect 87956 73392 88252 73412
rect 89956 72924 90252 72944
rect 90012 72922 90036 72924
rect 90092 72922 90116 72924
rect 90172 72922 90196 72924
rect 90034 72870 90036 72922
rect 90098 72870 90110 72922
rect 90172 72870 90174 72922
rect 90012 72868 90036 72870
rect 90092 72868 90116 72870
rect 90172 72868 90196 72870
rect 89956 72848 90252 72868
rect 87956 72380 88252 72400
rect 88012 72378 88036 72380
rect 88092 72378 88116 72380
rect 88172 72378 88196 72380
rect 88034 72326 88036 72378
rect 88098 72326 88110 72378
rect 88172 72326 88174 72378
rect 88012 72324 88036 72326
rect 88092 72324 88116 72326
rect 88172 72324 88196 72326
rect 87956 72304 88252 72324
rect 89956 71836 90252 71856
rect 90012 71834 90036 71836
rect 90092 71834 90116 71836
rect 90172 71834 90196 71836
rect 90034 71782 90036 71834
rect 90098 71782 90110 71834
rect 90172 71782 90174 71834
rect 90012 71780 90036 71782
rect 90092 71780 90116 71782
rect 90172 71780 90196 71782
rect 89956 71760 90252 71780
rect 87956 71292 88252 71312
rect 88012 71290 88036 71292
rect 88092 71290 88116 71292
rect 88172 71290 88196 71292
rect 88034 71238 88036 71290
rect 88098 71238 88110 71290
rect 88172 71238 88174 71290
rect 88012 71236 88036 71238
rect 88092 71236 88116 71238
rect 88172 71236 88196 71238
rect 87956 71216 88252 71236
rect 89956 70748 90252 70768
rect 90012 70746 90036 70748
rect 90092 70746 90116 70748
rect 90172 70746 90196 70748
rect 90034 70694 90036 70746
rect 90098 70694 90110 70746
rect 90172 70694 90174 70746
rect 90012 70692 90036 70694
rect 90092 70692 90116 70694
rect 90172 70692 90196 70694
rect 89956 70672 90252 70692
rect 87956 70204 88252 70224
rect 88012 70202 88036 70204
rect 88092 70202 88116 70204
rect 88172 70202 88196 70204
rect 88034 70150 88036 70202
rect 88098 70150 88110 70202
rect 88172 70150 88174 70202
rect 88012 70148 88036 70150
rect 88092 70148 88116 70150
rect 88172 70148 88196 70150
rect 87956 70128 88252 70148
rect 89956 69660 90252 69680
rect 90012 69658 90036 69660
rect 90092 69658 90116 69660
rect 90172 69658 90196 69660
rect 90034 69606 90036 69658
rect 90098 69606 90110 69658
rect 90172 69606 90174 69658
rect 90012 69604 90036 69606
rect 90092 69604 90116 69606
rect 90172 69604 90196 69606
rect 89956 69584 90252 69604
rect 87956 69116 88252 69136
rect 88012 69114 88036 69116
rect 88092 69114 88116 69116
rect 88172 69114 88196 69116
rect 88034 69062 88036 69114
rect 88098 69062 88110 69114
rect 88172 69062 88174 69114
rect 88012 69060 88036 69062
rect 88092 69060 88116 69062
rect 88172 69060 88196 69062
rect 87956 69040 88252 69060
rect 89956 68572 90252 68592
rect 90012 68570 90036 68572
rect 90092 68570 90116 68572
rect 90172 68570 90196 68572
rect 90034 68518 90036 68570
rect 90098 68518 90110 68570
rect 90172 68518 90174 68570
rect 90012 68516 90036 68518
rect 90092 68516 90116 68518
rect 90172 68516 90196 68518
rect 89956 68496 90252 68516
rect 87956 68028 88252 68048
rect 88012 68026 88036 68028
rect 88092 68026 88116 68028
rect 88172 68026 88196 68028
rect 88034 67974 88036 68026
rect 88098 67974 88110 68026
rect 88172 67974 88174 68026
rect 88012 67972 88036 67974
rect 88092 67972 88116 67974
rect 88172 67972 88196 67974
rect 87956 67952 88252 67972
rect 89956 67484 90252 67504
rect 90012 67482 90036 67484
rect 90092 67482 90116 67484
rect 90172 67482 90196 67484
rect 90034 67430 90036 67482
rect 90098 67430 90110 67482
rect 90172 67430 90174 67482
rect 90012 67428 90036 67430
rect 90092 67428 90116 67430
rect 90172 67428 90196 67430
rect 89956 67408 90252 67428
rect 87956 66940 88252 66960
rect 88012 66938 88036 66940
rect 88092 66938 88116 66940
rect 88172 66938 88196 66940
rect 88034 66886 88036 66938
rect 88098 66886 88110 66938
rect 88172 66886 88174 66938
rect 88012 66884 88036 66886
rect 88092 66884 88116 66886
rect 88172 66884 88196 66886
rect 87956 66864 88252 66884
rect 89956 66396 90252 66416
rect 90012 66394 90036 66396
rect 90092 66394 90116 66396
rect 90172 66394 90196 66396
rect 90034 66342 90036 66394
rect 90098 66342 90110 66394
rect 90172 66342 90174 66394
rect 90012 66340 90036 66342
rect 90092 66340 90116 66342
rect 90172 66340 90196 66342
rect 89956 66320 90252 66340
rect 87956 65852 88252 65872
rect 88012 65850 88036 65852
rect 88092 65850 88116 65852
rect 88172 65850 88196 65852
rect 88034 65798 88036 65850
rect 88098 65798 88110 65850
rect 88172 65798 88174 65850
rect 88012 65796 88036 65798
rect 88092 65796 88116 65798
rect 88172 65796 88196 65798
rect 87956 65776 88252 65796
rect 89956 65308 90252 65328
rect 90012 65306 90036 65308
rect 90092 65306 90116 65308
rect 90172 65306 90196 65308
rect 90034 65254 90036 65306
rect 90098 65254 90110 65306
rect 90172 65254 90174 65306
rect 90012 65252 90036 65254
rect 90092 65252 90116 65254
rect 90172 65252 90196 65254
rect 89956 65232 90252 65252
rect 87956 64764 88252 64784
rect 88012 64762 88036 64764
rect 88092 64762 88116 64764
rect 88172 64762 88196 64764
rect 88034 64710 88036 64762
rect 88098 64710 88110 64762
rect 88172 64710 88174 64762
rect 88012 64708 88036 64710
rect 88092 64708 88116 64710
rect 88172 64708 88196 64710
rect 87956 64688 88252 64708
rect 89956 64220 90252 64240
rect 90012 64218 90036 64220
rect 90092 64218 90116 64220
rect 90172 64218 90196 64220
rect 90034 64166 90036 64218
rect 90098 64166 90110 64218
rect 90172 64166 90174 64218
rect 90012 64164 90036 64166
rect 90092 64164 90116 64166
rect 90172 64164 90196 64166
rect 89956 64144 90252 64164
rect 87956 63676 88252 63696
rect 88012 63674 88036 63676
rect 88092 63674 88116 63676
rect 88172 63674 88196 63676
rect 88034 63622 88036 63674
rect 88098 63622 88110 63674
rect 88172 63622 88174 63674
rect 88012 63620 88036 63622
rect 88092 63620 88116 63622
rect 88172 63620 88196 63622
rect 87956 63600 88252 63620
rect 89956 63132 90252 63152
rect 90012 63130 90036 63132
rect 90092 63130 90116 63132
rect 90172 63130 90196 63132
rect 90034 63078 90036 63130
rect 90098 63078 90110 63130
rect 90172 63078 90174 63130
rect 90012 63076 90036 63078
rect 90092 63076 90116 63078
rect 90172 63076 90196 63078
rect 89956 63056 90252 63076
rect 87956 62588 88252 62608
rect 88012 62586 88036 62588
rect 88092 62586 88116 62588
rect 88172 62586 88196 62588
rect 88034 62534 88036 62586
rect 88098 62534 88110 62586
rect 88172 62534 88174 62586
rect 88012 62532 88036 62534
rect 88092 62532 88116 62534
rect 88172 62532 88196 62534
rect 87956 62512 88252 62532
rect 89956 62044 90252 62064
rect 90012 62042 90036 62044
rect 90092 62042 90116 62044
rect 90172 62042 90196 62044
rect 90034 61990 90036 62042
rect 90098 61990 90110 62042
rect 90172 61990 90174 62042
rect 90012 61988 90036 61990
rect 90092 61988 90116 61990
rect 90172 61988 90196 61990
rect 89956 61968 90252 61988
rect 87956 61500 88252 61520
rect 88012 61498 88036 61500
rect 88092 61498 88116 61500
rect 88172 61498 88196 61500
rect 88034 61446 88036 61498
rect 88098 61446 88110 61498
rect 88172 61446 88174 61498
rect 88012 61444 88036 61446
rect 88092 61444 88116 61446
rect 88172 61444 88196 61446
rect 87956 61424 88252 61444
rect 89956 60956 90252 60976
rect 90012 60954 90036 60956
rect 90092 60954 90116 60956
rect 90172 60954 90196 60956
rect 90034 60902 90036 60954
rect 90098 60902 90110 60954
rect 90172 60902 90174 60954
rect 90012 60900 90036 60902
rect 90092 60900 90116 60902
rect 90172 60900 90196 60902
rect 89956 60880 90252 60900
rect 87956 60412 88252 60432
rect 88012 60410 88036 60412
rect 88092 60410 88116 60412
rect 88172 60410 88196 60412
rect 88034 60358 88036 60410
rect 88098 60358 88110 60410
rect 88172 60358 88174 60410
rect 88012 60356 88036 60358
rect 88092 60356 88116 60358
rect 88172 60356 88196 60358
rect 87956 60336 88252 60356
rect 89956 59868 90252 59888
rect 90012 59866 90036 59868
rect 90092 59866 90116 59868
rect 90172 59866 90196 59868
rect 90034 59814 90036 59866
rect 90098 59814 90110 59866
rect 90172 59814 90174 59866
rect 90012 59812 90036 59814
rect 90092 59812 90116 59814
rect 90172 59812 90196 59814
rect 89956 59792 90252 59812
rect 87956 59324 88252 59344
rect 88012 59322 88036 59324
rect 88092 59322 88116 59324
rect 88172 59322 88196 59324
rect 88034 59270 88036 59322
rect 88098 59270 88110 59322
rect 88172 59270 88174 59322
rect 88012 59268 88036 59270
rect 88092 59268 88116 59270
rect 88172 59268 88196 59270
rect 87956 59248 88252 59268
rect 89956 58780 90252 58800
rect 90012 58778 90036 58780
rect 90092 58778 90116 58780
rect 90172 58778 90196 58780
rect 90034 58726 90036 58778
rect 90098 58726 90110 58778
rect 90172 58726 90174 58778
rect 90012 58724 90036 58726
rect 90092 58724 90116 58726
rect 90172 58724 90196 58726
rect 89956 58704 90252 58724
rect 87956 58236 88252 58256
rect 88012 58234 88036 58236
rect 88092 58234 88116 58236
rect 88172 58234 88196 58236
rect 88034 58182 88036 58234
rect 88098 58182 88110 58234
rect 88172 58182 88174 58234
rect 88012 58180 88036 58182
rect 88092 58180 88116 58182
rect 88172 58180 88196 58182
rect 87956 58160 88252 58180
rect 89956 57692 90252 57712
rect 90012 57690 90036 57692
rect 90092 57690 90116 57692
rect 90172 57690 90196 57692
rect 90034 57638 90036 57690
rect 90098 57638 90110 57690
rect 90172 57638 90174 57690
rect 90012 57636 90036 57638
rect 90092 57636 90116 57638
rect 90172 57636 90196 57638
rect 89956 57616 90252 57636
rect 87956 57148 88252 57168
rect 88012 57146 88036 57148
rect 88092 57146 88116 57148
rect 88172 57146 88196 57148
rect 88034 57094 88036 57146
rect 88098 57094 88110 57146
rect 88172 57094 88174 57146
rect 88012 57092 88036 57094
rect 88092 57092 88116 57094
rect 88172 57092 88196 57094
rect 87956 57072 88252 57092
rect 89956 56604 90252 56624
rect 90012 56602 90036 56604
rect 90092 56602 90116 56604
rect 90172 56602 90196 56604
rect 90034 56550 90036 56602
rect 90098 56550 90110 56602
rect 90172 56550 90174 56602
rect 90012 56548 90036 56550
rect 90092 56548 90116 56550
rect 90172 56548 90196 56550
rect 89956 56528 90252 56548
rect 87956 56060 88252 56080
rect 88012 56058 88036 56060
rect 88092 56058 88116 56060
rect 88172 56058 88196 56060
rect 88034 56006 88036 56058
rect 88098 56006 88110 56058
rect 88172 56006 88174 56058
rect 88012 56004 88036 56006
rect 88092 56004 88116 56006
rect 88172 56004 88196 56006
rect 87956 55984 88252 56004
rect 89956 55516 90252 55536
rect 90012 55514 90036 55516
rect 90092 55514 90116 55516
rect 90172 55514 90196 55516
rect 90034 55462 90036 55514
rect 90098 55462 90110 55514
rect 90172 55462 90174 55514
rect 90012 55460 90036 55462
rect 90092 55460 90116 55462
rect 90172 55460 90196 55462
rect 89956 55440 90252 55460
rect 87956 54972 88252 54992
rect 88012 54970 88036 54972
rect 88092 54970 88116 54972
rect 88172 54970 88196 54972
rect 88034 54918 88036 54970
rect 88098 54918 88110 54970
rect 88172 54918 88174 54970
rect 88012 54916 88036 54918
rect 88092 54916 88116 54918
rect 88172 54916 88196 54918
rect 87956 54896 88252 54916
rect 89956 54428 90252 54448
rect 90012 54426 90036 54428
rect 90092 54426 90116 54428
rect 90172 54426 90196 54428
rect 90034 54374 90036 54426
rect 90098 54374 90110 54426
rect 90172 54374 90174 54426
rect 90012 54372 90036 54374
rect 90092 54372 90116 54374
rect 90172 54372 90196 54374
rect 89956 54352 90252 54372
rect 87956 53884 88252 53904
rect 88012 53882 88036 53884
rect 88092 53882 88116 53884
rect 88172 53882 88196 53884
rect 88034 53830 88036 53882
rect 88098 53830 88110 53882
rect 88172 53830 88174 53882
rect 88012 53828 88036 53830
rect 88092 53828 88116 53830
rect 88172 53828 88196 53830
rect 87956 53808 88252 53828
rect 89956 53340 90252 53360
rect 90012 53338 90036 53340
rect 90092 53338 90116 53340
rect 90172 53338 90196 53340
rect 90034 53286 90036 53338
rect 90098 53286 90110 53338
rect 90172 53286 90174 53338
rect 90012 53284 90036 53286
rect 90092 53284 90116 53286
rect 90172 53284 90196 53286
rect 89956 53264 90252 53284
rect 87956 52796 88252 52816
rect 88012 52794 88036 52796
rect 88092 52794 88116 52796
rect 88172 52794 88196 52796
rect 88034 52742 88036 52794
rect 88098 52742 88110 52794
rect 88172 52742 88174 52794
rect 88012 52740 88036 52742
rect 88092 52740 88116 52742
rect 88172 52740 88196 52742
rect 87956 52720 88252 52740
rect 89956 52252 90252 52272
rect 90012 52250 90036 52252
rect 90092 52250 90116 52252
rect 90172 52250 90196 52252
rect 90034 52198 90036 52250
rect 90098 52198 90110 52250
rect 90172 52198 90174 52250
rect 90012 52196 90036 52198
rect 90092 52196 90116 52198
rect 90172 52196 90196 52198
rect 89956 52176 90252 52196
rect 87956 51708 88252 51728
rect 88012 51706 88036 51708
rect 88092 51706 88116 51708
rect 88172 51706 88196 51708
rect 88034 51654 88036 51706
rect 88098 51654 88110 51706
rect 88172 51654 88174 51706
rect 88012 51652 88036 51654
rect 88092 51652 88116 51654
rect 88172 51652 88196 51654
rect 87956 51632 88252 51652
rect 89956 51164 90252 51184
rect 90012 51162 90036 51164
rect 90092 51162 90116 51164
rect 90172 51162 90196 51164
rect 90034 51110 90036 51162
rect 90098 51110 90110 51162
rect 90172 51110 90174 51162
rect 90012 51108 90036 51110
rect 90092 51108 90116 51110
rect 90172 51108 90196 51110
rect 89956 51088 90252 51108
rect 87956 50620 88252 50640
rect 88012 50618 88036 50620
rect 88092 50618 88116 50620
rect 88172 50618 88196 50620
rect 88034 50566 88036 50618
rect 88098 50566 88110 50618
rect 88172 50566 88174 50618
rect 88012 50564 88036 50566
rect 88092 50564 88116 50566
rect 88172 50564 88196 50566
rect 87956 50544 88252 50564
rect 89956 50076 90252 50096
rect 90012 50074 90036 50076
rect 90092 50074 90116 50076
rect 90172 50074 90196 50076
rect 90034 50022 90036 50074
rect 90098 50022 90110 50074
rect 90172 50022 90174 50074
rect 90012 50020 90036 50022
rect 90092 50020 90116 50022
rect 90172 50020 90196 50022
rect 89956 50000 90252 50020
rect 87956 49532 88252 49552
rect 88012 49530 88036 49532
rect 88092 49530 88116 49532
rect 88172 49530 88196 49532
rect 88034 49478 88036 49530
rect 88098 49478 88110 49530
rect 88172 49478 88174 49530
rect 88012 49476 88036 49478
rect 88092 49476 88116 49478
rect 88172 49476 88196 49478
rect 87956 49456 88252 49476
rect 89956 48988 90252 49008
rect 90012 48986 90036 48988
rect 90092 48986 90116 48988
rect 90172 48986 90196 48988
rect 90034 48934 90036 48986
rect 90098 48934 90110 48986
rect 90172 48934 90174 48986
rect 90012 48932 90036 48934
rect 90092 48932 90116 48934
rect 90172 48932 90196 48934
rect 89956 48912 90252 48932
rect 87956 48444 88252 48464
rect 88012 48442 88036 48444
rect 88092 48442 88116 48444
rect 88172 48442 88196 48444
rect 88034 48390 88036 48442
rect 88098 48390 88110 48442
rect 88172 48390 88174 48442
rect 88012 48388 88036 48390
rect 88092 48388 88116 48390
rect 88172 48388 88196 48390
rect 87956 48368 88252 48388
rect 89956 47900 90252 47920
rect 90012 47898 90036 47900
rect 90092 47898 90116 47900
rect 90172 47898 90196 47900
rect 90034 47846 90036 47898
rect 90098 47846 90110 47898
rect 90172 47846 90174 47898
rect 90012 47844 90036 47846
rect 90092 47844 90116 47846
rect 90172 47844 90196 47846
rect 89956 47824 90252 47844
rect 87956 47356 88252 47376
rect 88012 47354 88036 47356
rect 88092 47354 88116 47356
rect 88172 47354 88196 47356
rect 88034 47302 88036 47354
rect 88098 47302 88110 47354
rect 88172 47302 88174 47354
rect 88012 47300 88036 47302
rect 88092 47300 88116 47302
rect 88172 47300 88196 47302
rect 87956 47280 88252 47300
rect 89956 46812 90252 46832
rect 90012 46810 90036 46812
rect 90092 46810 90116 46812
rect 90172 46810 90196 46812
rect 90034 46758 90036 46810
rect 90098 46758 90110 46810
rect 90172 46758 90174 46810
rect 90012 46756 90036 46758
rect 90092 46756 90116 46758
rect 90172 46756 90196 46758
rect 89956 46736 90252 46756
rect 87956 46268 88252 46288
rect 88012 46266 88036 46268
rect 88092 46266 88116 46268
rect 88172 46266 88196 46268
rect 88034 46214 88036 46266
rect 88098 46214 88110 46266
rect 88172 46214 88174 46266
rect 88012 46212 88036 46214
rect 88092 46212 88116 46214
rect 88172 46212 88196 46214
rect 87956 46192 88252 46212
rect 89956 45724 90252 45744
rect 90012 45722 90036 45724
rect 90092 45722 90116 45724
rect 90172 45722 90196 45724
rect 90034 45670 90036 45722
rect 90098 45670 90110 45722
rect 90172 45670 90174 45722
rect 90012 45668 90036 45670
rect 90092 45668 90116 45670
rect 90172 45668 90196 45670
rect 89956 45648 90252 45668
rect 87956 45180 88252 45200
rect 88012 45178 88036 45180
rect 88092 45178 88116 45180
rect 88172 45178 88196 45180
rect 88034 45126 88036 45178
rect 88098 45126 88110 45178
rect 88172 45126 88174 45178
rect 88012 45124 88036 45126
rect 88092 45124 88116 45126
rect 88172 45124 88196 45126
rect 87956 45104 88252 45124
rect 89956 44636 90252 44656
rect 90012 44634 90036 44636
rect 90092 44634 90116 44636
rect 90172 44634 90196 44636
rect 90034 44582 90036 44634
rect 90098 44582 90110 44634
rect 90172 44582 90174 44634
rect 90012 44580 90036 44582
rect 90092 44580 90116 44582
rect 90172 44580 90196 44582
rect 89956 44560 90252 44580
rect 87956 44092 88252 44112
rect 88012 44090 88036 44092
rect 88092 44090 88116 44092
rect 88172 44090 88196 44092
rect 88034 44038 88036 44090
rect 88098 44038 88110 44090
rect 88172 44038 88174 44090
rect 88012 44036 88036 44038
rect 88092 44036 88116 44038
rect 88172 44036 88196 44038
rect 87956 44016 88252 44036
rect 89956 43548 90252 43568
rect 90012 43546 90036 43548
rect 90092 43546 90116 43548
rect 90172 43546 90196 43548
rect 90034 43494 90036 43546
rect 90098 43494 90110 43546
rect 90172 43494 90174 43546
rect 90012 43492 90036 43494
rect 90092 43492 90116 43494
rect 90172 43492 90196 43494
rect 89956 43472 90252 43492
rect 87956 43004 88252 43024
rect 88012 43002 88036 43004
rect 88092 43002 88116 43004
rect 88172 43002 88196 43004
rect 88034 42950 88036 43002
rect 88098 42950 88110 43002
rect 88172 42950 88174 43002
rect 88012 42948 88036 42950
rect 88092 42948 88116 42950
rect 88172 42948 88196 42950
rect 87956 42928 88252 42948
rect 89956 42460 90252 42480
rect 90012 42458 90036 42460
rect 90092 42458 90116 42460
rect 90172 42458 90196 42460
rect 90034 42406 90036 42458
rect 90098 42406 90110 42458
rect 90172 42406 90174 42458
rect 90012 42404 90036 42406
rect 90092 42404 90116 42406
rect 90172 42404 90196 42406
rect 89956 42384 90252 42404
rect 87956 41916 88252 41936
rect 88012 41914 88036 41916
rect 88092 41914 88116 41916
rect 88172 41914 88196 41916
rect 88034 41862 88036 41914
rect 88098 41862 88110 41914
rect 88172 41862 88174 41914
rect 88012 41860 88036 41862
rect 88092 41860 88116 41862
rect 88172 41860 88196 41862
rect 87956 41840 88252 41860
rect 89956 41372 90252 41392
rect 90012 41370 90036 41372
rect 90092 41370 90116 41372
rect 90172 41370 90196 41372
rect 90034 41318 90036 41370
rect 90098 41318 90110 41370
rect 90172 41318 90174 41370
rect 90012 41316 90036 41318
rect 90092 41316 90116 41318
rect 90172 41316 90196 41318
rect 89956 41296 90252 41316
rect 87956 40828 88252 40848
rect 88012 40826 88036 40828
rect 88092 40826 88116 40828
rect 88172 40826 88196 40828
rect 88034 40774 88036 40826
rect 88098 40774 88110 40826
rect 88172 40774 88174 40826
rect 88012 40772 88036 40774
rect 88092 40772 88116 40774
rect 88172 40772 88196 40774
rect 87956 40752 88252 40772
rect 87880 40724 87932 40730
rect 87880 40666 87932 40672
rect 87878 40624 87934 40633
rect 87878 40559 87934 40568
rect 87892 40118 87920 40559
rect 89956 40284 90252 40304
rect 90012 40282 90036 40284
rect 90092 40282 90116 40284
rect 90172 40282 90196 40284
rect 90034 40230 90036 40282
rect 90098 40230 90110 40282
rect 90172 40230 90174 40282
rect 90012 40228 90036 40230
rect 90092 40228 90116 40230
rect 90172 40228 90196 40230
rect 89956 40208 90252 40228
rect 87880 40112 87932 40118
rect 87880 40054 87932 40060
rect 87956 39740 88252 39760
rect 88012 39738 88036 39740
rect 88092 39738 88116 39740
rect 88172 39738 88196 39740
rect 88034 39686 88036 39738
rect 88098 39686 88110 39738
rect 88172 39686 88174 39738
rect 88012 39684 88036 39686
rect 88092 39684 88116 39686
rect 88172 39684 88196 39686
rect 87956 39664 88252 39684
rect 89956 39196 90252 39216
rect 90012 39194 90036 39196
rect 90092 39194 90116 39196
rect 90172 39194 90196 39196
rect 90034 39142 90036 39194
rect 90098 39142 90110 39194
rect 90172 39142 90174 39194
rect 90012 39140 90036 39142
rect 90092 39140 90116 39142
rect 90172 39140 90196 39142
rect 89956 39120 90252 39140
rect 87956 38652 88252 38672
rect 88012 38650 88036 38652
rect 88092 38650 88116 38652
rect 88172 38650 88196 38652
rect 88034 38598 88036 38650
rect 88098 38598 88110 38650
rect 88172 38598 88174 38650
rect 88012 38596 88036 38598
rect 88092 38596 88116 38598
rect 88172 38596 88196 38598
rect 87956 38576 88252 38596
rect 89956 38108 90252 38128
rect 90012 38106 90036 38108
rect 90092 38106 90116 38108
rect 90172 38106 90196 38108
rect 90034 38054 90036 38106
rect 90098 38054 90110 38106
rect 90172 38054 90174 38106
rect 90012 38052 90036 38054
rect 90092 38052 90116 38054
rect 90172 38052 90196 38054
rect 89956 38032 90252 38052
rect 87956 37564 88252 37584
rect 88012 37562 88036 37564
rect 88092 37562 88116 37564
rect 88172 37562 88196 37564
rect 88034 37510 88036 37562
rect 88098 37510 88110 37562
rect 88172 37510 88174 37562
rect 88012 37508 88036 37510
rect 88092 37508 88116 37510
rect 88172 37508 88196 37510
rect 87956 37488 88252 37508
rect 89956 37020 90252 37040
rect 90012 37018 90036 37020
rect 90092 37018 90116 37020
rect 90172 37018 90196 37020
rect 90034 36966 90036 37018
rect 90098 36966 90110 37018
rect 90172 36966 90174 37018
rect 90012 36964 90036 36966
rect 90092 36964 90116 36966
rect 90172 36964 90196 36966
rect 89956 36944 90252 36964
rect 87956 36476 88252 36496
rect 88012 36474 88036 36476
rect 88092 36474 88116 36476
rect 88172 36474 88196 36476
rect 88034 36422 88036 36474
rect 88098 36422 88110 36474
rect 88172 36422 88174 36474
rect 88012 36420 88036 36422
rect 88092 36420 88116 36422
rect 88172 36420 88196 36422
rect 87956 36400 88252 36420
rect 89956 35932 90252 35952
rect 90012 35930 90036 35932
rect 90092 35930 90116 35932
rect 90172 35930 90196 35932
rect 90034 35878 90036 35930
rect 90098 35878 90110 35930
rect 90172 35878 90174 35930
rect 90012 35876 90036 35878
rect 90092 35876 90116 35878
rect 90172 35876 90196 35878
rect 89956 35856 90252 35876
rect 87956 35388 88252 35408
rect 88012 35386 88036 35388
rect 88092 35386 88116 35388
rect 88172 35386 88196 35388
rect 88034 35334 88036 35386
rect 88098 35334 88110 35386
rect 88172 35334 88174 35386
rect 88012 35332 88036 35334
rect 88092 35332 88116 35334
rect 88172 35332 88196 35334
rect 87956 35312 88252 35332
rect 89956 34844 90252 34864
rect 90012 34842 90036 34844
rect 90092 34842 90116 34844
rect 90172 34842 90196 34844
rect 90034 34790 90036 34842
rect 90098 34790 90110 34842
rect 90172 34790 90174 34842
rect 90012 34788 90036 34790
rect 90092 34788 90116 34790
rect 90172 34788 90196 34790
rect 89956 34768 90252 34788
rect 87956 34300 88252 34320
rect 88012 34298 88036 34300
rect 88092 34298 88116 34300
rect 88172 34298 88196 34300
rect 88034 34246 88036 34298
rect 88098 34246 88110 34298
rect 88172 34246 88174 34298
rect 88012 34244 88036 34246
rect 88092 34244 88116 34246
rect 88172 34244 88196 34246
rect 87956 34224 88252 34244
rect 89956 33756 90252 33776
rect 90012 33754 90036 33756
rect 90092 33754 90116 33756
rect 90172 33754 90196 33756
rect 90034 33702 90036 33754
rect 90098 33702 90110 33754
rect 90172 33702 90174 33754
rect 90012 33700 90036 33702
rect 90092 33700 90116 33702
rect 90172 33700 90196 33702
rect 89956 33680 90252 33700
rect 87956 33212 88252 33232
rect 88012 33210 88036 33212
rect 88092 33210 88116 33212
rect 88172 33210 88196 33212
rect 88034 33158 88036 33210
rect 88098 33158 88110 33210
rect 88172 33158 88174 33210
rect 88012 33156 88036 33158
rect 88092 33156 88116 33158
rect 88172 33156 88196 33158
rect 87956 33136 88252 33156
rect 89956 32668 90252 32688
rect 90012 32666 90036 32668
rect 90092 32666 90116 32668
rect 90172 32666 90196 32668
rect 90034 32614 90036 32666
rect 90098 32614 90110 32666
rect 90172 32614 90174 32666
rect 90012 32612 90036 32614
rect 90092 32612 90116 32614
rect 90172 32612 90196 32614
rect 89956 32592 90252 32612
rect 87956 32124 88252 32144
rect 88012 32122 88036 32124
rect 88092 32122 88116 32124
rect 88172 32122 88196 32124
rect 88034 32070 88036 32122
rect 88098 32070 88110 32122
rect 88172 32070 88174 32122
rect 88012 32068 88036 32070
rect 88092 32068 88116 32070
rect 88172 32068 88196 32070
rect 87956 32048 88252 32068
rect 89956 31580 90252 31600
rect 90012 31578 90036 31580
rect 90092 31578 90116 31580
rect 90172 31578 90196 31580
rect 90034 31526 90036 31578
rect 90098 31526 90110 31578
rect 90172 31526 90174 31578
rect 90012 31524 90036 31526
rect 90092 31524 90116 31526
rect 90172 31524 90196 31526
rect 89956 31504 90252 31524
rect 87956 31036 88252 31056
rect 88012 31034 88036 31036
rect 88092 31034 88116 31036
rect 88172 31034 88196 31036
rect 88034 30982 88036 31034
rect 88098 30982 88110 31034
rect 88172 30982 88174 31034
rect 88012 30980 88036 30982
rect 88092 30980 88116 30982
rect 88172 30980 88196 30982
rect 87956 30960 88252 30980
rect 89956 30492 90252 30512
rect 90012 30490 90036 30492
rect 90092 30490 90116 30492
rect 90172 30490 90196 30492
rect 90034 30438 90036 30490
rect 90098 30438 90110 30490
rect 90172 30438 90174 30490
rect 90012 30436 90036 30438
rect 90092 30436 90116 30438
rect 90172 30436 90196 30438
rect 89956 30416 90252 30436
rect 87956 29948 88252 29968
rect 88012 29946 88036 29948
rect 88092 29946 88116 29948
rect 88172 29946 88196 29948
rect 88034 29894 88036 29946
rect 88098 29894 88110 29946
rect 88172 29894 88174 29946
rect 88012 29892 88036 29894
rect 88092 29892 88116 29894
rect 88172 29892 88196 29894
rect 87956 29872 88252 29892
rect 89956 29404 90252 29424
rect 90012 29402 90036 29404
rect 90092 29402 90116 29404
rect 90172 29402 90196 29404
rect 90034 29350 90036 29402
rect 90098 29350 90110 29402
rect 90172 29350 90174 29402
rect 90012 29348 90036 29350
rect 90092 29348 90116 29350
rect 90172 29348 90196 29350
rect 89956 29328 90252 29348
rect 87956 28860 88252 28880
rect 88012 28858 88036 28860
rect 88092 28858 88116 28860
rect 88172 28858 88196 28860
rect 88034 28806 88036 28858
rect 88098 28806 88110 28858
rect 88172 28806 88174 28858
rect 88012 28804 88036 28806
rect 88092 28804 88116 28806
rect 88172 28804 88196 28806
rect 87956 28784 88252 28804
rect 89956 28316 90252 28336
rect 90012 28314 90036 28316
rect 90092 28314 90116 28316
rect 90172 28314 90196 28316
rect 90034 28262 90036 28314
rect 90098 28262 90110 28314
rect 90172 28262 90174 28314
rect 90012 28260 90036 28262
rect 90092 28260 90116 28262
rect 90172 28260 90196 28262
rect 89956 28240 90252 28260
rect 87956 27772 88252 27792
rect 88012 27770 88036 27772
rect 88092 27770 88116 27772
rect 88172 27770 88196 27772
rect 88034 27718 88036 27770
rect 88098 27718 88110 27770
rect 88172 27718 88174 27770
rect 88012 27716 88036 27718
rect 88092 27716 88116 27718
rect 88172 27716 88196 27718
rect 87956 27696 88252 27716
rect 89956 27228 90252 27248
rect 90012 27226 90036 27228
rect 90092 27226 90116 27228
rect 90172 27226 90196 27228
rect 90034 27174 90036 27226
rect 90098 27174 90110 27226
rect 90172 27174 90174 27226
rect 90012 27172 90036 27174
rect 90092 27172 90116 27174
rect 90172 27172 90196 27174
rect 89956 27152 90252 27172
rect 87956 26684 88252 26704
rect 88012 26682 88036 26684
rect 88092 26682 88116 26684
rect 88172 26682 88196 26684
rect 88034 26630 88036 26682
rect 88098 26630 88110 26682
rect 88172 26630 88174 26682
rect 88012 26628 88036 26630
rect 88092 26628 88116 26630
rect 88172 26628 88196 26630
rect 87956 26608 88252 26628
rect 89956 26140 90252 26160
rect 90012 26138 90036 26140
rect 90092 26138 90116 26140
rect 90172 26138 90196 26140
rect 90034 26086 90036 26138
rect 90098 26086 90110 26138
rect 90172 26086 90174 26138
rect 90012 26084 90036 26086
rect 90092 26084 90116 26086
rect 90172 26084 90196 26086
rect 89956 26064 90252 26084
rect 87956 25596 88252 25616
rect 88012 25594 88036 25596
rect 88092 25594 88116 25596
rect 88172 25594 88196 25596
rect 88034 25542 88036 25594
rect 88098 25542 88110 25594
rect 88172 25542 88174 25594
rect 88012 25540 88036 25542
rect 88092 25540 88116 25542
rect 88172 25540 88196 25542
rect 87956 25520 88252 25540
rect 89956 25052 90252 25072
rect 90012 25050 90036 25052
rect 90092 25050 90116 25052
rect 90172 25050 90196 25052
rect 90034 24998 90036 25050
rect 90098 24998 90110 25050
rect 90172 24998 90174 25050
rect 90012 24996 90036 24998
rect 90092 24996 90116 24998
rect 90172 24996 90196 24998
rect 89956 24976 90252 24996
rect 87956 24508 88252 24528
rect 88012 24506 88036 24508
rect 88092 24506 88116 24508
rect 88172 24506 88196 24508
rect 88034 24454 88036 24506
rect 88098 24454 88110 24506
rect 88172 24454 88174 24506
rect 88012 24452 88036 24454
rect 88092 24452 88116 24454
rect 88172 24452 88196 24454
rect 87956 24432 88252 24452
rect 89956 23964 90252 23984
rect 90012 23962 90036 23964
rect 90092 23962 90116 23964
rect 90172 23962 90196 23964
rect 90034 23910 90036 23962
rect 90098 23910 90110 23962
rect 90172 23910 90174 23962
rect 90012 23908 90036 23910
rect 90092 23908 90116 23910
rect 90172 23908 90196 23910
rect 89956 23888 90252 23908
rect 87956 23420 88252 23440
rect 88012 23418 88036 23420
rect 88092 23418 88116 23420
rect 88172 23418 88196 23420
rect 88034 23366 88036 23418
rect 88098 23366 88110 23418
rect 88172 23366 88174 23418
rect 88012 23364 88036 23366
rect 88092 23364 88116 23366
rect 88172 23364 88196 23366
rect 87956 23344 88252 23364
rect 89956 22876 90252 22896
rect 90012 22874 90036 22876
rect 90092 22874 90116 22876
rect 90172 22874 90196 22876
rect 90034 22822 90036 22874
rect 90098 22822 90110 22874
rect 90172 22822 90174 22874
rect 90012 22820 90036 22822
rect 90092 22820 90116 22822
rect 90172 22820 90196 22822
rect 89956 22800 90252 22820
rect 87956 22332 88252 22352
rect 88012 22330 88036 22332
rect 88092 22330 88116 22332
rect 88172 22330 88196 22332
rect 88034 22278 88036 22330
rect 88098 22278 88110 22330
rect 88172 22278 88174 22330
rect 88012 22276 88036 22278
rect 88092 22276 88116 22278
rect 88172 22276 88196 22278
rect 87956 22256 88252 22276
rect 89956 21788 90252 21808
rect 90012 21786 90036 21788
rect 90092 21786 90116 21788
rect 90172 21786 90196 21788
rect 90034 21734 90036 21786
rect 90098 21734 90110 21786
rect 90172 21734 90174 21786
rect 90012 21732 90036 21734
rect 90092 21732 90116 21734
rect 90172 21732 90196 21734
rect 89956 21712 90252 21732
rect 87956 21244 88252 21264
rect 88012 21242 88036 21244
rect 88092 21242 88116 21244
rect 88172 21242 88196 21244
rect 88034 21190 88036 21242
rect 88098 21190 88110 21242
rect 88172 21190 88174 21242
rect 88012 21188 88036 21190
rect 88092 21188 88116 21190
rect 88172 21188 88196 21190
rect 87956 21168 88252 21188
rect 87878 21040 87934 21049
rect 87878 20975 87934 20984
rect 87892 20806 87920 20975
rect 87880 20800 87932 20806
rect 87880 20742 87932 20748
rect 89956 20700 90252 20720
rect 90012 20698 90036 20700
rect 90092 20698 90116 20700
rect 90172 20698 90196 20700
rect 90034 20646 90036 20698
rect 90098 20646 90110 20698
rect 90172 20646 90174 20698
rect 90012 20644 90036 20646
rect 90092 20644 90116 20646
rect 90172 20644 90196 20646
rect 89956 20624 90252 20644
rect 87880 20596 87932 20602
rect 87880 20538 87932 20544
rect 87788 8084 87840 8090
rect 87616 4298 87644 8078
rect 87788 8026 87840 8032
rect 87892 7970 87920 20538
rect 87956 20156 88252 20176
rect 88012 20154 88036 20156
rect 88092 20154 88116 20156
rect 88172 20154 88196 20156
rect 88034 20102 88036 20154
rect 88098 20102 88110 20154
rect 88172 20102 88174 20154
rect 88012 20100 88036 20102
rect 88092 20100 88116 20102
rect 88172 20100 88196 20102
rect 87956 20080 88252 20100
rect 89956 19612 90252 19632
rect 90012 19610 90036 19612
rect 90092 19610 90116 19612
rect 90172 19610 90196 19612
rect 90034 19558 90036 19610
rect 90098 19558 90110 19610
rect 90172 19558 90174 19610
rect 90012 19556 90036 19558
rect 90092 19556 90116 19558
rect 90172 19556 90196 19558
rect 89956 19536 90252 19556
rect 87956 19068 88252 19088
rect 88012 19066 88036 19068
rect 88092 19066 88116 19068
rect 88172 19066 88196 19068
rect 88034 19014 88036 19066
rect 88098 19014 88110 19066
rect 88172 19014 88174 19066
rect 88012 19012 88036 19014
rect 88092 19012 88116 19014
rect 88172 19012 88196 19014
rect 87956 18992 88252 19012
rect 89956 18524 90252 18544
rect 90012 18522 90036 18524
rect 90092 18522 90116 18524
rect 90172 18522 90196 18524
rect 90034 18470 90036 18522
rect 90098 18470 90110 18522
rect 90172 18470 90174 18522
rect 90012 18468 90036 18470
rect 90092 18468 90116 18470
rect 90172 18468 90196 18470
rect 89956 18448 90252 18468
rect 87956 17980 88252 18000
rect 88012 17978 88036 17980
rect 88092 17978 88116 17980
rect 88172 17978 88196 17980
rect 88034 17926 88036 17978
rect 88098 17926 88110 17978
rect 88172 17926 88174 17978
rect 88012 17924 88036 17926
rect 88092 17924 88116 17926
rect 88172 17924 88196 17926
rect 87956 17904 88252 17924
rect 89956 17436 90252 17456
rect 90012 17434 90036 17436
rect 90092 17434 90116 17436
rect 90172 17434 90196 17436
rect 90034 17382 90036 17434
rect 90098 17382 90110 17434
rect 90172 17382 90174 17434
rect 90012 17380 90036 17382
rect 90092 17380 90116 17382
rect 90172 17380 90196 17382
rect 89956 17360 90252 17380
rect 87956 16892 88252 16912
rect 88012 16890 88036 16892
rect 88092 16890 88116 16892
rect 88172 16890 88196 16892
rect 88034 16838 88036 16890
rect 88098 16838 88110 16890
rect 88172 16838 88174 16890
rect 88012 16836 88036 16838
rect 88092 16836 88116 16838
rect 88172 16836 88196 16838
rect 87956 16816 88252 16836
rect 89956 16348 90252 16368
rect 90012 16346 90036 16348
rect 90092 16346 90116 16348
rect 90172 16346 90196 16348
rect 90034 16294 90036 16346
rect 90098 16294 90110 16346
rect 90172 16294 90174 16346
rect 90012 16292 90036 16294
rect 90092 16292 90116 16294
rect 90172 16292 90196 16294
rect 89956 16272 90252 16292
rect 87956 15804 88252 15824
rect 88012 15802 88036 15804
rect 88092 15802 88116 15804
rect 88172 15802 88196 15804
rect 88034 15750 88036 15802
rect 88098 15750 88110 15802
rect 88172 15750 88174 15802
rect 88012 15748 88036 15750
rect 88092 15748 88116 15750
rect 88172 15748 88196 15750
rect 87956 15728 88252 15748
rect 89956 15260 90252 15280
rect 90012 15258 90036 15260
rect 90092 15258 90116 15260
rect 90172 15258 90196 15260
rect 90034 15206 90036 15258
rect 90098 15206 90110 15258
rect 90172 15206 90174 15258
rect 90012 15204 90036 15206
rect 90092 15204 90116 15206
rect 90172 15204 90196 15206
rect 89956 15184 90252 15204
rect 87956 14716 88252 14736
rect 88012 14714 88036 14716
rect 88092 14714 88116 14716
rect 88172 14714 88196 14716
rect 88034 14662 88036 14714
rect 88098 14662 88110 14714
rect 88172 14662 88174 14714
rect 88012 14660 88036 14662
rect 88092 14660 88116 14662
rect 88172 14660 88196 14662
rect 87956 14640 88252 14660
rect 89956 14172 90252 14192
rect 90012 14170 90036 14172
rect 90092 14170 90116 14172
rect 90172 14170 90196 14172
rect 90034 14118 90036 14170
rect 90098 14118 90110 14170
rect 90172 14118 90174 14170
rect 90012 14116 90036 14118
rect 90092 14116 90116 14118
rect 90172 14116 90196 14118
rect 89956 14096 90252 14116
rect 87956 13628 88252 13648
rect 88012 13626 88036 13628
rect 88092 13626 88116 13628
rect 88172 13626 88196 13628
rect 88034 13574 88036 13626
rect 88098 13574 88110 13626
rect 88172 13574 88174 13626
rect 88012 13572 88036 13574
rect 88092 13572 88116 13574
rect 88172 13572 88196 13574
rect 87956 13552 88252 13572
rect 89956 13084 90252 13104
rect 90012 13082 90036 13084
rect 90092 13082 90116 13084
rect 90172 13082 90196 13084
rect 90034 13030 90036 13082
rect 90098 13030 90110 13082
rect 90172 13030 90174 13082
rect 90012 13028 90036 13030
rect 90092 13028 90116 13030
rect 90172 13028 90196 13030
rect 89956 13008 90252 13028
rect 87956 12540 88252 12560
rect 88012 12538 88036 12540
rect 88092 12538 88116 12540
rect 88172 12538 88196 12540
rect 88034 12486 88036 12538
rect 88098 12486 88110 12538
rect 88172 12486 88174 12538
rect 88012 12484 88036 12486
rect 88092 12484 88116 12486
rect 88172 12484 88196 12486
rect 87956 12464 88252 12484
rect 89956 11996 90252 12016
rect 90012 11994 90036 11996
rect 90092 11994 90116 11996
rect 90172 11994 90196 11996
rect 90034 11942 90036 11994
rect 90098 11942 90110 11994
rect 90172 11942 90174 11994
rect 90012 11940 90036 11942
rect 90092 11940 90116 11942
rect 90172 11940 90196 11942
rect 89956 11920 90252 11940
rect 87956 11452 88252 11472
rect 88012 11450 88036 11452
rect 88092 11450 88116 11452
rect 88172 11450 88196 11452
rect 88034 11398 88036 11450
rect 88098 11398 88110 11450
rect 88172 11398 88174 11450
rect 88012 11396 88036 11398
rect 88092 11396 88116 11398
rect 88172 11396 88196 11398
rect 87956 11376 88252 11396
rect 89956 10908 90252 10928
rect 90012 10906 90036 10908
rect 90092 10906 90116 10908
rect 90172 10906 90196 10908
rect 90034 10854 90036 10906
rect 90098 10854 90110 10906
rect 90172 10854 90174 10906
rect 90012 10852 90036 10854
rect 90092 10852 90116 10854
rect 90172 10852 90196 10854
rect 89956 10832 90252 10852
rect 87956 10364 88252 10384
rect 88012 10362 88036 10364
rect 88092 10362 88116 10364
rect 88172 10362 88196 10364
rect 88034 10310 88036 10362
rect 88098 10310 88110 10362
rect 88172 10310 88174 10362
rect 88012 10308 88036 10310
rect 88092 10308 88116 10310
rect 88172 10308 88196 10310
rect 87956 10288 88252 10308
rect 89956 9820 90252 9840
rect 90012 9818 90036 9820
rect 90092 9818 90116 9820
rect 90172 9818 90196 9820
rect 90034 9766 90036 9818
rect 90098 9766 90110 9818
rect 90172 9766 90174 9818
rect 90012 9764 90036 9766
rect 90092 9764 90116 9766
rect 90172 9764 90196 9766
rect 89956 9744 90252 9764
rect 87956 9276 88252 9296
rect 88012 9274 88036 9276
rect 88092 9274 88116 9276
rect 88172 9274 88196 9276
rect 88034 9222 88036 9274
rect 88098 9222 88110 9274
rect 88172 9222 88174 9274
rect 88012 9220 88036 9222
rect 88092 9220 88116 9222
rect 88172 9220 88196 9222
rect 87956 9200 88252 9220
rect 89956 8732 90252 8752
rect 90012 8730 90036 8732
rect 90092 8730 90116 8732
rect 90172 8730 90196 8732
rect 90034 8678 90036 8730
rect 90098 8678 90110 8730
rect 90172 8678 90174 8730
rect 90012 8676 90036 8678
rect 90092 8676 90116 8678
rect 90172 8676 90196 8678
rect 89956 8656 90252 8676
rect 87956 8188 88252 8208
rect 88012 8186 88036 8188
rect 88092 8186 88116 8188
rect 88172 8186 88196 8188
rect 88034 8134 88036 8186
rect 88098 8134 88110 8186
rect 88172 8134 88174 8186
rect 88012 8132 88036 8134
rect 88092 8132 88116 8134
rect 88172 8132 88196 8134
rect 87956 8112 88252 8132
rect 87708 7942 87920 7970
rect 87972 8016 88024 8022
rect 87972 7958 88024 7964
rect 87708 7410 87736 7942
rect 87878 7848 87934 7857
rect 87878 7783 87934 7792
rect 87788 7540 87840 7546
rect 87788 7482 87840 7488
rect 87696 7404 87748 7410
rect 87696 7346 87748 7352
rect 87696 7268 87748 7274
rect 87696 7210 87748 7216
rect 87708 4758 87736 7210
rect 87696 4752 87748 4758
rect 87696 4694 87748 4700
rect 87616 4270 87736 4298
rect 87602 4176 87658 4185
rect 87602 4111 87658 4120
rect 87616 2990 87644 4111
rect 87708 4078 87736 4270
rect 87696 4072 87748 4078
rect 87696 4014 87748 4020
rect 87604 2984 87656 2990
rect 87604 2926 87656 2932
rect 87512 2916 87564 2922
rect 87512 2858 87564 2864
rect 87800 2774 87828 7482
rect 87892 2938 87920 7783
rect 87984 7274 88012 7958
rect 89956 7644 90252 7664
rect 90012 7642 90036 7644
rect 90092 7642 90116 7644
rect 90172 7642 90196 7644
rect 90034 7590 90036 7642
rect 90098 7590 90110 7642
rect 90172 7590 90174 7642
rect 90012 7588 90036 7590
rect 90092 7588 90116 7590
rect 90172 7588 90196 7590
rect 89956 7568 90252 7588
rect 87972 7268 88024 7274
rect 87972 7210 88024 7216
rect 87956 7100 88252 7120
rect 88012 7098 88036 7100
rect 88092 7098 88116 7100
rect 88172 7098 88196 7100
rect 88034 7046 88036 7098
rect 88098 7046 88110 7098
rect 88172 7046 88174 7098
rect 88012 7044 88036 7046
rect 88092 7044 88116 7046
rect 88172 7044 88196 7046
rect 87956 7024 88252 7044
rect 89956 6556 90252 6576
rect 90012 6554 90036 6556
rect 90092 6554 90116 6556
rect 90172 6554 90196 6556
rect 90034 6502 90036 6554
rect 90098 6502 90110 6554
rect 90172 6502 90174 6554
rect 90012 6500 90036 6502
rect 90092 6500 90116 6502
rect 90172 6500 90196 6502
rect 89956 6480 90252 6500
rect 87956 6012 88252 6032
rect 88012 6010 88036 6012
rect 88092 6010 88116 6012
rect 88172 6010 88196 6012
rect 88034 5958 88036 6010
rect 88098 5958 88110 6010
rect 88172 5958 88174 6010
rect 88012 5956 88036 5958
rect 88092 5956 88116 5958
rect 88172 5956 88196 5958
rect 87956 5936 88252 5956
rect 89956 5468 90252 5488
rect 90012 5466 90036 5468
rect 90092 5466 90116 5468
rect 90172 5466 90196 5468
rect 90034 5414 90036 5466
rect 90098 5414 90110 5466
rect 90172 5414 90174 5466
rect 90012 5412 90036 5414
rect 90092 5412 90116 5414
rect 90172 5412 90196 5414
rect 89956 5392 90252 5412
rect 87956 4924 88252 4944
rect 88012 4922 88036 4924
rect 88092 4922 88116 4924
rect 88172 4922 88196 4924
rect 88034 4870 88036 4922
rect 88098 4870 88110 4922
rect 88172 4870 88174 4922
rect 88012 4868 88036 4870
rect 88092 4868 88116 4870
rect 88172 4868 88196 4870
rect 87956 4848 88252 4868
rect 87972 4752 88024 4758
rect 87972 4694 88024 4700
rect 87984 4010 88012 4694
rect 89956 4380 90252 4400
rect 90012 4378 90036 4380
rect 90092 4378 90116 4380
rect 90172 4378 90196 4380
rect 90034 4326 90036 4378
rect 90098 4326 90110 4378
rect 90172 4326 90174 4378
rect 90012 4324 90036 4326
rect 90092 4324 90116 4326
rect 90172 4324 90196 4326
rect 89956 4304 90252 4324
rect 87972 4004 88024 4010
rect 87972 3946 88024 3952
rect 87956 3836 88252 3856
rect 88012 3834 88036 3836
rect 88092 3834 88116 3836
rect 88172 3834 88196 3836
rect 88034 3782 88036 3834
rect 88098 3782 88110 3834
rect 88172 3782 88174 3834
rect 88012 3780 88036 3782
rect 88092 3780 88116 3782
rect 88172 3780 88196 3782
rect 87956 3760 88252 3780
rect 89956 3292 90252 3312
rect 90012 3290 90036 3292
rect 90092 3290 90116 3292
rect 90172 3290 90196 3292
rect 90034 3238 90036 3290
rect 90098 3238 90110 3290
rect 90172 3238 90174 3290
rect 90012 3236 90036 3238
rect 90092 3236 90116 3238
rect 90172 3236 90196 3238
rect 89956 3216 90252 3236
rect 87892 2910 88380 2938
rect 87800 2746 87920 2774
rect 87420 1760 87472 1766
rect 87420 1702 87472 1708
rect 87052 1692 87104 1698
rect 87052 1634 87104 1640
rect 87892 1630 87920 2746
rect 87956 2748 88252 2768
rect 88012 2746 88036 2748
rect 88092 2746 88116 2748
rect 88172 2746 88196 2748
rect 88034 2694 88036 2746
rect 88098 2694 88110 2746
rect 88172 2694 88174 2746
rect 88012 2692 88036 2694
rect 88092 2692 88116 2694
rect 88172 2692 88196 2694
rect 87956 2672 88252 2692
rect 88352 2530 88380 2910
rect 88260 2502 88380 2530
rect 87880 1624 87932 1630
rect 87880 1566 87932 1572
rect 88260 1494 88288 2502
rect 89956 2204 90252 2224
rect 90012 2202 90036 2204
rect 90092 2202 90116 2204
rect 90172 2202 90196 2204
rect 90034 2150 90036 2202
rect 90098 2150 90110 2202
rect 90172 2150 90174 2202
rect 90012 2148 90036 2150
rect 90092 2148 90116 2150
rect 90172 2148 90196 2150
rect 89956 2128 90252 2148
rect 88248 1488 88300 1494
rect 88248 1430 88300 1436
rect 86958 640 87014 649
rect 86958 575 87014 584
rect 86500 196 86552 202
rect 86500 138 86552 144
rect 24768 128 24820 134
rect 24768 70 24820 76
rect 86408 128 86460 134
rect 86408 70 86460 76
<< via2 >>
rect 1956 189338 2012 189340
rect 2036 189338 2092 189340
rect 2116 189338 2172 189340
rect 2196 189338 2252 189340
rect 1956 189286 1982 189338
rect 1982 189286 2012 189338
rect 2036 189286 2046 189338
rect 2046 189286 2092 189338
rect 2116 189286 2162 189338
rect 2162 189286 2172 189338
rect 2196 189286 2226 189338
rect 2226 189286 2252 189338
rect 1956 189284 2012 189286
rect 2036 189284 2092 189286
rect 2116 189284 2172 189286
rect 2196 189284 2252 189286
rect 85956 189338 86012 189340
rect 86036 189338 86092 189340
rect 86116 189338 86172 189340
rect 86196 189338 86252 189340
rect 85956 189286 85982 189338
rect 85982 189286 86012 189338
rect 86036 189286 86046 189338
rect 86046 189286 86092 189338
rect 86116 189286 86162 189338
rect 86162 189286 86172 189338
rect 86196 189286 86226 189338
rect 86226 189286 86252 189338
rect 85956 189284 86012 189286
rect 86036 189284 86092 189286
rect 86116 189284 86172 189286
rect 86196 189284 86252 189286
rect 89956 189338 90012 189340
rect 90036 189338 90092 189340
rect 90116 189338 90172 189340
rect 90196 189338 90252 189340
rect 89956 189286 89982 189338
rect 89982 189286 90012 189338
rect 90036 189286 90046 189338
rect 90046 189286 90092 189338
rect 90116 189286 90162 189338
rect 90162 189286 90172 189338
rect 90196 189286 90226 189338
rect 90226 189286 90252 189338
rect 89956 189284 90012 189286
rect 90036 189284 90092 189286
rect 90116 189284 90172 189286
rect 90196 189284 90252 189286
rect 75826 189100 75882 189136
rect 75826 189080 75828 189100
rect 75828 189080 75880 189100
rect 75880 189080 75882 189100
rect 3956 188794 4012 188796
rect 4036 188794 4092 188796
rect 4116 188794 4172 188796
rect 4196 188794 4252 188796
rect 3956 188742 3982 188794
rect 3982 188742 4012 188794
rect 4036 188742 4046 188794
rect 4046 188742 4092 188794
rect 4116 188742 4162 188794
rect 4162 188742 4172 188794
rect 4196 188742 4226 188794
rect 4226 188742 4252 188794
rect 3956 188740 4012 188742
rect 4036 188740 4092 188742
rect 4116 188740 4172 188742
rect 4196 188740 4252 188742
rect 1956 188250 2012 188252
rect 2036 188250 2092 188252
rect 2116 188250 2172 188252
rect 2196 188250 2252 188252
rect 1956 188198 1982 188250
rect 1982 188198 2012 188250
rect 2036 188198 2046 188250
rect 2046 188198 2092 188250
rect 2116 188198 2162 188250
rect 2162 188198 2172 188250
rect 2196 188198 2226 188250
rect 2226 188198 2252 188250
rect 1956 188196 2012 188198
rect 2036 188196 2092 188198
rect 2116 188196 2172 188198
rect 2196 188196 2252 188198
rect 3956 187706 4012 187708
rect 4036 187706 4092 187708
rect 4116 187706 4172 187708
rect 4196 187706 4252 187708
rect 3956 187654 3982 187706
rect 3982 187654 4012 187706
rect 4036 187654 4046 187706
rect 4046 187654 4092 187706
rect 4116 187654 4162 187706
rect 4162 187654 4172 187706
rect 4196 187654 4226 187706
rect 4226 187654 4252 187706
rect 3956 187652 4012 187654
rect 4036 187652 4092 187654
rect 4116 187652 4172 187654
rect 4196 187652 4252 187654
rect 1956 187162 2012 187164
rect 2036 187162 2092 187164
rect 2116 187162 2172 187164
rect 2196 187162 2252 187164
rect 1956 187110 1982 187162
rect 1982 187110 2012 187162
rect 2036 187110 2046 187162
rect 2046 187110 2092 187162
rect 2116 187110 2162 187162
rect 2162 187110 2172 187162
rect 2196 187110 2226 187162
rect 2226 187110 2252 187162
rect 1956 187108 2012 187110
rect 2036 187108 2092 187110
rect 2116 187108 2172 187110
rect 2196 187108 2252 187110
rect 87956 188794 88012 188796
rect 88036 188794 88092 188796
rect 88116 188794 88172 188796
rect 88196 188794 88252 188796
rect 87956 188742 87982 188794
rect 87982 188742 88012 188794
rect 88036 188742 88046 188794
rect 88046 188742 88092 188794
rect 88116 188742 88162 188794
rect 88162 188742 88172 188794
rect 88196 188742 88226 188794
rect 88226 188742 88252 188794
rect 87956 188740 88012 188742
rect 88036 188740 88092 188742
rect 88116 188740 88172 188742
rect 88196 188740 88252 188742
rect 85956 188250 86012 188252
rect 86036 188250 86092 188252
rect 86116 188250 86172 188252
rect 86196 188250 86252 188252
rect 85956 188198 85982 188250
rect 85982 188198 86012 188250
rect 86036 188198 86046 188250
rect 86046 188198 86092 188250
rect 86116 188198 86162 188250
rect 86162 188198 86172 188250
rect 86196 188198 86226 188250
rect 86226 188198 86252 188250
rect 85956 188196 86012 188198
rect 86036 188196 86092 188198
rect 86116 188196 86172 188198
rect 86196 188196 86252 188198
rect 89956 188250 90012 188252
rect 90036 188250 90092 188252
rect 90116 188250 90172 188252
rect 90196 188250 90252 188252
rect 89956 188198 89982 188250
rect 89982 188198 90012 188250
rect 90036 188198 90046 188250
rect 90046 188198 90092 188250
rect 90116 188198 90162 188250
rect 90162 188198 90172 188250
rect 90196 188198 90226 188250
rect 90226 188198 90252 188250
rect 89956 188196 90012 188198
rect 90036 188196 90092 188198
rect 90116 188196 90172 188198
rect 90196 188196 90252 188198
rect 87956 187706 88012 187708
rect 88036 187706 88092 187708
rect 88116 187706 88172 187708
rect 88196 187706 88252 187708
rect 87956 187654 87982 187706
rect 87982 187654 88012 187706
rect 88036 187654 88046 187706
rect 88046 187654 88092 187706
rect 88116 187654 88162 187706
rect 88162 187654 88172 187706
rect 88196 187654 88226 187706
rect 88226 187654 88252 187706
rect 87956 187652 88012 187654
rect 88036 187652 88092 187654
rect 88116 187652 88172 187654
rect 88196 187652 88252 187654
rect 79322 187040 79378 187096
rect 3956 186618 4012 186620
rect 4036 186618 4092 186620
rect 4116 186618 4172 186620
rect 4196 186618 4252 186620
rect 3956 186566 3982 186618
rect 3982 186566 4012 186618
rect 4036 186566 4046 186618
rect 4046 186566 4092 186618
rect 4116 186566 4162 186618
rect 4162 186566 4172 186618
rect 4196 186566 4226 186618
rect 4226 186566 4252 186618
rect 3956 186564 4012 186566
rect 4036 186564 4092 186566
rect 4116 186564 4172 186566
rect 4196 186564 4252 186566
rect 1956 186074 2012 186076
rect 2036 186074 2092 186076
rect 2116 186074 2172 186076
rect 2196 186074 2252 186076
rect 1956 186022 1982 186074
rect 1982 186022 2012 186074
rect 2036 186022 2046 186074
rect 2046 186022 2092 186074
rect 2116 186022 2162 186074
rect 2162 186022 2172 186074
rect 2196 186022 2226 186074
rect 2226 186022 2252 186074
rect 1956 186020 2012 186022
rect 2036 186020 2092 186022
rect 2116 186020 2172 186022
rect 2196 186020 2252 186022
rect 3956 185530 4012 185532
rect 4036 185530 4092 185532
rect 4116 185530 4172 185532
rect 4196 185530 4252 185532
rect 3956 185478 3982 185530
rect 3982 185478 4012 185530
rect 4036 185478 4046 185530
rect 4046 185478 4092 185530
rect 4116 185478 4162 185530
rect 4162 185478 4172 185530
rect 4196 185478 4226 185530
rect 4226 185478 4252 185530
rect 3956 185476 4012 185478
rect 4036 185476 4092 185478
rect 4116 185476 4172 185478
rect 4196 185476 4252 185478
rect 1956 184986 2012 184988
rect 2036 184986 2092 184988
rect 2116 184986 2172 184988
rect 2196 184986 2252 184988
rect 1956 184934 1982 184986
rect 1982 184934 2012 184986
rect 2036 184934 2046 184986
rect 2046 184934 2092 184986
rect 2116 184934 2162 184986
rect 2162 184934 2172 184986
rect 2196 184934 2226 184986
rect 2226 184934 2252 184986
rect 1956 184932 2012 184934
rect 2036 184932 2092 184934
rect 2116 184932 2172 184934
rect 2196 184932 2252 184934
rect 3956 184442 4012 184444
rect 4036 184442 4092 184444
rect 4116 184442 4172 184444
rect 4196 184442 4252 184444
rect 3956 184390 3982 184442
rect 3982 184390 4012 184442
rect 4036 184390 4046 184442
rect 4046 184390 4092 184442
rect 4116 184390 4162 184442
rect 4162 184390 4172 184442
rect 4196 184390 4226 184442
rect 4226 184390 4252 184442
rect 3956 184388 4012 184390
rect 4036 184388 4092 184390
rect 4116 184388 4172 184390
rect 4196 184388 4252 184390
rect 1956 183898 2012 183900
rect 2036 183898 2092 183900
rect 2116 183898 2172 183900
rect 2196 183898 2252 183900
rect 1956 183846 1982 183898
rect 1982 183846 2012 183898
rect 2036 183846 2046 183898
rect 2046 183846 2092 183898
rect 2116 183846 2162 183898
rect 2162 183846 2172 183898
rect 2196 183846 2226 183898
rect 2226 183846 2252 183898
rect 1956 183844 2012 183846
rect 2036 183844 2092 183846
rect 2116 183844 2172 183846
rect 2196 183844 2252 183846
rect 3956 183354 4012 183356
rect 4036 183354 4092 183356
rect 4116 183354 4172 183356
rect 4196 183354 4252 183356
rect 3956 183302 3982 183354
rect 3982 183302 4012 183354
rect 4036 183302 4046 183354
rect 4046 183302 4092 183354
rect 4116 183302 4162 183354
rect 4162 183302 4172 183354
rect 4196 183302 4226 183354
rect 4226 183302 4252 183354
rect 3956 183300 4012 183302
rect 4036 183300 4092 183302
rect 4116 183300 4172 183302
rect 4196 183300 4252 183302
rect 1956 182810 2012 182812
rect 2036 182810 2092 182812
rect 2116 182810 2172 182812
rect 2196 182810 2252 182812
rect 1956 182758 1982 182810
rect 1982 182758 2012 182810
rect 2036 182758 2046 182810
rect 2046 182758 2092 182810
rect 2116 182758 2162 182810
rect 2162 182758 2172 182810
rect 2196 182758 2226 182810
rect 2226 182758 2252 182810
rect 1956 182756 2012 182758
rect 2036 182756 2092 182758
rect 2116 182756 2172 182758
rect 2196 182756 2252 182758
rect 3956 182266 4012 182268
rect 4036 182266 4092 182268
rect 4116 182266 4172 182268
rect 4196 182266 4252 182268
rect 3956 182214 3982 182266
rect 3982 182214 4012 182266
rect 4036 182214 4046 182266
rect 4046 182214 4092 182266
rect 4116 182214 4162 182266
rect 4162 182214 4172 182266
rect 4196 182214 4226 182266
rect 4226 182214 4252 182266
rect 3956 182212 4012 182214
rect 4036 182212 4092 182214
rect 4116 182212 4172 182214
rect 4196 182212 4252 182214
rect 1956 181722 2012 181724
rect 2036 181722 2092 181724
rect 2116 181722 2172 181724
rect 2196 181722 2252 181724
rect 1956 181670 1982 181722
rect 1982 181670 2012 181722
rect 2036 181670 2046 181722
rect 2046 181670 2092 181722
rect 2116 181670 2162 181722
rect 2162 181670 2172 181722
rect 2196 181670 2226 181722
rect 2226 181670 2252 181722
rect 1956 181668 2012 181670
rect 2036 181668 2092 181670
rect 2116 181668 2172 181670
rect 2196 181668 2252 181670
rect 3956 181178 4012 181180
rect 4036 181178 4092 181180
rect 4116 181178 4172 181180
rect 4196 181178 4252 181180
rect 3956 181126 3982 181178
rect 3982 181126 4012 181178
rect 4036 181126 4046 181178
rect 4046 181126 4092 181178
rect 4116 181126 4162 181178
rect 4162 181126 4172 181178
rect 4196 181126 4226 181178
rect 4226 181126 4252 181178
rect 3956 181124 4012 181126
rect 4036 181124 4092 181126
rect 4116 181124 4172 181126
rect 4196 181124 4252 181126
rect 1956 180634 2012 180636
rect 2036 180634 2092 180636
rect 2116 180634 2172 180636
rect 2196 180634 2252 180636
rect 1956 180582 1982 180634
rect 1982 180582 2012 180634
rect 2036 180582 2046 180634
rect 2046 180582 2092 180634
rect 2116 180582 2162 180634
rect 2162 180582 2172 180634
rect 2196 180582 2226 180634
rect 2226 180582 2252 180634
rect 1956 180580 2012 180582
rect 2036 180580 2092 180582
rect 2116 180580 2172 180582
rect 2196 180580 2252 180582
rect 3956 180090 4012 180092
rect 4036 180090 4092 180092
rect 4116 180090 4172 180092
rect 4196 180090 4252 180092
rect 3956 180038 3982 180090
rect 3982 180038 4012 180090
rect 4036 180038 4046 180090
rect 4046 180038 4092 180090
rect 4116 180038 4162 180090
rect 4162 180038 4172 180090
rect 4196 180038 4226 180090
rect 4226 180038 4252 180090
rect 3956 180036 4012 180038
rect 4036 180036 4092 180038
rect 4116 180036 4172 180038
rect 4196 180036 4252 180038
rect 1956 179546 2012 179548
rect 2036 179546 2092 179548
rect 2116 179546 2172 179548
rect 2196 179546 2252 179548
rect 1956 179494 1982 179546
rect 1982 179494 2012 179546
rect 2036 179494 2046 179546
rect 2046 179494 2092 179546
rect 2116 179494 2162 179546
rect 2162 179494 2172 179546
rect 2196 179494 2226 179546
rect 2226 179494 2252 179546
rect 1956 179492 2012 179494
rect 2036 179492 2092 179494
rect 2116 179492 2172 179494
rect 2196 179492 2252 179494
rect 3956 179002 4012 179004
rect 4036 179002 4092 179004
rect 4116 179002 4172 179004
rect 4196 179002 4252 179004
rect 3956 178950 3982 179002
rect 3982 178950 4012 179002
rect 4036 178950 4046 179002
rect 4046 178950 4092 179002
rect 4116 178950 4162 179002
rect 4162 178950 4172 179002
rect 4196 178950 4226 179002
rect 4226 178950 4252 179002
rect 3956 178948 4012 178950
rect 4036 178948 4092 178950
rect 4116 178948 4172 178950
rect 4196 178948 4252 178950
rect 1956 178458 2012 178460
rect 2036 178458 2092 178460
rect 2116 178458 2172 178460
rect 2196 178458 2252 178460
rect 1956 178406 1982 178458
rect 1982 178406 2012 178458
rect 2036 178406 2046 178458
rect 2046 178406 2092 178458
rect 2116 178406 2162 178458
rect 2162 178406 2172 178458
rect 2196 178406 2226 178458
rect 2226 178406 2252 178458
rect 1956 178404 2012 178406
rect 2036 178404 2092 178406
rect 2116 178404 2172 178406
rect 2196 178404 2252 178406
rect 3956 177914 4012 177916
rect 4036 177914 4092 177916
rect 4116 177914 4172 177916
rect 4196 177914 4252 177916
rect 3956 177862 3982 177914
rect 3982 177862 4012 177914
rect 4036 177862 4046 177914
rect 4046 177862 4092 177914
rect 4116 177862 4162 177914
rect 4162 177862 4172 177914
rect 4196 177862 4226 177914
rect 4226 177862 4252 177914
rect 3956 177860 4012 177862
rect 4036 177860 4092 177862
rect 4116 177860 4172 177862
rect 4196 177860 4252 177862
rect 1956 177370 2012 177372
rect 2036 177370 2092 177372
rect 2116 177370 2172 177372
rect 2196 177370 2252 177372
rect 1956 177318 1982 177370
rect 1982 177318 2012 177370
rect 2036 177318 2046 177370
rect 2046 177318 2092 177370
rect 2116 177318 2162 177370
rect 2162 177318 2172 177370
rect 2196 177318 2226 177370
rect 2226 177318 2252 177370
rect 1956 177316 2012 177318
rect 2036 177316 2092 177318
rect 2116 177316 2172 177318
rect 2196 177316 2252 177318
rect 3956 176826 4012 176828
rect 4036 176826 4092 176828
rect 4116 176826 4172 176828
rect 4196 176826 4252 176828
rect 3956 176774 3982 176826
rect 3982 176774 4012 176826
rect 4036 176774 4046 176826
rect 4046 176774 4092 176826
rect 4116 176774 4162 176826
rect 4162 176774 4172 176826
rect 4196 176774 4226 176826
rect 4226 176774 4252 176826
rect 3956 176772 4012 176774
rect 4036 176772 4092 176774
rect 4116 176772 4172 176774
rect 4196 176772 4252 176774
rect 1956 176282 2012 176284
rect 2036 176282 2092 176284
rect 2116 176282 2172 176284
rect 2196 176282 2252 176284
rect 1956 176230 1982 176282
rect 1982 176230 2012 176282
rect 2036 176230 2046 176282
rect 2046 176230 2092 176282
rect 2116 176230 2162 176282
rect 2162 176230 2172 176282
rect 2196 176230 2226 176282
rect 2226 176230 2252 176282
rect 1956 176228 2012 176230
rect 2036 176228 2092 176230
rect 2116 176228 2172 176230
rect 2196 176228 2252 176230
rect 3956 175738 4012 175740
rect 4036 175738 4092 175740
rect 4116 175738 4172 175740
rect 4196 175738 4252 175740
rect 3956 175686 3982 175738
rect 3982 175686 4012 175738
rect 4036 175686 4046 175738
rect 4046 175686 4092 175738
rect 4116 175686 4162 175738
rect 4162 175686 4172 175738
rect 4196 175686 4226 175738
rect 4226 175686 4252 175738
rect 3956 175684 4012 175686
rect 4036 175684 4092 175686
rect 4116 175684 4172 175686
rect 4196 175684 4252 175686
rect 1956 175194 2012 175196
rect 2036 175194 2092 175196
rect 2116 175194 2172 175196
rect 2196 175194 2252 175196
rect 1956 175142 1982 175194
rect 1982 175142 2012 175194
rect 2036 175142 2046 175194
rect 2046 175142 2092 175194
rect 2116 175142 2162 175194
rect 2162 175142 2172 175194
rect 2196 175142 2226 175194
rect 2226 175142 2252 175194
rect 1956 175140 2012 175142
rect 2036 175140 2092 175142
rect 2116 175140 2172 175142
rect 2196 175140 2252 175142
rect 3956 174650 4012 174652
rect 4036 174650 4092 174652
rect 4116 174650 4172 174652
rect 4196 174650 4252 174652
rect 3956 174598 3982 174650
rect 3982 174598 4012 174650
rect 4036 174598 4046 174650
rect 4046 174598 4092 174650
rect 4116 174598 4162 174650
rect 4162 174598 4172 174650
rect 4196 174598 4226 174650
rect 4226 174598 4252 174650
rect 3956 174596 4012 174598
rect 4036 174596 4092 174598
rect 4116 174596 4172 174598
rect 4196 174596 4252 174598
rect 1956 174106 2012 174108
rect 2036 174106 2092 174108
rect 2116 174106 2172 174108
rect 2196 174106 2252 174108
rect 1956 174054 1982 174106
rect 1982 174054 2012 174106
rect 2036 174054 2046 174106
rect 2046 174054 2092 174106
rect 2116 174054 2162 174106
rect 2162 174054 2172 174106
rect 2196 174054 2226 174106
rect 2226 174054 2252 174106
rect 1956 174052 2012 174054
rect 2036 174052 2092 174054
rect 2116 174052 2172 174054
rect 2196 174052 2252 174054
rect 3956 173562 4012 173564
rect 4036 173562 4092 173564
rect 4116 173562 4172 173564
rect 4196 173562 4252 173564
rect 3956 173510 3982 173562
rect 3982 173510 4012 173562
rect 4036 173510 4046 173562
rect 4046 173510 4092 173562
rect 4116 173510 4162 173562
rect 4162 173510 4172 173562
rect 4196 173510 4226 173562
rect 4226 173510 4252 173562
rect 3956 173508 4012 173510
rect 4036 173508 4092 173510
rect 4116 173508 4172 173510
rect 4196 173508 4252 173510
rect 1956 173018 2012 173020
rect 2036 173018 2092 173020
rect 2116 173018 2172 173020
rect 2196 173018 2252 173020
rect 1956 172966 1982 173018
rect 1982 172966 2012 173018
rect 2036 172966 2046 173018
rect 2046 172966 2092 173018
rect 2116 172966 2162 173018
rect 2162 172966 2172 173018
rect 2196 172966 2226 173018
rect 2226 172966 2252 173018
rect 1956 172964 2012 172966
rect 2036 172964 2092 172966
rect 2116 172964 2172 172966
rect 2196 172964 2252 172966
rect 3956 172474 4012 172476
rect 4036 172474 4092 172476
rect 4116 172474 4172 172476
rect 4196 172474 4252 172476
rect 3956 172422 3982 172474
rect 3982 172422 4012 172474
rect 4036 172422 4046 172474
rect 4046 172422 4092 172474
rect 4116 172422 4162 172474
rect 4162 172422 4172 172474
rect 4196 172422 4226 172474
rect 4226 172422 4252 172474
rect 3956 172420 4012 172422
rect 4036 172420 4092 172422
rect 4116 172420 4172 172422
rect 4196 172420 4252 172422
rect 1956 171930 2012 171932
rect 2036 171930 2092 171932
rect 2116 171930 2172 171932
rect 2196 171930 2252 171932
rect 1956 171878 1982 171930
rect 1982 171878 2012 171930
rect 2036 171878 2046 171930
rect 2046 171878 2092 171930
rect 2116 171878 2162 171930
rect 2162 171878 2172 171930
rect 2196 171878 2226 171930
rect 2226 171878 2252 171930
rect 1956 171876 2012 171878
rect 2036 171876 2092 171878
rect 2116 171876 2172 171878
rect 2196 171876 2252 171878
rect 3956 171386 4012 171388
rect 4036 171386 4092 171388
rect 4116 171386 4172 171388
rect 4196 171386 4252 171388
rect 3956 171334 3982 171386
rect 3982 171334 4012 171386
rect 4036 171334 4046 171386
rect 4046 171334 4092 171386
rect 4116 171334 4162 171386
rect 4162 171334 4172 171386
rect 4196 171334 4226 171386
rect 4226 171334 4252 171386
rect 3956 171332 4012 171334
rect 4036 171332 4092 171334
rect 4116 171332 4172 171334
rect 4196 171332 4252 171334
rect 1956 170842 2012 170844
rect 2036 170842 2092 170844
rect 2116 170842 2172 170844
rect 2196 170842 2252 170844
rect 1956 170790 1982 170842
rect 1982 170790 2012 170842
rect 2036 170790 2046 170842
rect 2046 170790 2092 170842
rect 2116 170790 2162 170842
rect 2162 170790 2172 170842
rect 2196 170790 2226 170842
rect 2226 170790 2252 170842
rect 1956 170788 2012 170790
rect 2036 170788 2092 170790
rect 2116 170788 2172 170790
rect 2196 170788 2252 170790
rect 3956 170298 4012 170300
rect 4036 170298 4092 170300
rect 4116 170298 4172 170300
rect 4196 170298 4252 170300
rect 3956 170246 3982 170298
rect 3982 170246 4012 170298
rect 4036 170246 4046 170298
rect 4046 170246 4092 170298
rect 4116 170246 4162 170298
rect 4162 170246 4172 170298
rect 4196 170246 4226 170298
rect 4226 170246 4252 170298
rect 3956 170244 4012 170246
rect 4036 170244 4092 170246
rect 4116 170244 4172 170246
rect 4196 170244 4252 170246
rect 1956 169754 2012 169756
rect 2036 169754 2092 169756
rect 2116 169754 2172 169756
rect 2196 169754 2252 169756
rect 1956 169702 1982 169754
rect 1982 169702 2012 169754
rect 2036 169702 2046 169754
rect 2046 169702 2092 169754
rect 2116 169702 2162 169754
rect 2162 169702 2172 169754
rect 2196 169702 2226 169754
rect 2226 169702 2252 169754
rect 1956 169700 2012 169702
rect 2036 169700 2092 169702
rect 2116 169700 2172 169702
rect 2196 169700 2252 169702
rect 3956 169210 4012 169212
rect 4036 169210 4092 169212
rect 4116 169210 4172 169212
rect 4196 169210 4252 169212
rect 3956 169158 3982 169210
rect 3982 169158 4012 169210
rect 4036 169158 4046 169210
rect 4046 169158 4092 169210
rect 4116 169158 4162 169210
rect 4162 169158 4172 169210
rect 4196 169158 4226 169210
rect 4226 169158 4252 169210
rect 3956 169156 4012 169158
rect 4036 169156 4092 169158
rect 4116 169156 4172 169158
rect 4196 169156 4252 169158
rect 1956 168666 2012 168668
rect 2036 168666 2092 168668
rect 2116 168666 2172 168668
rect 2196 168666 2252 168668
rect 1956 168614 1982 168666
rect 1982 168614 2012 168666
rect 2036 168614 2046 168666
rect 2046 168614 2092 168666
rect 2116 168614 2162 168666
rect 2162 168614 2172 168666
rect 2196 168614 2226 168666
rect 2226 168614 2252 168666
rect 1956 168612 2012 168614
rect 2036 168612 2092 168614
rect 2116 168612 2172 168614
rect 2196 168612 2252 168614
rect 3956 168122 4012 168124
rect 4036 168122 4092 168124
rect 4116 168122 4172 168124
rect 4196 168122 4252 168124
rect 3956 168070 3982 168122
rect 3982 168070 4012 168122
rect 4036 168070 4046 168122
rect 4046 168070 4092 168122
rect 4116 168070 4162 168122
rect 4162 168070 4172 168122
rect 4196 168070 4226 168122
rect 4226 168070 4252 168122
rect 3956 168068 4012 168070
rect 4036 168068 4092 168070
rect 4116 168068 4172 168070
rect 4196 168068 4252 168070
rect 1956 167578 2012 167580
rect 2036 167578 2092 167580
rect 2116 167578 2172 167580
rect 2196 167578 2252 167580
rect 1956 167526 1982 167578
rect 1982 167526 2012 167578
rect 2036 167526 2046 167578
rect 2046 167526 2092 167578
rect 2116 167526 2162 167578
rect 2162 167526 2172 167578
rect 2196 167526 2226 167578
rect 2226 167526 2252 167578
rect 1956 167524 2012 167526
rect 2036 167524 2092 167526
rect 2116 167524 2172 167526
rect 2196 167524 2252 167526
rect 3956 167034 4012 167036
rect 4036 167034 4092 167036
rect 4116 167034 4172 167036
rect 4196 167034 4252 167036
rect 3956 166982 3982 167034
rect 3982 166982 4012 167034
rect 4036 166982 4046 167034
rect 4046 166982 4092 167034
rect 4116 166982 4162 167034
rect 4162 166982 4172 167034
rect 4196 166982 4226 167034
rect 4226 166982 4252 167034
rect 3956 166980 4012 166982
rect 4036 166980 4092 166982
rect 4116 166980 4172 166982
rect 4196 166980 4252 166982
rect 1956 166490 2012 166492
rect 2036 166490 2092 166492
rect 2116 166490 2172 166492
rect 2196 166490 2252 166492
rect 1956 166438 1982 166490
rect 1982 166438 2012 166490
rect 2036 166438 2046 166490
rect 2046 166438 2092 166490
rect 2116 166438 2162 166490
rect 2162 166438 2172 166490
rect 2196 166438 2226 166490
rect 2226 166438 2252 166490
rect 1956 166436 2012 166438
rect 2036 166436 2092 166438
rect 2116 166436 2172 166438
rect 2196 166436 2252 166438
rect 3956 165946 4012 165948
rect 4036 165946 4092 165948
rect 4116 165946 4172 165948
rect 4196 165946 4252 165948
rect 3956 165894 3982 165946
rect 3982 165894 4012 165946
rect 4036 165894 4046 165946
rect 4046 165894 4092 165946
rect 4116 165894 4162 165946
rect 4162 165894 4172 165946
rect 4196 165894 4226 165946
rect 4226 165894 4252 165946
rect 3956 165892 4012 165894
rect 4036 165892 4092 165894
rect 4116 165892 4172 165894
rect 4196 165892 4252 165894
rect 1956 165402 2012 165404
rect 2036 165402 2092 165404
rect 2116 165402 2172 165404
rect 2196 165402 2252 165404
rect 1956 165350 1982 165402
rect 1982 165350 2012 165402
rect 2036 165350 2046 165402
rect 2046 165350 2092 165402
rect 2116 165350 2162 165402
rect 2162 165350 2172 165402
rect 2196 165350 2226 165402
rect 2226 165350 2252 165402
rect 1956 165348 2012 165350
rect 2036 165348 2092 165350
rect 2116 165348 2172 165350
rect 2196 165348 2252 165350
rect 3956 164858 4012 164860
rect 4036 164858 4092 164860
rect 4116 164858 4172 164860
rect 4196 164858 4252 164860
rect 3956 164806 3982 164858
rect 3982 164806 4012 164858
rect 4036 164806 4046 164858
rect 4046 164806 4092 164858
rect 4116 164806 4162 164858
rect 4162 164806 4172 164858
rect 4196 164806 4226 164858
rect 4226 164806 4252 164858
rect 3956 164804 4012 164806
rect 4036 164804 4092 164806
rect 4116 164804 4172 164806
rect 4196 164804 4252 164806
rect 1956 164314 2012 164316
rect 2036 164314 2092 164316
rect 2116 164314 2172 164316
rect 2196 164314 2252 164316
rect 1956 164262 1982 164314
rect 1982 164262 2012 164314
rect 2036 164262 2046 164314
rect 2046 164262 2092 164314
rect 2116 164262 2162 164314
rect 2162 164262 2172 164314
rect 2196 164262 2226 164314
rect 2226 164262 2252 164314
rect 1956 164260 2012 164262
rect 2036 164260 2092 164262
rect 2116 164260 2172 164262
rect 2196 164260 2252 164262
rect 3956 163770 4012 163772
rect 4036 163770 4092 163772
rect 4116 163770 4172 163772
rect 4196 163770 4252 163772
rect 3956 163718 3982 163770
rect 3982 163718 4012 163770
rect 4036 163718 4046 163770
rect 4046 163718 4092 163770
rect 4116 163718 4162 163770
rect 4162 163718 4172 163770
rect 4196 163718 4226 163770
rect 4226 163718 4252 163770
rect 3956 163716 4012 163718
rect 4036 163716 4092 163718
rect 4116 163716 4172 163718
rect 4196 163716 4252 163718
rect 1956 163226 2012 163228
rect 2036 163226 2092 163228
rect 2116 163226 2172 163228
rect 2196 163226 2252 163228
rect 1956 163174 1982 163226
rect 1982 163174 2012 163226
rect 2036 163174 2046 163226
rect 2046 163174 2092 163226
rect 2116 163174 2162 163226
rect 2162 163174 2172 163226
rect 2196 163174 2226 163226
rect 2226 163174 2252 163226
rect 1956 163172 2012 163174
rect 2036 163172 2092 163174
rect 2116 163172 2172 163174
rect 2196 163172 2252 163174
rect 3956 162682 4012 162684
rect 4036 162682 4092 162684
rect 4116 162682 4172 162684
rect 4196 162682 4252 162684
rect 3956 162630 3982 162682
rect 3982 162630 4012 162682
rect 4036 162630 4046 162682
rect 4046 162630 4092 162682
rect 4116 162630 4162 162682
rect 4162 162630 4172 162682
rect 4196 162630 4226 162682
rect 4226 162630 4252 162682
rect 3956 162628 4012 162630
rect 4036 162628 4092 162630
rect 4116 162628 4172 162630
rect 4196 162628 4252 162630
rect 1956 162138 2012 162140
rect 2036 162138 2092 162140
rect 2116 162138 2172 162140
rect 2196 162138 2252 162140
rect 1956 162086 1982 162138
rect 1982 162086 2012 162138
rect 2036 162086 2046 162138
rect 2046 162086 2092 162138
rect 2116 162086 2162 162138
rect 2162 162086 2172 162138
rect 2196 162086 2226 162138
rect 2226 162086 2252 162138
rect 1956 162084 2012 162086
rect 2036 162084 2092 162086
rect 2116 162084 2172 162086
rect 2196 162084 2252 162086
rect 3956 161594 4012 161596
rect 4036 161594 4092 161596
rect 4116 161594 4172 161596
rect 4196 161594 4252 161596
rect 3956 161542 3982 161594
rect 3982 161542 4012 161594
rect 4036 161542 4046 161594
rect 4046 161542 4092 161594
rect 4116 161542 4162 161594
rect 4162 161542 4172 161594
rect 4196 161542 4226 161594
rect 4226 161542 4252 161594
rect 3956 161540 4012 161542
rect 4036 161540 4092 161542
rect 4116 161540 4172 161542
rect 4196 161540 4252 161542
rect 1956 161050 2012 161052
rect 2036 161050 2092 161052
rect 2116 161050 2172 161052
rect 2196 161050 2252 161052
rect 1956 160998 1982 161050
rect 1982 160998 2012 161050
rect 2036 160998 2046 161050
rect 2046 160998 2092 161050
rect 2116 160998 2162 161050
rect 2162 160998 2172 161050
rect 2196 160998 2226 161050
rect 2226 160998 2252 161050
rect 1956 160996 2012 160998
rect 2036 160996 2092 160998
rect 2116 160996 2172 160998
rect 2196 160996 2252 160998
rect 3956 160506 4012 160508
rect 4036 160506 4092 160508
rect 4116 160506 4172 160508
rect 4196 160506 4252 160508
rect 3956 160454 3982 160506
rect 3982 160454 4012 160506
rect 4036 160454 4046 160506
rect 4046 160454 4092 160506
rect 4116 160454 4162 160506
rect 4162 160454 4172 160506
rect 4196 160454 4226 160506
rect 4226 160454 4252 160506
rect 3956 160452 4012 160454
rect 4036 160452 4092 160454
rect 4116 160452 4172 160454
rect 4196 160452 4252 160454
rect 1956 159962 2012 159964
rect 2036 159962 2092 159964
rect 2116 159962 2172 159964
rect 2196 159962 2252 159964
rect 1956 159910 1982 159962
rect 1982 159910 2012 159962
rect 2036 159910 2046 159962
rect 2046 159910 2092 159962
rect 2116 159910 2162 159962
rect 2162 159910 2172 159962
rect 2196 159910 2226 159962
rect 2226 159910 2252 159962
rect 1956 159908 2012 159910
rect 2036 159908 2092 159910
rect 2116 159908 2172 159910
rect 2196 159908 2252 159910
rect 3956 159418 4012 159420
rect 4036 159418 4092 159420
rect 4116 159418 4172 159420
rect 4196 159418 4252 159420
rect 3956 159366 3982 159418
rect 3982 159366 4012 159418
rect 4036 159366 4046 159418
rect 4046 159366 4092 159418
rect 4116 159366 4162 159418
rect 4162 159366 4172 159418
rect 4196 159366 4226 159418
rect 4226 159366 4252 159418
rect 3956 159364 4012 159366
rect 4036 159364 4092 159366
rect 4116 159364 4172 159366
rect 4196 159364 4252 159366
rect 1956 158874 2012 158876
rect 2036 158874 2092 158876
rect 2116 158874 2172 158876
rect 2196 158874 2252 158876
rect 1956 158822 1982 158874
rect 1982 158822 2012 158874
rect 2036 158822 2046 158874
rect 2046 158822 2092 158874
rect 2116 158822 2162 158874
rect 2162 158822 2172 158874
rect 2196 158822 2226 158874
rect 2226 158822 2252 158874
rect 1956 158820 2012 158822
rect 2036 158820 2092 158822
rect 2116 158820 2172 158822
rect 2196 158820 2252 158822
rect 3956 158330 4012 158332
rect 4036 158330 4092 158332
rect 4116 158330 4172 158332
rect 4196 158330 4252 158332
rect 3956 158278 3982 158330
rect 3982 158278 4012 158330
rect 4036 158278 4046 158330
rect 4046 158278 4092 158330
rect 4116 158278 4162 158330
rect 4162 158278 4172 158330
rect 4196 158278 4226 158330
rect 4226 158278 4252 158330
rect 3956 158276 4012 158278
rect 4036 158276 4092 158278
rect 4116 158276 4172 158278
rect 4196 158276 4252 158278
rect 1956 157786 2012 157788
rect 2036 157786 2092 157788
rect 2116 157786 2172 157788
rect 2196 157786 2252 157788
rect 1956 157734 1982 157786
rect 1982 157734 2012 157786
rect 2036 157734 2046 157786
rect 2046 157734 2092 157786
rect 2116 157734 2162 157786
rect 2162 157734 2172 157786
rect 2196 157734 2226 157786
rect 2226 157734 2252 157786
rect 1956 157732 2012 157734
rect 2036 157732 2092 157734
rect 2116 157732 2172 157734
rect 2196 157732 2252 157734
rect 3956 157242 4012 157244
rect 4036 157242 4092 157244
rect 4116 157242 4172 157244
rect 4196 157242 4252 157244
rect 3956 157190 3982 157242
rect 3982 157190 4012 157242
rect 4036 157190 4046 157242
rect 4046 157190 4092 157242
rect 4116 157190 4162 157242
rect 4162 157190 4172 157242
rect 4196 157190 4226 157242
rect 4226 157190 4252 157242
rect 3956 157188 4012 157190
rect 4036 157188 4092 157190
rect 4116 157188 4172 157190
rect 4196 157188 4252 157190
rect 1956 156698 2012 156700
rect 2036 156698 2092 156700
rect 2116 156698 2172 156700
rect 2196 156698 2252 156700
rect 1956 156646 1982 156698
rect 1982 156646 2012 156698
rect 2036 156646 2046 156698
rect 2046 156646 2092 156698
rect 2116 156646 2162 156698
rect 2162 156646 2172 156698
rect 2196 156646 2226 156698
rect 2226 156646 2252 156698
rect 1956 156644 2012 156646
rect 2036 156644 2092 156646
rect 2116 156644 2172 156646
rect 2196 156644 2252 156646
rect 3956 156154 4012 156156
rect 4036 156154 4092 156156
rect 4116 156154 4172 156156
rect 4196 156154 4252 156156
rect 3956 156102 3982 156154
rect 3982 156102 4012 156154
rect 4036 156102 4046 156154
rect 4046 156102 4092 156154
rect 4116 156102 4162 156154
rect 4162 156102 4172 156154
rect 4196 156102 4226 156154
rect 4226 156102 4252 156154
rect 3956 156100 4012 156102
rect 4036 156100 4092 156102
rect 4116 156100 4172 156102
rect 4196 156100 4252 156102
rect 1956 155610 2012 155612
rect 2036 155610 2092 155612
rect 2116 155610 2172 155612
rect 2196 155610 2252 155612
rect 1956 155558 1982 155610
rect 1982 155558 2012 155610
rect 2036 155558 2046 155610
rect 2046 155558 2092 155610
rect 2116 155558 2162 155610
rect 2162 155558 2172 155610
rect 2196 155558 2226 155610
rect 2226 155558 2252 155610
rect 1956 155556 2012 155558
rect 2036 155556 2092 155558
rect 2116 155556 2172 155558
rect 2196 155556 2252 155558
rect 3956 155066 4012 155068
rect 4036 155066 4092 155068
rect 4116 155066 4172 155068
rect 4196 155066 4252 155068
rect 3956 155014 3982 155066
rect 3982 155014 4012 155066
rect 4036 155014 4046 155066
rect 4046 155014 4092 155066
rect 4116 155014 4162 155066
rect 4162 155014 4172 155066
rect 4196 155014 4226 155066
rect 4226 155014 4252 155066
rect 3956 155012 4012 155014
rect 4036 155012 4092 155014
rect 4116 155012 4172 155014
rect 4196 155012 4252 155014
rect 1956 154522 2012 154524
rect 2036 154522 2092 154524
rect 2116 154522 2172 154524
rect 2196 154522 2252 154524
rect 1956 154470 1982 154522
rect 1982 154470 2012 154522
rect 2036 154470 2046 154522
rect 2046 154470 2092 154522
rect 2116 154470 2162 154522
rect 2162 154470 2172 154522
rect 2196 154470 2226 154522
rect 2226 154470 2252 154522
rect 1956 154468 2012 154470
rect 2036 154468 2092 154470
rect 2116 154468 2172 154470
rect 2196 154468 2252 154470
rect 3956 153978 4012 153980
rect 4036 153978 4092 153980
rect 4116 153978 4172 153980
rect 4196 153978 4252 153980
rect 3956 153926 3982 153978
rect 3982 153926 4012 153978
rect 4036 153926 4046 153978
rect 4046 153926 4092 153978
rect 4116 153926 4162 153978
rect 4162 153926 4172 153978
rect 4196 153926 4226 153978
rect 4226 153926 4252 153978
rect 3956 153924 4012 153926
rect 4036 153924 4092 153926
rect 4116 153924 4172 153926
rect 4196 153924 4252 153926
rect 1956 153434 2012 153436
rect 2036 153434 2092 153436
rect 2116 153434 2172 153436
rect 2196 153434 2252 153436
rect 1956 153382 1982 153434
rect 1982 153382 2012 153434
rect 2036 153382 2046 153434
rect 2046 153382 2092 153434
rect 2116 153382 2162 153434
rect 2162 153382 2172 153434
rect 2196 153382 2226 153434
rect 2226 153382 2252 153434
rect 1956 153380 2012 153382
rect 2036 153380 2092 153382
rect 2116 153380 2172 153382
rect 2196 153380 2252 153382
rect 3956 152890 4012 152892
rect 4036 152890 4092 152892
rect 4116 152890 4172 152892
rect 4196 152890 4252 152892
rect 3956 152838 3982 152890
rect 3982 152838 4012 152890
rect 4036 152838 4046 152890
rect 4046 152838 4092 152890
rect 4116 152838 4162 152890
rect 4162 152838 4172 152890
rect 4196 152838 4226 152890
rect 4226 152838 4252 152890
rect 3956 152836 4012 152838
rect 4036 152836 4092 152838
rect 4116 152836 4172 152838
rect 4196 152836 4252 152838
rect 1956 152346 2012 152348
rect 2036 152346 2092 152348
rect 2116 152346 2172 152348
rect 2196 152346 2252 152348
rect 1956 152294 1982 152346
rect 1982 152294 2012 152346
rect 2036 152294 2046 152346
rect 2046 152294 2092 152346
rect 2116 152294 2162 152346
rect 2162 152294 2172 152346
rect 2196 152294 2226 152346
rect 2226 152294 2252 152346
rect 1956 152292 2012 152294
rect 2036 152292 2092 152294
rect 2116 152292 2172 152294
rect 2196 152292 2252 152294
rect 3956 151802 4012 151804
rect 4036 151802 4092 151804
rect 4116 151802 4172 151804
rect 4196 151802 4252 151804
rect 3956 151750 3982 151802
rect 3982 151750 4012 151802
rect 4036 151750 4046 151802
rect 4046 151750 4092 151802
rect 4116 151750 4162 151802
rect 4162 151750 4172 151802
rect 4196 151750 4226 151802
rect 4226 151750 4252 151802
rect 3956 151748 4012 151750
rect 4036 151748 4092 151750
rect 4116 151748 4172 151750
rect 4196 151748 4252 151750
rect 1956 151258 2012 151260
rect 2036 151258 2092 151260
rect 2116 151258 2172 151260
rect 2196 151258 2252 151260
rect 1956 151206 1982 151258
rect 1982 151206 2012 151258
rect 2036 151206 2046 151258
rect 2046 151206 2092 151258
rect 2116 151206 2162 151258
rect 2162 151206 2172 151258
rect 2196 151206 2226 151258
rect 2226 151206 2252 151258
rect 1956 151204 2012 151206
rect 2036 151204 2092 151206
rect 2116 151204 2172 151206
rect 2196 151204 2252 151206
rect 3956 150714 4012 150716
rect 4036 150714 4092 150716
rect 4116 150714 4172 150716
rect 4196 150714 4252 150716
rect 3956 150662 3982 150714
rect 3982 150662 4012 150714
rect 4036 150662 4046 150714
rect 4046 150662 4092 150714
rect 4116 150662 4162 150714
rect 4162 150662 4172 150714
rect 4196 150662 4226 150714
rect 4226 150662 4252 150714
rect 3956 150660 4012 150662
rect 4036 150660 4092 150662
rect 4116 150660 4172 150662
rect 4196 150660 4252 150662
rect 1956 150170 2012 150172
rect 2036 150170 2092 150172
rect 2116 150170 2172 150172
rect 2196 150170 2252 150172
rect 1956 150118 1982 150170
rect 1982 150118 2012 150170
rect 2036 150118 2046 150170
rect 2046 150118 2092 150170
rect 2116 150118 2162 150170
rect 2162 150118 2172 150170
rect 2196 150118 2226 150170
rect 2226 150118 2252 150170
rect 1956 150116 2012 150118
rect 2036 150116 2092 150118
rect 2116 150116 2172 150118
rect 2196 150116 2252 150118
rect 3956 149626 4012 149628
rect 4036 149626 4092 149628
rect 4116 149626 4172 149628
rect 4196 149626 4252 149628
rect 3956 149574 3982 149626
rect 3982 149574 4012 149626
rect 4036 149574 4046 149626
rect 4046 149574 4092 149626
rect 4116 149574 4162 149626
rect 4162 149574 4172 149626
rect 4196 149574 4226 149626
rect 4226 149574 4252 149626
rect 3956 149572 4012 149574
rect 4036 149572 4092 149574
rect 4116 149572 4172 149574
rect 4196 149572 4252 149574
rect 1956 149082 2012 149084
rect 2036 149082 2092 149084
rect 2116 149082 2172 149084
rect 2196 149082 2252 149084
rect 1956 149030 1982 149082
rect 1982 149030 2012 149082
rect 2036 149030 2046 149082
rect 2046 149030 2092 149082
rect 2116 149030 2162 149082
rect 2162 149030 2172 149082
rect 2196 149030 2226 149082
rect 2226 149030 2252 149082
rect 1956 149028 2012 149030
rect 2036 149028 2092 149030
rect 2116 149028 2172 149030
rect 2196 149028 2252 149030
rect 3956 148538 4012 148540
rect 4036 148538 4092 148540
rect 4116 148538 4172 148540
rect 4196 148538 4252 148540
rect 3956 148486 3982 148538
rect 3982 148486 4012 148538
rect 4036 148486 4046 148538
rect 4046 148486 4092 148538
rect 4116 148486 4162 148538
rect 4162 148486 4172 148538
rect 4196 148486 4226 148538
rect 4226 148486 4252 148538
rect 3956 148484 4012 148486
rect 4036 148484 4092 148486
rect 4116 148484 4172 148486
rect 4196 148484 4252 148486
rect 1956 147994 2012 147996
rect 2036 147994 2092 147996
rect 2116 147994 2172 147996
rect 2196 147994 2252 147996
rect 1956 147942 1982 147994
rect 1982 147942 2012 147994
rect 2036 147942 2046 147994
rect 2046 147942 2092 147994
rect 2116 147942 2162 147994
rect 2162 147942 2172 147994
rect 2196 147942 2226 147994
rect 2226 147942 2252 147994
rect 1956 147940 2012 147942
rect 2036 147940 2092 147942
rect 2116 147940 2172 147942
rect 2196 147940 2252 147942
rect 3956 147450 4012 147452
rect 4036 147450 4092 147452
rect 4116 147450 4172 147452
rect 4196 147450 4252 147452
rect 3956 147398 3982 147450
rect 3982 147398 4012 147450
rect 4036 147398 4046 147450
rect 4046 147398 4092 147450
rect 4116 147398 4162 147450
rect 4162 147398 4172 147450
rect 4196 147398 4226 147450
rect 4226 147398 4252 147450
rect 3956 147396 4012 147398
rect 4036 147396 4092 147398
rect 4116 147396 4172 147398
rect 4196 147396 4252 147398
rect 1956 146906 2012 146908
rect 2036 146906 2092 146908
rect 2116 146906 2172 146908
rect 2196 146906 2252 146908
rect 1956 146854 1982 146906
rect 1982 146854 2012 146906
rect 2036 146854 2046 146906
rect 2046 146854 2092 146906
rect 2116 146854 2162 146906
rect 2162 146854 2172 146906
rect 2196 146854 2226 146906
rect 2226 146854 2252 146906
rect 1956 146852 2012 146854
rect 2036 146852 2092 146854
rect 2116 146852 2172 146854
rect 2196 146852 2252 146854
rect 3956 146362 4012 146364
rect 4036 146362 4092 146364
rect 4116 146362 4172 146364
rect 4196 146362 4252 146364
rect 3956 146310 3982 146362
rect 3982 146310 4012 146362
rect 4036 146310 4046 146362
rect 4046 146310 4092 146362
rect 4116 146310 4162 146362
rect 4162 146310 4172 146362
rect 4196 146310 4226 146362
rect 4226 146310 4252 146362
rect 3956 146308 4012 146310
rect 4036 146308 4092 146310
rect 4116 146308 4172 146310
rect 4196 146308 4252 146310
rect 1956 145818 2012 145820
rect 2036 145818 2092 145820
rect 2116 145818 2172 145820
rect 2196 145818 2252 145820
rect 1956 145766 1982 145818
rect 1982 145766 2012 145818
rect 2036 145766 2046 145818
rect 2046 145766 2092 145818
rect 2116 145766 2162 145818
rect 2162 145766 2172 145818
rect 2196 145766 2226 145818
rect 2226 145766 2252 145818
rect 1956 145764 2012 145766
rect 2036 145764 2092 145766
rect 2116 145764 2172 145766
rect 2196 145764 2252 145766
rect 3956 145274 4012 145276
rect 4036 145274 4092 145276
rect 4116 145274 4172 145276
rect 4196 145274 4252 145276
rect 3956 145222 3982 145274
rect 3982 145222 4012 145274
rect 4036 145222 4046 145274
rect 4046 145222 4092 145274
rect 4116 145222 4162 145274
rect 4162 145222 4172 145274
rect 4196 145222 4226 145274
rect 4226 145222 4252 145274
rect 3956 145220 4012 145222
rect 4036 145220 4092 145222
rect 4116 145220 4172 145222
rect 4196 145220 4252 145222
rect 1956 144730 2012 144732
rect 2036 144730 2092 144732
rect 2116 144730 2172 144732
rect 2196 144730 2252 144732
rect 1956 144678 1982 144730
rect 1982 144678 2012 144730
rect 2036 144678 2046 144730
rect 2046 144678 2092 144730
rect 2116 144678 2162 144730
rect 2162 144678 2172 144730
rect 2196 144678 2226 144730
rect 2226 144678 2252 144730
rect 1956 144676 2012 144678
rect 2036 144676 2092 144678
rect 2116 144676 2172 144678
rect 2196 144676 2252 144678
rect 3956 144186 4012 144188
rect 4036 144186 4092 144188
rect 4116 144186 4172 144188
rect 4196 144186 4252 144188
rect 3956 144134 3982 144186
rect 3982 144134 4012 144186
rect 4036 144134 4046 144186
rect 4046 144134 4092 144186
rect 4116 144134 4162 144186
rect 4162 144134 4172 144186
rect 4196 144134 4226 144186
rect 4226 144134 4252 144186
rect 3956 144132 4012 144134
rect 4036 144132 4092 144134
rect 4116 144132 4172 144134
rect 4196 144132 4252 144134
rect 1956 143642 2012 143644
rect 2036 143642 2092 143644
rect 2116 143642 2172 143644
rect 2196 143642 2252 143644
rect 1956 143590 1982 143642
rect 1982 143590 2012 143642
rect 2036 143590 2046 143642
rect 2046 143590 2092 143642
rect 2116 143590 2162 143642
rect 2162 143590 2172 143642
rect 2196 143590 2226 143642
rect 2226 143590 2252 143642
rect 1956 143588 2012 143590
rect 2036 143588 2092 143590
rect 2116 143588 2172 143590
rect 2196 143588 2252 143590
rect 3956 143098 4012 143100
rect 4036 143098 4092 143100
rect 4116 143098 4172 143100
rect 4196 143098 4252 143100
rect 3956 143046 3982 143098
rect 3982 143046 4012 143098
rect 4036 143046 4046 143098
rect 4046 143046 4092 143098
rect 4116 143046 4162 143098
rect 4162 143046 4172 143098
rect 4196 143046 4226 143098
rect 4226 143046 4252 143098
rect 3956 143044 4012 143046
rect 4036 143044 4092 143046
rect 4116 143044 4172 143046
rect 4196 143044 4252 143046
rect 1956 142554 2012 142556
rect 2036 142554 2092 142556
rect 2116 142554 2172 142556
rect 2196 142554 2252 142556
rect 1956 142502 1982 142554
rect 1982 142502 2012 142554
rect 2036 142502 2046 142554
rect 2046 142502 2092 142554
rect 2116 142502 2162 142554
rect 2162 142502 2172 142554
rect 2196 142502 2226 142554
rect 2226 142502 2252 142554
rect 1956 142500 2012 142502
rect 2036 142500 2092 142502
rect 2116 142500 2172 142502
rect 2196 142500 2252 142502
rect 3956 142010 4012 142012
rect 4036 142010 4092 142012
rect 4116 142010 4172 142012
rect 4196 142010 4252 142012
rect 3956 141958 3982 142010
rect 3982 141958 4012 142010
rect 4036 141958 4046 142010
rect 4046 141958 4092 142010
rect 4116 141958 4162 142010
rect 4162 141958 4172 142010
rect 4196 141958 4226 142010
rect 4226 141958 4252 142010
rect 3956 141956 4012 141958
rect 4036 141956 4092 141958
rect 4116 141956 4172 141958
rect 4196 141956 4252 141958
rect 1956 141466 2012 141468
rect 2036 141466 2092 141468
rect 2116 141466 2172 141468
rect 2196 141466 2252 141468
rect 1956 141414 1982 141466
rect 1982 141414 2012 141466
rect 2036 141414 2046 141466
rect 2046 141414 2092 141466
rect 2116 141414 2162 141466
rect 2162 141414 2172 141466
rect 2196 141414 2226 141466
rect 2226 141414 2252 141466
rect 1956 141412 2012 141414
rect 2036 141412 2092 141414
rect 2116 141412 2172 141414
rect 2196 141412 2252 141414
rect 3956 140922 4012 140924
rect 4036 140922 4092 140924
rect 4116 140922 4172 140924
rect 4196 140922 4252 140924
rect 3956 140870 3982 140922
rect 3982 140870 4012 140922
rect 4036 140870 4046 140922
rect 4046 140870 4092 140922
rect 4116 140870 4162 140922
rect 4162 140870 4172 140922
rect 4196 140870 4226 140922
rect 4226 140870 4252 140922
rect 3956 140868 4012 140870
rect 4036 140868 4092 140870
rect 4116 140868 4172 140870
rect 4196 140868 4252 140870
rect 1956 140378 2012 140380
rect 2036 140378 2092 140380
rect 2116 140378 2172 140380
rect 2196 140378 2252 140380
rect 1956 140326 1982 140378
rect 1982 140326 2012 140378
rect 2036 140326 2046 140378
rect 2046 140326 2092 140378
rect 2116 140326 2162 140378
rect 2162 140326 2172 140378
rect 2196 140326 2226 140378
rect 2226 140326 2252 140378
rect 1956 140324 2012 140326
rect 2036 140324 2092 140326
rect 2116 140324 2172 140326
rect 2196 140324 2252 140326
rect 3956 139834 4012 139836
rect 4036 139834 4092 139836
rect 4116 139834 4172 139836
rect 4196 139834 4252 139836
rect 3956 139782 3982 139834
rect 3982 139782 4012 139834
rect 4036 139782 4046 139834
rect 4046 139782 4092 139834
rect 4116 139782 4162 139834
rect 4162 139782 4172 139834
rect 4196 139782 4226 139834
rect 4226 139782 4252 139834
rect 3956 139780 4012 139782
rect 4036 139780 4092 139782
rect 4116 139780 4172 139782
rect 4196 139780 4252 139782
rect 1956 139290 2012 139292
rect 2036 139290 2092 139292
rect 2116 139290 2172 139292
rect 2196 139290 2252 139292
rect 1956 139238 1982 139290
rect 1982 139238 2012 139290
rect 2036 139238 2046 139290
rect 2046 139238 2092 139290
rect 2116 139238 2162 139290
rect 2162 139238 2172 139290
rect 2196 139238 2226 139290
rect 2226 139238 2252 139290
rect 1956 139236 2012 139238
rect 2036 139236 2092 139238
rect 2116 139236 2172 139238
rect 2196 139236 2252 139238
rect 3956 138746 4012 138748
rect 4036 138746 4092 138748
rect 4116 138746 4172 138748
rect 4196 138746 4252 138748
rect 3956 138694 3982 138746
rect 3982 138694 4012 138746
rect 4036 138694 4046 138746
rect 4046 138694 4092 138746
rect 4116 138694 4162 138746
rect 4162 138694 4172 138746
rect 4196 138694 4226 138746
rect 4226 138694 4252 138746
rect 3956 138692 4012 138694
rect 4036 138692 4092 138694
rect 4116 138692 4172 138694
rect 4196 138692 4252 138694
rect 1956 138202 2012 138204
rect 2036 138202 2092 138204
rect 2116 138202 2172 138204
rect 2196 138202 2252 138204
rect 1956 138150 1982 138202
rect 1982 138150 2012 138202
rect 2036 138150 2046 138202
rect 2046 138150 2092 138202
rect 2116 138150 2162 138202
rect 2162 138150 2172 138202
rect 2196 138150 2226 138202
rect 2226 138150 2252 138202
rect 1956 138148 2012 138150
rect 2036 138148 2092 138150
rect 2116 138148 2172 138150
rect 2196 138148 2252 138150
rect 3956 137658 4012 137660
rect 4036 137658 4092 137660
rect 4116 137658 4172 137660
rect 4196 137658 4252 137660
rect 3956 137606 3982 137658
rect 3982 137606 4012 137658
rect 4036 137606 4046 137658
rect 4046 137606 4092 137658
rect 4116 137606 4162 137658
rect 4162 137606 4172 137658
rect 4196 137606 4226 137658
rect 4226 137606 4252 137658
rect 3956 137604 4012 137606
rect 4036 137604 4092 137606
rect 4116 137604 4172 137606
rect 4196 137604 4252 137606
rect 1956 137114 2012 137116
rect 2036 137114 2092 137116
rect 2116 137114 2172 137116
rect 2196 137114 2252 137116
rect 1956 137062 1982 137114
rect 1982 137062 2012 137114
rect 2036 137062 2046 137114
rect 2046 137062 2092 137114
rect 2116 137062 2162 137114
rect 2162 137062 2172 137114
rect 2196 137062 2226 137114
rect 2226 137062 2252 137114
rect 1956 137060 2012 137062
rect 2036 137060 2092 137062
rect 2116 137060 2172 137062
rect 2196 137060 2252 137062
rect 3956 136570 4012 136572
rect 4036 136570 4092 136572
rect 4116 136570 4172 136572
rect 4196 136570 4252 136572
rect 3956 136518 3982 136570
rect 3982 136518 4012 136570
rect 4036 136518 4046 136570
rect 4046 136518 4092 136570
rect 4116 136518 4162 136570
rect 4162 136518 4172 136570
rect 4196 136518 4226 136570
rect 4226 136518 4252 136570
rect 3956 136516 4012 136518
rect 4036 136516 4092 136518
rect 4116 136516 4172 136518
rect 4196 136516 4252 136518
rect 1956 136026 2012 136028
rect 2036 136026 2092 136028
rect 2116 136026 2172 136028
rect 2196 136026 2252 136028
rect 1956 135974 1982 136026
rect 1982 135974 2012 136026
rect 2036 135974 2046 136026
rect 2046 135974 2092 136026
rect 2116 135974 2162 136026
rect 2162 135974 2172 136026
rect 2196 135974 2226 136026
rect 2226 135974 2252 136026
rect 1956 135972 2012 135974
rect 2036 135972 2092 135974
rect 2116 135972 2172 135974
rect 2196 135972 2252 135974
rect 3956 135482 4012 135484
rect 4036 135482 4092 135484
rect 4116 135482 4172 135484
rect 4196 135482 4252 135484
rect 3956 135430 3982 135482
rect 3982 135430 4012 135482
rect 4036 135430 4046 135482
rect 4046 135430 4092 135482
rect 4116 135430 4162 135482
rect 4162 135430 4172 135482
rect 4196 135430 4226 135482
rect 4226 135430 4252 135482
rect 3956 135428 4012 135430
rect 4036 135428 4092 135430
rect 4116 135428 4172 135430
rect 4196 135428 4252 135430
rect 1956 134938 2012 134940
rect 2036 134938 2092 134940
rect 2116 134938 2172 134940
rect 2196 134938 2252 134940
rect 1956 134886 1982 134938
rect 1982 134886 2012 134938
rect 2036 134886 2046 134938
rect 2046 134886 2092 134938
rect 2116 134886 2162 134938
rect 2162 134886 2172 134938
rect 2196 134886 2226 134938
rect 2226 134886 2252 134938
rect 1956 134884 2012 134886
rect 2036 134884 2092 134886
rect 2116 134884 2172 134886
rect 2196 134884 2252 134886
rect 3956 134394 4012 134396
rect 4036 134394 4092 134396
rect 4116 134394 4172 134396
rect 4196 134394 4252 134396
rect 3956 134342 3982 134394
rect 3982 134342 4012 134394
rect 4036 134342 4046 134394
rect 4046 134342 4092 134394
rect 4116 134342 4162 134394
rect 4162 134342 4172 134394
rect 4196 134342 4226 134394
rect 4226 134342 4252 134394
rect 3956 134340 4012 134342
rect 4036 134340 4092 134342
rect 4116 134340 4172 134342
rect 4196 134340 4252 134342
rect 1956 133850 2012 133852
rect 2036 133850 2092 133852
rect 2116 133850 2172 133852
rect 2196 133850 2252 133852
rect 1956 133798 1982 133850
rect 1982 133798 2012 133850
rect 2036 133798 2046 133850
rect 2046 133798 2092 133850
rect 2116 133798 2162 133850
rect 2162 133798 2172 133850
rect 2196 133798 2226 133850
rect 2226 133798 2252 133850
rect 1956 133796 2012 133798
rect 2036 133796 2092 133798
rect 2116 133796 2172 133798
rect 2196 133796 2252 133798
rect 3956 133306 4012 133308
rect 4036 133306 4092 133308
rect 4116 133306 4172 133308
rect 4196 133306 4252 133308
rect 3956 133254 3982 133306
rect 3982 133254 4012 133306
rect 4036 133254 4046 133306
rect 4046 133254 4092 133306
rect 4116 133254 4162 133306
rect 4162 133254 4172 133306
rect 4196 133254 4226 133306
rect 4226 133254 4252 133306
rect 3956 133252 4012 133254
rect 4036 133252 4092 133254
rect 4116 133252 4172 133254
rect 4196 133252 4252 133254
rect 1956 132762 2012 132764
rect 2036 132762 2092 132764
rect 2116 132762 2172 132764
rect 2196 132762 2252 132764
rect 1956 132710 1982 132762
rect 1982 132710 2012 132762
rect 2036 132710 2046 132762
rect 2046 132710 2092 132762
rect 2116 132710 2162 132762
rect 2162 132710 2172 132762
rect 2196 132710 2226 132762
rect 2226 132710 2252 132762
rect 1956 132708 2012 132710
rect 2036 132708 2092 132710
rect 2116 132708 2172 132710
rect 2196 132708 2252 132710
rect 3956 132218 4012 132220
rect 4036 132218 4092 132220
rect 4116 132218 4172 132220
rect 4196 132218 4252 132220
rect 3956 132166 3982 132218
rect 3982 132166 4012 132218
rect 4036 132166 4046 132218
rect 4046 132166 4092 132218
rect 4116 132166 4162 132218
rect 4162 132166 4172 132218
rect 4196 132166 4226 132218
rect 4226 132166 4252 132218
rect 3956 132164 4012 132166
rect 4036 132164 4092 132166
rect 4116 132164 4172 132166
rect 4196 132164 4252 132166
rect 1956 131674 2012 131676
rect 2036 131674 2092 131676
rect 2116 131674 2172 131676
rect 2196 131674 2252 131676
rect 1956 131622 1982 131674
rect 1982 131622 2012 131674
rect 2036 131622 2046 131674
rect 2046 131622 2092 131674
rect 2116 131622 2162 131674
rect 2162 131622 2172 131674
rect 2196 131622 2226 131674
rect 2226 131622 2252 131674
rect 1956 131620 2012 131622
rect 2036 131620 2092 131622
rect 2116 131620 2172 131622
rect 2196 131620 2252 131622
rect 3956 131130 4012 131132
rect 4036 131130 4092 131132
rect 4116 131130 4172 131132
rect 4196 131130 4252 131132
rect 3956 131078 3982 131130
rect 3982 131078 4012 131130
rect 4036 131078 4046 131130
rect 4046 131078 4092 131130
rect 4116 131078 4162 131130
rect 4162 131078 4172 131130
rect 4196 131078 4226 131130
rect 4226 131078 4252 131130
rect 3956 131076 4012 131078
rect 4036 131076 4092 131078
rect 4116 131076 4172 131078
rect 4196 131076 4252 131078
rect 1956 130586 2012 130588
rect 2036 130586 2092 130588
rect 2116 130586 2172 130588
rect 2196 130586 2252 130588
rect 1956 130534 1982 130586
rect 1982 130534 2012 130586
rect 2036 130534 2046 130586
rect 2046 130534 2092 130586
rect 2116 130534 2162 130586
rect 2162 130534 2172 130586
rect 2196 130534 2226 130586
rect 2226 130534 2252 130586
rect 1956 130532 2012 130534
rect 2036 130532 2092 130534
rect 2116 130532 2172 130534
rect 2196 130532 2252 130534
rect 3956 130042 4012 130044
rect 4036 130042 4092 130044
rect 4116 130042 4172 130044
rect 4196 130042 4252 130044
rect 3956 129990 3982 130042
rect 3982 129990 4012 130042
rect 4036 129990 4046 130042
rect 4046 129990 4092 130042
rect 4116 129990 4162 130042
rect 4162 129990 4172 130042
rect 4196 129990 4226 130042
rect 4226 129990 4252 130042
rect 3956 129988 4012 129990
rect 4036 129988 4092 129990
rect 4116 129988 4172 129990
rect 4196 129988 4252 129990
rect 1956 129498 2012 129500
rect 2036 129498 2092 129500
rect 2116 129498 2172 129500
rect 2196 129498 2252 129500
rect 1956 129446 1982 129498
rect 1982 129446 2012 129498
rect 2036 129446 2046 129498
rect 2046 129446 2092 129498
rect 2116 129446 2162 129498
rect 2162 129446 2172 129498
rect 2196 129446 2226 129498
rect 2226 129446 2252 129498
rect 1956 129444 2012 129446
rect 2036 129444 2092 129446
rect 2116 129444 2172 129446
rect 2196 129444 2252 129446
rect 3956 128954 4012 128956
rect 4036 128954 4092 128956
rect 4116 128954 4172 128956
rect 4196 128954 4252 128956
rect 3956 128902 3982 128954
rect 3982 128902 4012 128954
rect 4036 128902 4046 128954
rect 4046 128902 4092 128954
rect 4116 128902 4162 128954
rect 4162 128902 4172 128954
rect 4196 128902 4226 128954
rect 4226 128902 4252 128954
rect 3956 128900 4012 128902
rect 4036 128900 4092 128902
rect 4116 128900 4172 128902
rect 4196 128900 4252 128902
rect 1956 128410 2012 128412
rect 2036 128410 2092 128412
rect 2116 128410 2172 128412
rect 2196 128410 2252 128412
rect 1956 128358 1982 128410
rect 1982 128358 2012 128410
rect 2036 128358 2046 128410
rect 2046 128358 2092 128410
rect 2116 128358 2162 128410
rect 2162 128358 2172 128410
rect 2196 128358 2226 128410
rect 2226 128358 2252 128410
rect 1956 128356 2012 128358
rect 2036 128356 2092 128358
rect 2116 128356 2172 128358
rect 2196 128356 2252 128358
rect 3956 127866 4012 127868
rect 4036 127866 4092 127868
rect 4116 127866 4172 127868
rect 4196 127866 4252 127868
rect 3956 127814 3982 127866
rect 3982 127814 4012 127866
rect 4036 127814 4046 127866
rect 4046 127814 4092 127866
rect 4116 127814 4162 127866
rect 4162 127814 4172 127866
rect 4196 127814 4226 127866
rect 4226 127814 4252 127866
rect 3956 127812 4012 127814
rect 4036 127812 4092 127814
rect 4116 127812 4172 127814
rect 4196 127812 4252 127814
rect 1956 127322 2012 127324
rect 2036 127322 2092 127324
rect 2116 127322 2172 127324
rect 2196 127322 2252 127324
rect 1956 127270 1982 127322
rect 1982 127270 2012 127322
rect 2036 127270 2046 127322
rect 2046 127270 2092 127322
rect 2116 127270 2162 127322
rect 2162 127270 2172 127322
rect 2196 127270 2226 127322
rect 2226 127270 2252 127322
rect 1956 127268 2012 127270
rect 2036 127268 2092 127270
rect 2116 127268 2172 127270
rect 2196 127268 2252 127270
rect 3956 126778 4012 126780
rect 4036 126778 4092 126780
rect 4116 126778 4172 126780
rect 4196 126778 4252 126780
rect 3956 126726 3982 126778
rect 3982 126726 4012 126778
rect 4036 126726 4046 126778
rect 4046 126726 4092 126778
rect 4116 126726 4162 126778
rect 4162 126726 4172 126778
rect 4196 126726 4226 126778
rect 4226 126726 4252 126778
rect 3956 126724 4012 126726
rect 4036 126724 4092 126726
rect 4116 126724 4172 126726
rect 4196 126724 4252 126726
rect 1956 126234 2012 126236
rect 2036 126234 2092 126236
rect 2116 126234 2172 126236
rect 2196 126234 2252 126236
rect 1956 126182 1982 126234
rect 1982 126182 2012 126234
rect 2036 126182 2046 126234
rect 2046 126182 2092 126234
rect 2116 126182 2162 126234
rect 2162 126182 2172 126234
rect 2196 126182 2226 126234
rect 2226 126182 2252 126234
rect 1956 126180 2012 126182
rect 2036 126180 2092 126182
rect 2116 126180 2172 126182
rect 2196 126180 2252 126182
rect 3956 125690 4012 125692
rect 4036 125690 4092 125692
rect 4116 125690 4172 125692
rect 4196 125690 4252 125692
rect 3956 125638 3982 125690
rect 3982 125638 4012 125690
rect 4036 125638 4046 125690
rect 4046 125638 4092 125690
rect 4116 125638 4162 125690
rect 4162 125638 4172 125690
rect 4196 125638 4226 125690
rect 4226 125638 4252 125690
rect 3956 125636 4012 125638
rect 4036 125636 4092 125638
rect 4116 125636 4172 125638
rect 4196 125636 4252 125638
rect 1956 125146 2012 125148
rect 2036 125146 2092 125148
rect 2116 125146 2172 125148
rect 2196 125146 2252 125148
rect 1956 125094 1982 125146
rect 1982 125094 2012 125146
rect 2036 125094 2046 125146
rect 2046 125094 2092 125146
rect 2116 125094 2162 125146
rect 2162 125094 2172 125146
rect 2196 125094 2226 125146
rect 2226 125094 2252 125146
rect 1956 125092 2012 125094
rect 2036 125092 2092 125094
rect 2116 125092 2172 125094
rect 2196 125092 2252 125094
rect 3956 124602 4012 124604
rect 4036 124602 4092 124604
rect 4116 124602 4172 124604
rect 4196 124602 4252 124604
rect 3956 124550 3982 124602
rect 3982 124550 4012 124602
rect 4036 124550 4046 124602
rect 4046 124550 4092 124602
rect 4116 124550 4162 124602
rect 4162 124550 4172 124602
rect 4196 124550 4226 124602
rect 4226 124550 4252 124602
rect 3956 124548 4012 124550
rect 4036 124548 4092 124550
rect 4116 124548 4172 124550
rect 4196 124548 4252 124550
rect 1956 124058 2012 124060
rect 2036 124058 2092 124060
rect 2116 124058 2172 124060
rect 2196 124058 2252 124060
rect 1956 124006 1982 124058
rect 1982 124006 2012 124058
rect 2036 124006 2046 124058
rect 2046 124006 2092 124058
rect 2116 124006 2162 124058
rect 2162 124006 2172 124058
rect 2196 124006 2226 124058
rect 2226 124006 2252 124058
rect 1956 124004 2012 124006
rect 2036 124004 2092 124006
rect 2116 124004 2172 124006
rect 2196 124004 2252 124006
rect 3956 123514 4012 123516
rect 4036 123514 4092 123516
rect 4116 123514 4172 123516
rect 4196 123514 4252 123516
rect 3956 123462 3982 123514
rect 3982 123462 4012 123514
rect 4036 123462 4046 123514
rect 4046 123462 4092 123514
rect 4116 123462 4162 123514
rect 4162 123462 4172 123514
rect 4196 123462 4226 123514
rect 4226 123462 4252 123514
rect 3956 123460 4012 123462
rect 4036 123460 4092 123462
rect 4116 123460 4172 123462
rect 4196 123460 4252 123462
rect 1956 122970 2012 122972
rect 2036 122970 2092 122972
rect 2116 122970 2172 122972
rect 2196 122970 2252 122972
rect 1956 122918 1982 122970
rect 1982 122918 2012 122970
rect 2036 122918 2046 122970
rect 2046 122918 2092 122970
rect 2116 122918 2162 122970
rect 2162 122918 2172 122970
rect 2196 122918 2226 122970
rect 2226 122918 2252 122970
rect 1956 122916 2012 122918
rect 2036 122916 2092 122918
rect 2116 122916 2172 122918
rect 2196 122916 2252 122918
rect 3956 122426 4012 122428
rect 4036 122426 4092 122428
rect 4116 122426 4172 122428
rect 4196 122426 4252 122428
rect 3956 122374 3982 122426
rect 3982 122374 4012 122426
rect 4036 122374 4046 122426
rect 4046 122374 4092 122426
rect 4116 122374 4162 122426
rect 4162 122374 4172 122426
rect 4196 122374 4226 122426
rect 4226 122374 4252 122426
rect 3956 122372 4012 122374
rect 4036 122372 4092 122374
rect 4116 122372 4172 122374
rect 4196 122372 4252 122374
rect 1956 121882 2012 121884
rect 2036 121882 2092 121884
rect 2116 121882 2172 121884
rect 2196 121882 2252 121884
rect 1956 121830 1982 121882
rect 1982 121830 2012 121882
rect 2036 121830 2046 121882
rect 2046 121830 2092 121882
rect 2116 121830 2162 121882
rect 2162 121830 2172 121882
rect 2196 121830 2226 121882
rect 2226 121830 2252 121882
rect 1956 121828 2012 121830
rect 2036 121828 2092 121830
rect 2116 121828 2172 121830
rect 2196 121828 2252 121830
rect 3956 121338 4012 121340
rect 4036 121338 4092 121340
rect 4116 121338 4172 121340
rect 4196 121338 4252 121340
rect 3956 121286 3982 121338
rect 3982 121286 4012 121338
rect 4036 121286 4046 121338
rect 4046 121286 4092 121338
rect 4116 121286 4162 121338
rect 4162 121286 4172 121338
rect 4196 121286 4226 121338
rect 4226 121286 4252 121338
rect 3956 121284 4012 121286
rect 4036 121284 4092 121286
rect 4116 121284 4172 121286
rect 4196 121284 4252 121286
rect 1956 120794 2012 120796
rect 2036 120794 2092 120796
rect 2116 120794 2172 120796
rect 2196 120794 2252 120796
rect 1956 120742 1982 120794
rect 1982 120742 2012 120794
rect 2036 120742 2046 120794
rect 2046 120742 2092 120794
rect 2116 120742 2162 120794
rect 2162 120742 2172 120794
rect 2196 120742 2226 120794
rect 2226 120742 2252 120794
rect 1956 120740 2012 120742
rect 2036 120740 2092 120742
rect 2116 120740 2172 120742
rect 2196 120740 2252 120742
rect 3956 120250 4012 120252
rect 4036 120250 4092 120252
rect 4116 120250 4172 120252
rect 4196 120250 4252 120252
rect 3956 120198 3982 120250
rect 3982 120198 4012 120250
rect 4036 120198 4046 120250
rect 4046 120198 4092 120250
rect 4116 120198 4162 120250
rect 4162 120198 4172 120250
rect 4196 120198 4226 120250
rect 4226 120198 4252 120250
rect 3956 120196 4012 120198
rect 4036 120196 4092 120198
rect 4116 120196 4172 120198
rect 4196 120196 4252 120198
rect 1956 119706 2012 119708
rect 2036 119706 2092 119708
rect 2116 119706 2172 119708
rect 2196 119706 2252 119708
rect 1956 119654 1982 119706
rect 1982 119654 2012 119706
rect 2036 119654 2046 119706
rect 2046 119654 2092 119706
rect 2116 119654 2162 119706
rect 2162 119654 2172 119706
rect 2196 119654 2226 119706
rect 2226 119654 2252 119706
rect 1956 119652 2012 119654
rect 2036 119652 2092 119654
rect 2116 119652 2172 119654
rect 2196 119652 2252 119654
rect 3956 119162 4012 119164
rect 4036 119162 4092 119164
rect 4116 119162 4172 119164
rect 4196 119162 4252 119164
rect 3956 119110 3982 119162
rect 3982 119110 4012 119162
rect 4036 119110 4046 119162
rect 4046 119110 4092 119162
rect 4116 119110 4162 119162
rect 4162 119110 4172 119162
rect 4196 119110 4226 119162
rect 4226 119110 4252 119162
rect 3956 119108 4012 119110
rect 4036 119108 4092 119110
rect 4116 119108 4172 119110
rect 4196 119108 4252 119110
rect 1956 118618 2012 118620
rect 2036 118618 2092 118620
rect 2116 118618 2172 118620
rect 2196 118618 2252 118620
rect 1956 118566 1982 118618
rect 1982 118566 2012 118618
rect 2036 118566 2046 118618
rect 2046 118566 2092 118618
rect 2116 118566 2162 118618
rect 2162 118566 2172 118618
rect 2196 118566 2226 118618
rect 2226 118566 2252 118618
rect 1956 118564 2012 118566
rect 2036 118564 2092 118566
rect 2116 118564 2172 118566
rect 2196 118564 2252 118566
rect 3956 118074 4012 118076
rect 4036 118074 4092 118076
rect 4116 118074 4172 118076
rect 4196 118074 4252 118076
rect 3956 118022 3982 118074
rect 3982 118022 4012 118074
rect 4036 118022 4046 118074
rect 4046 118022 4092 118074
rect 4116 118022 4162 118074
rect 4162 118022 4172 118074
rect 4196 118022 4226 118074
rect 4226 118022 4252 118074
rect 3956 118020 4012 118022
rect 4036 118020 4092 118022
rect 4116 118020 4172 118022
rect 4196 118020 4252 118022
rect 1956 117530 2012 117532
rect 2036 117530 2092 117532
rect 2116 117530 2172 117532
rect 2196 117530 2252 117532
rect 1956 117478 1982 117530
rect 1982 117478 2012 117530
rect 2036 117478 2046 117530
rect 2046 117478 2092 117530
rect 2116 117478 2162 117530
rect 2162 117478 2172 117530
rect 2196 117478 2226 117530
rect 2226 117478 2252 117530
rect 1956 117476 2012 117478
rect 2036 117476 2092 117478
rect 2116 117476 2172 117478
rect 2196 117476 2252 117478
rect 3956 116986 4012 116988
rect 4036 116986 4092 116988
rect 4116 116986 4172 116988
rect 4196 116986 4252 116988
rect 3956 116934 3982 116986
rect 3982 116934 4012 116986
rect 4036 116934 4046 116986
rect 4046 116934 4092 116986
rect 4116 116934 4162 116986
rect 4162 116934 4172 116986
rect 4196 116934 4226 116986
rect 4226 116934 4252 116986
rect 3956 116932 4012 116934
rect 4036 116932 4092 116934
rect 4116 116932 4172 116934
rect 4196 116932 4252 116934
rect 1956 116442 2012 116444
rect 2036 116442 2092 116444
rect 2116 116442 2172 116444
rect 2196 116442 2252 116444
rect 1956 116390 1982 116442
rect 1982 116390 2012 116442
rect 2036 116390 2046 116442
rect 2046 116390 2092 116442
rect 2116 116390 2162 116442
rect 2162 116390 2172 116442
rect 2196 116390 2226 116442
rect 2226 116390 2252 116442
rect 1956 116388 2012 116390
rect 2036 116388 2092 116390
rect 2116 116388 2172 116390
rect 2196 116388 2252 116390
rect 3956 115898 4012 115900
rect 4036 115898 4092 115900
rect 4116 115898 4172 115900
rect 4196 115898 4252 115900
rect 3956 115846 3982 115898
rect 3982 115846 4012 115898
rect 4036 115846 4046 115898
rect 4046 115846 4092 115898
rect 4116 115846 4162 115898
rect 4162 115846 4172 115898
rect 4196 115846 4226 115898
rect 4226 115846 4252 115898
rect 3956 115844 4012 115846
rect 4036 115844 4092 115846
rect 4116 115844 4172 115846
rect 4196 115844 4252 115846
rect 1956 115354 2012 115356
rect 2036 115354 2092 115356
rect 2116 115354 2172 115356
rect 2196 115354 2252 115356
rect 1956 115302 1982 115354
rect 1982 115302 2012 115354
rect 2036 115302 2046 115354
rect 2046 115302 2092 115354
rect 2116 115302 2162 115354
rect 2162 115302 2172 115354
rect 2196 115302 2226 115354
rect 2226 115302 2252 115354
rect 1956 115300 2012 115302
rect 2036 115300 2092 115302
rect 2116 115300 2172 115302
rect 2196 115300 2252 115302
rect 3956 114810 4012 114812
rect 4036 114810 4092 114812
rect 4116 114810 4172 114812
rect 4196 114810 4252 114812
rect 3956 114758 3982 114810
rect 3982 114758 4012 114810
rect 4036 114758 4046 114810
rect 4046 114758 4092 114810
rect 4116 114758 4162 114810
rect 4162 114758 4172 114810
rect 4196 114758 4226 114810
rect 4226 114758 4252 114810
rect 3956 114756 4012 114758
rect 4036 114756 4092 114758
rect 4116 114756 4172 114758
rect 4196 114756 4252 114758
rect 1956 114266 2012 114268
rect 2036 114266 2092 114268
rect 2116 114266 2172 114268
rect 2196 114266 2252 114268
rect 1956 114214 1982 114266
rect 1982 114214 2012 114266
rect 2036 114214 2046 114266
rect 2046 114214 2092 114266
rect 2116 114214 2162 114266
rect 2162 114214 2172 114266
rect 2196 114214 2226 114266
rect 2226 114214 2252 114266
rect 1956 114212 2012 114214
rect 2036 114212 2092 114214
rect 2116 114212 2172 114214
rect 2196 114212 2252 114214
rect 3956 113722 4012 113724
rect 4036 113722 4092 113724
rect 4116 113722 4172 113724
rect 4196 113722 4252 113724
rect 3956 113670 3982 113722
rect 3982 113670 4012 113722
rect 4036 113670 4046 113722
rect 4046 113670 4092 113722
rect 4116 113670 4162 113722
rect 4162 113670 4172 113722
rect 4196 113670 4226 113722
rect 4226 113670 4252 113722
rect 3956 113668 4012 113670
rect 4036 113668 4092 113670
rect 4116 113668 4172 113670
rect 4196 113668 4252 113670
rect 1956 113178 2012 113180
rect 2036 113178 2092 113180
rect 2116 113178 2172 113180
rect 2196 113178 2252 113180
rect 1956 113126 1982 113178
rect 1982 113126 2012 113178
rect 2036 113126 2046 113178
rect 2046 113126 2092 113178
rect 2116 113126 2162 113178
rect 2162 113126 2172 113178
rect 2196 113126 2226 113178
rect 2226 113126 2252 113178
rect 1956 113124 2012 113126
rect 2036 113124 2092 113126
rect 2116 113124 2172 113126
rect 2196 113124 2252 113126
rect 3956 112634 4012 112636
rect 4036 112634 4092 112636
rect 4116 112634 4172 112636
rect 4196 112634 4252 112636
rect 3956 112582 3982 112634
rect 3982 112582 4012 112634
rect 4036 112582 4046 112634
rect 4046 112582 4092 112634
rect 4116 112582 4162 112634
rect 4162 112582 4172 112634
rect 4196 112582 4226 112634
rect 4226 112582 4252 112634
rect 3956 112580 4012 112582
rect 4036 112580 4092 112582
rect 4116 112580 4172 112582
rect 4196 112580 4252 112582
rect 1956 112090 2012 112092
rect 2036 112090 2092 112092
rect 2116 112090 2172 112092
rect 2196 112090 2252 112092
rect 1956 112038 1982 112090
rect 1982 112038 2012 112090
rect 2036 112038 2046 112090
rect 2046 112038 2092 112090
rect 2116 112038 2162 112090
rect 2162 112038 2172 112090
rect 2196 112038 2226 112090
rect 2226 112038 2252 112090
rect 1956 112036 2012 112038
rect 2036 112036 2092 112038
rect 2116 112036 2172 112038
rect 2196 112036 2252 112038
rect 3956 111546 4012 111548
rect 4036 111546 4092 111548
rect 4116 111546 4172 111548
rect 4196 111546 4252 111548
rect 3956 111494 3982 111546
rect 3982 111494 4012 111546
rect 4036 111494 4046 111546
rect 4046 111494 4092 111546
rect 4116 111494 4162 111546
rect 4162 111494 4172 111546
rect 4196 111494 4226 111546
rect 4226 111494 4252 111546
rect 3956 111492 4012 111494
rect 4036 111492 4092 111494
rect 4116 111492 4172 111494
rect 4196 111492 4252 111494
rect 1956 111002 2012 111004
rect 2036 111002 2092 111004
rect 2116 111002 2172 111004
rect 2196 111002 2252 111004
rect 1956 110950 1982 111002
rect 1982 110950 2012 111002
rect 2036 110950 2046 111002
rect 2046 110950 2092 111002
rect 2116 110950 2162 111002
rect 2162 110950 2172 111002
rect 2196 110950 2226 111002
rect 2226 110950 2252 111002
rect 1956 110948 2012 110950
rect 2036 110948 2092 110950
rect 2116 110948 2172 110950
rect 2196 110948 2252 110950
rect 3956 110458 4012 110460
rect 4036 110458 4092 110460
rect 4116 110458 4172 110460
rect 4196 110458 4252 110460
rect 3956 110406 3982 110458
rect 3982 110406 4012 110458
rect 4036 110406 4046 110458
rect 4046 110406 4092 110458
rect 4116 110406 4162 110458
rect 4162 110406 4172 110458
rect 4196 110406 4226 110458
rect 4226 110406 4252 110458
rect 3956 110404 4012 110406
rect 4036 110404 4092 110406
rect 4116 110404 4172 110406
rect 4196 110404 4252 110406
rect 1956 109914 2012 109916
rect 2036 109914 2092 109916
rect 2116 109914 2172 109916
rect 2196 109914 2252 109916
rect 1956 109862 1982 109914
rect 1982 109862 2012 109914
rect 2036 109862 2046 109914
rect 2046 109862 2092 109914
rect 2116 109862 2162 109914
rect 2162 109862 2172 109914
rect 2196 109862 2226 109914
rect 2226 109862 2252 109914
rect 1956 109860 2012 109862
rect 2036 109860 2092 109862
rect 2116 109860 2172 109862
rect 2196 109860 2252 109862
rect 3956 109370 4012 109372
rect 4036 109370 4092 109372
rect 4116 109370 4172 109372
rect 4196 109370 4252 109372
rect 3956 109318 3982 109370
rect 3982 109318 4012 109370
rect 4036 109318 4046 109370
rect 4046 109318 4092 109370
rect 4116 109318 4162 109370
rect 4162 109318 4172 109370
rect 4196 109318 4226 109370
rect 4226 109318 4252 109370
rect 3956 109316 4012 109318
rect 4036 109316 4092 109318
rect 4116 109316 4172 109318
rect 4196 109316 4252 109318
rect 1956 108826 2012 108828
rect 2036 108826 2092 108828
rect 2116 108826 2172 108828
rect 2196 108826 2252 108828
rect 1956 108774 1982 108826
rect 1982 108774 2012 108826
rect 2036 108774 2046 108826
rect 2046 108774 2092 108826
rect 2116 108774 2162 108826
rect 2162 108774 2172 108826
rect 2196 108774 2226 108826
rect 2226 108774 2252 108826
rect 1956 108772 2012 108774
rect 2036 108772 2092 108774
rect 2116 108772 2172 108774
rect 2196 108772 2252 108774
rect 3956 108282 4012 108284
rect 4036 108282 4092 108284
rect 4116 108282 4172 108284
rect 4196 108282 4252 108284
rect 3956 108230 3982 108282
rect 3982 108230 4012 108282
rect 4036 108230 4046 108282
rect 4046 108230 4092 108282
rect 4116 108230 4162 108282
rect 4162 108230 4172 108282
rect 4196 108230 4226 108282
rect 4226 108230 4252 108282
rect 3956 108228 4012 108230
rect 4036 108228 4092 108230
rect 4116 108228 4172 108230
rect 4196 108228 4252 108230
rect 1956 107738 2012 107740
rect 2036 107738 2092 107740
rect 2116 107738 2172 107740
rect 2196 107738 2252 107740
rect 1956 107686 1982 107738
rect 1982 107686 2012 107738
rect 2036 107686 2046 107738
rect 2046 107686 2092 107738
rect 2116 107686 2162 107738
rect 2162 107686 2172 107738
rect 2196 107686 2226 107738
rect 2226 107686 2252 107738
rect 1956 107684 2012 107686
rect 2036 107684 2092 107686
rect 2116 107684 2172 107686
rect 2196 107684 2252 107686
rect 3956 107194 4012 107196
rect 4036 107194 4092 107196
rect 4116 107194 4172 107196
rect 4196 107194 4252 107196
rect 3956 107142 3982 107194
rect 3982 107142 4012 107194
rect 4036 107142 4046 107194
rect 4046 107142 4092 107194
rect 4116 107142 4162 107194
rect 4162 107142 4172 107194
rect 4196 107142 4226 107194
rect 4226 107142 4252 107194
rect 3956 107140 4012 107142
rect 4036 107140 4092 107142
rect 4116 107140 4172 107142
rect 4196 107140 4252 107142
rect 1956 106650 2012 106652
rect 2036 106650 2092 106652
rect 2116 106650 2172 106652
rect 2196 106650 2252 106652
rect 1956 106598 1982 106650
rect 1982 106598 2012 106650
rect 2036 106598 2046 106650
rect 2046 106598 2092 106650
rect 2116 106598 2162 106650
rect 2162 106598 2172 106650
rect 2196 106598 2226 106650
rect 2226 106598 2252 106650
rect 1956 106596 2012 106598
rect 2036 106596 2092 106598
rect 2116 106596 2172 106598
rect 2196 106596 2252 106598
rect 3956 106106 4012 106108
rect 4036 106106 4092 106108
rect 4116 106106 4172 106108
rect 4196 106106 4252 106108
rect 3956 106054 3982 106106
rect 3982 106054 4012 106106
rect 4036 106054 4046 106106
rect 4046 106054 4092 106106
rect 4116 106054 4162 106106
rect 4162 106054 4172 106106
rect 4196 106054 4226 106106
rect 4226 106054 4252 106106
rect 3956 106052 4012 106054
rect 4036 106052 4092 106054
rect 4116 106052 4172 106054
rect 4196 106052 4252 106054
rect 84382 186224 84438 186280
rect 4802 182980 4858 183016
rect 4802 182960 4804 182980
rect 4804 182960 4856 182980
rect 4856 182960 4858 182980
rect 5170 182960 5226 183016
rect 4802 181892 4858 181928
rect 4802 181872 4804 181892
rect 4804 181872 4856 181892
rect 4856 181872 4858 181892
rect 4618 180140 4620 180160
rect 4620 180140 4672 180160
rect 4672 180140 4674 180160
rect 4618 180104 4674 180140
rect 4526 179052 4528 179072
rect 4528 179052 4580 179072
rect 4580 179052 4582 179072
rect 4526 179016 4582 179052
rect 4710 176976 4766 177032
rect 1956 105562 2012 105564
rect 2036 105562 2092 105564
rect 2116 105562 2172 105564
rect 2196 105562 2252 105564
rect 1956 105510 1982 105562
rect 1982 105510 2012 105562
rect 2036 105510 2046 105562
rect 2046 105510 2092 105562
rect 2116 105510 2162 105562
rect 2162 105510 2172 105562
rect 2196 105510 2226 105562
rect 2226 105510 2252 105562
rect 1956 105508 2012 105510
rect 2036 105508 2092 105510
rect 2116 105508 2172 105510
rect 2196 105508 2252 105510
rect 3956 105018 4012 105020
rect 4036 105018 4092 105020
rect 4116 105018 4172 105020
rect 4196 105018 4252 105020
rect 3956 104966 3982 105018
rect 3982 104966 4012 105018
rect 4036 104966 4046 105018
rect 4046 104966 4092 105018
rect 4116 104966 4162 105018
rect 4162 104966 4172 105018
rect 4196 104966 4226 105018
rect 4226 104966 4252 105018
rect 3956 104964 4012 104966
rect 4036 104964 4092 104966
rect 4116 104964 4172 104966
rect 4196 104964 4252 104966
rect 1956 104474 2012 104476
rect 2036 104474 2092 104476
rect 2116 104474 2172 104476
rect 2196 104474 2252 104476
rect 1956 104422 1982 104474
rect 1982 104422 2012 104474
rect 2036 104422 2046 104474
rect 2046 104422 2092 104474
rect 2116 104422 2162 104474
rect 2162 104422 2172 104474
rect 2196 104422 2226 104474
rect 2226 104422 2252 104474
rect 1956 104420 2012 104422
rect 2036 104420 2092 104422
rect 2116 104420 2172 104422
rect 2196 104420 2252 104422
rect 3956 103930 4012 103932
rect 4036 103930 4092 103932
rect 4116 103930 4172 103932
rect 4196 103930 4252 103932
rect 3956 103878 3982 103930
rect 3982 103878 4012 103930
rect 4036 103878 4046 103930
rect 4046 103878 4092 103930
rect 4116 103878 4162 103930
rect 4162 103878 4172 103930
rect 4196 103878 4226 103930
rect 4226 103878 4252 103930
rect 3956 103876 4012 103878
rect 4036 103876 4092 103878
rect 4116 103876 4172 103878
rect 4196 103876 4252 103878
rect 1956 103386 2012 103388
rect 2036 103386 2092 103388
rect 2116 103386 2172 103388
rect 2196 103386 2252 103388
rect 1956 103334 1982 103386
rect 1982 103334 2012 103386
rect 2036 103334 2046 103386
rect 2046 103334 2092 103386
rect 2116 103334 2162 103386
rect 2162 103334 2172 103386
rect 2196 103334 2226 103386
rect 2226 103334 2252 103386
rect 1956 103332 2012 103334
rect 2036 103332 2092 103334
rect 2116 103332 2172 103334
rect 2196 103332 2252 103334
rect 3956 102842 4012 102844
rect 4036 102842 4092 102844
rect 4116 102842 4172 102844
rect 4196 102842 4252 102844
rect 3956 102790 3982 102842
rect 3982 102790 4012 102842
rect 4036 102790 4046 102842
rect 4046 102790 4092 102842
rect 4116 102790 4162 102842
rect 4162 102790 4172 102842
rect 4196 102790 4226 102842
rect 4226 102790 4252 102842
rect 3956 102788 4012 102790
rect 4036 102788 4092 102790
rect 4116 102788 4172 102790
rect 4196 102788 4252 102790
rect 1956 102298 2012 102300
rect 2036 102298 2092 102300
rect 2116 102298 2172 102300
rect 2196 102298 2252 102300
rect 1956 102246 1982 102298
rect 1982 102246 2012 102298
rect 2036 102246 2046 102298
rect 2046 102246 2092 102298
rect 2116 102246 2162 102298
rect 2162 102246 2172 102298
rect 2196 102246 2226 102298
rect 2226 102246 2252 102298
rect 1956 102244 2012 102246
rect 2036 102244 2092 102246
rect 2116 102244 2172 102246
rect 2196 102244 2252 102246
rect 3956 101754 4012 101756
rect 4036 101754 4092 101756
rect 4116 101754 4172 101756
rect 4196 101754 4252 101756
rect 3956 101702 3982 101754
rect 3982 101702 4012 101754
rect 4036 101702 4046 101754
rect 4046 101702 4092 101754
rect 4116 101702 4162 101754
rect 4162 101702 4172 101754
rect 4196 101702 4226 101754
rect 4226 101702 4252 101754
rect 3956 101700 4012 101702
rect 4036 101700 4092 101702
rect 4116 101700 4172 101702
rect 4196 101700 4252 101702
rect 1956 101210 2012 101212
rect 2036 101210 2092 101212
rect 2116 101210 2172 101212
rect 2196 101210 2252 101212
rect 1956 101158 1982 101210
rect 1982 101158 2012 101210
rect 2036 101158 2046 101210
rect 2046 101158 2092 101210
rect 2116 101158 2162 101210
rect 2162 101158 2172 101210
rect 2196 101158 2226 101210
rect 2226 101158 2252 101210
rect 1956 101156 2012 101158
rect 2036 101156 2092 101158
rect 2116 101156 2172 101158
rect 2196 101156 2252 101158
rect 3956 100666 4012 100668
rect 4036 100666 4092 100668
rect 4116 100666 4172 100668
rect 4196 100666 4252 100668
rect 3956 100614 3982 100666
rect 3982 100614 4012 100666
rect 4036 100614 4046 100666
rect 4046 100614 4092 100666
rect 4116 100614 4162 100666
rect 4162 100614 4172 100666
rect 4196 100614 4226 100666
rect 4226 100614 4252 100666
rect 3956 100612 4012 100614
rect 4036 100612 4092 100614
rect 4116 100612 4172 100614
rect 4196 100612 4252 100614
rect 1956 100122 2012 100124
rect 2036 100122 2092 100124
rect 2116 100122 2172 100124
rect 2196 100122 2252 100124
rect 1956 100070 1982 100122
rect 1982 100070 2012 100122
rect 2036 100070 2046 100122
rect 2046 100070 2092 100122
rect 2116 100070 2162 100122
rect 2162 100070 2172 100122
rect 2196 100070 2226 100122
rect 2226 100070 2252 100122
rect 1956 100068 2012 100070
rect 2036 100068 2092 100070
rect 2116 100068 2172 100070
rect 2196 100068 2252 100070
rect 3956 99578 4012 99580
rect 4036 99578 4092 99580
rect 4116 99578 4172 99580
rect 4196 99578 4252 99580
rect 3956 99526 3982 99578
rect 3982 99526 4012 99578
rect 4036 99526 4046 99578
rect 4046 99526 4092 99578
rect 4116 99526 4162 99578
rect 4162 99526 4172 99578
rect 4196 99526 4226 99578
rect 4226 99526 4252 99578
rect 3956 99524 4012 99526
rect 4036 99524 4092 99526
rect 4116 99524 4172 99526
rect 4196 99524 4252 99526
rect 1956 99034 2012 99036
rect 2036 99034 2092 99036
rect 2116 99034 2172 99036
rect 2196 99034 2252 99036
rect 1956 98982 1982 99034
rect 1982 98982 2012 99034
rect 2036 98982 2046 99034
rect 2046 98982 2092 99034
rect 2116 98982 2162 99034
rect 2162 98982 2172 99034
rect 2196 98982 2226 99034
rect 2226 98982 2252 99034
rect 1956 98980 2012 98982
rect 2036 98980 2092 98982
rect 2116 98980 2172 98982
rect 2196 98980 2252 98982
rect 3956 98490 4012 98492
rect 4036 98490 4092 98492
rect 4116 98490 4172 98492
rect 4196 98490 4252 98492
rect 3956 98438 3982 98490
rect 3982 98438 4012 98490
rect 4036 98438 4046 98490
rect 4046 98438 4092 98490
rect 4116 98438 4162 98490
rect 4162 98438 4172 98490
rect 4196 98438 4226 98490
rect 4226 98438 4252 98490
rect 3956 98436 4012 98438
rect 4036 98436 4092 98438
rect 4116 98436 4172 98438
rect 4196 98436 4252 98438
rect 1956 97946 2012 97948
rect 2036 97946 2092 97948
rect 2116 97946 2172 97948
rect 2196 97946 2252 97948
rect 1956 97894 1982 97946
rect 1982 97894 2012 97946
rect 2036 97894 2046 97946
rect 2046 97894 2092 97946
rect 2116 97894 2162 97946
rect 2162 97894 2172 97946
rect 2196 97894 2226 97946
rect 2226 97894 2252 97946
rect 1956 97892 2012 97894
rect 2036 97892 2092 97894
rect 2116 97892 2172 97894
rect 2196 97892 2252 97894
rect 1956 96858 2012 96860
rect 2036 96858 2092 96860
rect 2116 96858 2172 96860
rect 2196 96858 2252 96860
rect 1956 96806 1982 96858
rect 1982 96806 2012 96858
rect 2036 96806 2046 96858
rect 2046 96806 2092 96858
rect 2116 96806 2162 96858
rect 2162 96806 2172 96858
rect 2196 96806 2226 96858
rect 2226 96806 2252 96858
rect 1956 96804 2012 96806
rect 2036 96804 2092 96806
rect 2116 96804 2172 96806
rect 2196 96804 2252 96806
rect 1956 95770 2012 95772
rect 2036 95770 2092 95772
rect 2116 95770 2172 95772
rect 2196 95770 2252 95772
rect 1956 95718 1982 95770
rect 1982 95718 2012 95770
rect 2036 95718 2046 95770
rect 2046 95718 2092 95770
rect 2116 95718 2162 95770
rect 2162 95718 2172 95770
rect 2196 95718 2226 95770
rect 2226 95718 2252 95770
rect 1956 95716 2012 95718
rect 2036 95716 2092 95718
rect 2116 95716 2172 95718
rect 2196 95716 2252 95718
rect 1956 94682 2012 94684
rect 2036 94682 2092 94684
rect 2116 94682 2172 94684
rect 2196 94682 2252 94684
rect 1956 94630 1982 94682
rect 1982 94630 2012 94682
rect 2036 94630 2046 94682
rect 2046 94630 2092 94682
rect 2116 94630 2162 94682
rect 2162 94630 2172 94682
rect 2196 94630 2226 94682
rect 2226 94630 2252 94682
rect 1956 94628 2012 94630
rect 2036 94628 2092 94630
rect 2116 94628 2172 94630
rect 2196 94628 2252 94630
rect 1956 93594 2012 93596
rect 2036 93594 2092 93596
rect 2116 93594 2172 93596
rect 2196 93594 2252 93596
rect 1956 93542 1982 93594
rect 1982 93542 2012 93594
rect 2036 93542 2046 93594
rect 2046 93542 2092 93594
rect 2116 93542 2162 93594
rect 2162 93542 2172 93594
rect 2196 93542 2226 93594
rect 2226 93542 2252 93594
rect 1956 93540 2012 93542
rect 2036 93540 2092 93542
rect 2116 93540 2172 93542
rect 2196 93540 2252 93542
rect 1956 92506 2012 92508
rect 2036 92506 2092 92508
rect 2116 92506 2172 92508
rect 2196 92506 2252 92508
rect 1956 92454 1982 92506
rect 1982 92454 2012 92506
rect 2036 92454 2046 92506
rect 2046 92454 2092 92506
rect 2116 92454 2162 92506
rect 2162 92454 2172 92506
rect 2196 92454 2226 92506
rect 2226 92454 2252 92506
rect 1956 92452 2012 92454
rect 2036 92452 2092 92454
rect 2116 92452 2172 92454
rect 2196 92452 2252 92454
rect 1956 91418 2012 91420
rect 2036 91418 2092 91420
rect 2116 91418 2172 91420
rect 2196 91418 2252 91420
rect 1956 91366 1982 91418
rect 1982 91366 2012 91418
rect 2036 91366 2046 91418
rect 2046 91366 2092 91418
rect 2116 91366 2162 91418
rect 2162 91366 2172 91418
rect 2196 91366 2226 91418
rect 2226 91366 2252 91418
rect 1956 91364 2012 91366
rect 2036 91364 2092 91366
rect 2116 91364 2172 91366
rect 2196 91364 2252 91366
rect 1956 90330 2012 90332
rect 2036 90330 2092 90332
rect 2116 90330 2172 90332
rect 2196 90330 2252 90332
rect 1956 90278 1982 90330
rect 1982 90278 2012 90330
rect 2036 90278 2046 90330
rect 2046 90278 2092 90330
rect 2116 90278 2162 90330
rect 2162 90278 2172 90330
rect 2196 90278 2226 90330
rect 2226 90278 2252 90330
rect 1956 90276 2012 90278
rect 2036 90276 2092 90278
rect 2116 90276 2172 90278
rect 2196 90276 2252 90278
rect 1956 89242 2012 89244
rect 2036 89242 2092 89244
rect 2116 89242 2172 89244
rect 2196 89242 2252 89244
rect 1956 89190 1982 89242
rect 1982 89190 2012 89242
rect 2036 89190 2046 89242
rect 2046 89190 2092 89242
rect 2116 89190 2162 89242
rect 2162 89190 2172 89242
rect 2196 89190 2226 89242
rect 2226 89190 2252 89242
rect 1956 89188 2012 89190
rect 2036 89188 2092 89190
rect 2116 89188 2172 89190
rect 2196 89188 2252 89190
rect 1956 88154 2012 88156
rect 2036 88154 2092 88156
rect 2116 88154 2172 88156
rect 2196 88154 2252 88156
rect 1956 88102 1982 88154
rect 1982 88102 2012 88154
rect 2036 88102 2046 88154
rect 2046 88102 2092 88154
rect 2116 88102 2162 88154
rect 2162 88102 2172 88154
rect 2196 88102 2226 88154
rect 2226 88102 2252 88154
rect 1956 88100 2012 88102
rect 2036 88100 2092 88102
rect 2116 88100 2172 88102
rect 2196 88100 2252 88102
rect 1956 87066 2012 87068
rect 2036 87066 2092 87068
rect 2116 87066 2172 87068
rect 2196 87066 2252 87068
rect 1956 87014 1982 87066
rect 1982 87014 2012 87066
rect 2036 87014 2046 87066
rect 2046 87014 2092 87066
rect 2116 87014 2162 87066
rect 2162 87014 2172 87066
rect 2196 87014 2226 87066
rect 2226 87014 2252 87066
rect 1956 87012 2012 87014
rect 2036 87012 2092 87014
rect 2116 87012 2172 87014
rect 2196 87012 2252 87014
rect 1956 85978 2012 85980
rect 2036 85978 2092 85980
rect 2116 85978 2172 85980
rect 2196 85978 2252 85980
rect 1956 85926 1982 85978
rect 1982 85926 2012 85978
rect 2036 85926 2046 85978
rect 2046 85926 2092 85978
rect 2116 85926 2162 85978
rect 2162 85926 2172 85978
rect 2196 85926 2226 85978
rect 2226 85926 2252 85978
rect 1956 85924 2012 85926
rect 2036 85924 2092 85926
rect 2116 85924 2172 85926
rect 2196 85924 2252 85926
rect 1956 84890 2012 84892
rect 2036 84890 2092 84892
rect 2116 84890 2172 84892
rect 2196 84890 2252 84892
rect 1956 84838 1982 84890
rect 1982 84838 2012 84890
rect 2036 84838 2046 84890
rect 2046 84838 2092 84890
rect 2116 84838 2162 84890
rect 2162 84838 2172 84890
rect 2196 84838 2226 84890
rect 2226 84838 2252 84890
rect 1956 84836 2012 84838
rect 2036 84836 2092 84838
rect 2116 84836 2172 84838
rect 2196 84836 2252 84838
rect 3956 97402 4012 97404
rect 4036 97402 4092 97404
rect 4116 97402 4172 97404
rect 4196 97402 4252 97404
rect 3956 97350 3982 97402
rect 3982 97350 4012 97402
rect 4036 97350 4046 97402
rect 4046 97350 4092 97402
rect 4116 97350 4162 97402
rect 4162 97350 4172 97402
rect 4196 97350 4226 97402
rect 4226 97350 4252 97402
rect 3956 97348 4012 97350
rect 4036 97348 4092 97350
rect 4116 97348 4172 97350
rect 4196 97348 4252 97350
rect 1956 83802 2012 83804
rect 2036 83802 2092 83804
rect 2116 83802 2172 83804
rect 2196 83802 2252 83804
rect 1956 83750 1982 83802
rect 1982 83750 2012 83802
rect 2036 83750 2046 83802
rect 2046 83750 2092 83802
rect 2116 83750 2162 83802
rect 2162 83750 2172 83802
rect 2196 83750 2226 83802
rect 2226 83750 2252 83802
rect 1956 83748 2012 83750
rect 2036 83748 2092 83750
rect 2116 83748 2172 83750
rect 2196 83748 2252 83750
rect 1956 82714 2012 82716
rect 2036 82714 2092 82716
rect 2116 82714 2172 82716
rect 2196 82714 2252 82716
rect 1956 82662 1982 82714
rect 1982 82662 2012 82714
rect 2036 82662 2046 82714
rect 2046 82662 2092 82714
rect 2116 82662 2162 82714
rect 2162 82662 2172 82714
rect 2196 82662 2226 82714
rect 2226 82662 2252 82714
rect 1956 82660 2012 82662
rect 2036 82660 2092 82662
rect 2116 82660 2172 82662
rect 2196 82660 2252 82662
rect 1956 81626 2012 81628
rect 2036 81626 2092 81628
rect 2116 81626 2172 81628
rect 2196 81626 2252 81628
rect 1956 81574 1982 81626
rect 1982 81574 2012 81626
rect 2036 81574 2046 81626
rect 2046 81574 2092 81626
rect 2116 81574 2162 81626
rect 2162 81574 2172 81626
rect 2196 81574 2226 81626
rect 2226 81574 2252 81626
rect 1956 81572 2012 81574
rect 2036 81572 2092 81574
rect 2116 81572 2172 81574
rect 2196 81572 2252 81574
rect 1956 80538 2012 80540
rect 2036 80538 2092 80540
rect 2116 80538 2172 80540
rect 2196 80538 2252 80540
rect 1956 80486 1982 80538
rect 1982 80486 2012 80538
rect 2036 80486 2046 80538
rect 2046 80486 2092 80538
rect 2116 80486 2162 80538
rect 2162 80486 2172 80538
rect 2196 80486 2226 80538
rect 2226 80486 2252 80538
rect 1956 80484 2012 80486
rect 2036 80484 2092 80486
rect 2116 80484 2172 80486
rect 2196 80484 2252 80486
rect 1956 79450 2012 79452
rect 2036 79450 2092 79452
rect 2116 79450 2172 79452
rect 2196 79450 2252 79452
rect 1956 79398 1982 79450
rect 1982 79398 2012 79450
rect 2036 79398 2046 79450
rect 2046 79398 2092 79450
rect 2116 79398 2162 79450
rect 2162 79398 2172 79450
rect 2196 79398 2226 79450
rect 2226 79398 2252 79450
rect 1956 79396 2012 79398
rect 2036 79396 2092 79398
rect 2116 79396 2172 79398
rect 2196 79396 2252 79398
rect 1956 78362 2012 78364
rect 2036 78362 2092 78364
rect 2116 78362 2172 78364
rect 2196 78362 2252 78364
rect 1956 78310 1982 78362
rect 1982 78310 2012 78362
rect 2036 78310 2046 78362
rect 2046 78310 2092 78362
rect 2116 78310 2162 78362
rect 2162 78310 2172 78362
rect 2196 78310 2226 78362
rect 2226 78310 2252 78362
rect 1956 78308 2012 78310
rect 2036 78308 2092 78310
rect 2116 78308 2172 78310
rect 2196 78308 2252 78310
rect 1956 77274 2012 77276
rect 2036 77274 2092 77276
rect 2116 77274 2172 77276
rect 2196 77274 2252 77276
rect 1956 77222 1982 77274
rect 1982 77222 2012 77274
rect 2036 77222 2046 77274
rect 2046 77222 2092 77274
rect 2116 77222 2162 77274
rect 2162 77222 2172 77274
rect 2196 77222 2226 77274
rect 2226 77222 2252 77274
rect 1956 77220 2012 77222
rect 2036 77220 2092 77222
rect 2116 77220 2172 77222
rect 2196 77220 2252 77222
rect 1956 76186 2012 76188
rect 2036 76186 2092 76188
rect 2116 76186 2172 76188
rect 2196 76186 2252 76188
rect 1956 76134 1982 76186
rect 1982 76134 2012 76186
rect 2036 76134 2046 76186
rect 2046 76134 2092 76186
rect 2116 76134 2162 76186
rect 2162 76134 2172 76186
rect 2196 76134 2226 76186
rect 2226 76134 2252 76186
rect 1956 76132 2012 76134
rect 2036 76132 2092 76134
rect 2116 76132 2172 76134
rect 2196 76132 2252 76134
rect 1956 75098 2012 75100
rect 2036 75098 2092 75100
rect 2116 75098 2172 75100
rect 2196 75098 2252 75100
rect 1956 75046 1982 75098
rect 1982 75046 2012 75098
rect 2036 75046 2046 75098
rect 2046 75046 2092 75098
rect 2116 75046 2162 75098
rect 2162 75046 2172 75098
rect 2196 75046 2226 75098
rect 2226 75046 2252 75098
rect 1956 75044 2012 75046
rect 2036 75044 2092 75046
rect 2116 75044 2172 75046
rect 2196 75044 2252 75046
rect 1956 74010 2012 74012
rect 2036 74010 2092 74012
rect 2116 74010 2172 74012
rect 2196 74010 2252 74012
rect 1956 73958 1982 74010
rect 1982 73958 2012 74010
rect 2036 73958 2046 74010
rect 2046 73958 2092 74010
rect 2116 73958 2162 74010
rect 2162 73958 2172 74010
rect 2196 73958 2226 74010
rect 2226 73958 2252 74010
rect 1956 73956 2012 73958
rect 2036 73956 2092 73958
rect 2116 73956 2172 73958
rect 2196 73956 2252 73958
rect 1956 72922 2012 72924
rect 2036 72922 2092 72924
rect 2116 72922 2172 72924
rect 2196 72922 2252 72924
rect 1956 72870 1982 72922
rect 1982 72870 2012 72922
rect 2036 72870 2046 72922
rect 2046 72870 2092 72922
rect 2116 72870 2162 72922
rect 2162 72870 2172 72922
rect 2196 72870 2226 72922
rect 2226 72870 2252 72922
rect 1956 72868 2012 72870
rect 2036 72868 2092 72870
rect 2116 72868 2172 72870
rect 2196 72868 2252 72870
rect 1956 71834 2012 71836
rect 2036 71834 2092 71836
rect 2116 71834 2172 71836
rect 2196 71834 2252 71836
rect 1956 71782 1982 71834
rect 1982 71782 2012 71834
rect 2036 71782 2046 71834
rect 2046 71782 2092 71834
rect 2116 71782 2162 71834
rect 2162 71782 2172 71834
rect 2196 71782 2226 71834
rect 2226 71782 2252 71834
rect 1956 71780 2012 71782
rect 2036 71780 2092 71782
rect 2116 71780 2172 71782
rect 2196 71780 2252 71782
rect 1956 70746 2012 70748
rect 2036 70746 2092 70748
rect 2116 70746 2172 70748
rect 2196 70746 2252 70748
rect 1956 70694 1982 70746
rect 1982 70694 2012 70746
rect 2036 70694 2046 70746
rect 2046 70694 2092 70746
rect 2116 70694 2162 70746
rect 2162 70694 2172 70746
rect 2196 70694 2226 70746
rect 2226 70694 2252 70746
rect 1956 70692 2012 70694
rect 2036 70692 2092 70694
rect 2116 70692 2172 70694
rect 2196 70692 2252 70694
rect 1956 69658 2012 69660
rect 2036 69658 2092 69660
rect 2116 69658 2172 69660
rect 2196 69658 2252 69660
rect 1956 69606 1982 69658
rect 1982 69606 2012 69658
rect 2036 69606 2046 69658
rect 2046 69606 2092 69658
rect 2116 69606 2162 69658
rect 2162 69606 2172 69658
rect 2196 69606 2226 69658
rect 2226 69606 2252 69658
rect 1956 69604 2012 69606
rect 2036 69604 2092 69606
rect 2116 69604 2172 69606
rect 2196 69604 2252 69606
rect 1956 68570 2012 68572
rect 2036 68570 2092 68572
rect 2116 68570 2172 68572
rect 2196 68570 2252 68572
rect 1956 68518 1982 68570
rect 1982 68518 2012 68570
rect 2036 68518 2046 68570
rect 2046 68518 2092 68570
rect 2116 68518 2162 68570
rect 2162 68518 2172 68570
rect 2196 68518 2226 68570
rect 2226 68518 2252 68570
rect 1956 68516 2012 68518
rect 2036 68516 2092 68518
rect 2116 68516 2172 68518
rect 2196 68516 2252 68518
rect 1956 67482 2012 67484
rect 2036 67482 2092 67484
rect 2116 67482 2172 67484
rect 2196 67482 2252 67484
rect 1956 67430 1982 67482
rect 1982 67430 2012 67482
rect 2036 67430 2046 67482
rect 2046 67430 2092 67482
rect 2116 67430 2162 67482
rect 2162 67430 2172 67482
rect 2196 67430 2226 67482
rect 2226 67430 2252 67482
rect 1956 67428 2012 67430
rect 2036 67428 2092 67430
rect 2116 67428 2172 67430
rect 2196 67428 2252 67430
rect 1956 66394 2012 66396
rect 2036 66394 2092 66396
rect 2116 66394 2172 66396
rect 2196 66394 2252 66396
rect 1956 66342 1982 66394
rect 1982 66342 2012 66394
rect 2036 66342 2046 66394
rect 2046 66342 2092 66394
rect 2116 66342 2162 66394
rect 2162 66342 2172 66394
rect 2196 66342 2226 66394
rect 2226 66342 2252 66394
rect 1956 66340 2012 66342
rect 2036 66340 2092 66342
rect 2116 66340 2172 66342
rect 2196 66340 2252 66342
rect 1956 65306 2012 65308
rect 2036 65306 2092 65308
rect 2116 65306 2172 65308
rect 2196 65306 2252 65308
rect 1956 65254 1982 65306
rect 1982 65254 2012 65306
rect 2036 65254 2046 65306
rect 2046 65254 2092 65306
rect 2116 65254 2162 65306
rect 2162 65254 2172 65306
rect 2196 65254 2226 65306
rect 2226 65254 2252 65306
rect 1956 65252 2012 65254
rect 2036 65252 2092 65254
rect 2116 65252 2172 65254
rect 2196 65252 2252 65254
rect 1956 64218 2012 64220
rect 2036 64218 2092 64220
rect 2116 64218 2172 64220
rect 2196 64218 2252 64220
rect 1956 64166 1982 64218
rect 1982 64166 2012 64218
rect 2036 64166 2046 64218
rect 2046 64166 2092 64218
rect 2116 64166 2162 64218
rect 2162 64166 2172 64218
rect 2196 64166 2226 64218
rect 2226 64166 2252 64218
rect 1956 64164 2012 64166
rect 2036 64164 2092 64166
rect 2116 64164 2172 64166
rect 2196 64164 2252 64166
rect 1956 63130 2012 63132
rect 2036 63130 2092 63132
rect 2116 63130 2172 63132
rect 2196 63130 2252 63132
rect 1956 63078 1982 63130
rect 1982 63078 2012 63130
rect 2036 63078 2046 63130
rect 2046 63078 2092 63130
rect 2116 63078 2162 63130
rect 2162 63078 2172 63130
rect 2196 63078 2226 63130
rect 2226 63078 2252 63130
rect 1956 63076 2012 63078
rect 2036 63076 2092 63078
rect 2116 63076 2172 63078
rect 2196 63076 2252 63078
rect 1956 62042 2012 62044
rect 2036 62042 2092 62044
rect 2116 62042 2172 62044
rect 2196 62042 2252 62044
rect 1956 61990 1982 62042
rect 1982 61990 2012 62042
rect 2036 61990 2046 62042
rect 2046 61990 2092 62042
rect 2116 61990 2162 62042
rect 2162 61990 2172 62042
rect 2196 61990 2226 62042
rect 2226 61990 2252 62042
rect 1956 61988 2012 61990
rect 2036 61988 2092 61990
rect 2116 61988 2172 61990
rect 2196 61988 2252 61990
rect 1956 60954 2012 60956
rect 2036 60954 2092 60956
rect 2116 60954 2172 60956
rect 2196 60954 2252 60956
rect 1956 60902 1982 60954
rect 1982 60902 2012 60954
rect 2036 60902 2046 60954
rect 2046 60902 2092 60954
rect 2116 60902 2162 60954
rect 2162 60902 2172 60954
rect 2196 60902 2226 60954
rect 2226 60902 2252 60954
rect 1956 60900 2012 60902
rect 2036 60900 2092 60902
rect 2116 60900 2172 60902
rect 2196 60900 2252 60902
rect 1956 59866 2012 59868
rect 2036 59866 2092 59868
rect 2116 59866 2172 59868
rect 2196 59866 2252 59868
rect 1956 59814 1982 59866
rect 1982 59814 2012 59866
rect 2036 59814 2046 59866
rect 2046 59814 2092 59866
rect 2116 59814 2162 59866
rect 2162 59814 2172 59866
rect 2196 59814 2226 59866
rect 2226 59814 2252 59866
rect 1956 59812 2012 59814
rect 2036 59812 2092 59814
rect 2116 59812 2172 59814
rect 2196 59812 2252 59814
rect 1956 58778 2012 58780
rect 2036 58778 2092 58780
rect 2116 58778 2172 58780
rect 2196 58778 2252 58780
rect 1956 58726 1982 58778
rect 1982 58726 2012 58778
rect 2036 58726 2046 58778
rect 2046 58726 2092 58778
rect 2116 58726 2162 58778
rect 2162 58726 2172 58778
rect 2196 58726 2226 58778
rect 2226 58726 2252 58778
rect 1956 58724 2012 58726
rect 2036 58724 2092 58726
rect 2116 58724 2172 58726
rect 2196 58724 2252 58726
rect 1956 57690 2012 57692
rect 2036 57690 2092 57692
rect 2116 57690 2172 57692
rect 2196 57690 2252 57692
rect 1956 57638 1982 57690
rect 1982 57638 2012 57690
rect 2036 57638 2046 57690
rect 2046 57638 2092 57690
rect 2116 57638 2162 57690
rect 2162 57638 2172 57690
rect 2196 57638 2226 57690
rect 2226 57638 2252 57690
rect 1956 57636 2012 57638
rect 2036 57636 2092 57638
rect 2116 57636 2172 57638
rect 2196 57636 2252 57638
rect 1956 56602 2012 56604
rect 2036 56602 2092 56604
rect 2116 56602 2172 56604
rect 2196 56602 2252 56604
rect 1956 56550 1982 56602
rect 1982 56550 2012 56602
rect 2036 56550 2046 56602
rect 2046 56550 2092 56602
rect 2116 56550 2162 56602
rect 2162 56550 2172 56602
rect 2196 56550 2226 56602
rect 2226 56550 2252 56602
rect 1956 56548 2012 56550
rect 2036 56548 2092 56550
rect 2116 56548 2172 56550
rect 2196 56548 2252 56550
rect 1956 55514 2012 55516
rect 2036 55514 2092 55516
rect 2116 55514 2172 55516
rect 2196 55514 2252 55516
rect 1956 55462 1982 55514
rect 1982 55462 2012 55514
rect 2036 55462 2046 55514
rect 2046 55462 2092 55514
rect 2116 55462 2162 55514
rect 2162 55462 2172 55514
rect 2196 55462 2226 55514
rect 2226 55462 2252 55514
rect 1956 55460 2012 55462
rect 2036 55460 2092 55462
rect 2116 55460 2172 55462
rect 2196 55460 2252 55462
rect 1956 54426 2012 54428
rect 2036 54426 2092 54428
rect 2116 54426 2172 54428
rect 2196 54426 2252 54428
rect 1956 54374 1982 54426
rect 1982 54374 2012 54426
rect 2036 54374 2046 54426
rect 2046 54374 2092 54426
rect 2116 54374 2162 54426
rect 2162 54374 2172 54426
rect 2196 54374 2226 54426
rect 2226 54374 2252 54426
rect 1956 54372 2012 54374
rect 2036 54372 2092 54374
rect 2116 54372 2172 54374
rect 2196 54372 2252 54374
rect 1956 53338 2012 53340
rect 2036 53338 2092 53340
rect 2116 53338 2172 53340
rect 2196 53338 2252 53340
rect 1956 53286 1982 53338
rect 1982 53286 2012 53338
rect 2036 53286 2046 53338
rect 2046 53286 2092 53338
rect 2116 53286 2162 53338
rect 2162 53286 2172 53338
rect 2196 53286 2226 53338
rect 2226 53286 2252 53338
rect 1956 53284 2012 53286
rect 2036 53284 2092 53286
rect 2116 53284 2172 53286
rect 2196 53284 2252 53286
rect 1956 52250 2012 52252
rect 2036 52250 2092 52252
rect 2116 52250 2172 52252
rect 2196 52250 2252 52252
rect 1956 52198 1982 52250
rect 1982 52198 2012 52250
rect 2036 52198 2046 52250
rect 2046 52198 2092 52250
rect 2116 52198 2162 52250
rect 2162 52198 2172 52250
rect 2196 52198 2226 52250
rect 2226 52198 2252 52250
rect 1956 52196 2012 52198
rect 2036 52196 2092 52198
rect 2116 52196 2172 52198
rect 2196 52196 2252 52198
rect 1956 51162 2012 51164
rect 2036 51162 2092 51164
rect 2116 51162 2172 51164
rect 2196 51162 2252 51164
rect 1956 51110 1982 51162
rect 1982 51110 2012 51162
rect 2036 51110 2046 51162
rect 2046 51110 2092 51162
rect 2116 51110 2162 51162
rect 2162 51110 2172 51162
rect 2196 51110 2226 51162
rect 2226 51110 2252 51162
rect 1956 51108 2012 51110
rect 2036 51108 2092 51110
rect 2116 51108 2172 51110
rect 2196 51108 2252 51110
rect 1956 50074 2012 50076
rect 2036 50074 2092 50076
rect 2116 50074 2172 50076
rect 2196 50074 2252 50076
rect 1956 50022 1982 50074
rect 1982 50022 2012 50074
rect 2036 50022 2046 50074
rect 2046 50022 2092 50074
rect 2116 50022 2162 50074
rect 2162 50022 2172 50074
rect 2196 50022 2226 50074
rect 2226 50022 2252 50074
rect 1956 50020 2012 50022
rect 2036 50020 2092 50022
rect 2116 50020 2172 50022
rect 2196 50020 2252 50022
rect 1956 48986 2012 48988
rect 2036 48986 2092 48988
rect 2116 48986 2172 48988
rect 2196 48986 2252 48988
rect 1956 48934 1982 48986
rect 1982 48934 2012 48986
rect 2036 48934 2046 48986
rect 2046 48934 2092 48986
rect 2116 48934 2162 48986
rect 2162 48934 2172 48986
rect 2196 48934 2226 48986
rect 2226 48934 2252 48986
rect 1956 48932 2012 48934
rect 2036 48932 2092 48934
rect 2116 48932 2172 48934
rect 2196 48932 2252 48934
rect 1956 47898 2012 47900
rect 2036 47898 2092 47900
rect 2116 47898 2172 47900
rect 2196 47898 2252 47900
rect 1956 47846 1982 47898
rect 1982 47846 2012 47898
rect 2036 47846 2046 47898
rect 2046 47846 2092 47898
rect 2116 47846 2162 47898
rect 2162 47846 2172 47898
rect 2196 47846 2226 47898
rect 2226 47846 2252 47898
rect 1956 47844 2012 47846
rect 2036 47844 2092 47846
rect 2116 47844 2172 47846
rect 2196 47844 2252 47846
rect 1956 46810 2012 46812
rect 2036 46810 2092 46812
rect 2116 46810 2172 46812
rect 2196 46810 2252 46812
rect 1956 46758 1982 46810
rect 1982 46758 2012 46810
rect 2036 46758 2046 46810
rect 2046 46758 2092 46810
rect 2116 46758 2162 46810
rect 2162 46758 2172 46810
rect 2196 46758 2226 46810
rect 2226 46758 2252 46810
rect 1956 46756 2012 46758
rect 2036 46756 2092 46758
rect 2116 46756 2172 46758
rect 2196 46756 2252 46758
rect 1956 45722 2012 45724
rect 2036 45722 2092 45724
rect 2116 45722 2172 45724
rect 2196 45722 2252 45724
rect 1956 45670 1982 45722
rect 1982 45670 2012 45722
rect 2036 45670 2046 45722
rect 2046 45670 2092 45722
rect 2116 45670 2162 45722
rect 2162 45670 2172 45722
rect 2196 45670 2226 45722
rect 2226 45670 2252 45722
rect 1956 45668 2012 45670
rect 2036 45668 2092 45670
rect 2116 45668 2172 45670
rect 2196 45668 2252 45670
rect 1956 44634 2012 44636
rect 2036 44634 2092 44636
rect 2116 44634 2172 44636
rect 2196 44634 2252 44636
rect 1956 44582 1982 44634
rect 1982 44582 2012 44634
rect 2036 44582 2046 44634
rect 2046 44582 2092 44634
rect 2116 44582 2162 44634
rect 2162 44582 2172 44634
rect 2196 44582 2226 44634
rect 2226 44582 2252 44634
rect 1956 44580 2012 44582
rect 2036 44580 2092 44582
rect 2116 44580 2172 44582
rect 2196 44580 2252 44582
rect 1956 43546 2012 43548
rect 2036 43546 2092 43548
rect 2116 43546 2172 43548
rect 2196 43546 2252 43548
rect 1956 43494 1982 43546
rect 1982 43494 2012 43546
rect 2036 43494 2046 43546
rect 2046 43494 2092 43546
rect 2116 43494 2162 43546
rect 2162 43494 2172 43546
rect 2196 43494 2226 43546
rect 2226 43494 2252 43546
rect 1956 43492 2012 43494
rect 2036 43492 2092 43494
rect 2116 43492 2172 43494
rect 2196 43492 2252 43494
rect 1956 42458 2012 42460
rect 2036 42458 2092 42460
rect 2116 42458 2172 42460
rect 2196 42458 2252 42460
rect 1956 42406 1982 42458
rect 1982 42406 2012 42458
rect 2036 42406 2046 42458
rect 2046 42406 2092 42458
rect 2116 42406 2162 42458
rect 2162 42406 2172 42458
rect 2196 42406 2226 42458
rect 2226 42406 2252 42458
rect 1956 42404 2012 42406
rect 2036 42404 2092 42406
rect 2116 42404 2172 42406
rect 2196 42404 2252 42406
rect 1956 41370 2012 41372
rect 2036 41370 2092 41372
rect 2116 41370 2172 41372
rect 2196 41370 2252 41372
rect 1956 41318 1982 41370
rect 1982 41318 2012 41370
rect 2036 41318 2046 41370
rect 2046 41318 2092 41370
rect 2116 41318 2162 41370
rect 2162 41318 2172 41370
rect 2196 41318 2226 41370
rect 2226 41318 2252 41370
rect 1956 41316 2012 41318
rect 2036 41316 2092 41318
rect 2116 41316 2172 41318
rect 2196 41316 2252 41318
rect 1956 40282 2012 40284
rect 2036 40282 2092 40284
rect 2116 40282 2172 40284
rect 2196 40282 2252 40284
rect 1956 40230 1982 40282
rect 1982 40230 2012 40282
rect 2036 40230 2046 40282
rect 2046 40230 2092 40282
rect 2116 40230 2162 40282
rect 2162 40230 2172 40282
rect 2196 40230 2226 40282
rect 2226 40230 2252 40282
rect 1956 40228 2012 40230
rect 2036 40228 2092 40230
rect 2116 40228 2172 40230
rect 2196 40228 2252 40230
rect 1956 39194 2012 39196
rect 2036 39194 2092 39196
rect 2116 39194 2172 39196
rect 2196 39194 2252 39196
rect 1956 39142 1982 39194
rect 1982 39142 2012 39194
rect 2036 39142 2046 39194
rect 2046 39142 2092 39194
rect 2116 39142 2162 39194
rect 2162 39142 2172 39194
rect 2196 39142 2226 39194
rect 2226 39142 2252 39194
rect 1956 39140 2012 39142
rect 2036 39140 2092 39142
rect 2116 39140 2172 39142
rect 2196 39140 2252 39142
rect 1956 38106 2012 38108
rect 2036 38106 2092 38108
rect 2116 38106 2172 38108
rect 2196 38106 2252 38108
rect 1956 38054 1982 38106
rect 1982 38054 2012 38106
rect 2036 38054 2046 38106
rect 2046 38054 2092 38106
rect 2116 38054 2162 38106
rect 2162 38054 2172 38106
rect 2196 38054 2226 38106
rect 2226 38054 2252 38106
rect 1956 38052 2012 38054
rect 2036 38052 2092 38054
rect 2116 38052 2172 38054
rect 2196 38052 2252 38054
rect 1956 37018 2012 37020
rect 2036 37018 2092 37020
rect 2116 37018 2172 37020
rect 2196 37018 2252 37020
rect 1956 36966 1982 37018
rect 1982 36966 2012 37018
rect 2036 36966 2046 37018
rect 2046 36966 2092 37018
rect 2116 36966 2162 37018
rect 2162 36966 2172 37018
rect 2196 36966 2226 37018
rect 2226 36966 2252 37018
rect 1956 36964 2012 36966
rect 2036 36964 2092 36966
rect 2116 36964 2172 36966
rect 2196 36964 2252 36966
rect 1956 35930 2012 35932
rect 2036 35930 2092 35932
rect 2116 35930 2172 35932
rect 2196 35930 2252 35932
rect 1956 35878 1982 35930
rect 1982 35878 2012 35930
rect 2036 35878 2046 35930
rect 2046 35878 2092 35930
rect 2116 35878 2162 35930
rect 2162 35878 2172 35930
rect 2196 35878 2226 35930
rect 2226 35878 2252 35930
rect 1956 35876 2012 35878
rect 2036 35876 2092 35878
rect 2116 35876 2172 35878
rect 2196 35876 2252 35878
rect 1956 34842 2012 34844
rect 2036 34842 2092 34844
rect 2116 34842 2172 34844
rect 2196 34842 2252 34844
rect 1956 34790 1982 34842
rect 1982 34790 2012 34842
rect 2036 34790 2046 34842
rect 2046 34790 2092 34842
rect 2116 34790 2162 34842
rect 2162 34790 2172 34842
rect 2196 34790 2226 34842
rect 2226 34790 2252 34842
rect 1956 34788 2012 34790
rect 2036 34788 2092 34790
rect 2116 34788 2172 34790
rect 2196 34788 2252 34790
rect 1956 33754 2012 33756
rect 2036 33754 2092 33756
rect 2116 33754 2172 33756
rect 2196 33754 2252 33756
rect 1956 33702 1982 33754
rect 1982 33702 2012 33754
rect 2036 33702 2046 33754
rect 2046 33702 2092 33754
rect 2116 33702 2162 33754
rect 2162 33702 2172 33754
rect 2196 33702 2226 33754
rect 2226 33702 2252 33754
rect 1956 33700 2012 33702
rect 2036 33700 2092 33702
rect 2116 33700 2172 33702
rect 2196 33700 2252 33702
rect 1956 32666 2012 32668
rect 2036 32666 2092 32668
rect 2116 32666 2172 32668
rect 2196 32666 2252 32668
rect 1956 32614 1982 32666
rect 1982 32614 2012 32666
rect 2036 32614 2046 32666
rect 2046 32614 2092 32666
rect 2116 32614 2162 32666
rect 2162 32614 2172 32666
rect 2196 32614 2226 32666
rect 2226 32614 2252 32666
rect 1956 32612 2012 32614
rect 2036 32612 2092 32614
rect 2116 32612 2172 32614
rect 2196 32612 2252 32614
rect 1956 31578 2012 31580
rect 2036 31578 2092 31580
rect 2116 31578 2172 31580
rect 2196 31578 2252 31580
rect 1956 31526 1982 31578
rect 1982 31526 2012 31578
rect 2036 31526 2046 31578
rect 2046 31526 2092 31578
rect 2116 31526 2162 31578
rect 2162 31526 2172 31578
rect 2196 31526 2226 31578
rect 2226 31526 2252 31578
rect 1956 31524 2012 31526
rect 2036 31524 2092 31526
rect 2116 31524 2172 31526
rect 2196 31524 2252 31526
rect 1956 30490 2012 30492
rect 2036 30490 2092 30492
rect 2116 30490 2172 30492
rect 2196 30490 2252 30492
rect 1956 30438 1982 30490
rect 1982 30438 2012 30490
rect 2036 30438 2046 30490
rect 2046 30438 2092 30490
rect 2116 30438 2162 30490
rect 2162 30438 2172 30490
rect 2196 30438 2226 30490
rect 2226 30438 2252 30490
rect 1956 30436 2012 30438
rect 2036 30436 2092 30438
rect 2116 30436 2172 30438
rect 2196 30436 2252 30438
rect 1956 29402 2012 29404
rect 2036 29402 2092 29404
rect 2116 29402 2172 29404
rect 2196 29402 2252 29404
rect 1956 29350 1982 29402
rect 1982 29350 2012 29402
rect 2036 29350 2046 29402
rect 2046 29350 2092 29402
rect 2116 29350 2162 29402
rect 2162 29350 2172 29402
rect 2196 29350 2226 29402
rect 2226 29350 2252 29402
rect 1956 29348 2012 29350
rect 2036 29348 2092 29350
rect 2116 29348 2172 29350
rect 2196 29348 2252 29350
rect 1956 28314 2012 28316
rect 2036 28314 2092 28316
rect 2116 28314 2172 28316
rect 2196 28314 2252 28316
rect 1956 28262 1982 28314
rect 1982 28262 2012 28314
rect 2036 28262 2046 28314
rect 2046 28262 2092 28314
rect 2116 28262 2162 28314
rect 2162 28262 2172 28314
rect 2196 28262 2226 28314
rect 2226 28262 2252 28314
rect 1956 28260 2012 28262
rect 2036 28260 2092 28262
rect 2116 28260 2172 28262
rect 2196 28260 2252 28262
rect 1956 27226 2012 27228
rect 2036 27226 2092 27228
rect 2116 27226 2172 27228
rect 2196 27226 2252 27228
rect 1956 27174 1982 27226
rect 1982 27174 2012 27226
rect 2036 27174 2046 27226
rect 2046 27174 2092 27226
rect 2116 27174 2162 27226
rect 2162 27174 2172 27226
rect 2196 27174 2226 27226
rect 2226 27174 2252 27226
rect 1956 27172 2012 27174
rect 2036 27172 2092 27174
rect 2116 27172 2172 27174
rect 2196 27172 2252 27174
rect 1956 26138 2012 26140
rect 2036 26138 2092 26140
rect 2116 26138 2172 26140
rect 2196 26138 2252 26140
rect 1956 26086 1982 26138
rect 1982 26086 2012 26138
rect 2036 26086 2046 26138
rect 2046 26086 2092 26138
rect 2116 26086 2162 26138
rect 2162 26086 2172 26138
rect 2196 26086 2226 26138
rect 2226 26086 2252 26138
rect 1956 26084 2012 26086
rect 2036 26084 2092 26086
rect 2116 26084 2172 26086
rect 2196 26084 2252 26086
rect 1956 25050 2012 25052
rect 2036 25050 2092 25052
rect 2116 25050 2172 25052
rect 2196 25050 2252 25052
rect 1956 24998 1982 25050
rect 1982 24998 2012 25050
rect 2036 24998 2046 25050
rect 2046 24998 2092 25050
rect 2116 24998 2162 25050
rect 2162 24998 2172 25050
rect 2196 24998 2226 25050
rect 2226 24998 2252 25050
rect 1956 24996 2012 24998
rect 2036 24996 2092 24998
rect 2116 24996 2172 24998
rect 2196 24996 2252 24998
rect 1956 23962 2012 23964
rect 2036 23962 2092 23964
rect 2116 23962 2172 23964
rect 2196 23962 2252 23964
rect 1956 23910 1982 23962
rect 1982 23910 2012 23962
rect 2036 23910 2046 23962
rect 2046 23910 2092 23962
rect 2116 23910 2162 23962
rect 2162 23910 2172 23962
rect 2196 23910 2226 23962
rect 2226 23910 2252 23962
rect 1956 23908 2012 23910
rect 2036 23908 2092 23910
rect 2116 23908 2172 23910
rect 2196 23908 2252 23910
rect 1956 22874 2012 22876
rect 2036 22874 2092 22876
rect 2116 22874 2172 22876
rect 2196 22874 2252 22876
rect 1956 22822 1982 22874
rect 1982 22822 2012 22874
rect 2036 22822 2046 22874
rect 2046 22822 2092 22874
rect 2116 22822 2162 22874
rect 2162 22822 2172 22874
rect 2196 22822 2226 22874
rect 2226 22822 2252 22874
rect 1956 22820 2012 22822
rect 2036 22820 2092 22822
rect 2116 22820 2172 22822
rect 2196 22820 2252 22822
rect 1956 21786 2012 21788
rect 2036 21786 2092 21788
rect 2116 21786 2172 21788
rect 2196 21786 2252 21788
rect 1956 21734 1982 21786
rect 1982 21734 2012 21786
rect 2036 21734 2046 21786
rect 2046 21734 2092 21786
rect 2116 21734 2162 21786
rect 2162 21734 2172 21786
rect 2196 21734 2226 21786
rect 2226 21734 2252 21786
rect 1956 21732 2012 21734
rect 2036 21732 2092 21734
rect 2116 21732 2172 21734
rect 2196 21732 2252 21734
rect 1956 20698 2012 20700
rect 2036 20698 2092 20700
rect 2116 20698 2172 20700
rect 2196 20698 2252 20700
rect 1956 20646 1982 20698
rect 1982 20646 2012 20698
rect 2036 20646 2046 20698
rect 2046 20646 2092 20698
rect 2116 20646 2162 20698
rect 2162 20646 2172 20698
rect 2196 20646 2226 20698
rect 2226 20646 2252 20698
rect 1956 20644 2012 20646
rect 2036 20644 2092 20646
rect 2116 20644 2172 20646
rect 2196 20644 2252 20646
rect 1956 19610 2012 19612
rect 2036 19610 2092 19612
rect 2116 19610 2172 19612
rect 2196 19610 2252 19612
rect 1956 19558 1982 19610
rect 1982 19558 2012 19610
rect 2036 19558 2046 19610
rect 2046 19558 2092 19610
rect 2116 19558 2162 19610
rect 2162 19558 2172 19610
rect 2196 19558 2226 19610
rect 2226 19558 2252 19610
rect 1956 19556 2012 19558
rect 2036 19556 2092 19558
rect 2116 19556 2172 19558
rect 2196 19556 2252 19558
rect 1956 18522 2012 18524
rect 2036 18522 2092 18524
rect 2116 18522 2172 18524
rect 2196 18522 2252 18524
rect 1956 18470 1982 18522
rect 1982 18470 2012 18522
rect 2036 18470 2046 18522
rect 2046 18470 2092 18522
rect 2116 18470 2162 18522
rect 2162 18470 2172 18522
rect 2196 18470 2226 18522
rect 2226 18470 2252 18522
rect 1956 18468 2012 18470
rect 2036 18468 2092 18470
rect 2116 18468 2172 18470
rect 2196 18468 2252 18470
rect 1956 17434 2012 17436
rect 2036 17434 2092 17436
rect 2116 17434 2172 17436
rect 2196 17434 2252 17436
rect 1956 17382 1982 17434
rect 1982 17382 2012 17434
rect 2036 17382 2046 17434
rect 2046 17382 2092 17434
rect 2116 17382 2162 17434
rect 2162 17382 2172 17434
rect 2196 17382 2226 17434
rect 2226 17382 2252 17434
rect 1956 17380 2012 17382
rect 2036 17380 2092 17382
rect 2116 17380 2172 17382
rect 2196 17380 2252 17382
rect 1956 16346 2012 16348
rect 2036 16346 2092 16348
rect 2116 16346 2172 16348
rect 2196 16346 2252 16348
rect 1956 16294 1982 16346
rect 1982 16294 2012 16346
rect 2036 16294 2046 16346
rect 2046 16294 2092 16346
rect 2116 16294 2162 16346
rect 2162 16294 2172 16346
rect 2196 16294 2226 16346
rect 2226 16294 2252 16346
rect 1956 16292 2012 16294
rect 2036 16292 2092 16294
rect 2116 16292 2172 16294
rect 2196 16292 2252 16294
rect 1956 15258 2012 15260
rect 2036 15258 2092 15260
rect 2116 15258 2172 15260
rect 2196 15258 2252 15260
rect 1956 15206 1982 15258
rect 1982 15206 2012 15258
rect 2036 15206 2046 15258
rect 2046 15206 2092 15258
rect 2116 15206 2162 15258
rect 2162 15206 2172 15258
rect 2196 15206 2226 15258
rect 2226 15206 2252 15258
rect 1956 15204 2012 15206
rect 2036 15204 2092 15206
rect 2116 15204 2172 15206
rect 2196 15204 2252 15206
rect 1956 14170 2012 14172
rect 2036 14170 2092 14172
rect 2116 14170 2172 14172
rect 2196 14170 2252 14172
rect 1956 14118 1982 14170
rect 1982 14118 2012 14170
rect 2036 14118 2046 14170
rect 2046 14118 2092 14170
rect 2116 14118 2162 14170
rect 2162 14118 2172 14170
rect 2196 14118 2226 14170
rect 2226 14118 2252 14170
rect 1956 14116 2012 14118
rect 2036 14116 2092 14118
rect 2116 14116 2172 14118
rect 2196 14116 2252 14118
rect 1956 13082 2012 13084
rect 2036 13082 2092 13084
rect 2116 13082 2172 13084
rect 2196 13082 2252 13084
rect 1956 13030 1982 13082
rect 1982 13030 2012 13082
rect 2036 13030 2046 13082
rect 2046 13030 2092 13082
rect 2116 13030 2162 13082
rect 2162 13030 2172 13082
rect 2196 13030 2226 13082
rect 2226 13030 2252 13082
rect 1956 13028 2012 13030
rect 2036 13028 2092 13030
rect 2116 13028 2172 13030
rect 2196 13028 2252 13030
rect 1956 11994 2012 11996
rect 2036 11994 2092 11996
rect 2116 11994 2172 11996
rect 2196 11994 2252 11996
rect 1956 11942 1982 11994
rect 1982 11942 2012 11994
rect 2036 11942 2046 11994
rect 2046 11942 2092 11994
rect 2116 11942 2162 11994
rect 2162 11942 2172 11994
rect 2196 11942 2226 11994
rect 2226 11942 2252 11994
rect 1956 11940 2012 11942
rect 2036 11940 2092 11942
rect 2116 11940 2172 11942
rect 2196 11940 2252 11942
rect 1956 10906 2012 10908
rect 2036 10906 2092 10908
rect 2116 10906 2172 10908
rect 2196 10906 2252 10908
rect 1956 10854 1982 10906
rect 1982 10854 2012 10906
rect 2036 10854 2046 10906
rect 2046 10854 2092 10906
rect 2116 10854 2162 10906
rect 2162 10854 2172 10906
rect 2196 10854 2226 10906
rect 2226 10854 2252 10906
rect 1956 10852 2012 10854
rect 2036 10852 2092 10854
rect 2116 10852 2172 10854
rect 2196 10852 2252 10854
rect 1956 9818 2012 9820
rect 2036 9818 2092 9820
rect 2116 9818 2172 9820
rect 2196 9818 2252 9820
rect 1956 9766 1982 9818
rect 1982 9766 2012 9818
rect 2036 9766 2046 9818
rect 2046 9766 2092 9818
rect 2116 9766 2162 9818
rect 2162 9766 2172 9818
rect 2196 9766 2226 9818
rect 2226 9766 2252 9818
rect 1956 9764 2012 9766
rect 2036 9764 2092 9766
rect 2116 9764 2172 9766
rect 2196 9764 2252 9766
rect 1956 8730 2012 8732
rect 2036 8730 2092 8732
rect 2116 8730 2172 8732
rect 2196 8730 2252 8732
rect 1956 8678 1982 8730
rect 1982 8678 2012 8730
rect 2036 8678 2046 8730
rect 2046 8678 2092 8730
rect 2116 8678 2162 8730
rect 2162 8678 2172 8730
rect 2196 8678 2226 8730
rect 2226 8678 2252 8730
rect 1956 8676 2012 8678
rect 2036 8676 2092 8678
rect 2116 8676 2172 8678
rect 2196 8676 2252 8678
rect 1956 7642 2012 7644
rect 2036 7642 2092 7644
rect 2116 7642 2172 7644
rect 2196 7642 2252 7644
rect 1956 7590 1982 7642
rect 1982 7590 2012 7642
rect 2036 7590 2046 7642
rect 2046 7590 2092 7642
rect 2116 7590 2162 7642
rect 2162 7590 2172 7642
rect 2196 7590 2226 7642
rect 2226 7590 2252 7642
rect 1956 7588 2012 7590
rect 2036 7588 2092 7590
rect 2116 7588 2172 7590
rect 2196 7588 2252 7590
rect 1956 6554 2012 6556
rect 2036 6554 2092 6556
rect 2116 6554 2172 6556
rect 2196 6554 2252 6556
rect 1956 6502 1982 6554
rect 1982 6502 2012 6554
rect 2036 6502 2046 6554
rect 2046 6502 2092 6554
rect 2116 6502 2162 6554
rect 2162 6502 2172 6554
rect 2196 6502 2226 6554
rect 2226 6502 2252 6554
rect 1956 6500 2012 6502
rect 2036 6500 2092 6502
rect 2116 6500 2172 6502
rect 2196 6500 2252 6502
rect 1956 5466 2012 5468
rect 2036 5466 2092 5468
rect 2116 5466 2172 5468
rect 2196 5466 2252 5468
rect 1956 5414 1982 5466
rect 1982 5414 2012 5466
rect 2036 5414 2046 5466
rect 2046 5414 2092 5466
rect 2116 5414 2162 5466
rect 2162 5414 2172 5466
rect 2196 5414 2226 5466
rect 2226 5414 2252 5466
rect 1956 5412 2012 5414
rect 2036 5412 2092 5414
rect 2116 5412 2172 5414
rect 2196 5412 2252 5414
rect 1956 4378 2012 4380
rect 2036 4378 2092 4380
rect 2116 4378 2172 4380
rect 2196 4378 2252 4380
rect 1956 4326 1982 4378
rect 1982 4326 2012 4378
rect 2036 4326 2046 4378
rect 2046 4326 2092 4378
rect 2116 4326 2162 4378
rect 2162 4326 2172 4378
rect 2196 4326 2226 4378
rect 2226 4326 2252 4378
rect 1956 4324 2012 4326
rect 2036 4324 2092 4326
rect 2116 4324 2172 4326
rect 2196 4324 2252 4326
rect 1956 3290 2012 3292
rect 2036 3290 2092 3292
rect 2116 3290 2172 3292
rect 2196 3290 2252 3292
rect 1956 3238 1982 3290
rect 1982 3238 2012 3290
rect 2036 3238 2046 3290
rect 2046 3238 2092 3290
rect 2116 3238 2162 3290
rect 2162 3238 2172 3290
rect 2196 3238 2226 3290
rect 2226 3238 2252 3290
rect 1956 3236 2012 3238
rect 2036 3236 2092 3238
rect 2116 3236 2172 3238
rect 2196 3236 2252 3238
rect 3956 96314 4012 96316
rect 4036 96314 4092 96316
rect 4116 96314 4172 96316
rect 4196 96314 4252 96316
rect 3956 96262 3982 96314
rect 3982 96262 4012 96314
rect 4036 96262 4046 96314
rect 4046 96262 4092 96314
rect 4116 96262 4162 96314
rect 4162 96262 4172 96314
rect 4196 96262 4226 96314
rect 4226 96262 4252 96314
rect 3956 96260 4012 96262
rect 4036 96260 4092 96262
rect 4116 96260 4172 96262
rect 4196 96260 4252 96262
rect 3514 3304 3570 3360
rect 3956 95226 4012 95228
rect 4036 95226 4092 95228
rect 4116 95226 4172 95228
rect 4196 95226 4252 95228
rect 3956 95174 3982 95226
rect 3982 95174 4012 95226
rect 4036 95174 4046 95226
rect 4046 95174 4092 95226
rect 4116 95174 4162 95226
rect 4162 95174 4172 95226
rect 4196 95174 4226 95226
rect 4226 95174 4252 95226
rect 3956 95172 4012 95174
rect 4036 95172 4092 95174
rect 4116 95172 4172 95174
rect 4196 95172 4252 95174
rect 3956 94138 4012 94140
rect 4036 94138 4092 94140
rect 4116 94138 4172 94140
rect 4196 94138 4252 94140
rect 3956 94086 3982 94138
rect 3982 94086 4012 94138
rect 4036 94086 4046 94138
rect 4046 94086 4092 94138
rect 4116 94086 4162 94138
rect 4162 94086 4172 94138
rect 4196 94086 4226 94138
rect 4226 94086 4252 94138
rect 3956 94084 4012 94086
rect 4036 94084 4092 94086
rect 4116 94084 4172 94086
rect 4196 94084 4252 94086
rect 3956 93050 4012 93052
rect 4036 93050 4092 93052
rect 4116 93050 4172 93052
rect 4196 93050 4252 93052
rect 3956 92998 3982 93050
rect 3982 92998 4012 93050
rect 4036 92998 4046 93050
rect 4046 92998 4092 93050
rect 4116 92998 4162 93050
rect 4162 92998 4172 93050
rect 4196 92998 4226 93050
rect 4226 92998 4252 93050
rect 3956 92996 4012 92998
rect 4036 92996 4092 92998
rect 4116 92996 4172 92998
rect 4196 92996 4252 92998
rect 3956 91962 4012 91964
rect 4036 91962 4092 91964
rect 4116 91962 4172 91964
rect 4196 91962 4252 91964
rect 3956 91910 3982 91962
rect 3982 91910 4012 91962
rect 4036 91910 4046 91962
rect 4046 91910 4092 91962
rect 4116 91910 4162 91962
rect 4162 91910 4172 91962
rect 4196 91910 4226 91962
rect 4226 91910 4252 91962
rect 3956 91908 4012 91910
rect 4036 91908 4092 91910
rect 4116 91908 4172 91910
rect 4196 91908 4252 91910
rect 3956 90874 4012 90876
rect 4036 90874 4092 90876
rect 4116 90874 4172 90876
rect 4196 90874 4252 90876
rect 3956 90822 3982 90874
rect 3982 90822 4012 90874
rect 4036 90822 4046 90874
rect 4046 90822 4092 90874
rect 4116 90822 4162 90874
rect 4162 90822 4172 90874
rect 4196 90822 4226 90874
rect 4226 90822 4252 90874
rect 3956 90820 4012 90822
rect 4036 90820 4092 90822
rect 4116 90820 4172 90822
rect 4196 90820 4252 90822
rect 4434 93472 4490 93528
rect 3956 89786 4012 89788
rect 4036 89786 4092 89788
rect 4116 89786 4172 89788
rect 4196 89786 4252 89788
rect 3956 89734 3982 89786
rect 3982 89734 4012 89786
rect 4036 89734 4046 89786
rect 4046 89734 4092 89786
rect 4116 89734 4162 89786
rect 4162 89734 4172 89786
rect 4196 89734 4226 89786
rect 4226 89734 4252 89786
rect 3956 89732 4012 89734
rect 4036 89732 4092 89734
rect 4116 89732 4172 89734
rect 4196 89732 4252 89734
rect 3956 88698 4012 88700
rect 4036 88698 4092 88700
rect 4116 88698 4172 88700
rect 4196 88698 4252 88700
rect 3956 88646 3982 88698
rect 3982 88646 4012 88698
rect 4036 88646 4046 88698
rect 4046 88646 4092 88698
rect 4116 88646 4162 88698
rect 4162 88646 4172 88698
rect 4196 88646 4226 88698
rect 4226 88646 4252 88698
rect 3956 88644 4012 88646
rect 4036 88644 4092 88646
rect 4116 88644 4172 88646
rect 4196 88644 4252 88646
rect 3956 87610 4012 87612
rect 4036 87610 4092 87612
rect 4116 87610 4172 87612
rect 4196 87610 4252 87612
rect 3956 87558 3982 87610
rect 3982 87558 4012 87610
rect 4036 87558 4046 87610
rect 4046 87558 4092 87610
rect 4116 87558 4162 87610
rect 4162 87558 4172 87610
rect 4196 87558 4226 87610
rect 4226 87558 4252 87610
rect 3956 87556 4012 87558
rect 4036 87556 4092 87558
rect 4116 87556 4172 87558
rect 4196 87556 4252 87558
rect 3956 86522 4012 86524
rect 4036 86522 4092 86524
rect 4116 86522 4172 86524
rect 4196 86522 4252 86524
rect 3956 86470 3982 86522
rect 3982 86470 4012 86522
rect 4036 86470 4046 86522
rect 4046 86470 4092 86522
rect 4116 86470 4162 86522
rect 4162 86470 4172 86522
rect 4196 86470 4226 86522
rect 4226 86470 4252 86522
rect 3956 86468 4012 86470
rect 4036 86468 4092 86470
rect 4116 86468 4172 86470
rect 4196 86468 4252 86470
rect 3956 85434 4012 85436
rect 4036 85434 4092 85436
rect 4116 85434 4172 85436
rect 4196 85434 4252 85436
rect 3956 85382 3982 85434
rect 3982 85382 4012 85434
rect 4036 85382 4046 85434
rect 4046 85382 4092 85434
rect 4116 85382 4162 85434
rect 4162 85382 4172 85434
rect 4196 85382 4226 85434
rect 4226 85382 4252 85434
rect 3956 85380 4012 85382
rect 4036 85380 4092 85382
rect 4116 85380 4172 85382
rect 4196 85380 4252 85382
rect 3956 84346 4012 84348
rect 4036 84346 4092 84348
rect 4116 84346 4172 84348
rect 4196 84346 4252 84348
rect 3956 84294 3982 84346
rect 3982 84294 4012 84346
rect 4036 84294 4046 84346
rect 4046 84294 4092 84346
rect 4116 84294 4162 84346
rect 4162 84294 4172 84346
rect 4196 84294 4226 84346
rect 4226 84294 4252 84346
rect 3956 84292 4012 84294
rect 4036 84292 4092 84294
rect 4116 84292 4172 84294
rect 4196 84292 4252 84294
rect 3956 83258 4012 83260
rect 4036 83258 4092 83260
rect 4116 83258 4172 83260
rect 4196 83258 4252 83260
rect 3956 83206 3982 83258
rect 3982 83206 4012 83258
rect 4036 83206 4046 83258
rect 4046 83206 4092 83258
rect 4116 83206 4162 83258
rect 4162 83206 4172 83258
rect 4196 83206 4226 83258
rect 4226 83206 4252 83258
rect 3956 83204 4012 83206
rect 4036 83204 4092 83206
rect 4116 83204 4172 83206
rect 4196 83204 4252 83206
rect 3956 82170 4012 82172
rect 4036 82170 4092 82172
rect 4116 82170 4172 82172
rect 4196 82170 4252 82172
rect 3956 82118 3982 82170
rect 3982 82118 4012 82170
rect 4036 82118 4046 82170
rect 4046 82118 4092 82170
rect 4116 82118 4162 82170
rect 4162 82118 4172 82170
rect 4196 82118 4226 82170
rect 4226 82118 4252 82170
rect 3956 82116 4012 82118
rect 4036 82116 4092 82118
rect 4116 82116 4172 82118
rect 4196 82116 4252 82118
rect 3956 81082 4012 81084
rect 4036 81082 4092 81084
rect 4116 81082 4172 81084
rect 4196 81082 4252 81084
rect 3956 81030 3982 81082
rect 3982 81030 4012 81082
rect 4036 81030 4046 81082
rect 4046 81030 4092 81082
rect 4116 81030 4162 81082
rect 4162 81030 4172 81082
rect 4196 81030 4226 81082
rect 4226 81030 4252 81082
rect 3956 81028 4012 81030
rect 4036 81028 4092 81030
rect 4116 81028 4172 81030
rect 4196 81028 4252 81030
rect 3956 79994 4012 79996
rect 4036 79994 4092 79996
rect 4116 79994 4172 79996
rect 4196 79994 4252 79996
rect 3956 79942 3982 79994
rect 3982 79942 4012 79994
rect 4036 79942 4046 79994
rect 4046 79942 4092 79994
rect 4116 79942 4162 79994
rect 4162 79942 4172 79994
rect 4196 79942 4226 79994
rect 4226 79942 4252 79994
rect 3956 79940 4012 79942
rect 4036 79940 4092 79942
rect 4116 79940 4172 79942
rect 4196 79940 4252 79942
rect 3956 78906 4012 78908
rect 4036 78906 4092 78908
rect 4116 78906 4172 78908
rect 4196 78906 4252 78908
rect 3956 78854 3982 78906
rect 3982 78854 4012 78906
rect 4036 78854 4046 78906
rect 4046 78854 4092 78906
rect 4116 78854 4162 78906
rect 4162 78854 4172 78906
rect 4196 78854 4226 78906
rect 4226 78854 4252 78906
rect 3956 78852 4012 78854
rect 4036 78852 4092 78854
rect 4116 78852 4172 78854
rect 4196 78852 4252 78854
rect 3956 77818 4012 77820
rect 4036 77818 4092 77820
rect 4116 77818 4172 77820
rect 4196 77818 4252 77820
rect 3956 77766 3982 77818
rect 3982 77766 4012 77818
rect 4036 77766 4046 77818
rect 4046 77766 4092 77818
rect 4116 77766 4162 77818
rect 4162 77766 4172 77818
rect 4196 77766 4226 77818
rect 4226 77766 4252 77818
rect 3956 77764 4012 77766
rect 4036 77764 4092 77766
rect 4116 77764 4172 77766
rect 4196 77764 4252 77766
rect 3956 76730 4012 76732
rect 4036 76730 4092 76732
rect 4116 76730 4172 76732
rect 4196 76730 4252 76732
rect 3956 76678 3982 76730
rect 3982 76678 4012 76730
rect 4036 76678 4046 76730
rect 4046 76678 4092 76730
rect 4116 76678 4162 76730
rect 4162 76678 4172 76730
rect 4196 76678 4226 76730
rect 4226 76678 4252 76730
rect 3956 76676 4012 76678
rect 4036 76676 4092 76678
rect 4116 76676 4172 76678
rect 4196 76676 4252 76678
rect 3956 75642 4012 75644
rect 4036 75642 4092 75644
rect 4116 75642 4172 75644
rect 4196 75642 4252 75644
rect 3956 75590 3982 75642
rect 3982 75590 4012 75642
rect 4036 75590 4046 75642
rect 4046 75590 4092 75642
rect 4116 75590 4162 75642
rect 4162 75590 4172 75642
rect 4196 75590 4226 75642
rect 4226 75590 4252 75642
rect 3956 75588 4012 75590
rect 4036 75588 4092 75590
rect 4116 75588 4172 75590
rect 4196 75588 4252 75590
rect 3956 74554 4012 74556
rect 4036 74554 4092 74556
rect 4116 74554 4172 74556
rect 4196 74554 4252 74556
rect 3956 74502 3982 74554
rect 3982 74502 4012 74554
rect 4036 74502 4046 74554
rect 4046 74502 4092 74554
rect 4116 74502 4162 74554
rect 4162 74502 4172 74554
rect 4196 74502 4226 74554
rect 4226 74502 4252 74554
rect 3956 74500 4012 74502
rect 4036 74500 4092 74502
rect 4116 74500 4172 74502
rect 4196 74500 4252 74502
rect 3956 73466 4012 73468
rect 4036 73466 4092 73468
rect 4116 73466 4172 73468
rect 4196 73466 4252 73468
rect 3956 73414 3982 73466
rect 3982 73414 4012 73466
rect 4036 73414 4046 73466
rect 4046 73414 4092 73466
rect 4116 73414 4162 73466
rect 4162 73414 4172 73466
rect 4196 73414 4226 73466
rect 4226 73414 4252 73466
rect 3956 73412 4012 73414
rect 4036 73412 4092 73414
rect 4116 73412 4172 73414
rect 4196 73412 4252 73414
rect 3956 72378 4012 72380
rect 4036 72378 4092 72380
rect 4116 72378 4172 72380
rect 4196 72378 4252 72380
rect 3956 72326 3982 72378
rect 3982 72326 4012 72378
rect 4036 72326 4046 72378
rect 4046 72326 4092 72378
rect 4116 72326 4162 72378
rect 4162 72326 4172 72378
rect 4196 72326 4226 72378
rect 4226 72326 4252 72378
rect 3956 72324 4012 72326
rect 4036 72324 4092 72326
rect 4116 72324 4172 72326
rect 4196 72324 4252 72326
rect 3956 71290 4012 71292
rect 4036 71290 4092 71292
rect 4116 71290 4172 71292
rect 4196 71290 4252 71292
rect 3956 71238 3982 71290
rect 3982 71238 4012 71290
rect 4036 71238 4046 71290
rect 4046 71238 4092 71290
rect 4116 71238 4162 71290
rect 4162 71238 4172 71290
rect 4196 71238 4226 71290
rect 4226 71238 4252 71290
rect 3956 71236 4012 71238
rect 4036 71236 4092 71238
rect 4116 71236 4172 71238
rect 4196 71236 4252 71238
rect 3956 70202 4012 70204
rect 4036 70202 4092 70204
rect 4116 70202 4172 70204
rect 4196 70202 4252 70204
rect 3956 70150 3982 70202
rect 3982 70150 4012 70202
rect 4036 70150 4046 70202
rect 4046 70150 4092 70202
rect 4116 70150 4162 70202
rect 4162 70150 4172 70202
rect 4196 70150 4226 70202
rect 4226 70150 4252 70202
rect 3956 70148 4012 70150
rect 4036 70148 4092 70150
rect 4116 70148 4172 70150
rect 4196 70148 4252 70150
rect 3956 69114 4012 69116
rect 4036 69114 4092 69116
rect 4116 69114 4172 69116
rect 4196 69114 4252 69116
rect 3956 69062 3982 69114
rect 3982 69062 4012 69114
rect 4036 69062 4046 69114
rect 4046 69062 4092 69114
rect 4116 69062 4162 69114
rect 4162 69062 4172 69114
rect 4196 69062 4226 69114
rect 4226 69062 4252 69114
rect 3956 69060 4012 69062
rect 4036 69060 4092 69062
rect 4116 69060 4172 69062
rect 4196 69060 4252 69062
rect 3956 68026 4012 68028
rect 4036 68026 4092 68028
rect 4116 68026 4172 68028
rect 4196 68026 4252 68028
rect 3956 67974 3982 68026
rect 3982 67974 4012 68026
rect 4036 67974 4046 68026
rect 4046 67974 4092 68026
rect 4116 67974 4162 68026
rect 4162 67974 4172 68026
rect 4196 67974 4226 68026
rect 4226 67974 4252 68026
rect 3956 67972 4012 67974
rect 4036 67972 4092 67974
rect 4116 67972 4172 67974
rect 4196 67972 4252 67974
rect 3956 66938 4012 66940
rect 4036 66938 4092 66940
rect 4116 66938 4172 66940
rect 4196 66938 4252 66940
rect 3956 66886 3982 66938
rect 3982 66886 4012 66938
rect 4036 66886 4046 66938
rect 4046 66886 4092 66938
rect 4116 66886 4162 66938
rect 4162 66886 4172 66938
rect 4196 66886 4226 66938
rect 4226 66886 4252 66938
rect 3956 66884 4012 66886
rect 4036 66884 4092 66886
rect 4116 66884 4172 66886
rect 4196 66884 4252 66886
rect 3956 65850 4012 65852
rect 4036 65850 4092 65852
rect 4116 65850 4172 65852
rect 4196 65850 4252 65852
rect 3956 65798 3982 65850
rect 3982 65798 4012 65850
rect 4036 65798 4046 65850
rect 4046 65798 4092 65850
rect 4116 65798 4162 65850
rect 4162 65798 4172 65850
rect 4196 65798 4226 65850
rect 4226 65798 4252 65850
rect 3956 65796 4012 65798
rect 4036 65796 4092 65798
rect 4116 65796 4172 65798
rect 4196 65796 4252 65798
rect 3956 64762 4012 64764
rect 4036 64762 4092 64764
rect 4116 64762 4172 64764
rect 4196 64762 4252 64764
rect 3956 64710 3982 64762
rect 3982 64710 4012 64762
rect 4036 64710 4046 64762
rect 4046 64710 4092 64762
rect 4116 64710 4162 64762
rect 4162 64710 4172 64762
rect 4196 64710 4226 64762
rect 4226 64710 4252 64762
rect 3956 64708 4012 64710
rect 4036 64708 4092 64710
rect 4116 64708 4172 64710
rect 4196 64708 4252 64710
rect 3956 63674 4012 63676
rect 4036 63674 4092 63676
rect 4116 63674 4172 63676
rect 4196 63674 4252 63676
rect 3956 63622 3982 63674
rect 3982 63622 4012 63674
rect 4036 63622 4046 63674
rect 4046 63622 4092 63674
rect 4116 63622 4162 63674
rect 4162 63622 4172 63674
rect 4196 63622 4226 63674
rect 4226 63622 4252 63674
rect 3956 63620 4012 63622
rect 4036 63620 4092 63622
rect 4116 63620 4172 63622
rect 4196 63620 4252 63622
rect 3956 62586 4012 62588
rect 4036 62586 4092 62588
rect 4116 62586 4172 62588
rect 4196 62586 4252 62588
rect 3956 62534 3982 62586
rect 3982 62534 4012 62586
rect 4036 62534 4046 62586
rect 4046 62534 4092 62586
rect 4116 62534 4162 62586
rect 4162 62534 4172 62586
rect 4196 62534 4226 62586
rect 4226 62534 4252 62586
rect 3956 62532 4012 62534
rect 4036 62532 4092 62534
rect 4116 62532 4172 62534
rect 4196 62532 4252 62534
rect 3956 61498 4012 61500
rect 4036 61498 4092 61500
rect 4116 61498 4172 61500
rect 4196 61498 4252 61500
rect 3956 61446 3982 61498
rect 3982 61446 4012 61498
rect 4036 61446 4046 61498
rect 4046 61446 4092 61498
rect 4116 61446 4162 61498
rect 4162 61446 4172 61498
rect 4196 61446 4226 61498
rect 4226 61446 4252 61498
rect 3956 61444 4012 61446
rect 4036 61444 4092 61446
rect 4116 61444 4172 61446
rect 4196 61444 4252 61446
rect 3956 60410 4012 60412
rect 4036 60410 4092 60412
rect 4116 60410 4172 60412
rect 4196 60410 4252 60412
rect 3956 60358 3982 60410
rect 3982 60358 4012 60410
rect 4036 60358 4046 60410
rect 4046 60358 4092 60410
rect 4116 60358 4162 60410
rect 4162 60358 4172 60410
rect 4196 60358 4226 60410
rect 4226 60358 4252 60410
rect 3956 60356 4012 60358
rect 4036 60356 4092 60358
rect 4116 60356 4172 60358
rect 4196 60356 4252 60358
rect 3956 59322 4012 59324
rect 4036 59322 4092 59324
rect 4116 59322 4172 59324
rect 4196 59322 4252 59324
rect 3956 59270 3982 59322
rect 3982 59270 4012 59322
rect 4036 59270 4046 59322
rect 4046 59270 4092 59322
rect 4116 59270 4162 59322
rect 4162 59270 4172 59322
rect 4196 59270 4226 59322
rect 4226 59270 4252 59322
rect 3956 59268 4012 59270
rect 4036 59268 4092 59270
rect 4116 59268 4172 59270
rect 4196 59268 4252 59270
rect 3956 58234 4012 58236
rect 4036 58234 4092 58236
rect 4116 58234 4172 58236
rect 4196 58234 4252 58236
rect 3956 58182 3982 58234
rect 3982 58182 4012 58234
rect 4036 58182 4046 58234
rect 4046 58182 4092 58234
rect 4116 58182 4162 58234
rect 4162 58182 4172 58234
rect 4196 58182 4226 58234
rect 4226 58182 4252 58234
rect 3956 58180 4012 58182
rect 4036 58180 4092 58182
rect 4116 58180 4172 58182
rect 4196 58180 4252 58182
rect 3956 57146 4012 57148
rect 4036 57146 4092 57148
rect 4116 57146 4172 57148
rect 4196 57146 4252 57148
rect 3956 57094 3982 57146
rect 3982 57094 4012 57146
rect 4036 57094 4046 57146
rect 4046 57094 4092 57146
rect 4116 57094 4162 57146
rect 4162 57094 4172 57146
rect 4196 57094 4226 57146
rect 4226 57094 4252 57146
rect 3956 57092 4012 57094
rect 4036 57092 4092 57094
rect 4116 57092 4172 57094
rect 4196 57092 4252 57094
rect 3956 56058 4012 56060
rect 4036 56058 4092 56060
rect 4116 56058 4172 56060
rect 4196 56058 4252 56060
rect 3956 56006 3982 56058
rect 3982 56006 4012 56058
rect 4036 56006 4046 56058
rect 4046 56006 4092 56058
rect 4116 56006 4162 56058
rect 4162 56006 4172 56058
rect 4196 56006 4226 56058
rect 4226 56006 4252 56058
rect 3956 56004 4012 56006
rect 4036 56004 4092 56006
rect 4116 56004 4172 56006
rect 4196 56004 4252 56006
rect 3956 54970 4012 54972
rect 4036 54970 4092 54972
rect 4116 54970 4172 54972
rect 4196 54970 4252 54972
rect 3956 54918 3982 54970
rect 3982 54918 4012 54970
rect 4036 54918 4046 54970
rect 4046 54918 4092 54970
rect 4116 54918 4162 54970
rect 4162 54918 4172 54970
rect 4196 54918 4226 54970
rect 4226 54918 4252 54970
rect 3956 54916 4012 54918
rect 4036 54916 4092 54918
rect 4116 54916 4172 54918
rect 4196 54916 4252 54918
rect 3956 53882 4012 53884
rect 4036 53882 4092 53884
rect 4116 53882 4172 53884
rect 4196 53882 4252 53884
rect 3956 53830 3982 53882
rect 3982 53830 4012 53882
rect 4036 53830 4046 53882
rect 4046 53830 4092 53882
rect 4116 53830 4162 53882
rect 4162 53830 4172 53882
rect 4196 53830 4226 53882
rect 4226 53830 4252 53882
rect 3956 53828 4012 53830
rect 4036 53828 4092 53830
rect 4116 53828 4172 53830
rect 4196 53828 4252 53830
rect 3956 52794 4012 52796
rect 4036 52794 4092 52796
rect 4116 52794 4172 52796
rect 4196 52794 4252 52796
rect 3956 52742 3982 52794
rect 3982 52742 4012 52794
rect 4036 52742 4046 52794
rect 4046 52742 4092 52794
rect 4116 52742 4162 52794
rect 4162 52742 4172 52794
rect 4196 52742 4226 52794
rect 4226 52742 4252 52794
rect 3956 52740 4012 52742
rect 4036 52740 4092 52742
rect 4116 52740 4172 52742
rect 4196 52740 4252 52742
rect 3956 51706 4012 51708
rect 4036 51706 4092 51708
rect 4116 51706 4172 51708
rect 4196 51706 4252 51708
rect 3956 51654 3982 51706
rect 3982 51654 4012 51706
rect 4036 51654 4046 51706
rect 4046 51654 4092 51706
rect 4116 51654 4162 51706
rect 4162 51654 4172 51706
rect 4196 51654 4226 51706
rect 4226 51654 4252 51706
rect 3956 51652 4012 51654
rect 4036 51652 4092 51654
rect 4116 51652 4172 51654
rect 4196 51652 4252 51654
rect 3956 50618 4012 50620
rect 4036 50618 4092 50620
rect 4116 50618 4172 50620
rect 4196 50618 4252 50620
rect 3956 50566 3982 50618
rect 3982 50566 4012 50618
rect 4036 50566 4046 50618
rect 4046 50566 4092 50618
rect 4116 50566 4162 50618
rect 4162 50566 4172 50618
rect 4196 50566 4226 50618
rect 4226 50566 4252 50618
rect 3956 50564 4012 50566
rect 4036 50564 4092 50566
rect 4116 50564 4172 50566
rect 4196 50564 4252 50566
rect 3956 49530 4012 49532
rect 4036 49530 4092 49532
rect 4116 49530 4172 49532
rect 4196 49530 4252 49532
rect 3956 49478 3982 49530
rect 3982 49478 4012 49530
rect 4036 49478 4046 49530
rect 4046 49478 4092 49530
rect 4116 49478 4162 49530
rect 4162 49478 4172 49530
rect 4196 49478 4226 49530
rect 4226 49478 4252 49530
rect 3956 49476 4012 49478
rect 4036 49476 4092 49478
rect 4116 49476 4172 49478
rect 4196 49476 4252 49478
rect 3956 48442 4012 48444
rect 4036 48442 4092 48444
rect 4116 48442 4172 48444
rect 4196 48442 4252 48444
rect 3956 48390 3982 48442
rect 3982 48390 4012 48442
rect 4036 48390 4046 48442
rect 4046 48390 4092 48442
rect 4116 48390 4162 48442
rect 4162 48390 4172 48442
rect 4196 48390 4226 48442
rect 4226 48390 4252 48442
rect 3956 48388 4012 48390
rect 4036 48388 4092 48390
rect 4116 48388 4172 48390
rect 4196 48388 4252 48390
rect 3956 47354 4012 47356
rect 4036 47354 4092 47356
rect 4116 47354 4172 47356
rect 4196 47354 4252 47356
rect 3956 47302 3982 47354
rect 3982 47302 4012 47354
rect 4036 47302 4046 47354
rect 4046 47302 4092 47354
rect 4116 47302 4162 47354
rect 4162 47302 4172 47354
rect 4196 47302 4226 47354
rect 4226 47302 4252 47354
rect 3956 47300 4012 47302
rect 4036 47300 4092 47302
rect 4116 47300 4172 47302
rect 4196 47300 4252 47302
rect 3956 46266 4012 46268
rect 4036 46266 4092 46268
rect 4116 46266 4172 46268
rect 4196 46266 4252 46268
rect 3956 46214 3982 46266
rect 3982 46214 4012 46266
rect 4036 46214 4046 46266
rect 4046 46214 4092 46266
rect 4116 46214 4162 46266
rect 4162 46214 4172 46266
rect 4196 46214 4226 46266
rect 4226 46214 4252 46266
rect 3956 46212 4012 46214
rect 4036 46212 4092 46214
rect 4116 46212 4172 46214
rect 4196 46212 4252 46214
rect 3956 45178 4012 45180
rect 4036 45178 4092 45180
rect 4116 45178 4172 45180
rect 4196 45178 4252 45180
rect 3956 45126 3982 45178
rect 3982 45126 4012 45178
rect 4036 45126 4046 45178
rect 4046 45126 4092 45178
rect 4116 45126 4162 45178
rect 4162 45126 4172 45178
rect 4196 45126 4226 45178
rect 4226 45126 4252 45178
rect 3956 45124 4012 45126
rect 4036 45124 4092 45126
rect 4116 45124 4172 45126
rect 4196 45124 4252 45126
rect 3956 44090 4012 44092
rect 4036 44090 4092 44092
rect 4116 44090 4172 44092
rect 4196 44090 4252 44092
rect 3956 44038 3982 44090
rect 3982 44038 4012 44090
rect 4036 44038 4046 44090
rect 4046 44038 4092 44090
rect 4116 44038 4162 44090
rect 4162 44038 4172 44090
rect 4196 44038 4226 44090
rect 4226 44038 4252 44090
rect 3956 44036 4012 44038
rect 4036 44036 4092 44038
rect 4116 44036 4172 44038
rect 4196 44036 4252 44038
rect 3956 43002 4012 43004
rect 4036 43002 4092 43004
rect 4116 43002 4172 43004
rect 4196 43002 4252 43004
rect 3956 42950 3982 43002
rect 3982 42950 4012 43002
rect 4036 42950 4046 43002
rect 4046 42950 4092 43002
rect 4116 42950 4162 43002
rect 4162 42950 4172 43002
rect 4196 42950 4226 43002
rect 4226 42950 4252 43002
rect 3956 42948 4012 42950
rect 4036 42948 4092 42950
rect 4116 42948 4172 42950
rect 4196 42948 4252 42950
rect 3956 41914 4012 41916
rect 4036 41914 4092 41916
rect 4116 41914 4172 41916
rect 4196 41914 4252 41916
rect 3956 41862 3982 41914
rect 3982 41862 4012 41914
rect 4036 41862 4046 41914
rect 4046 41862 4092 41914
rect 4116 41862 4162 41914
rect 4162 41862 4172 41914
rect 4196 41862 4226 41914
rect 4226 41862 4252 41914
rect 3956 41860 4012 41862
rect 4036 41860 4092 41862
rect 4116 41860 4172 41862
rect 4196 41860 4252 41862
rect 3956 40826 4012 40828
rect 4036 40826 4092 40828
rect 4116 40826 4172 40828
rect 4196 40826 4252 40828
rect 3956 40774 3982 40826
rect 3982 40774 4012 40826
rect 4036 40774 4046 40826
rect 4046 40774 4092 40826
rect 4116 40774 4162 40826
rect 4162 40774 4172 40826
rect 4196 40774 4226 40826
rect 4226 40774 4252 40826
rect 3956 40772 4012 40774
rect 4036 40772 4092 40774
rect 4116 40772 4172 40774
rect 4196 40772 4252 40774
rect 3956 39738 4012 39740
rect 4036 39738 4092 39740
rect 4116 39738 4172 39740
rect 4196 39738 4252 39740
rect 3956 39686 3982 39738
rect 3982 39686 4012 39738
rect 4036 39686 4046 39738
rect 4046 39686 4092 39738
rect 4116 39686 4162 39738
rect 4162 39686 4172 39738
rect 4196 39686 4226 39738
rect 4226 39686 4252 39738
rect 3956 39684 4012 39686
rect 4036 39684 4092 39686
rect 4116 39684 4172 39686
rect 4196 39684 4252 39686
rect 3956 38650 4012 38652
rect 4036 38650 4092 38652
rect 4116 38650 4172 38652
rect 4196 38650 4252 38652
rect 3956 38598 3982 38650
rect 3982 38598 4012 38650
rect 4036 38598 4046 38650
rect 4046 38598 4092 38650
rect 4116 38598 4162 38650
rect 4162 38598 4172 38650
rect 4196 38598 4226 38650
rect 4226 38598 4252 38650
rect 3956 38596 4012 38598
rect 4036 38596 4092 38598
rect 4116 38596 4172 38598
rect 4196 38596 4252 38598
rect 3956 37562 4012 37564
rect 4036 37562 4092 37564
rect 4116 37562 4172 37564
rect 4196 37562 4252 37564
rect 3956 37510 3982 37562
rect 3982 37510 4012 37562
rect 4036 37510 4046 37562
rect 4046 37510 4092 37562
rect 4116 37510 4162 37562
rect 4162 37510 4172 37562
rect 4196 37510 4226 37562
rect 4226 37510 4252 37562
rect 3956 37508 4012 37510
rect 4036 37508 4092 37510
rect 4116 37508 4172 37510
rect 4196 37508 4252 37510
rect 3956 36474 4012 36476
rect 4036 36474 4092 36476
rect 4116 36474 4172 36476
rect 4196 36474 4252 36476
rect 3956 36422 3982 36474
rect 3982 36422 4012 36474
rect 4036 36422 4046 36474
rect 4046 36422 4092 36474
rect 4116 36422 4162 36474
rect 4162 36422 4172 36474
rect 4196 36422 4226 36474
rect 4226 36422 4252 36474
rect 3956 36420 4012 36422
rect 4036 36420 4092 36422
rect 4116 36420 4172 36422
rect 4196 36420 4252 36422
rect 3956 35386 4012 35388
rect 4036 35386 4092 35388
rect 4116 35386 4172 35388
rect 4196 35386 4252 35388
rect 3956 35334 3982 35386
rect 3982 35334 4012 35386
rect 4036 35334 4046 35386
rect 4046 35334 4092 35386
rect 4116 35334 4162 35386
rect 4162 35334 4172 35386
rect 4196 35334 4226 35386
rect 4226 35334 4252 35386
rect 3956 35332 4012 35334
rect 4036 35332 4092 35334
rect 4116 35332 4172 35334
rect 4196 35332 4252 35334
rect 3956 34298 4012 34300
rect 4036 34298 4092 34300
rect 4116 34298 4172 34300
rect 4196 34298 4252 34300
rect 3956 34246 3982 34298
rect 3982 34246 4012 34298
rect 4036 34246 4046 34298
rect 4046 34246 4092 34298
rect 4116 34246 4162 34298
rect 4162 34246 4172 34298
rect 4196 34246 4226 34298
rect 4226 34246 4252 34298
rect 3956 34244 4012 34246
rect 4036 34244 4092 34246
rect 4116 34244 4172 34246
rect 4196 34244 4252 34246
rect 3956 33210 4012 33212
rect 4036 33210 4092 33212
rect 4116 33210 4172 33212
rect 4196 33210 4252 33212
rect 3956 33158 3982 33210
rect 3982 33158 4012 33210
rect 4036 33158 4046 33210
rect 4046 33158 4092 33210
rect 4116 33158 4162 33210
rect 4162 33158 4172 33210
rect 4196 33158 4226 33210
rect 4226 33158 4252 33210
rect 3956 33156 4012 33158
rect 4036 33156 4092 33158
rect 4116 33156 4172 33158
rect 4196 33156 4252 33158
rect 3956 32122 4012 32124
rect 4036 32122 4092 32124
rect 4116 32122 4172 32124
rect 4196 32122 4252 32124
rect 3956 32070 3982 32122
rect 3982 32070 4012 32122
rect 4036 32070 4046 32122
rect 4046 32070 4092 32122
rect 4116 32070 4162 32122
rect 4162 32070 4172 32122
rect 4196 32070 4226 32122
rect 4226 32070 4252 32122
rect 3956 32068 4012 32070
rect 4036 32068 4092 32070
rect 4116 32068 4172 32070
rect 4196 32068 4252 32070
rect 3956 31034 4012 31036
rect 4036 31034 4092 31036
rect 4116 31034 4172 31036
rect 4196 31034 4252 31036
rect 3956 30982 3982 31034
rect 3982 30982 4012 31034
rect 4036 30982 4046 31034
rect 4046 30982 4092 31034
rect 4116 30982 4162 31034
rect 4162 30982 4172 31034
rect 4196 30982 4226 31034
rect 4226 30982 4252 31034
rect 3956 30980 4012 30982
rect 4036 30980 4092 30982
rect 4116 30980 4172 30982
rect 4196 30980 4252 30982
rect 3956 29946 4012 29948
rect 4036 29946 4092 29948
rect 4116 29946 4172 29948
rect 4196 29946 4252 29948
rect 3956 29894 3982 29946
rect 3982 29894 4012 29946
rect 4036 29894 4046 29946
rect 4046 29894 4092 29946
rect 4116 29894 4162 29946
rect 4162 29894 4172 29946
rect 4196 29894 4226 29946
rect 4226 29894 4252 29946
rect 3956 29892 4012 29894
rect 4036 29892 4092 29894
rect 4116 29892 4172 29894
rect 4196 29892 4252 29894
rect 3956 28858 4012 28860
rect 4036 28858 4092 28860
rect 4116 28858 4172 28860
rect 4196 28858 4252 28860
rect 3956 28806 3982 28858
rect 3982 28806 4012 28858
rect 4036 28806 4046 28858
rect 4046 28806 4092 28858
rect 4116 28806 4162 28858
rect 4162 28806 4172 28858
rect 4196 28806 4226 28858
rect 4226 28806 4252 28858
rect 3956 28804 4012 28806
rect 4036 28804 4092 28806
rect 4116 28804 4172 28806
rect 4196 28804 4252 28806
rect 3956 27770 4012 27772
rect 4036 27770 4092 27772
rect 4116 27770 4172 27772
rect 4196 27770 4252 27772
rect 3956 27718 3982 27770
rect 3982 27718 4012 27770
rect 4036 27718 4046 27770
rect 4046 27718 4092 27770
rect 4116 27718 4162 27770
rect 4162 27718 4172 27770
rect 4196 27718 4226 27770
rect 4226 27718 4252 27770
rect 3956 27716 4012 27718
rect 4036 27716 4092 27718
rect 4116 27716 4172 27718
rect 4196 27716 4252 27718
rect 3956 26682 4012 26684
rect 4036 26682 4092 26684
rect 4116 26682 4172 26684
rect 4196 26682 4252 26684
rect 3956 26630 3982 26682
rect 3982 26630 4012 26682
rect 4036 26630 4046 26682
rect 4046 26630 4092 26682
rect 4116 26630 4162 26682
rect 4162 26630 4172 26682
rect 4196 26630 4226 26682
rect 4226 26630 4252 26682
rect 3956 26628 4012 26630
rect 4036 26628 4092 26630
rect 4116 26628 4172 26630
rect 4196 26628 4252 26630
rect 3956 25594 4012 25596
rect 4036 25594 4092 25596
rect 4116 25594 4172 25596
rect 4196 25594 4252 25596
rect 3956 25542 3982 25594
rect 3982 25542 4012 25594
rect 4036 25542 4046 25594
rect 4046 25542 4092 25594
rect 4116 25542 4162 25594
rect 4162 25542 4172 25594
rect 4196 25542 4226 25594
rect 4226 25542 4252 25594
rect 3956 25540 4012 25542
rect 4036 25540 4092 25542
rect 4116 25540 4172 25542
rect 4196 25540 4252 25542
rect 3956 24506 4012 24508
rect 4036 24506 4092 24508
rect 4116 24506 4172 24508
rect 4196 24506 4252 24508
rect 3956 24454 3982 24506
rect 3982 24454 4012 24506
rect 4036 24454 4046 24506
rect 4046 24454 4092 24506
rect 4116 24454 4162 24506
rect 4162 24454 4172 24506
rect 4196 24454 4226 24506
rect 4226 24454 4252 24506
rect 3956 24452 4012 24454
rect 4036 24452 4092 24454
rect 4116 24452 4172 24454
rect 4196 24452 4252 24454
rect 3956 23418 4012 23420
rect 4036 23418 4092 23420
rect 4116 23418 4172 23420
rect 4196 23418 4252 23420
rect 3956 23366 3982 23418
rect 3982 23366 4012 23418
rect 4036 23366 4046 23418
rect 4046 23366 4092 23418
rect 4116 23366 4162 23418
rect 4162 23366 4172 23418
rect 4196 23366 4226 23418
rect 4226 23366 4252 23418
rect 3956 23364 4012 23366
rect 4036 23364 4092 23366
rect 4116 23364 4172 23366
rect 4196 23364 4252 23366
rect 3956 22330 4012 22332
rect 4036 22330 4092 22332
rect 4116 22330 4172 22332
rect 4196 22330 4252 22332
rect 3956 22278 3982 22330
rect 3982 22278 4012 22330
rect 4036 22278 4046 22330
rect 4046 22278 4092 22330
rect 4116 22278 4162 22330
rect 4162 22278 4172 22330
rect 4196 22278 4226 22330
rect 4226 22278 4252 22330
rect 3956 22276 4012 22278
rect 4036 22276 4092 22278
rect 4116 22276 4172 22278
rect 4196 22276 4252 22278
rect 3956 21242 4012 21244
rect 4036 21242 4092 21244
rect 4116 21242 4172 21244
rect 4196 21242 4252 21244
rect 3956 21190 3982 21242
rect 3982 21190 4012 21242
rect 4036 21190 4046 21242
rect 4046 21190 4092 21242
rect 4116 21190 4162 21242
rect 4162 21190 4172 21242
rect 4196 21190 4226 21242
rect 4226 21190 4252 21242
rect 3956 21188 4012 21190
rect 4036 21188 4092 21190
rect 4116 21188 4172 21190
rect 4196 21188 4252 21190
rect 3956 20154 4012 20156
rect 4036 20154 4092 20156
rect 4116 20154 4172 20156
rect 4196 20154 4252 20156
rect 3956 20102 3982 20154
rect 3982 20102 4012 20154
rect 4036 20102 4046 20154
rect 4046 20102 4092 20154
rect 4116 20102 4162 20154
rect 4162 20102 4172 20154
rect 4196 20102 4226 20154
rect 4226 20102 4252 20154
rect 3956 20100 4012 20102
rect 4036 20100 4092 20102
rect 4116 20100 4172 20102
rect 4196 20100 4252 20102
rect 3956 19066 4012 19068
rect 4036 19066 4092 19068
rect 4116 19066 4172 19068
rect 4196 19066 4252 19068
rect 3956 19014 3982 19066
rect 3982 19014 4012 19066
rect 4036 19014 4046 19066
rect 4046 19014 4092 19066
rect 4116 19014 4162 19066
rect 4162 19014 4172 19066
rect 4196 19014 4226 19066
rect 4226 19014 4252 19066
rect 3956 19012 4012 19014
rect 4036 19012 4092 19014
rect 4116 19012 4172 19014
rect 4196 19012 4252 19014
rect 3956 17978 4012 17980
rect 4036 17978 4092 17980
rect 4116 17978 4172 17980
rect 4196 17978 4252 17980
rect 3956 17926 3982 17978
rect 3982 17926 4012 17978
rect 4036 17926 4046 17978
rect 4046 17926 4092 17978
rect 4116 17926 4162 17978
rect 4162 17926 4172 17978
rect 4196 17926 4226 17978
rect 4226 17926 4252 17978
rect 3956 17924 4012 17926
rect 4036 17924 4092 17926
rect 4116 17924 4172 17926
rect 4196 17924 4252 17926
rect 3956 16890 4012 16892
rect 4036 16890 4092 16892
rect 4116 16890 4172 16892
rect 4196 16890 4252 16892
rect 3956 16838 3982 16890
rect 3982 16838 4012 16890
rect 4036 16838 4046 16890
rect 4046 16838 4092 16890
rect 4116 16838 4162 16890
rect 4162 16838 4172 16890
rect 4196 16838 4226 16890
rect 4226 16838 4252 16890
rect 3956 16836 4012 16838
rect 4036 16836 4092 16838
rect 4116 16836 4172 16838
rect 4196 16836 4252 16838
rect 3956 15802 4012 15804
rect 4036 15802 4092 15804
rect 4116 15802 4172 15804
rect 4196 15802 4252 15804
rect 3956 15750 3982 15802
rect 3982 15750 4012 15802
rect 4036 15750 4046 15802
rect 4046 15750 4092 15802
rect 4116 15750 4162 15802
rect 4162 15750 4172 15802
rect 4196 15750 4226 15802
rect 4226 15750 4252 15802
rect 3956 15748 4012 15750
rect 4036 15748 4092 15750
rect 4116 15748 4172 15750
rect 4196 15748 4252 15750
rect 3956 14714 4012 14716
rect 4036 14714 4092 14716
rect 4116 14714 4172 14716
rect 4196 14714 4252 14716
rect 3956 14662 3982 14714
rect 3982 14662 4012 14714
rect 4036 14662 4046 14714
rect 4046 14662 4092 14714
rect 4116 14662 4162 14714
rect 4162 14662 4172 14714
rect 4196 14662 4226 14714
rect 4226 14662 4252 14714
rect 3956 14660 4012 14662
rect 4036 14660 4092 14662
rect 4116 14660 4172 14662
rect 4196 14660 4252 14662
rect 3956 13626 4012 13628
rect 4036 13626 4092 13628
rect 4116 13626 4172 13628
rect 4196 13626 4252 13628
rect 3956 13574 3982 13626
rect 3982 13574 4012 13626
rect 4036 13574 4046 13626
rect 4046 13574 4092 13626
rect 4116 13574 4162 13626
rect 4162 13574 4172 13626
rect 4196 13574 4226 13626
rect 4226 13574 4252 13626
rect 3956 13572 4012 13574
rect 4036 13572 4092 13574
rect 4116 13572 4172 13574
rect 4196 13572 4252 13574
rect 3956 12538 4012 12540
rect 4036 12538 4092 12540
rect 4116 12538 4172 12540
rect 4196 12538 4252 12540
rect 3956 12486 3982 12538
rect 3982 12486 4012 12538
rect 4036 12486 4046 12538
rect 4046 12486 4092 12538
rect 4116 12486 4162 12538
rect 4162 12486 4172 12538
rect 4196 12486 4226 12538
rect 4226 12486 4252 12538
rect 3956 12484 4012 12486
rect 4036 12484 4092 12486
rect 4116 12484 4172 12486
rect 4196 12484 4252 12486
rect 3956 11450 4012 11452
rect 4036 11450 4092 11452
rect 4116 11450 4172 11452
rect 4196 11450 4252 11452
rect 3956 11398 3982 11450
rect 3982 11398 4012 11450
rect 4036 11398 4046 11450
rect 4046 11398 4092 11450
rect 4116 11398 4162 11450
rect 4162 11398 4172 11450
rect 4196 11398 4226 11450
rect 4226 11398 4252 11450
rect 3956 11396 4012 11398
rect 4036 11396 4092 11398
rect 4116 11396 4172 11398
rect 4196 11396 4252 11398
rect 3956 10362 4012 10364
rect 4036 10362 4092 10364
rect 4116 10362 4172 10364
rect 4196 10362 4252 10364
rect 3956 10310 3982 10362
rect 3982 10310 4012 10362
rect 4036 10310 4046 10362
rect 4046 10310 4092 10362
rect 4116 10310 4162 10362
rect 4162 10310 4172 10362
rect 4196 10310 4226 10362
rect 4226 10310 4252 10362
rect 3956 10308 4012 10310
rect 4036 10308 4092 10310
rect 4116 10308 4172 10310
rect 4196 10308 4252 10310
rect 3956 9274 4012 9276
rect 4036 9274 4092 9276
rect 4116 9274 4172 9276
rect 4196 9274 4252 9276
rect 3956 9222 3982 9274
rect 3982 9222 4012 9274
rect 4036 9222 4046 9274
rect 4046 9222 4092 9274
rect 4116 9222 4162 9274
rect 4162 9222 4172 9274
rect 4196 9222 4226 9274
rect 4226 9222 4252 9274
rect 3956 9220 4012 9222
rect 4036 9220 4092 9222
rect 4116 9220 4172 9222
rect 4196 9220 4252 9222
rect 3956 8186 4012 8188
rect 4036 8186 4092 8188
rect 4116 8186 4172 8188
rect 4196 8186 4252 8188
rect 3956 8134 3982 8186
rect 3982 8134 4012 8186
rect 4036 8134 4046 8186
rect 4046 8134 4092 8186
rect 4116 8134 4162 8186
rect 4162 8134 4172 8186
rect 4196 8134 4226 8186
rect 4226 8134 4252 8186
rect 3956 8132 4012 8134
rect 4036 8132 4092 8134
rect 4116 8132 4172 8134
rect 4196 8132 4252 8134
rect 3956 7098 4012 7100
rect 4036 7098 4092 7100
rect 4116 7098 4172 7100
rect 4196 7098 4252 7100
rect 3956 7046 3982 7098
rect 3982 7046 4012 7098
rect 4036 7046 4046 7098
rect 4046 7046 4092 7098
rect 4116 7046 4162 7098
rect 4162 7046 4172 7098
rect 4196 7046 4226 7098
rect 4226 7046 4252 7098
rect 3956 7044 4012 7046
rect 4036 7044 4092 7046
rect 4116 7044 4172 7046
rect 4196 7044 4252 7046
rect 3956 6010 4012 6012
rect 4036 6010 4092 6012
rect 4116 6010 4172 6012
rect 4196 6010 4252 6012
rect 3956 5958 3982 6010
rect 3982 5958 4012 6010
rect 4036 5958 4046 6010
rect 4046 5958 4092 6010
rect 4116 5958 4162 6010
rect 4162 5958 4172 6010
rect 4196 5958 4226 6010
rect 4226 5958 4252 6010
rect 3956 5956 4012 5958
rect 4036 5956 4092 5958
rect 4116 5956 4172 5958
rect 4196 5956 4252 5958
rect 3956 4922 4012 4924
rect 4036 4922 4092 4924
rect 4116 4922 4172 4924
rect 4196 4922 4252 4924
rect 3956 4870 3982 4922
rect 3982 4870 4012 4922
rect 4036 4870 4046 4922
rect 4046 4870 4092 4922
rect 4116 4870 4162 4922
rect 4162 4870 4172 4922
rect 4196 4870 4226 4922
rect 4226 4870 4252 4922
rect 3956 4868 4012 4870
rect 4036 4868 4092 4870
rect 4116 4868 4172 4870
rect 4196 4868 4252 4870
rect 3606 2896 3662 2952
rect 1956 2202 2012 2204
rect 2036 2202 2092 2204
rect 2116 2202 2172 2204
rect 2196 2202 2252 2204
rect 1956 2150 1982 2202
rect 1982 2150 2012 2202
rect 2036 2150 2046 2202
rect 2046 2150 2092 2202
rect 2116 2150 2162 2202
rect 2162 2150 2172 2202
rect 2196 2150 2226 2202
rect 2226 2150 2252 2202
rect 1956 2148 2012 2150
rect 2036 2148 2092 2150
rect 2116 2148 2172 2150
rect 2196 2148 2252 2150
rect 3790 3032 3846 3088
rect 3956 3834 4012 3836
rect 4036 3834 4092 3836
rect 4116 3834 4172 3836
rect 4196 3834 4252 3836
rect 3956 3782 3982 3834
rect 3982 3782 4012 3834
rect 4036 3782 4046 3834
rect 4046 3782 4092 3834
rect 4116 3782 4162 3834
rect 4162 3782 4172 3834
rect 4196 3782 4226 3834
rect 4226 3782 4252 3834
rect 3956 3780 4012 3782
rect 4036 3780 4092 3782
rect 4116 3780 4172 3782
rect 4196 3780 4252 3782
rect 4434 10124 4490 10160
rect 4434 10104 4436 10124
rect 4436 10104 4488 10124
rect 4488 10104 4490 10124
rect 4342 3168 4398 3224
rect 3956 2746 4012 2748
rect 4036 2746 4092 2748
rect 4116 2746 4172 2748
rect 4196 2746 4252 2748
rect 3956 2694 3982 2746
rect 3982 2694 4012 2746
rect 4036 2694 4046 2746
rect 4046 2694 4092 2746
rect 4116 2694 4162 2746
rect 4162 2694 4172 2746
rect 4196 2694 4226 2746
rect 4226 2694 4252 2746
rect 3956 2692 4012 2694
rect 4036 2692 4092 2694
rect 4116 2692 4172 2694
rect 4196 2692 4252 2694
rect 4802 176180 4858 176216
rect 4802 176160 4804 176180
rect 4804 176160 4856 176180
rect 4856 176160 4858 176180
rect 4802 174548 4858 174584
rect 4802 174528 4804 174548
rect 4804 174528 4856 174548
rect 4856 174528 4858 174548
rect 4710 92384 4766 92440
rect 4710 91024 4766 91080
rect 4710 89256 4766 89312
rect 5262 176160 5318 176216
rect 5262 174528 5318 174584
rect 5446 121488 5502 121544
rect 5354 116612 5410 116648
rect 5354 116592 5356 116612
rect 5356 116592 5408 116612
rect 5408 116592 5410 116612
rect 5446 114980 5502 115016
rect 5446 114960 5448 114980
rect 5448 114960 5500 114980
rect 5500 114960 5502 114980
rect 5078 91024 5134 91080
rect 5170 89392 5226 89448
rect 4802 89020 4804 89040
rect 4804 89020 4856 89040
rect 4856 89020 4858 89040
rect 4802 88984 4858 89020
rect 4802 88848 4858 88904
rect 4710 86672 4766 86728
rect 4710 85176 4766 85232
rect 4802 83308 4804 83328
rect 4804 83308 4856 83328
rect 4856 83308 4858 83328
rect 4802 83272 4858 83308
rect 4802 82220 4804 82240
rect 4804 82220 4856 82240
rect 4856 82220 4858 82240
rect 4802 82184 4858 82220
rect 4802 80436 4858 80472
rect 4802 80416 4804 80436
rect 4804 80416 4856 80436
rect 4856 80416 4858 80436
rect 4710 22380 4712 22400
rect 4712 22380 4764 22400
rect 4764 22380 4766 22400
rect 4710 22344 4766 22380
rect 4618 3168 4674 3224
rect 4802 20868 4858 20904
rect 4802 20848 4804 20868
rect 4804 20848 4856 20868
rect 4856 20848 4858 20868
rect 5078 89120 5134 89176
rect 4986 87760 5042 87816
rect 5262 88712 5318 88768
rect 5170 86264 5226 86320
rect 5170 82184 5226 82240
rect 5262 80416 5318 80472
rect 4802 3884 4804 3904
rect 4804 3884 4856 3904
rect 4856 3884 4858 3904
rect 4802 3848 4858 3884
rect 4894 3032 4950 3088
rect 5354 2760 5410 2816
rect 5722 96872 5778 96928
rect 6182 96872 6238 96928
rect 5906 96736 5962 96792
rect 5814 96600 5870 96656
rect 5906 3304 5962 3360
rect 5722 3032 5778 3088
rect 5630 2896 5686 2952
rect 6366 96736 6422 96792
rect 21914 97180 21916 97200
rect 21916 97180 21968 97200
rect 21968 97180 21970 97200
rect 21914 97144 21970 97180
rect 22650 97144 22706 97200
rect 14646 97028 14702 97064
rect 14646 97008 14648 97028
rect 14648 97008 14700 97028
rect 14700 97008 14702 97028
rect 17130 97028 17186 97064
rect 17130 97008 17132 97028
rect 17132 97008 17184 97028
rect 17184 97008 17186 97028
rect 18050 97044 18052 97064
rect 18052 97044 18104 97064
rect 18104 97044 18106 97064
rect 18050 97008 18106 97044
rect 78954 97144 79010 97200
rect 24306 97008 24362 97064
rect 25410 97008 25466 97064
rect 30102 97008 30158 97064
rect 32034 97008 32090 97064
rect 33138 97008 33194 97064
rect 77390 97008 77446 97064
rect 78678 97008 78734 97064
rect 54850 96872 54906 96928
rect 60462 96872 60518 96928
rect 60646 96872 60702 96928
rect 16486 96484 16542 96520
rect 16486 96464 16488 96484
rect 16488 96464 16540 96484
rect 16540 96464 16542 96484
rect 15750 96348 15806 96384
rect 15750 96328 15752 96348
rect 15752 96328 15804 96348
rect 15804 96328 15806 96348
rect 9586 96212 9642 96248
rect 9586 96192 9588 96212
rect 9588 96192 9640 96212
rect 9640 96192 9642 96212
rect 6550 2896 6606 2952
rect 53746 96600 53802 96656
rect 22098 96192 22154 96248
rect 27986 96192 28042 96248
rect 29182 96192 29238 96248
rect 20994 96056 21050 96112
rect 26790 96056 26846 96112
rect 24582 95240 24638 95296
rect 12806 95104 12862 95160
rect 19338 95124 19394 95160
rect 19338 95104 19340 95124
rect 19340 95104 19392 95124
rect 19392 95104 19394 95124
rect 24766 95140 24768 95160
rect 24768 95140 24820 95160
rect 24820 95140 24822 95160
rect 24766 95104 24822 95140
rect 25962 95104 26018 95160
rect 23386 94968 23442 95024
rect 31482 96056 31538 96112
rect 34978 96056 35034 96112
rect 46846 96328 46902 96384
rect 50342 96328 50398 96384
rect 51170 96328 51226 96384
rect 39578 95920 39634 95976
rect 38474 95784 38530 95840
rect 41970 96192 42026 96248
rect 44178 96192 44234 96248
rect 37830 95240 37886 95296
rect 41142 95240 41198 95296
rect 38566 95104 38622 95160
rect 44086 95104 44142 95160
rect 20626 94852 20682 94888
rect 20626 94832 20628 94852
rect 20628 94832 20680 94852
rect 20680 94832 20682 94852
rect 30286 94988 30342 95024
rect 30286 94968 30288 94988
rect 30288 94968 30340 94988
rect 30340 94968 30342 94988
rect 31666 94968 31722 95024
rect 37278 94580 37334 94616
rect 37278 94560 37280 94580
rect 37280 94560 37332 94580
rect 37332 94560 37334 94580
rect 42706 94424 42762 94480
rect 45374 95260 45430 95296
rect 45374 95240 45376 95260
rect 45376 95240 45428 95260
rect 45428 95240 45430 95260
rect 45190 95104 45246 95160
rect 45558 95104 45614 95160
rect 46662 95104 46718 95160
rect 47950 95240 48006 95296
rect 48226 95240 48282 95296
rect 48134 95104 48190 95160
rect 45098 94424 45154 94480
rect 50802 95104 50858 95160
rect 49882 94424 49938 94480
rect 50158 94424 50214 94480
rect 50158 94152 50214 94208
rect 50986 94016 51042 94072
rect 57610 96600 57666 96656
rect 57886 96600 57942 96656
rect 58070 96600 58126 96656
rect 59542 96600 59598 96656
rect 59726 96600 59782 96656
rect 59910 96600 59966 96656
rect 60462 96600 60518 96656
rect 40866 93608 40922 93664
rect 42614 93608 42670 93664
rect 44086 93608 44142 93664
rect 46662 93608 46718 93664
rect 47950 93608 48006 93664
rect 48778 93628 48834 93664
rect 48778 93608 48780 93628
rect 48780 93608 48832 93628
rect 48832 93608 48834 93628
rect 40866 93336 40922 93392
rect 40590 93200 40646 93256
rect 32862 92812 32918 92848
rect 32862 92792 32864 92812
rect 32864 92792 32916 92812
rect 32916 92792 32918 92812
rect 34150 92812 34206 92848
rect 34150 92792 34152 92812
rect 34152 92792 34204 92812
rect 34204 92792 34206 92812
rect 35254 92792 35310 92848
rect 49054 93608 49110 93664
rect 49606 93608 49662 93664
rect 49974 93608 50030 93664
rect 50618 93608 50674 93664
rect 51262 93608 51318 93664
rect 51446 93608 51502 93664
rect 52182 93608 52238 93664
rect 52550 93608 52606 93664
rect 53286 93608 53342 93664
rect 53746 93608 53802 93664
rect 54022 93608 54078 93664
rect 54206 93628 54262 93664
rect 54206 93608 54208 93628
rect 54208 93608 54260 93628
rect 54260 93608 54262 93628
rect 54574 93608 54630 93664
rect 54942 93608 54998 93664
rect 61566 96736 61622 96792
rect 61750 96736 61806 96792
rect 61934 96736 61990 96792
rect 77114 96872 77170 96928
rect 76930 96600 76986 96656
rect 77114 96600 77170 96656
rect 79506 96736 79562 96792
rect 80150 97144 80206 97200
rect 79230 96600 79286 96656
rect 82174 96600 82230 96656
rect 80150 96328 80206 96384
rect 74630 95920 74686 95976
rect 74814 95920 74870 95976
rect 74814 95648 74870 95704
rect 79506 96056 79562 96112
rect 79690 96056 79746 96112
rect 76838 95956 76840 95976
rect 76840 95956 76892 95976
rect 76892 95956 76894 95976
rect 76838 95920 76894 95956
rect 77022 95920 77078 95976
rect 75182 95512 75238 95568
rect 76102 95512 76158 95568
rect 63958 95240 64014 95296
rect 64142 95276 64144 95296
rect 64144 95276 64196 95296
rect 64196 95276 64198 95296
rect 64142 95240 64198 95276
rect 64326 95240 64382 95296
rect 79506 95376 79562 95432
rect 80242 95920 80298 95976
rect 80518 96192 80574 96248
rect 80426 95920 80482 95976
rect 79506 94968 79562 95024
rect 80058 94968 80114 95024
rect 79230 94016 79286 94072
rect 80518 94968 80574 95024
rect 81438 94968 81494 95024
rect 82542 153992 82598 154048
rect 82542 132232 82598 132288
rect 82634 114280 82690 114336
rect 82450 95648 82506 95704
rect 82634 96736 82690 96792
rect 82818 97552 82874 97608
rect 82910 96736 82966 96792
rect 82174 94560 82230 94616
rect 82358 94560 82414 94616
rect 79506 93880 79562 93936
rect 77022 93608 77078 93664
rect 77298 93608 77354 93664
rect 79046 93608 79102 93664
rect 79506 93336 79562 93392
rect 77482 93064 77538 93120
rect 77666 93064 77722 93120
rect 82634 93744 82690 93800
rect 36726 92828 36728 92848
rect 36728 92828 36780 92848
rect 36780 92828 36782 92848
rect 36726 92792 36782 92828
rect 38382 92792 38438 92848
rect 39946 92792 40002 92848
rect 40590 92792 40646 92848
rect 77666 92792 77722 92848
rect 82082 92792 82138 92848
rect 83278 97008 83334 97064
rect 83554 96056 83610 96112
rect 83370 95784 83426 95840
rect 82910 94968 82966 95024
rect 82726 92928 82782 92984
rect 82450 55256 82506 55312
rect 82450 45464 82506 45520
rect 82450 16632 82506 16688
rect 8114 2624 8170 2680
rect 15290 2624 15346 2680
rect 20718 2624 20774 2680
rect 22650 2508 22706 2544
rect 22650 2488 22652 2508
rect 22652 2488 22704 2508
rect 22704 2488 22706 2508
rect 47766 3168 47822 3224
rect 48686 3168 48742 3224
rect 48686 2896 48742 2952
rect 49974 2896 50030 2952
rect 25042 2624 25098 2680
rect 9770 2216 9826 2272
rect 13910 2216 13966 2272
rect 16302 2216 16358 2272
rect 22098 2216 22154 2272
rect 24122 2216 24178 2272
rect 32678 2216 32734 2272
rect 36174 2216 36230 2272
rect 37462 2236 37518 2272
rect 37462 2216 37464 2236
rect 37464 2216 37516 2236
rect 37516 2216 37518 2236
rect 32770 2080 32826 2136
rect 33966 2100 34022 2136
rect 36266 2116 36268 2136
rect 36268 2116 36320 2136
rect 36320 2116 36322 2136
rect 33966 2080 33968 2100
rect 33968 2080 34020 2100
rect 34020 2080 34022 2100
rect 36266 2080 36322 2116
rect 29090 1964 29146 2000
rect 29090 1944 29092 1964
rect 29092 1944 29144 1964
rect 29144 1944 29146 1964
rect 30470 1964 30526 2000
rect 30470 1944 30472 1964
rect 30472 1944 30524 1964
rect 30524 1944 30526 1964
rect 31666 1944 31722 2000
rect 17498 1808 17554 1864
rect 21086 1808 21142 1864
rect 22282 1808 22338 1864
rect 25778 1828 25834 1864
rect 25778 1808 25780 1828
rect 25780 1808 25832 1828
rect 25832 1808 25834 1828
rect 9770 1400 9826 1456
rect 26974 1808 27030 1864
rect 28170 1808 28226 1864
rect 12438 1300 12440 1320
rect 12440 1300 12492 1320
rect 12492 1300 12494 1320
rect 12438 1264 12494 1300
rect 19246 1264 19302 1320
rect 30286 1264 30342 1320
rect 35530 1300 35532 1320
rect 35532 1300 35584 1320
rect 35584 1300 35586 1320
rect 35530 1264 35586 1300
rect 39854 1264 39910 1320
rect 17958 1128 18014 1184
rect 19338 1128 19394 1184
rect 28998 1128 29054 1184
rect 34518 1128 34574 1184
rect 39946 1148 40002 1184
rect 39946 1128 39948 1148
rect 39948 1128 40000 1148
rect 40000 1128 40002 1148
rect 24766 992 24822 1048
rect 30378 1012 30434 1048
rect 30378 992 30380 1012
rect 30380 992 30432 1012
rect 30432 992 30434 1012
rect 41326 1012 41382 1048
rect 41326 992 41328 1012
rect 41328 992 41380 1012
rect 41380 992 41382 1012
rect 44914 1284 44970 1320
rect 48226 1300 48228 1320
rect 48228 1300 48280 1320
rect 48280 1300 48282 1320
rect 44914 1264 44916 1284
rect 44916 1264 44968 1284
rect 44968 1264 44970 1284
rect 48226 1264 48282 1300
rect 53470 2896 53526 2952
rect 84106 169904 84162 169960
rect 84106 164056 84162 164112
rect 84014 96192 84070 96248
rect 83738 95104 83794 95160
rect 51354 2252 51356 2272
rect 51356 2252 51408 2272
rect 51408 2252 51410 2272
rect 51354 2216 51410 2252
rect 52550 2216 52606 2272
rect 52366 1128 52422 1184
rect 42706 992 42762 1048
rect 46754 992 46810 1048
rect 49606 992 49662 1048
rect 27618 856 27674 912
rect 42798 856 42854 912
rect 44086 876 44142 912
rect 44086 856 44088 876
rect 44088 856 44140 876
rect 44140 856 44142 876
rect 24766 720 24822 776
rect 33138 740 33194 776
rect 33138 720 33140 740
rect 33140 720 33192 740
rect 33192 720 33194 740
rect 20626 196 20682 232
rect 20626 176 20628 196
rect 20628 176 20680 196
rect 20680 176 20682 196
rect 46846 856 46902 912
rect 50986 720 51042 776
rect 54666 992 54722 1048
rect 53746 468 53802 504
rect 53746 448 53748 468
rect 53748 448 53800 468
rect 53800 448 53802 468
rect 55034 720 55090 776
rect 55126 448 55182 504
rect 83002 2916 83058 2952
rect 83002 2896 83004 2916
rect 83004 2896 83056 2916
rect 83056 2896 83058 2916
rect 82910 2760 82966 2816
rect 83186 3168 83242 3224
rect 83186 2760 83242 2816
rect 85956 187162 86012 187164
rect 86036 187162 86092 187164
rect 86116 187162 86172 187164
rect 86196 187162 86252 187164
rect 85956 187110 85982 187162
rect 85982 187110 86012 187162
rect 86036 187110 86046 187162
rect 86046 187110 86092 187162
rect 86116 187110 86162 187162
rect 86162 187110 86172 187162
rect 86196 187110 86226 187162
rect 86226 187110 86252 187162
rect 85956 187108 86012 187110
rect 86036 187108 86092 187110
rect 86116 187108 86172 187110
rect 86196 187108 86252 187110
rect 89956 187162 90012 187164
rect 90036 187162 90092 187164
rect 90116 187162 90172 187164
rect 90196 187162 90252 187164
rect 89956 187110 89982 187162
rect 89982 187110 90012 187162
rect 90036 187110 90046 187162
rect 90046 187110 90092 187162
rect 90116 187110 90162 187162
rect 90162 187110 90172 187162
rect 90196 187110 90226 187162
rect 90226 187110 90252 187162
rect 89956 187108 90012 187110
rect 90036 187108 90092 187110
rect 90116 187108 90172 187110
rect 90196 187108 90252 187110
rect 87956 186618 88012 186620
rect 88036 186618 88092 186620
rect 88116 186618 88172 186620
rect 88196 186618 88252 186620
rect 87956 186566 87982 186618
rect 87982 186566 88012 186618
rect 88036 186566 88046 186618
rect 88046 186566 88092 186618
rect 88116 186566 88162 186618
rect 88162 186566 88172 186618
rect 88196 186566 88226 186618
rect 88226 186566 88252 186618
rect 87956 186564 88012 186566
rect 88036 186564 88092 186566
rect 88116 186564 88172 186566
rect 88196 186564 88252 186566
rect 85956 186074 86012 186076
rect 86036 186074 86092 186076
rect 86116 186074 86172 186076
rect 86196 186074 86252 186076
rect 85956 186022 85982 186074
rect 85982 186022 86012 186074
rect 86036 186022 86046 186074
rect 86046 186022 86092 186074
rect 86116 186022 86162 186074
rect 86162 186022 86172 186074
rect 86196 186022 86226 186074
rect 86226 186022 86252 186074
rect 85956 186020 86012 186022
rect 86036 186020 86092 186022
rect 86116 186020 86172 186022
rect 86196 186020 86252 186022
rect 89956 186074 90012 186076
rect 90036 186074 90092 186076
rect 90116 186074 90172 186076
rect 90196 186074 90252 186076
rect 89956 186022 89982 186074
rect 89982 186022 90012 186074
rect 90036 186022 90046 186074
rect 90046 186022 90092 186074
rect 90116 186022 90162 186074
rect 90162 186022 90172 186074
rect 90196 186022 90226 186074
rect 90226 186022 90252 186074
rect 89956 186020 90012 186022
rect 90036 186020 90092 186022
rect 90116 186020 90172 186022
rect 90196 186020 90252 186022
rect 87956 185530 88012 185532
rect 88036 185530 88092 185532
rect 88116 185530 88172 185532
rect 88196 185530 88252 185532
rect 87956 185478 87982 185530
rect 87982 185478 88012 185530
rect 88036 185478 88046 185530
rect 88046 185478 88092 185530
rect 88116 185478 88162 185530
rect 88162 185478 88172 185530
rect 88196 185478 88226 185530
rect 88226 185478 88252 185530
rect 87956 185476 88012 185478
rect 88036 185476 88092 185478
rect 88116 185476 88172 185478
rect 88196 185476 88252 185478
rect 85956 184986 86012 184988
rect 86036 184986 86092 184988
rect 86116 184986 86172 184988
rect 86196 184986 86252 184988
rect 85956 184934 85982 184986
rect 85982 184934 86012 184986
rect 86036 184934 86046 184986
rect 86046 184934 86092 184986
rect 86116 184934 86162 184986
rect 86162 184934 86172 184986
rect 86196 184934 86226 184986
rect 86226 184934 86252 184986
rect 85956 184932 86012 184934
rect 86036 184932 86092 184934
rect 86116 184932 86172 184934
rect 86196 184932 86252 184934
rect 89956 184986 90012 184988
rect 90036 184986 90092 184988
rect 90116 184986 90172 184988
rect 90196 184986 90252 184988
rect 89956 184934 89982 184986
rect 89982 184934 90012 184986
rect 90036 184934 90046 184986
rect 90046 184934 90092 184986
rect 90116 184934 90162 184986
rect 90162 184934 90172 184986
rect 90196 184934 90226 184986
rect 90226 184934 90252 184986
rect 89956 184932 90012 184934
rect 90036 184932 90092 184934
rect 90116 184932 90172 184934
rect 90196 184932 90252 184934
rect 87956 184442 88012 184444
rect 88036 184442 88092 184444
rect 88116 184442 88172 184444
rect 88196 184442 88252 184444
rect 87956 184390 87982 184442
rect 87982 184390 88012 184442
rect 88036 184390 88046 184442
rect 88046 184390 88092 184442
rect 88116 184390 88162 184442
rect 88162 184390 88172 184442
rect 88196 184390 88226 184442
rect 88226 184390 88252 184442
rect 87956 184388 88012 184390
rect 88036 184388 88092 184390
rect 88116 184388 88172 184390
rect 88196 184388 88252 184390
rect 85956 183898 86012 183900
rect 86036 183898 86092 183900
rect 86116 183898 86172 183900
rect 86196 183898 86252 183900
rect 85956 183846 85982 183898
rect 85982 183846 86012 183898
rect 86036 183846 86046 183898
rect 86046 183846 86092 183898
rect 86116 183846 86162 183898
rect 86162 183846 86172 183898
rect 86196 183846 86226 183898
rect 86226 183846 86252 183898
rect 85956 183844 86012 183846
rect 86036 183844 86092 183846
rect 86116 183844 86172 183846
rect 86196 183844 86252 183846
rect 89956 183898 90012 183900
rect 90036 183898 90092 183900
rect 90116 183898 90172 183900
rect 90196 183898 90252 183900
rect 89956 183846 89982 183898
rect 89982 183846 90012 183898
rect 90036 183846 90046 183898
rect 90046 183846 90092 183898
rect 90116 183846 90162 183898
rect 90162 183846 90172 183898
rect 90196 183846 90226 183898
rect 90226 183846 90252 183898
rect 89956 183844 90012 183846
rect 90036 183844 90092 183846
rect 90116 183844 90172 183846
rect 90196 183844 90252 183846
rect 87956 183354 88012 183356
rect 88036 183354 88092 183356
rect 88116 183354 88172 183356
rect 88196 183354 88252 183356
rect 87956 183302 87982 183354
rect 87982 183302 88012 183354
rect 88036 183302 88046 183354
rect 88046 183302 88092 183354
rect 88116 183302 88162 183354
rect 88162 183302 88172 183354
rect 88196 183302 88226 183354
rect 88226 183302 88252 183354
rect 87956 183300 88012 183302
rect 88036 183300 88092 183302
rect 88116 183300 88172 183302
rect 88196 183300 88252 183302
rect 85956 182810 86012 182812
rect 86036 182810 86092 182812
rect 86116 182810 86172 182812
rect 86196 182810 86252 182812
rect 85956 182758 85982 182810
rect 85982 182758 86012 182810
rect 86036 182758 86046 182810
rect 86046 182758 86092 182810
rect 86116 182758 86162 182810
rect 86162 182758 86172 182810
rect 86196 182758 86226 182810
rect 86226 182758 86252 182810
rect 85956 182756 86012 182758
rect 86036 182756 86092 182758
rect 86116 182756 86172 182758
rect 86196 182756 86252 182758
rect 89956 182810 90012 182812
rect 90036 182810 90092 182812
rect 90116 182810 90172 182812
rect 90196 182810 90252 182812
rect 89956 182758 89982 182810
rect 89982 182758 90012 182810
rect 90036 182758 90046 182810
rect 90046 182758 90092 182810
rect 90116 182758 90162 182810
rect 90162 182758 90172 182810
rect 90196 182758 90226 182810
rect 90226 182758 90252 182810
rect 89956 182756 90012 182758
rect 90036 182756 90092 182758
rect 90116 182756 90172 182758
rect 90196 182756 90252 182758
rect 87956 182266 88012 182268
rect 88036 182266 88092 182268
rect 88116 182266 88172 182268
rect 88196 182266 88252 182268
rect 87956 182214 87982 182266
rect 87982 182214 88012 182266
rect 88036 182214 88046 182266
rect 88046 182214 88092 182266
rect 88116 182214 88162 182266
rect 88162 182214 88172 182266
rect 88196 182214 88226 182266
rect 88226 182214 88252 182266
rect 87956 182212 88012 182214
rect 88036 182212 88092 182214
rect 88116 182212 88172 182214
rect 88196 182212 88252 182214
rect 85956 181722 86012 181724
rect 86036 181722 86092 181724
rect 86116 181722 86172 181724
rect 86196 181722 86252 181724
rect 85956 181670 85982 181722
rect 85982 181670 86012 181722
rect 86036 181670 86046 181722
rect 86046 181670 86092 181722
rect 86116 181670 86162 181722
rect 86162 181670 86172 181722
rect 86196 181670 86226 181722
rect 86226 181670 86252 181722
rect 85956 181668 86012 181670
rect 86036 181668 86092 181670
rect 86116 181668 86172 181670
rect 86196 181668 86252 181670
rect 89956 181722 90012 181724
rect 90036 181722 90092 181724
rect 90116 181722 90172 181724
rect 90196 181722 90252 181724
rect 89956 181670 89982 181722
rect 89982 181670 90012 181722
rect 90036 181670 90046 181722
rect 90046 181670 90092 181722
rect 90116 181670 90162 181722
rect 90162 181670 90172 181722
rect 90196 181670 90226 181722
rect 90226 181670 90252 181722
rect 89956 181668 90012 181670
rect 90036 181668 90092 181670
rect 90116 181668 90172 181670
rect 90196 181668 90252 181670
rect 87694 181464 87750 181520
rect 87956 181178 88012 181180
rect 88036 181178 88092 181180
rect 88116 181178 88172 181180
rect 88196 181178 88252 181180
rect 87956 181126 87982 181178
rect 87982 181126 88012 181178
rect 88036 181126 88046 181178
rect 88046 181126 88092 181178
rect 88116 181126 88162 181178
rect 88162 181126 88172 181178
rect 88196 181126 88226 181178
rect 88226 181126 88252 181178
rect 87956 181124 88012 181126
rect 88036 181124 88092 181126
rect 88116 181124 88172 181126
rect 88196 181124 88252 181126
rect 85956 180634 86012 180636
rect 86036 180634 86092 180636
rect 86116 180634 86172 180636
rect 86196 180634 86252 180636
rect 85956 180582 85982 180634
rect 85982 180582 86012 180634
rect 86036 180582 86046 180634
rect 86046 180582 86092 180634
rect 86116 180582 86162 180634
rect 86162 180582 86172 180634
rect 86196 180582 86226 180634
rect 86226 180582 86252 180634
rect 85956 180580 86012 180582
rect 86036 180580 86092 180582
rect 86116 180580 86172 180582
rect 86196 180580 86252 180582
rect 89956 180634 90012 180636
rect 90036 180634 90092 180636
rect 90116 180634 90172 180636
rect 90196 180634 90252 180636
rect 89956 180582 89982 180634
rect 89982 180582 90012 180634
rect 90036 180582 90046 180634
rect 90046 180582 90092 180634
rect 90116 180582 90162 180634
rect 90162 180582 90172 180634
rect 90196 180582 90226 180634
rect 90226 180582 90252 180634
rect 89956 180580 90012 180582
rect 90036 180580 90092 180582
rect 90116 180580 90172 180582
rect 90196 180580 90252 180582
rect 87956 180090 88012 180092
rect 88036 180090 88092 180092
rect 88116 180090 88172 180092
rect 88196 180090 88252 180092
rect 87956 180038 87982 180090
rect 87982 180038 88012 180090
rect 88036 180038 88046 180090
rect 88046 180038 88092 180090
rect 88116 180038 88162 180090
rect 88162 180038 88172 180090
rect 88196 180038 88226 180090
rect 88226 180038 88252 180090
rect 87956 180036 88012 180038
rect 88036 180036 88092 180038
rect 88116 180036 88172 180038
rect 88196 180036 88252 180038
rect 85956 179546 86012 179548
rect 86036 179546 86092 179548
rect 86116 179546 86172 179548
rect 86196 179546 86252 179548
rect 85956 179494 85982 179546
rect 85982 179494 86012 179546
rect 86036 179494 86046 179546
rect 86046 179494 86092 179546
rect 86116 179494 86162 179546
rect 86162 179494 86172 179546
rect 86196 179494 86226 179546
rect 86226 179494 86252 179546
rect 85956 179492 86012 179494
rect 86036 179492 86092 179494
rect 86116 179492 86172 179494
rect 86196 179492 86252 179494
rect 89956 179546 90012 179548
rect 90036 179546 90092 179548
rect 90116 179546 90172 179548
rect 90196 179546 90252 179548
rect 89956 179494 89982 179546
rect 89982 179494 90012 179546
rect 90036 179494 90046 179546
rect 90046 179494 90092 179546
rect 90116 179494 90162 179546
rect 90162 179494 90172 179546
rect 90196 179494 90226 179546
rect 90226 179494 90252 179546
rect 89956 179492 90012 179494
rect 90036 179492 90092 179494
rect 90116 179492 90172 179494
rect 90196 179492 90252 179494
rect 87956 179002 88012 179004
rect 88036 179002 88092 179004
rect 88116 179002 88172 179004
rect 88196 179002 88252 179004
rect 87956 178950 87982 179002
rect 87982 178950 88012 179002
rect 88036 178950 88046 179002
rect 88046 178950 88092 179002
rect 88116 178950 88162 179002
rect 88162 178950 88172 179002
rect 88196 178950 88226 179002
rect 88226 178950 88252 179002
rect 87956 178948 88012 178950
rect 88036 178948 88092 178950
rect 88116 178948 88172 178950
rect 88196 178948 88252 178950
rect 85956 178458 86012 178460
rect 86036 178458 86092 178460
rect 86116 178458 86172 178460
rect 86196 178458 86252 178460
rect 85956 178406 85982 178458
rect 85982 178406 86012 178458
rect 86036 178406 86046 178458
rect 86046 178406 86092 178458
rect 86116 178406 86162 178458
rect 86162 178406 86172 178458
rect 86196 178406 86226 178458
rect 86226 178406 86252 178458
rect 85956 178404 86012 178406
rect 86036 178404 86092 178406
rect 86116 178404 86172 178406
rect 86196 178404 86252 178406
rect 89956 178458 90012 178460
rect 90036 178458 90092 178460
rect 90116 178458 90172 178460
rect 90196 178458 90252 178460
rect 89956 178406 89982 178458
rect 89982 178406 90012 178458
rect 90036 178406 90046 178458
rect 90046 178406 90092 178458
rect 90116 178406 90162 178458
rect 90162 178406 90172 178458
rect 90196 178406 90226 178458
rect 90226 178406 90252 178458
rect 89956 178404 90012 178406
rect 90036 178404 90092 178406
rect 90116 178404 90172 178406
rect 90196 178404 90252 178406
rect 87956 177914 88012 177916
rect 88036 177914 88092 177916
rect 88116 177914 88172 177916
rect 88196 177914 88252 177916
rect 87956 177862 87982 177914
rect 87982 177862 88012 177914
rect 88036 177862 88046 177914
rect 88046 177862 88092 177914
rect 88116 177862 88162 177914
rect 88162 177862 88172 177914
rect 88196 177862 88226 177914
rect 88226 177862 88252 177914
rect 87956 177860 88012 177862
rect 88036 177860 88092 177862
rect 88116 177860 88172 177862
rect 88196 177860 88252 177862
rect 87786 177656 87842 177712
rect 85956 177370 86012 177372
rect 86036 177370 86092 177372
rect 86116 177370 86172 177372
rect 86196 177370 86252 177372
rect 85956 177318 85982 177370
rect 85982 177318 86012 177370
rect 86036 177318 86046 177370
rect 86046 177318 86092 177370
rect 86116 177318 86162 177370
rect 86162 177318 86172 177370
rect 86196 177318 86226 177370
rect 86226 177318 86252 177370
rect 85956 177316 86012 177318
rect 86036 177316 86092 177318
rect 86116 177316 86172 177318
rect 86196 177316 86252 177318
rect 85956 176282 86012 176284
rect 86036 176282 86092 176284
rect 86116 176282 86172 176284
rect 86196 176282 86252 176284
rect 85956 176230 85982 176282
rect 85982 176230 86012 176282
rect 86036 176230 86046 176282
rect 86046 176230 86092 176282
rect 86116 176230 86162 176282
rect 86162 176230 86172 176282
rect 86196 176230 86226 176282
rect 86226 176230 86252 176282
rect 85956 176228 86012 176230
rect 86036 176228 86092 176230
rect 86116 176228 86172 176230
rect 86196 176228 86252 176230
rect 85956 175194 86012 175196
rect 86036 175194 86092 175196
rect 86116 175194 86172 175196
rect 86196 175194 86252 175196
rect 85956 175142 85982 175194
rect 85982 175142 86012 175194
rect 86036 175142 86046 175194
rect 86046 175142 86092 175194
rect 86116 175142 86162 175194
rect 86162 175142 86172 175194
rect 86196 175142 86226 175194
rect 86226 175142 86252 175194
rect 85956 175140 86012 175142
rect 86036 175140 86092 175142
rect 86116 175140 86172 175142
rect 86196 175140 86252 175142
rect 87418 174256 87474 174312
rect 85956 174106 86012 174108
rect 86036 174106 86092 174108
rect 86116 174106 86172 174108
rect 86196 174106 86252 174108
rect 85956 174054 85982 174106
rect 85982 174054 86012 174106
rect 86036 174054 86046 174106
rect 86046 174054 86092 174106
rect 86116 174054 86162 174106
rect 86162 174054 86172 174106
rect 86196 174054 86226 174106
rect 86226 174054 86252 174106
rect 85956 174052 86012 174054
rect 86036 174052 86092 174054
rect 86116 174052 86172 174054
rect 86196 174052 86252 174054
rect 87602 173168 87658 173224
rect 85956 173018 86012 173020
rect 86036 173018 86092 173020
rect 86116 173018 86172 173020
rect 86196 173018 86252 173020
rect 85956 172966 85982 173018
rect 85982 172966 86012 173018
rect 86036 172966 86046 173018
rect 86046 172966 86092 173018
rect 86116 172966 86162 173018
rect 86162 172966 86172 173018
rect 86196 172966 86226 173018
rect 86226 172966 86252 173018
rect 85956 172964 86012 172966
rect 86036 172964 86092 172966
rect 86116 172964 86172 172966
rect 86196 172964 86252 172966
rect 85956 171930 86012 171932
rect 86036 171930 86092 171932
rect 86116 171930 86172 171932
rect 86196 171930 86252 171932
rect 85956 171878 85982 171930
rect 85982 171878 86012 171930
rect 86036 171878 86046 171930
rect 86046 171878 86092 171930
rect 86116 171878 86162 171930
rect 86162 171878 86172 171930
rect 86196 171878 86226 171930
rect 86226 171878 86252 171930
rect 85956 171876 86012 171878
rect 86036 171876 86092 171878
rect 86116 171876 86172 171878
rect 86196 171876 86252 171878
rect 85956 170842 86012 170844
rect 86036 170842 86092 170844
rect 86116 170842 86172 170844
rect 86196 170842 86252 170844
rect 85956 170790 85982 170842
rect 85982 170790 86012 170842
rect 86036 170790 86046 170842
rect 86046 170790 86092 170842
rect 86116 170790 86162 170842
rect 86162 170790 86172 170842
rect 86196 170790 86226 170842
rect 86226 170790 86252 170842
rect 85956 170788 86012 170790
rect 86036 170788 86092 170790
rect 86116 170788 86172 170790
rect 86196 170788 86252 170790
rect 85956 169754 86012 169756
rect 86036 169754 86092 169756
rect 86116 169754 86172 169756
rect 86196 169754 86252 169756
rect 85956 169702 85982 169754
rect 85982 169702 86012 169754
rect 86036 169702 86046 169754
rect 86046 169702 86092 169754
rect 86116 169702 86162 169754
rect 86162 169702 86172 169754
rect 86196 169702 86226 169754
rect 86226 169702 86252 169754
rect 85956 169700 86012 169702
rect 86036 169700 86092 169702
rect 86116 169700 86172 169702
rect 86196 169700 86252 169702
rect 85956 168666 86012 168668
rect 86036 168666 86092 168668
rect 86116 168666 86172 168668
rect 86196 168666 86252 168668
rect 85956 168614 85982 168666
rect 85982 168614 86012 168666
rect 86036 168614 86046 168666
rect 86046 168614 86092 168666
rect 86116 168614 86162 168666
rect 86162 168614 86172 168666
rect 86196 168614 86226 168666
rect 86226 168614 86252 168666
rect 85956 168612 86012 168614
rect 86036 168612 86092 168614
rect 86116 168612 86172 168614
rect 86196 168612 86252 168614
rect 87050 168272 87106 168328
rect 85956 167578 86012 167580
rect 86036 167578 86092 167580
rect 86116 167578 86172 167580
rect 86196 167578 86252 167580
rect 85956 167526 85982 167578
rect 85982 167526 86012 167578
rect 86036 167526 86046 167578
rect 86046 167526 86092 167578
rect 86116 167526 86162 167578
rect 86162 167526 86172 167578
rect 86196 167526 86226 167578
rect 86226 167526 86252 167578
rect 85956 167524 86012 167526
rect 86036 167524 86092 167526
rect 86116 167524 86172 167526
rect 86196 167524 86252 167526
rect 85956 166490 86012 166492
rect 86036 166490 86092 166492
rect 86116 166490 86172 166492
rect 86196 166490 86252 166492
rect 85956 166438 85982 166490
rect 85982 166438 86012 166490
rect 86036 166438 86046 166490
rect 86046 166438 86092 166490
rect 86116 166438 86162 166490
rect 86162 166438 86172 166490
rect 86196 166438 86226 166490
rect 86226 166438 86252 166490
rect 85956 166436 86012 166438
rect 86036 166436 86092 166438
rect 86116 166436 86172 166438
rect 86196 166436 86252 166438
rect 87510 165688 87566 165744
rect 85956 165402 86012 165404
rect 86036 165402 86092 165404
rect 86116 165402 86172 165404
rect 86196 165402 86252 165404
rect 85956 165350 85982 165402
rect 85982 165350 86012 165402
rect 86036 165350 86046 165402
rect 86046 165350 86092 165402
rect 86116 165350 86162 165402
rect 86162 165350 86172 165402
rect 86196 165350 86226 165402
rect 86226 165350 86252 165402
rect 85956 165348 86012 165350
rect 86036 165348 86092 165350
rect 86116 165348 86172 165350
rect 86196 165348 86252 165350
rect 85956 164314 86012 164316
rect 86036 164314 86092 164316
rect 86116 164314 86172 164316
rect 86196 164314 86252 164316
rect 85956 164262 85982 164314
rect 85982 164262 86012 164314
rect 86036 164262 86046 164314
rect 86046 164262 86092 164314
rect 86116 164262 86162 164314
rect 86162 164262 86172 164314
rect 86196 164262 86226 164314
rect 86226 164262 86252 164314
rect 85956 164260 86012 164262
rect 86036 164260 86092 164262
rect 86116 164260 86172 164262
rect 86196 164260 86252 164262
rect 85956 163226 86012 163228
rect 86036 163226 86092 163228
rect 86116 163226 86172 163228
rect 86196 163226 86252 163228
rect 85956 163174 85982 163226
rect 85982 163174 86012 163226
rect 86036 163174 86046 163226
rect 86046 163174 86092 163226
rect 86116 163174 86162 163226
rect 86162 163174 86172 163226
rect 86196 163174 86226 163226
rect 86226 163174 86252 163226
rect 85956 163172 86012 163174
rect 86036 163172 86092 163174
rect 86116 163172 86172 163174
rect 86196 163172 86252 163174
rect 85956 162138 86012 162140
rect 86036 162138 86092 162140
rect 86116 162138 86172 162140
rect 86196 162138 86252 162140
rect 85956 162086 85982 162138
rect 85982 162086 86012 162138
rect 86036 162086 86046 162138
rect 86046 162086 86092 162138
rect 86116 162086 86162 162138
rect 86162 162086 86172 162138
rect 86196 162086 86226 162138
rect 86226 162086 86252 162138
rect 85956 162084 86012 162086
rect 86036 162084 86092 162086
rect 86116 162084 86172 162086
rect 86196 162084 86252 162086
rect 85118 161744 85174 161800
rect 85956 161050 86012 161052
rect 86036 161050 86092 161052
rect 86116 161050 86172 161052
rect 86196 161050 86252 161052
rect 85956 160998 85982 161050
rect 85982 160998 86012 161050
rect 86036 160998 86046 161050
rect 86046 160998 86092 161050
rect 86116 160998 86162 161050
rect 86162 160998 86172 161050
rect 86196 160998 86226 161050
rect 86226 160998 86252 161050
rect 85956 160996 86012 160998
rect 86036 160996 86092 160998
rect 86116 160996 86172 160998
rect 86196 160996 86252 160998
rect 85956 159962 86012 159964
rect 86036 159962 86092 159964
rect 86116 159962 86172 159964
rect 86196 159962 86252 159964
rect 85956 159910 85982 159962
rect 85982 159910 86012 159962
rect 86036 159910 86046 159962
rect 86046 159910 86092 159962
rect 86116 159910 86162 159962
rect 86162 159910 86172 159962
rect 86196 159910 86226 159962
rect 86226 159910 86252 159962
rect 85956 159908 86012 159910
rect 86036 159908 86092 159910
rect 86116 159908 86172 159910
rect 86196 159908 86252 159910
rect 87418 159704 87474 159760
rect 85956 158874 86012 158876
rect 86036 158874 86092 158876
rect 86116 158874 86172 158876
rect 86196 158874 86252 158876
rect 85956 158822 85982 158874
rect 85982 158822 86012 158874
rect 86036 158822 86046 158874
rect 86046 158822 86092 158874
rect 86116 158822 86162 158874
rect 86162 158822 86172 158874
rect 86196 158822 86226 158874
rect 86226 158822 86252 158874
rect 85956 158820 86012 158822
rect 86036 158820 86092 158822
rect 86116 158820 86172 158822
rect 86196 158820 86252 158822
rect 86590 158480 86646 158536
rect 85956 157786 86012 157788
rect 86036 157786 86092 157788
rect 86116 157786 86172 157788
rect 86196 157786 86252 157788
rect 85956 157734 85982 157786
rect 85982 157734 86012 157786
rect 86036 157734 86046 157786
rect 86046 157734 86092 157786
rect 86116 157734 86162 157786
rect 86162 157734 86172 157786
rect 86196 157734 86226 157786
rect 86226 157734 86252 157786
rect 85956 157732 86012 157734
rect 86036 157732 86092 157734
rect 86116 157732 86172 157734
rect 86196 157732 86252 157734
rect 85956 156698 86012 156700
rect 86036 156698 86092 156700
rect 86116 156698 86172 156700
rect 86196 156698 86252 156700
rect 85956 156646 85982 156698
rect 85982 156646 86012 156698
rect 86036 156646 86046 156698
rect 86046 156646 86092 156698
rect 86116 156646 86162 156698
rect 86162 156646 86172 156698
rect 86196 156646 86226 156698
rect 86226 156646 86252 156698
rect 85956 156644 86012 156646
rect 86036 156644 86092 156646
rect 86116 156644 86172 156646
rect 86196 156644 86252 156646
rect 85956 155610 86012 155612
rect 86036 155610 86092 155612
rect 86116 155610 86172 155612
rect 86196 155610 86252 155612
rect 85956 155558 85982 155610
rect 85982 155558 86012 155610
rect 86036 155558 86046 155610
rect 86046 155558 86092 155610
rect 86116 155558 86162 155610
rect 86162 155558 86172 155610
rect 86196 155558 86226 155610
rect 86226 155558 86252 155610
rect 85956 155556 86012 155558
rect 86036 155556 86092 155558
rect 86116 155556 86172 155558
rect 86196 155556 86252 155558
rect 85956 154522 86012 154524
rect 86036 154522 86092 154524
rect 86116 154522 86172 154524
rect 86196 154522 86252 154524
rect 85956 154470 85982 154522
rect 85982 154470 86012 154522
rect 86036 154470 86046 154522
rect 86046 154470 86092 154522
rect 86116 154470 86162 154522
rect 86162 154470 86172 154522
rect 86196 154470 86226 154522
rect 86226 154470 86252 154522
rect 85956 154468 86012 154470
rect 86036 154468 86092 154470
rect 86116 154468 86172 154470
rect 86196 154468 86252 154470
rect 85956 153434 86012 153436
rect 86036 153434 86092 153436
rect 86116 153434 86172 153436
rect 86196 153434 86252 153436
rect 85956 153382 85982 153434
rect 85982 153382 86012 153434
rect 86036 153382 86046 153434
rect 86046 153382 86092 153434
rect 86116 153382 86162 153434
rect 86162 153382 86172 153434
rect 86196 153382 86226 153434
rect 86226 153382 86252 153434
rect 85956 153380 86012 153382
rect 86036 153380 86092 153382
rect 86116 153380 86172 153382
rect 86196 153380 86252 153382
rect 85956 152346 86012 152348
rect 86036 152346 86092 152348
rect 86116 152346 86172 152348
rect 86196 152346 86252 152348
rect 85956 152294 85982 152346
rect 85982 152294 86012 152346
rect 86036 152294 86046 152346
rect 86046 152294 86092 152346
rect 86116 152294 86162 152346
rect 86162 152294 86172 152346
rect 86196 152294 86226 152346
rect 86226 152294 86252 152346
rect 85956 152292 86012 152294
rect 86036 152292 86092 152294
rect 86116 152292 86172 152294
rect 86196 152292 86252 152294
rect 85956 151258 86012 151260
rect 86036 151258 86092 151260
rect 86116 151258 86172 151260
rect 86196 151258 86252 151260
rect 85956 151206 85982 151258
rect 85982 151206 86012 151258
rect 86036 151206 86046 151258
rect 86046 151206 86092 151258
rect 86116 151206 86162 151258
rect 86162 151206 86172 151258
rect 86196 151206 86226 151258
rect 86226 151206 86252 151258
rect 85956 151204 86012 151206
rect 86036 151204 86092 151206
rect 86116 151204 86172 151206
rect 86196 151204 86252 151206
rect 85956 150170 86012 150172
rect 86036 150170 86092 150172
rect 86116 150170 86172 150172
rect 86196 150170 86252 150172
rect 85956 150118 85982 150170
rect 85982 150118 86012 150170
rect 86036 150118 86046 150170
rect 86046 150118 86092 150170
rect 86116 150118 86162 150170
rect 86162 150118 86172 150170
rect 86196 150118 86226 150170
rect 86226 150118 86252 150170
rect 85956 150116 86012 150118
rect 86036 150116 86092 150118
rect 86116 150116 86172 150118
rect 86196 150116 86252 150118
rect 85956 149082 86012 149084
rect 86036 149082 86092 149084
rect 86116 149082 86172 149084
rect 86196 149082 86252 149084
rect 85956 149030 85982 149082
rect 85982 149030 86012 149082
rect 86036 149030 86046 149082
rect 86046 149030 86092 149082
rect 86116 149030 86162 149082
rect 86162 149030 86172 149082
rect 86196 149030 86226 149082
rect 86226 149030 86252 149082
rect 85956 149028 86012 149030
rect 86036 149028 86092 149030
rect 86116 149028 86172 149030
rect 86196 149028 86252 149030
rect 85956 147994 86012 147996
rect 86036 147994 86092 147996
rect 86116 147994 86172 147996
rect 86196 147994 86252 147996
rect 85956 147942 85982 147994
rect 85982 147942 86012 147994
rect 86036 147942 86046 147994
rect 86046 147942 86092 147994
rect 86116 147942 86162 147994
rect 86162 147942 86172 147994
rect 86196 147942 86226 147994
rect 86226 147942 86252 147994
rect 85956 147940 86012 147942
rect 86036 147940 86092 147942
rect 86116 147940 86172 147942
rect 86196 147940 86252 147942
rect 85956 146906 86012 146908
rect 86036 146906 86092 146908
rect 86116 146906 86172 146908
rect 86196 146906 86252 146908
rect 85956 146854 85982 146906
rect 85982 146854 86012 146906
rect 86036 146854 86046 146906
rect 86046 146854 86092 146906
rect 86116 146854 86162 146906
rect 86162 146854 86172 146906
rect 86196 146854 86226 146906
rect 86226 146854 86252 146906
rect 85956 146852 86012 146854
rect 86036 146852 86092 146854
rect 86116 146852 86172 146854
rect 86196 146852 86252 146854
rect 85956 145818 86012 145820
rect 86036 145818 86092 145820
rect 86116 145818 86172 145820
rect 86196 145818 86252 145820
rect 85956 145766 85982 145818
rect 85982 145766 86012 145818
rect 86036 145766 86046 145818
rect 86046 145766 86092 145818
rect 86116 145766 86162 145818
rect 86162 145766 86172 145818
rect 86196 145766 86226 145818
rect 86226 145766 86252 145818
rect 85956 145764 86012 145766
rect 86036 145764 86092 145766
rect 86116 145764 86172 145766
rect 86196 145764 86252 145766
rect 84566 125740 84568 125760
rect 84568 125740 84620 125760
rect 84620 125740 84622 125760
rect 84566 125704 84622 125740
rect 84474 124072 84530 124128
rect 84382 122984 84438 123040
rect 84474 120944 84530 121000
rect 84382 118224 84438 118280
rect 84198 99456 84254 99512
rect 84106 94696 84162 94752
rect 84014 94424 84070 94480
rect 83462 3032 83518 3088
rect 83554 1536 83610 1592
rect 84290 24404 84346 24440
rect 84290 24384 84292 24404
rect 84292 24384 84344 24404
rect 84344 24384 84346 24404
rect 84290 23316 84346 23352
rect 84290 23296 84292 23316
rect 84292 23296 84344 23316
rect 84344 23296 84346 23316
rect 84566 120128 84622 120184
rect 84566 117272 84622 117328
rect 84566 93200 84622 93256
rect 84566 28872 84622 28928
rect 84566 27548 84568 27568
rect 84568 27548 84620 27568
rect 84620 27548 84622 27568
rect 84566 27512 84622 27548
rect 84566 26152 84622 26208
rect 85956 144730 86012 144732
rect 86036 144730 86092 144732
rect 86116 144730 86172 144732
rect 86196 144730 86252 144732
rect 85956 144678 85982 144730
rect 85982 144678 86012 144730
rect 86036 144678 86046 144730
rect 86046 144678 86092 144730
rect 86116 144678 86162 144730
rect 86162 144678 86172 144730
rect 86196 144678 86226 144730
rect 86226 144678 86252 144730
rect 85956 144676 86012 144678
rect 86036 144676 86092 144678
rect 86116 144676 86172 144678
rect 86196 144676 86252 144678
rect 85486 118360 85542 118416
rect 85118 99456 85174 99512
rect 85118 99320 85174 99376
rect 84750 97416 84806 97472
rect 85026 97416 85082 97472
rect 85670 104080 85726 104136
rect 85956 143642 86012 143644
rect 86036 143642 86092 143644
rect 86116 143642 86172 143644
rect 86196 143642 86252 143644
rect 85956 143590 85982 143642
rect 85982 143590 86012 143642
rect 86036 143590 86046 143642
rect 86046 143590 86092 143642
rect 86116 143590 86162 143642
rect 86162 143590 86172 143642
rect 86196 143590 86226 143642
rect 86226 143590 86252 143642
rect 85956 143588 86012 143590
rect 86036 143588 86092 143590
rect 86116 143588 86172 143590
rect 86196 143588 86252 143590
rect 85956 142554 86012 142556
rect 86036 142554 86092 142556
rect 86116 142554 86172 142556
rect 86196 142554 86252 142556
rect 85956 142502 85982 142554
rect 85982 142502 86012 142554
rect 86036 142502 86046 142554
rect 86046 142502 86092 142554
rect 86116 142502 86162 142554
rect 86162 142502 86172 142554
rect 86196 142502 86226 142554
rect 86226 142502 86252 142554
rect 85956 142500 86012 142502
rect 86036 142500 86092 142502
rect 86116 142500 86172 142502
rect 86196 142500 86252 142502
rect 85956 141466 86012 141468
rect 86036 141466 86092 141468
rect 86116 141466 86172 141468
rect 86196 141466 86252 141468
rect 85956 141414 85982 141466
rect 85982 141414 86012 141466
rect 86036 141414 86046 141466
rect 86046 141414 86092 141466
rect 86116 141414 86162 141466
rect 86162 141414 86172 141466
rect 86196 141414 86226 141466
rect 86226 141414 86252 141466
rect 85956 141412 86012 141414
rect 86036 141412 86092 141414
rect 86116 141412 86172 141414
rect 86196 141412 86252 141414
rect 85956 140378 86012 140380
rect 86036 140378 86092 140380
rect 86116 140378 86172 140380
rect 86196 140378 86252 140380
rect 85956 140326 85982 140378
rect 85982 140326 86012 140378
rect 86036 140326 86046 140378
rect 86046 140326 86092 140378
rect 86116 140326 86162 140378
rect 86162 140326 86172 140378
rect 86196 140326 86226 140378
rect 86226 140326 86252 140378
rect 85956 140324 86012 140326
rect 86036 140324 86092 140326
rect 86116 140324 86172 140326
rect 86196 140324 86252 140326
rect 85956 139290 86012 139292
rect 86036 139290 86092 139292
rect 86116 139290 86172 139292
rect 86196 139290 86252 139292
rect 85956 139238 85982 139290
rect 85982 139238 86012 139290
rect 86036 139238 86046 139290
rect 86046 139238 86092 139290
rect 86116 139238 86162 139290
rect 86162 139238 86172 139290
rect 86196 139238 86226 139290
rect 86226 139238 86252 139290
rect 85956 139236 86012 139238
rect 86036 139236 86092 139238
rect 86116 139236 86172 139238
rect 86196 139236 86252 139238
rect 85956 138202 86012 138204
rect 86036 138202 86092 138204
rect 86116 138202 86172 138204
rect 86196 138202 86252 138204
rect 85956 138150 85982 138202
rect 85982 138150 86012 138202
rect 86036 138150 86046 138202
rect 86046 138150 86092 138202
rect 86116 138150 86162 138202
rect 86162 138150 86172 138202
rect 86196 138150 86226 138202
rect 86226 138150 86252 138202
rect 85956 138148 86012 138150
rect 86036 138148 86092 138150
rect 86116 138148 86172 138150
rect 86196 138148 86252 138150
rect 86498 137808 86554 137864
rect 85956 137114 86012 137116
rect 86036 137114 86092 137116
rect 86116 137114 86172 137116
rect 86196 137114 86252 137116
rect 85956 137062 85982 137114
rect 85982 137062 86012 137114
rect 86036 137062 86046 137114
rect 86046 137062 86092 137114
rect 86116 137062 86162 137114
rect 86162 137062 86172 137114
rect 86196 137062 86226 137114
rect 86226 137062 86252 137114
rect 85956 137060 86012 137062
rect 86036 137060 86092 137062
rect 86116 137060 86172 137062
rect 86196 137060 86252 137062
rect 86314 136312 86370 136368
rect 85956 136026 86012 136028
rect 86036 136026 86092 136028
rect 86116 136026 86172 136028
rect 86196 136026 86252 136028
rect 85956 135974 85982 136026
rect 85982 135974 86012 136026
rect 86036 135974 86046 136026
rect 86046 135974 86092 136026
rect 86116 135974 86162 136026
rect 86162 135974 86172 136026
rect 86196 135974 86226 136026
rect 86226 135974 86252 136026
rect 85956 135972 86012 135974
rect 86036 135972 86092 135974
rect 86116 135972 86172 135974
rect 86196 135972 86252 135974
rect 85956 134938 86012 134940
rect 86036 134938 86092 134940
rect 86116 134938 86172 134940
rect 86196 134938 86252 134940
rect 85956 134886 85982 134938
rect 85982 134886 86012 134938
rect 86036 134886 86046 134938
rect 86046 134886 86092 134938
rect 86116 134886 86162 134938
rect 86162 134886 86172 134938
rect 86196 134886 86226 134938
rect 86226 134886 86252 134938
rect 85956 134884 86012 134886
rect 86036 134884 86092 134886
rect 86116 134884 86172 134886
rect 86196 134884 86252 134886
rect 85956 133850 86012 133852
rect 86036 133850 86092 133852
rect 86116 133850 86172 133852
rect 86196 133850 86252 133852
rect 85956 133798 85982 133850
rect 85982 133798 86012 133850
rect 86036 133798 86046 133850
rect 86046 133798 86092 133850
rect 86116 133798 86162 133850
rect 86162 133798 86172 133850
rect 86196 133798 86226 133850
rect 86226 133798 86252 133850
rect 85956 133796 86012 133798
rect 86036 133796 86092 133798
rect 86116 133796 86172 133798
rect 86196 133796 86252 133798
rect 85956 132762 86012 132764
rect 86036 132762 86092 132764
rect 86116 132762 86172 132764
rect 86196 132762 86252 132764
rect 85956 132710 85982 132762
rect 85982 132710 86012 132762
rect 86036 132710 86046 132762
rect 86046 132710 86092 132762
rect 86116 132710 86162 132762
rect 86162 132710 86172 132762
rect 86196 132710 86226 132762
rect 86226 132710 86252 132762
rect 85956 132708 86012 132710
rect 86036 132708 86092 132710
rect 86116 132708 86172 132710
rect 86196 132708 86252 132710
rect 85956 131674 86012 131676
rect 86036 131674 86092 131676
rect 86116 131674 86172 131676
rect 86196 131674 86252 131676
rect 85956 131622 85982 131674
rect 85982 131622 86012 131674
rect 86036 131622 86046 131674
rect 86046 131622 86092 131674
rect 86116 131622 86162 131674
rect 86162 131622 86172 131674
rect 86196 131622 86226 131674
rect 86226 131622 86252 131674
rect 85956 131620 86012 131622
rect 86036 131620 86092 131622
rect 86116 131620 86172 131622
rect 86196 131620 86252 131622
rect 85956 130586 86012 130588
rect 86036 130586 86092 130588
rect 86116 130586 86172 130588
rect 86196 130586 86252 130588
rect 85956 130534 85982 130586
rect 85982 130534 86012 130586
rect 86036 130534 86046 130586
rect 86046 130534 86092 130586
rect 86116 130534 86162 130586
rect 86162 130534 86172 130586
rect 86196 130534 86226 130586
rect 86226 130534 86252 130586
rect 85956 130532 86012 130534
rect 86036 130532 86092 130534
rect 86116 130532 86172 130534
rect 86196 130532 86252 130534
rect 85956 129498 86012 129500
rect 86036 129498 86092 129500
rect 86116 129498 86172 129500
rect 86196 129498 86252 129500
rect 85956 129446 85982 129498
rect 85982 129446 86012 129498
rect 86036 129446 86046 129498
rect 86046 129446 86092 129498
rect 86116 129446 86162 129498
rect 86162 129446 86172 129498
rect 86196 129446 86226 129498
rect 86226 129446 86252 129498
rect 85956 129444 86012 129446
rect 86036 129444 86092 129446
rect 86116 129444 86172 129446
rect 86196 129444 86252 129446
rect 85956 128410 86012 128412
rect 86036 128410 86092 128412
rect 86116 128410 86172 128412
rect 86196 128410 86252 128412
rect 85956 128358 85982 128410
rect 85982 128358 86012 128410
rect 86036 128358 86046 128410
rect 86046 128358 86092 128410
rect 86116 128358 86162 128410
rect 86162 128358 86172 128410
rect 86196 128358 86226 128410
rect 86226 128358 86252 128410
rect 85956 128356 86012 128358
rect 86036 128356 86092 128358
rect 86116 128356 86172 128358
rect 86196 128356 86252 128358
rect 85956 127322 86012 127324
rect 86036 127322 86092 127324
rect 86116 127322 86172 127324
rect 86196 127322 86252 127324
rect 85956 127270 85982 127322
rect 85982 127270 86012 127322
rect 86036 127270 86046 127322
rect 86046 127270 86092 127322
rect 86116 127270 86162 127322
rect 86162 127270 86172 127322
rect 86196 127270 86226 127322
rect 86226 127270 86252 127322
rect 85956 127268 86012 127270
rect 86036 127268 86092 127270
rect 86116 127268 86172 127270
rect 86196 127268 86252 127270
rect 85956 126234 86012 126236
rect 86036 126234 86092 126236
rect 86116 126234 86172 126236
rect 86196 126234 86252 126236
rect 85956 126182 85982 126234
rect 85982 126182 86012 126234
rect 86036 126182 86046 126234
rect 86046 126182 86092 126234
rect 86116 126182 86162 126234
rect 86162 126182 86172 126234
rect 86196 126182 86226 126234
rect 86226 126182 86252 126234
rect 85956 126180 86012 126182
rect 86036 126180 86092 126182
rect 86116 126180 86172 126182
rect 86196 126180 86252 126182
rect 85956 125146 86012 125148
rect 86036 125146 86092 125148
rect 86116 125146 86172 125148
rect 86196 125146 86252 125148
rect 85956 125094 85982 125146
rect 85982 125094 86012 125146
rect 86036 125094 86046 125146
rect 86046 125094 86092 125146
rect 86116 125094 86162 125146
rect 86162 125094 86172 125146
rect 86196 125094 86226 125146
rect 86226 125094 86252 125146
rect 85956 125092 86012 125094
rect 86036 125092 86092 125094
rect 86116 125092 86172 125094
rect 86196 125092 86252 125094
rect 85956 124058 86012 124060
rect 86036 124058 86092 124060
rect 86116 124058 86172 124060
rect 86196 124058 86252 124060
rect 85956 124006 85982 124058
rect 85982 124006 86012 124058
rect 86036 124006 86046 124058
rect 86046 124006 86092 124058
rect 86116 124006 86162 124058
rect 86162 124006 86172 124058
rect 86196 124006 86226 124058
rect 86226 124006 86252 124058
rect 85956 124004 86012 124006
rect 86036 124004 86092 124006
rect 86116 124004 86172 124006
rect 86196 124004 86252 124006
rect 85956 122970 86012 122972
rect 86036 122970 86092 122972
rect 86116 122970 86172 122972
rect 86196 122970 86252 122972
rect 85956 122918 85982 122970
rect 85982 122918 86012 122970
rect 86036 122918 86046 122970
rect 86046 122918 86092 122970
rect 86116 122918 86162 122970
rect 86162 122918 86172 122970
rect 86196 122918 86226 122970
rect 86226 122918 86252 122970
rect 85956 122916 86012 122918
rect 86036 122916 86092 122918
rect 86116 122916 86172 122918
rect 86196 122916 86252 122918
rect 86406 135224 86462 135280
rect 85956 121882 86012 121884
rect 86036 121882 86092 121884
rect 86116 121882 86172 121884
rect 86196 121882 86252 121884
rect 85956 121830 85982 121882
rect 85982 121830 86012 121882
rect 86036 121830 86046 121882
rect 86046 121830 86092 121882
rect 86116 121830 86162 121882
rect 86162 121830 86172 121882
rect 86196 121830 86226 121882
rect 86226 121830 86252 121882
rect 85956 121828 86012 121830
rect 86036 121828 86092 121830
rect 86116 121828 86172 121830
rect 86196 121828 86252 121830
rect 85956 120794 86012 120796
rect 86036 120794 86092 120796
rect 86116 120794 86172 120796
rect 86196 120794 86252 120796
rect 85956 120742 85982 120794
rect 85982 120742 86012 120794
rect 86036 120742 86046 120794
rect 86046 120742 86092 120794
rect 86116 120742 86162 120794
rect 86162 120742 86172 120794
rect 86196 120742 86226 120794
rect 86226 120742 86252 120794
rect 85956 120740 86012 120742
rect 86036 120740 86092 120742
rect 86116 120740 86172 120742
rect 86196 120740 86252 120742
rect 85956 119706 86012 119708
rect 86036 119706 86092 119708
rect 86116 119706 86172 119708
rect 86196 119706 86252 119708
rect 85956 119654 85982 119706
rect 85982 119654 86012 119706
rect 86036 119654 86046 119706
rect 86046 119654 86092 119706
rect 86116 119654 86162 119706
rect 86162 119654 86172 119706
rect 86196 119654 86226 119706
rect 86226 119654 86252 119706
rect 85956 119652 86012 119654
rect 86036 119652 86092 119654
rect 86116 119652 86172 119654
rect 86196 119652 86252 119654
rect 85956 118618 86012 118620
rect 86036 118618 86092 118620
rect 86116 118618 86172 118620
rect 86196 118618 86252 118620
rect 85956 118566 85982 118618
rect 85982 118566 86012 118618
rect 86036 118566 86046 118618
rect 86046 118566 86092 118618
rect 86116 118566 86162 118618
rect 86162 118566 86172 118618
rect 86196 118566 86226 118618
rect 86226 118566 86252 118618
rect 85956 118564 86012 118566
rect 86036 118564 86092 118566
rect 86116 118564 86172 118566
rect 86196 118564 86252 118566
rect 85956 117530 86012 117532
rect 86036 117530 86092 117532
rect 86116 117530 86172 117532
rect 86196 117530 86252 117532
rect 85956 117478 85982 117530
rect 85982 117478 86012 117530
rect 86036 117478 86046 117530
rect 86046 117478 86092 117530
rect 86116 117478 86162 117530
rect 86162 117478 86172 117530
rect 86196 117478 86226 117530
rect 86226 117478 86252 117530
rect 85956 117476 86012 117478
rect 86036 117476 86092 117478
rect 86116 117476 86172 117478
rect 86196 117476 86252 117478
rect 85956 116442 86012 116444
rect 86036 116442 86092 116444
rect 86116 116442 86172 116444
rect 86196 116442 86252 116444
rect 85956 116390 85982 116442
rect 85982 116390 86012 116442
rect 86036 116390 86046 116442
rect 86046 116390 86092 116442
rect 86116 116390 86162 116442
rect 86162 116390 86172 116442
rect 86196 116390 86226 116442
rect 86226 116390 86252 116442
rect 85956 116388 86012 116390
rect 86036 116388 86092 116390
rect 86116 116388 86172 116390
rect 86196 116388 86252 116390
rect 86314 116048 86370 116104
rect 85956 115354 86012 115356
rect 86036 115354 86092 115356
rect 86116 115354 86172 115356
rect 86196 115354 86252 115356
rect 85956 115302 85982 115354
rect 85982 115302 86012 115354
rect 86036 115302 86046 115354
rect 86046 115302 86092 115354
rect 86116 115302 86162 115354
rect 86162 115302 86172 115354
rect 86196 115302 86226 115354
rect 86226 115302 86252 115354
rect 85956 115300 86012 115302
rect 86036 115300 86092 115302
rect 86116 115300 86172 115302
rect 86196 115300 86252 115302
rect 85956 114266 86012 114268
rect 86036 114266 86092 114268
rect 86116 114266 86172 114268
rect 86196 114266 86252 114268
rect 85956 114214 85982 114266
rect 85982 114214 86012 114266
rect 86036 114214 86046 114266
rect 86046 114214 86092 114266
rect 86116 114214 86162 114266
rect 86162 114214 86172 114266
rect 86196 114214 86226 114266
rect 86226 114214 86252 114266
rect 85956 114212 86012 114214
rect 86036 114212 86092 114214
rect 86116 114212 86172 114214
rect 86196 114212 86252 114214
rect 85956 113178 86012 113180
rect 86036 113178 86092 113180
rect 86116 113178 86172 113180
rect 86196 113178 86252 113180
rect 85956 113126 85982 113178
rect 85982 113126 86012 113178
rect 86036 113126 86046 113178
rect 86046 113126 86092 113178
rect 86116 113126 86162 113178
rect 86162 113126 86172 113178
rect 86196 113126 86226 113178
rect 86226 113126 86252 113178
rect 85956 113124 86012 113126
rect 86036 113124 86092 113126
rect 86116 113124 86172 113126
rect 86196 113124 86252 113126
rect 85956 112090 86012 112092
rect 86036 112090 86092 112092
rect 86116 112090 86172 112092
rect 86196 112090 86252 112092
rect 85956 112038 85982 112090
rect 85982 112038 86012 112090
rect 86036 112038 86046 112090
rect 86046 112038 86092 112090
rect 86116 112038 86162 112090
rect 86162 112038 86172 112090
rect 86196 112038 86226 112090
rect 86226 112038 86252 112090
rect 85956 112036 86012 112038
rect 86036 112036 86092 112038
rect 86116 112036 86172 112038
rect 86196 112036 86252 112038
rect 85956 111002 86012 111004
rect 86036 111002 86092 111004
rect 86116 111002 86172 111004
rect 86196 111002 86252 111004
rect 85956 110950 85982 111002
rect 85982 110950 86012 111002
rect 86036 110950 86046 111002
rect 86046 110950 86092 111002
rect 86116 110950 86162 111002
rect 86162 110950 86172 111002
rect 86196 110950 86226 111002
rect 86226 110950 86252 111002
rect 85956 110948 86012 110950
rect 86036 110948 86092 110950
rect 86116 110948 86172 110950
rect 86196 110948 86252 110950
rect 85956 109914 86012 109916
rect 86036 109914 86092 109916
rect 86116 109914 86172 109916
rect 86196 109914 86252 109916
rect 85956 109862 85982 109914
rect 85982 109862 86012 109914
rect 86036 109862 86046 109914
rect 86046 109862 86092 109914
rect 86116 109862 86162 109914
rect 86162 109862 86172 109914
rect 86196 109862 86226 109914
rect 86226 109862 86252 109914
rect 85956 109860 86012 109862
rect 86036 109860 86092 109862
rect 86116 109860 86172 109862
rect 86196 109860 86252 109862
rect 85956 108826 86012 108828
rect 86036 108826 86092 108828
rect 86116 108826 86172 108828
rect 86196 108826 86252 108828
rect 85956 108774 85982 108826
rect 85982 108774 86012 108826
rect 86036 108774 86046 108826
rect 86046 108774 86092 108826
rect 86116 108774 86162 108826
rect 86162 108774 86172 108826
rect 86196 108774 86226 108826
rect 86226 108774 86252 108826
rect 85956 108772 86012 108774
rect 86036 108772 86092 108774
rect 86116 108772 86172 108774
rect 86196 108772 86252 108774
rect 85956 107738 86012 107740
rect 86036 107738 86092 107740
rect 86116 107738 86172 107740
rect 86196 107738 86252 107740
rect 85956 107686 85982 107738
rect 85982 107686 86012 107738
rect 86036 107686 86046 107738
rect 86046 107686 86092 107738
rect 86116 107686 86162 107738
rect 86162 107686 86172 107738
rect 86196 107686 86226 107738
rect 86226 107686 86252 107738
rect 85956 107684 86012 107686
rect 86036 107684 86092 107686
rect 86116 107684 86172 107686
rect 86196 107684 86252 107686
rect 85956 106650 86012 106652
rect 86036 106650 86092 106652
rect 86116 106650 86172 106652
rect 86196 106650 86252 106652
rect 85956 106598 85982 106650
rect 85982 106598 86012 106650
rect 86036 106598 86046 106650
rect 86046 106598 86092 106650
rect 86116 106598 86162 106650
rect 86162 106598 86172 106650
rect 86196 106598 86226 106650
rect 86226 106598 86252 106650
rect 85956 106596 86012 106598
rect 86036 106596 86092 106598
rect 86116 106596 86172 106598
rect 86196 106596 86252 106598
rect 86498 113464 86554 113520
rect 85956 105562 86012 105564
rect 86036 105562 86092 105564
rect 86116 105562 86172 105564
rect 86196 105562 86252 105564
rect 85956 105510 85982 105562
rect 85982 105510 86012 105562
rect 86036 105510 86046 105562
rect 86046 105510 86092 105562
rect 86116 105510 86162 105562
rect 86162 105510 86172 105562
rect 86196 105510 86226 105562
rect 86226 105510 86252 105562
rect 85956 105508 86012 105510
rect 86036 105508 86092 105510
rect 86116 105508 86172 105510
rect 86196 105508 86252 105510
rect 85956 104474 86012 104476
rect 86036 104474 86092 104476
rect 86116 104474 86172 104476
rect 86196 104474 86252 104476
rect 85956 104422 85982 104474
rect 85982 104422 86012 104474
rect 86036 104422 86046 104474
rect 86046 104422 86092 104474
rect 86116 104422 86162 104474
rect 86162 104422 86172 104474
rect 86196 104422 86226 104474
rect 86226 104422 86252 104474
rect 85956 104420 86012 104422
rect 86036 104420 86092 104422
rect 86116 104420 86172 104422
rect 86196 104420 86252 104422
rect 86406 106256 86462 106312
rect 85956 103386 86012 103388
rect 86036 103386 86092 103388
rect 86116 103386 86172 103388
rect 86196 103386 86252 103388
rect 85956 103334 85982 103386
rect 85982 103334 86012 103386
rect 86036 103334 86046 103386
rect 86046 103334 86092 103386
rect 86116 103334 86162 103386
rect 86162 103334 86172 103386
rect 86196 103334 86226 103386
rect 86226 103334 86252 103386
rect 85956 103332 86012 103334
rect 86036 103332 86092 103334
rect 86116 103332 86172 103334
rect 86196 103332 86252 103334
rect 85956 102298 86012 102300
rect 86036 102298 86092 102300
rect 86116 102298 86172 102300
rect 86196 102298 86252 102300
rect 85956 102246 85982 102298
rect 85982 102246 86012 102298
rect 86036 102246 86046 102298
rect 86046 102246 86092 102298
rect 86116 102246 86162 102298
rect 86162 102246 86172 102298
rect 86196 102246 86226 102298
rect 86226 102246 86252 102298
rect 85956 102244 86012 102246
rect 86036 102244 86092 102246
rect 86116 102244 86172 102246
rect 86196 102244 86252 102246
rect 85956 101210 86012 101212
rect 86036 101210 86092 101212
rect 86116 101210 86172 101212
rect 86196 101210 86252 101212
rect 85956 101158 85982 101210
rect 85982 101158 86012 101210
rect 86036 101158 86046 101210
rect 86046 101158 86092 101210
rect 86116 101158 86162 101210
rect 86162 101158 86172 101210
rect 86196 101158 86226 101210
rect 86226 101158 86252 101210
rect 85956 101156 86012 101158
rect 86036 101156 86092 101158
rect 86116 101156 86172 101158
rect 86196 101156 86252 101158
rect 85956 100122 86012 100124
rect 86036 100122 86092 100124
rect 86116 100122 86172 100124
rect 86196 100122 86252 100124
rect 85956 100070 85982 100122
rect 85982 100070 86012 100122
rect 86036 100070 86046 100122
rect 86046 100070 86092 100122
rect 86116 100070 86162 100122
rect 86162 100070 86172 100122
rect 86196 100070 86226 100122
rect 86226 100070 86252 100122
rect 85956 100068 86012 100070
rect 86036 100068 86092 100070
rect 86116 100068 86172 100070
rect 86196 100068 86252 100070
rect 85394 99048 85450 99104
rect 84934 94424 84990 94480
rect 85578 95376 85634 95432
rect 85118 93608 85174 93664
rect 85026 93472 85082 93528
rect 85026 85312 85082 85368
rect 84750 32020 84806 32056
rect 84750 32000 84752 32020
rect 84752 32000 84804 32020
rect 84804 32000 84806 32020
rect 84750 30268 84752 30288
rect 84752 30268 84804 30288
rect 84804 30268 84806 30288
rect 84750 30232 84806 30268
rect 85026 84904 85082 84960
rect 85026 84632 85082 84688
rect 85394 85040 85450 85096
rect 85578 92012 85580 92032
rect 85580 92012 85632 92032
rect 85632 92012 85634 92032
rect 85578 91976 85634 92012
rect 85956 99034 86012 99036
rect 86036 99034 86092 99036
rect 86116 99034 86172 99036
rect 86196 99034 86252 99036
rect 85956 98982 85982 99034
rect 85982 98982 86012 99034
rect 86036 98982 86046 99034
rect 86046 98982 86092 99034
rect 86116 98982 86162 99034
rect 86162 98982 86172 99034
rect 86196 98982 86226 99034
rect 86226 98982 86252 99034
rect 85956 98980 86012 98982
rect 86036 98980 86092 98982
rect 86116 98980 86172 98982
rect 86196 98980 86252 98982
rect 85956 97946 86012 97948
rect 86036 97946 86092 97948
rect 86116 97946 86172 97948
rect 86196 97946 86252 97948
rect 85956 97894 85982 97946
rect 85982 97894 86012 97946
rect 86036 97894 86046 97946
rect 86046 97894 86092 97946
rect 86116 97894 86162 97946
rect 86162 97894 86172 97946
rect 86196 97894 86226 97946
rect 86226 97894 86252 97946
rect 85956 97892 86012 97894
rect 86036 97892 86092 97894
rect 86116 97892 86172 97894
rect 86196 97892 86252 97894
rect 85956 96858 86012 96860
rect 86036 96858 86092 96860
rect 86116 96858 86172 96860
rect 86196 96858 86252 96860
rect 85956 96806 85982 96858
rect 85982 96806 86012 96858
rect 86036 96806 86046 96858
rect 86046 96806 86092 96858
rect 86116 96806 86162 96858
rect 86162 96806 86172 96858
rect 86196 96806 86226 96858
rect 86226 96806 86252 96858
rect 85956 96804 86012 96806
rect 86036 96804 86092 96806
rect 86116 96804 86172 96806
rect 86196 96804 86252 96806
rect 85956 95770 86012 95772
rect 86036 95770 86092 95772
rect 86116 95770 86172 95772
rect 86196 95770 86252 95772
rect 85956 95718 85982 95770
rect 85982 95718 86012 95770
rect 86036 95718 86046 95770
rect 86046 95718 86092 95770
rect 86116 95718 86162 95770
rect 86162 95718 86172 95770
rect 86196 95718 86226 95770
rect 86226 95718 86252 95770
rect 85956 95716 86012 95718
rect 86036 95716 86092 95718
rect 86116 95716 86172 95718
rect 86196 95716 86252 95718
rect 87326 156984 87382 157040
rect 87142 154808 87198 154864
rect 86774 152496 86830 152552
rect 86682 151000 86738 151056
rect 86682 104624 86738 104680
rect 86590 101360 86646 101416
rect 86498 99320 86554 99376
rect 85956 94682 86012 94684
rect 86036 94682 86092 94684
rect 86116 94682 86172 94684
rect 86196 94682 86252 94684
rect 85956 94630 85982 94682
rect 85982 94630 86012 94682
rect 86036 94630 86046 94682
rect 86046 94630 86092 94682
rect 86116 94630 86162 94682
rect 86162 94630 86172 94682
rect 86196 94630 86226 94682
rect 86226 94630 86252 94682
rect 85956 94628 86012 94630
rect 86036 94628 86092 94630
rect 86116 94628 86172 94630
rect 86196 94628 86252 94630
rect 85956 93594 86012 93596
rect 86036 93594 86092 93596
rect 86116 93594 86172 93596
rect 86196 93594 86252 93596
rect 85956 93542 85982 93594
rect 85982 93542 86012 93594
rect 86036 93542 86046 93594
rect 86046 93542 86092 93594
rect 86116 93542 86162 93594
rect 86162 93542 86172 93594
rect 86196 93542 86226 93594
rect 86226 93542 86252 93594
rect 85956 93540 86012 93542
rect 86036 93540 86092 93542
rect 86116 93540 86172 93542
rect 86196 93540 86252 93542
rect 85956 92506 86012 92508
rect 86036 92506 86092 92508
rect 86116 92506 86172 92508
rect 86196 92506 86252 92508
rect 85956 92454 85982 92506
rect 85982 92454 86012 92506
rect 86036 92454 86046 92506
rect 86046 92454 86092 92506
rect 86116 92454 86162 92506
rect 86162 92454 86172 92506
rect 86196 92454 86226 92506
rect 86226 92454 86252 92506
rect 85956 92452 86012 92454
rect 86036 92452 86092 92454
rect 86116 92452 86172 92454
rect 86196 92452 86252 92454
rect 85956 91418 86012 91420
rect 86036 91418 86092 91420
rect 86116 91418 86172 91420
rect 86196 91418 86252 91420
rect 85956 91366 85982 91418
rect 85982 91366 86012 91418
rect 86036 91366 86046 91418
rect 86046 91366 86092 91418
rect 86116 91366 86162 91418
rect 86162 91366 86172 91418
rect 86196 91366 86226 91418
rect 86226 91366 86252 91418
rect 85956 91364 86012 91366
rect 86036 91364 86092 91366
rect 86116 91364 86172 91366
rect 86196 91364 86252 91366
rect 85956 90330 86012 90332
rect 86036 90330 86092 90332
rect 86116 90330 86172 90332
rect 86196 90330 86252 90332
rect 85956 90278 85982 90330
rect 85982 90278 86012 90330
rect 86036 90278 86046 90330
rect 86046 90278 86092 90330
rect 86116 90278 86162 90330
rect 86162 90278 86172 90330
rect 86196 90278 86226 90330
rect 86226 90278 86252 90330
rect 85956 90276 86012 90278
rect 86036 90276 86092 90278
rect 86116 90276 86172 90278
rect 86196 90276 86252 90278
rect 85956 89242 86012 89244
rect 86036 89242 86092 89244
rect 86116 89242 86172 89244
rect 86196 89242 86252 89244
rect 85956 89190 85982 89242
rect 85982 89190 86012 89242
rect 86036 89190 86046 89242
rect 86046 89190 86092 89242
rect 86116 89190 86162 89242
rect 86162 89190 86172 89242
rect 86196 89190 86226 89242
rect 86226 89190 86252 89242
rect 85956 89188 86012 89190
rect 86036 89188 86092 89190
rect 86116 89188 86172 89190
rect 86196 89188 86252 89190
rect 85956 88154 86012 88156
rect 86036 88154 86092 88156
rect 86116 88154 86172 88156
rect 86196 88154 86252 88156
rect 85956 88102 85982 88154
rect 85982 88102 86012 88154
rect 86036 88102 86046 88154
rect 86046 88102 86092 88154
rect 86116 88102 86162 88154
rect 86162 88102 86172 88154
rect 86196 88102 86226 88154
rect 86226 88102 86252 88154
rect 85956 88100 86012 88102
rect 86036 88100 86092 88102
rect 86116 88100 86172 88102
rect 86196 88100 86252 88102
rect 85956 87066 86012 87068
rect 86036 87066 86092 87068
rect 86116 87066 86172 87068
rect 86196 87066 86252 87068
rect 85956 87014 85982 87066
rect 85982 87014 86012 87066
rect 86036 87014 86046 87066
rect 86046 87014 86092 87066
rect 86116 87014 86162 87066
rect 86162 87014 86172 87066
rect 86196 87014 86226 87066
rect 86226 87014 86252 87066
rect 85956 87012 86012 87014
rect 86036 87012 86092 87014
rect 86116 87012 86172 87014
rect 86196 87012 86252 87014
rect 85956 85978 86012 85980
rect 86036 85978 86092 85980
rect 86116 85978 86172 85980
rect 86196 85978 86252 85980
rect 85956 85926 85982 85978
rect 85982 85926 86012 85978
rect 86036 85926 86046 85978
rect 86046 85926 86092 85978
rect 86116 85926 86162 85978
rect 86162 85926 86172 85978
rect 86196 85926 86226 85978
rect 86226 85926 86252 85978
rect 85956 85924 86012 85926
rect 86036 85924 86092 85926
rect 86116 85924 86172 85926
rect 86196 85924 86252 85926
rect 85956 84890 86012 84892
rect 86036 84890 86092 84892
rect 86116 84890 86172 84892
rect 86196 84890 86252 84892
rect 85956 84838 85982 84890
rect 85982 84838 86012 84890
rect 86036 84838 86046 84890
rect 86046 84838 86092 84890
rect 86116 84838 86162 84890
rect 86162 84838 86172 84890
rect 86196 84838 86226 84890
rect 86226 84838 86252 84890
rect 85956 84836 86012 84838
rect 86036 84836 86092 84838
rect 86116 84836 86172 84838
rect 86196 84836 86252 84838
rect 85956 83802 86012 83804
rect 86036 83802 86092 83804
rect 86116 83802 86172 83804
rect 86196 83802 86252 83804
rect 85956 83750 85982 83802
rect 85982 83750 86012 83802
rect 86036 83750 86046 83802
rect 86046 83750 86092 83802
rect 86116 83750 86162 83802
rect 86162 83750 86172 83802
rect 86196 83750 86226 83802
rect 86226 83750 86252 83802
rect 85956 83748 86012 83750
rect 86036 83748 86092 83750
rect 86116 83748 86172 83750
rect 86196 83748 86252 83750
rect 85956 82714 86012 82716
rect 86036 82714 86092 82716
rect 86116 82714 86172 82716
rect 86196 82714 86252 82716
rect 85956 82662 85982 82714
rect 85982 82662 86012 82714
rect 86036 82662 86046 82714
rect 86046 82662 86092 82714
rect 86116 82662 86162 82714
rect 86162 82662 86172 82714
rect 86196 82662 86226 82714
rect 86226 82662 86252 82714
rect 85956 82660 86012 82662
rect 86036 82660 86092 82662
rect 86116 82660 86172 82662
rect 86196 82660 86252 82662
rect 85956 81626 86012 81628
rect 86036 81626 86092 81628
rect 86116 81626 86172 81628
rect 86196 81626 86252 81628
rect 85956 81574 85982 81626
rect 85982 81574 86012 81626
rect 86036 81574 86046 81626
rect 86046 81574 86092 81626
rect 86116 81574 86162 81626
rect 86162 81574 86172 81626
rect 86196 81574 86226 81626
rect 86226 81574 86252 81626
rect 85956 81572 86012 81574
rect 86036 81572 86092 81574
rect 86116 81572 86172 81574
rect 86196 81572 86252 81574
rect 85956 80538 86012 80540
rect 86036 80538 86092 80540
rect 86116 80538 86172 80540
rect 86196 80538 86252 80540
rect 85956 80486 85982 80538
rect 85982 80486 86012 80538
rect 86036 80486 86046 80538
rect 86046 80486 86092 80538
rect 86116 80486 86162 80538
rect 86162 80486 86172 80538
rect 86196 80486 86226 80538
rect 86226 80486 86252 80538
rect 85956 80484 86012 80486
rect 86036 80484 86092 80486
rect 86116 80484 86172 80486
rect 86196 80484 86252 80486
rect 85956 79450 86012 79452
rect 86036 79450 86092 79452
rect 86116 79450 86172 79452
rect 86196 79450 86252 79452
rect 85956 79398 85982 79450
rect 85982 79398 86012 79450
rect 86036 79398 86046 79450
rect 86046 79398 86092 79450
rect 86116 79398 86162 79450
rect 86162 79398 86172 79450
rect 86196 79398 86226 79450
rect 86226 79398 86252 79450
rect 85956 79396 86012 79398
rect 86036 79396 86092 79398
rect 86116 79396 86172 79398
rect 86196 79396 86252 79398
rect 85956 78362 86012 78364
rect 86036 78362 86092 78364
rect 86116 78362 86172 78364
rect 86196 78362 86252 78364
rect 85956 78310 85982 78362
rect 85982 78310 86012 78362
rect 86036 78310 86046 78362
rect 86046 78310 86092 78362
rect 86116 78310 86162 78362
rect 86162 78310 86172 78362
rect 86196 78310 86226 78362
rect 86226 78310 86252 78362
rect 85956 78308 86012 78310
rect 86036 78308 86092 78310
rect 86116 78308 86172 78310
rect 86196 78308 86252 78310
rect 85956 77274 86012 77276
rect 86036 77274 86092 77276
rect 86116 77274 86172 77276
rect 86196 77274 86252 77276
rect 85956 77222 85982 77274
rect 85982 77222 86012 77274
rect 86036 77222 86046 77274
rect 86046 77222 86092 77274
rect 86116 77222 86162 77274
rect 86162 77222 86172 77274
rect 86196 77222 86226 77274
rect 86226 77222 86252 77274
rect 85956 77220 86012 77222
rect 86036 77220 86092 77222
rect 86116 77220 86172 77222
rect 86196 77220 86252 77222
rect 85956 76186 86012 76188
rect 86036 76186 86092 76188
rect 86116 76186 86172 76188
rect 86196 76186 86252 76188
rect 85956 76134 85982 76186
rect 85982 76134 86012 76186
rect 86036 76134 86046 76186
rect 86046 76134 86092 76186
rect 86116 76134 86162 76186
rect 86162 76134 86172 76186
rect 86196 76134 86226 76186
rect 86226 76134 86252 76186
rect 85956 76132 86012 76134
rect 86036 76132 86092 76134
rect 86116 76132 86172 76134
rect 86196 76132 86252 76134
rect 85956 75098 86012 75100
rect 86036 75098 86092 75100
rect 86116 75098 86172 75100
rect 86196 75098 86252 75100
rect 85956 75046 85982 75098
rect 85982 75046 86012 75098
rect 86036 75046 86046 75098
rect 86046 75046 86092 75098
rect 86116 75046 86162 75098
rect 86162 75046 86172 75098
rect 86196 75046 86226 75098
rect 86226 75046 86252 75098
rect 85956 75044 86012 75046
rect 86036 75044 86092 75046
rect 86116 75044 86172 75046
rect 86196 75044 86252 75046
rect 85956 74010 86012 74012
rect 86036 74010 86092 74012
rect 86116 74010 86172 74012
rect 86196 74010 86252 74012
rect 85956 73958 85982 74010
rect 85982 73958 86012 74010
rect 86036 73958 86046 74010
rect 86046 73958 86092 74010
rect 86116 73958 86162 74010
rect 86162 73958 86172 74010
rect 86196 73958 86226 74010
rect 86226 73958 86252 74010
rect 85956 73956 86012 73958
rect 86036 73956 86092 73958
rect 86116 73956 86172 73958
rect 86196 73956 86252 73958
rect 85956 72922 86012 72924
rect 86036 72922 86092 72924
rect 86116 72922 86172 72924
rect 86196 72922 86252 72924
rect 85956 72870 85982 72922
rect 85982 72870 86012 72922
rect 86036 72870 86046 72922
rect 86046 72870 86092 72922
rect 86116 72870 86162 72922
rect 86162 72870 86172 72922
rect 86196 72870 86226 72922
rect 86226 72870 86252 72922
rect 85956 72868 86012 72870
rect 86036 72868 86092 72870
rect 86116 72868 86172 72870
rect 86196 72868 86252 72870
rect 85956 71834 86012 71836
rect 86036 71834 86092 71836
rect 86116 71834 86172 71836
rect 86196 71834 86252 71836
rect 85956 71782 85982 71834
rect 85982 71782 86012 71834
rect 86036 71782 86046 71834
rect 86046 71782 86092 71834
rect 86116 71782 86162 71834
rect 86162 71782 86172 71834
rect 86196 71782 86226 71834
rect 86226 71782 86252 71834
rect 85956 71780 86012 71782
rect 86036 71780 86092 71782
rect 86116 71780 86172 71782
rect 86196 71780 86252 71782
rect 85956 70746 86012 70748
rect 86036 70746 86092 70748
rect 86116 70746 86172 70748
rect 86196 70746 86252 70748
rect 85956 70694 85982 70746
rect 85982 70694 86012 70746
rect 86036 70694 86046 70746
rect 86046 70694 86092 70746
rect 86116 70694 86162 70746
rect 86162 70694 86172 70746
rect 86196 70694 86226 70746
rect 86226 70694 86252 70746
rect 85956 70692 86012 70694
rect 86036 70692 86092 70694
rect 86116 70692 86172 70694
rect 86196 70692 86252 70694
rect 85956 69658 86012 69660
rect 86036 69658 86092 69660
rect 86116 69658 86172 69660
rect 86196 69658 86252 69660
rect 85956 69606 85982 69658
rect 85982 69606 86012 69658
rect 86036 69606 86046 69658
rect 86046 69606 86092 69658
rect 86116 69606 86162 69658
rect 86162 69606 86172 69658
rect 86196 69606 86226 69658
rect 86226 69606 86252 69658
rect 85956 69604 86012 69606
rect 86036 69604 86092 69606
rect 86116 69604 86172 69606
rect 86196 69604 86252 69606
rect 85956 68570 86012 68572
rect 86036 68570 86092 68572
rect 86116 68570 86172 68572
rect 86196 68570 86252 68572
rect 85956 68518 85982 68570
rect 85982 68518 86012 68570
rect 86036 68518 86046 68570
rect 86046 68518 86092 68570
rect 86116 68518 86162 68570
rect 86162 68518 86172 68570
rect 86196 68518 86226 68570
rect 86226 68518 86252 68570
rect 85956 68516 86012 68518
rect 86036 68516 86092 68518
rect 86116 68516 86172 68518
rect 86196 68516 86252 68518
rect 85956 67482 86012 67484
rect 86036 67482 86092 67484
rect 86116 67482 86172 67484
rect 86196 67482 86252 67484
rect 85956 67430 85982 67482
rect 85982 67430 86012 67482
rect 86036 67430 86046 67482
rect 86046 67430 86092 67482
rect 86116 67430 86162 67482
rect 86162 67430 86172 67482
rect 86196 67430 86226 67482
rect 86226 67430 86252 67482
rect 85956 67428 86012 67430
rect 86036 67428 86092 67430
rect 86116 67428 86172 67430
rect 86196 67428 86252 67430
rect 85956 66394 86012 66396
rect 86036 66394 86092 66396
rect 86116 66394 86172 66396
rect 86196 66394 86252 66396
rect 85956 66342 85982 66394
rect 85982 66342 86012 66394
rect 86036 66342 86046 66394
rect 86046 66342 86092 66394
rect 86116 66342 86162 66394
rect 86162 66342 86172 66394
rect 86196 66342 86226 66394
rect 86226 66342 86252 66394
rect 85956 66340 86012 66342
rect 86036 66340 86092 66342
rect 86116 66340 86172 66342
rect 86196 66340 86252 66342
rect 85956 65306 86012 65308
rect 86036 65306 86092 65308
rect 86116 65306 86172 65308
rect 86196 65306 86252 65308
rect 85956 65254 85982 65306
rect 85982 65254 86012 65306
rect 86036 65254 86046 65306
rect 86046 65254 86092 65306
rect 86116 65254 86162 65306
rect 86162 65254 86172 65306
rect 86196 65254 86226 65306
rect 86226 65254 86252 65306
rect 85956 65252 86012 65254
rect 86036 65252 86092 65254
rect 86116 65252 86172 65254
rect 86196 65252 86252 65254
rect 85956 64218 86012 64220
rect 86036 64218 86092 64220
rect 86116 64218 86172 64220
rect 86196 64218 86252 64220
rect 85956 64166 85982 64218
rect 85982 64166 86012 64218
rect 86036 64166 86046 64218
rect 86046 64166 86092 64218
rect 86116 64166 86162 64218
rect 86162 64166 86172 64218
rect 86196 64166 86226 64218
rect 86226 64166 86252 64218
rect 85956 64164 86012 64166
rect 86036 64164 86092 64166
rect 86116 64164 86172 64166
rect 86196 64164 86252 64166
rect 85956 63130 86012 63132
rect 86036 63130 86092 63132
rect 86116 63130 86172 63132
rect 86196 63130 86252 63132
rect 85956 63078 85982 63130
rect 85982 63078 86012 63130
rect 86036 63078 86046 63130
rect 86046 63078 86092 63130
rect 86116 63078 86162 63130
rect 86162 63078 86172 63130
rect 86196 63078 86226 63130
rect 86226 63078 86252 63130
rect 85956 63076 86012 63078
rect 86036 63076 86092 63078
rect 86116 63076 86172 63078
rect 86196 63076 86252 63078
rect 85956 62042 86012 62044
rect 86036 62042 86092 62044
rect 86116 62042 86172 62044
rect 86196 62042 86252 62044
rect 85956 61990 85982 62042
rect 85982 61990 86012 62042
rect 86036 61990 86046 62042
rect 86046 61990 86092 62042
rect 86116 61990 86162 62042
rect 86162 61990 86172 62042
rect 86196 61990 86226 62042
rect 86226 61990 86252 62042
rect 85956 61988 86012 61990
rect 86036 61988 86092 61990
rect 86116 61988 86172 61990
rect 86196 61988 86252 61990
rect 85956 60954 86012 60956
rect 86036 60954 86092 60956
rect 86116 60954 86172 60956
rect 86196 60954 86252 60956
rect 85956 60902 85982 60954
rect 85982 60902 86012 60954
rect 86036 60902 86046 60954
rect 86046 60902 86092 60954
rect 86116 60902 86162 60954
rect 86162 60902 86172 60954
rect 86196 60902 86226 60954
rect 86226 60902 86252 60954
rect 85956 60900 86012 60902
rect 86036 60900 86092 60902
rect 86116 60900 86172 60902
rect 86196 60900 86252 60902
rect 85956 59866 86012 59868
rect 86036 59866 86092 59868
rect 86116 59866 86172 59868
rect 86196 59866 86252 59868
rect 85956 59814 85982 59866
rect 85982 59814 86012 59866
rect 86036 59814 86046 59866
rect 86046 59814 86092 59866
rect 86116 59814 86162 59866
rect 86162 59814 86172 59866
rect 86196 59814 86226 59866
rect 86226 59814 86252 59866
rect 85956 59812 86012 59814
rect 86036 59812 86092 59814
rect 86116 59812 86172 59814
rect 86196 59812 86252 59814
rect 85956 58778 86012 58780
rect 86036 58778 86092 58780
rect 86116 58778 86172 58780
rect 86196 58778 86252 58780
rect 85956 58726 85982 58778
rect 85982 58726 86012 58778
rect 86036 58726 86046 58778
rect 86046 58726 86092 58778
rect 86116 58726 86162 58778
rect 86162 58726 86172 58778
rect 86196 58726 86226 58778
rect 86226 58726 86252 58778
rect 85956 58724 86012 58726
rect 86036 58724 86092 58726
rect 86116 58724 86172 58726
rect 86196 58724 86252 58726
rect 85956 57690 86012 57692
rect 86036 57690 86092 57692
rect 86116 57690 86172 57692
rect 86196 57690 86252 57692
rect 85956 57638 85982 57690
rect 85982 57638 86012 57690
rect 86036 57638 86046 57690
rect 86046 57638 86092 57690
rect 86116 57638 86162 57690
rect 86162 57638 86172 57690
rect 86196 57638 86226 57690
rect 86226 57638 86252 57690
rect 85956 57636 86012 57638
rect 86036 57636 86092 57638
rect 86116 57636 86172 57638
rect 86196 57636 86252 57638
rect 85956 56602 86012 56604
rect 86036 56602 86092 56604
rect 86116 56602 86172 56604
rect 86196 56602 86252 56604
rect 85956 56550 85982 56602
rect 85982 56550 86012 56602
rect 86036 56550 86046 56602
rect 86046 56550 86092 56602
rect 86116 56550 86162 56602
rect 86162 56550 86172 56602
rect 86196 56550 86226 56602
rect 86226 56550 86252 56602
rect 85956 56548 86012 56550
rect 86036 56548 86092 56550
rect 86116 56548 86172 56550
rect 86196 56548 86252 56550
rect 85956 55514 86012 55516
rect 86036 55514 86092 55516
rect 86116 55514 86172 55516
rect 86196 55514 86252 55516
rect 85956 55462 85982 55514
rect 85982 55462 86012 55514
rect 86036 55462 86046 55514
rect 86046 55462 86092 55514
rect 86116 55462 86162 55514
rect 86162 55462 86172 55514
rect 86196 55462 86226 55514
rect 86226 55462 86252 55514
rect 85956 55460 86012 55462
rect 86036 55460 86092 55462
rect 86116 55460 86172 55462
rect 86196 55460 86252 55462
rect 85956 54426 86012 54428
rect 86036 54426 86092 54428
rect 86116 54426 86172 54428
rect 86196 54426 86252 54428
rect 85956 54374 85982 54426
rect 85982 54374 86012 54426
rect 86036 54374 86046 54426
rect 86046 54374 86092 54426
rect 86116 54374 86162 54426
rect 86162 54374 86172 54426
rect 86196 54374 86226 54426
rect 86226 54374 86252 54426
rect 85956 54372 86012 54374
rect 86036 54372 86092 54374
rect 86116 54372 86172 54374
rect 86196 54372 86252 54374
rect 85956 53338 86012 53340
rect 86036 53338 86092 53340
rect 86116 53338 86172 53340
rect 86196 53338 86252 53340
rect 85956 53286 85982 53338
rect 85982 53286 86012 53338
rect 86036 53286 86046 53338
rect 86046 53286 86092 53338
rect 86116 53286 86162 53338
rect 86162 53286 86172 53338
rect 86196 53286 86226 53338
rect 86226 53286 86252 53338
rect 85956 53284 86012 53286
rect 86036 53284 86092 53286
rect 86116 53284 86172 53286
rect 86196 53284 86252 53286
rect 85956 52250 86012 52252
rect 86036 52250 86092 52252
rect 86116 52250 86172 52252
rect 86196 52250 86252 52252
rect 85956 52198 85982 52250
rect 85982 52198 86012 52250
rect 86036 52198 86046 52250
rect 86046 52198 86092 52250
rect 86116 52198 86162 52250
rect 86162 52198 86172 52250
rect 86196 52198 86226 52250
rect 86226 52198 86252 52250
rect 85956 52196 86012 52198
rect 86036 52196 86092 52198
rect 86116 52196 86172 52198
rect 86196 52196 86252 52198
rect 85956 51162 86012 51164
rect 86036 51162 86092 51164
rect 86116 51162 86172 51164
rect 86196 51162 86252 51164
rect 85956 51110 85982 51162
rect 85982 51110 86012 51162
rect 86036 51110 86046 51162
rect 86046 51110 86092 51162
rect 86116 51110 86162 51162
rect 86162 51110 86172 51162
rect 86196 51110 86226 51162
rect 86226 51110 86252 51162
rect 85956 51108 86012 51110
rect 86036 51108 86092 51110
rect 86116 51108 86172 51110
rect 86196 51108 86252 51110
rect 85956 50074 86012 50076
rect 86036 50074 86092 50076
rect 86116 50074 86172 50076
rect 86196 50074 86252 50076
rect 85956 50022 85982 50074
rect 85982 50022 86012 50074
rect 86036 50022 86046 50074
rect 86046 50022 86092 50074
rect 86116 50022 86162 50074
rect 86162 50022 86172 50074
rect 86196 50022 86226 50074
rect 86226 50022 86252 50074
rect 85956 50020 86012 50022
rect 86036 50020 86092 50022
rect 86116 50020 86172 50022
rect 86196 50020 86252 50022
rect 85956 48986 86012 48988
rect 86036 48986 86092 48988
rect 86116 48986 86172 48988
rect 86196 48986 86252 48988
rect 85956 48934 85982 48986
rect 85982 48934 86012 48986
rect 86036 48934 86046 48986
rect 86046 48934 86092 48986
rect 86116 48934 86162 48986
rect 86162 48934 86172 48986
rect 86196 48934 86226 48986
rect 86226 48934 86252 48986
rect 85956 48932 86012 48934
rect 86036 48932 86092 48934
rect 86116 48932 86172 48934
rect 86196 48932 86252 48934
rect 85956 47898 86012 47900
rect 86036 47898 86092 47900
rect 86116 47898 86172 47900
rect 86196 47898 86252 47900
rect 85956 47846 85982 47898
rect 85982 47846 86012 47898
rect 86036 47846 86046 47898
rect 86046 47846 86092 47898
rect 86116 47846 86162 47898
rect 86162 47846 86172 47898
rect 86196 47846 86226 47898
rect 86226 47846 86252 47898
rect 85956 47844 86012 47846
rect 86036 47844 86092 47846
rect 86116 47844 86172 47846
rect 86196 47844 86252 47846
rect 85956 46810 86012 46812
rect 86036 46810 86092 46812
rect 86116 46810 86172 46812
rect 86196 46810 86252 46812
rect 85956 46758 85982 46810
rect 85982 46758 86012 46810
rect 86036 46758 86046 46810
rect 86046 46758 86092 46810
rect 86116 46758 86162 46810
rect 86162 46758 86172 46810
rect 86196 46758 86226 46810
rect 86226 46758 86252 46810
rect 85956 46756 86012 46758
rect 86036 46756 86092 46758
rect 86116 46756 86172 46758
rect 86196 46756 86252 46758
rect 85956 45722 86012 45724
rect 86036 45722 86092 45724
rect 86116 45722 86172 45724
rect 86196 45722 86252 45724
rect 85956 45670 85982 45722
rect 85982 45670 86012 45722
rect 86036 45670 86046 45722
rect 86046 45670 86092 45722
rect 86116 45670 86162 45722
rect 86162 45670 86172 45722
rect 86196 45670 86226 45722
rect 86226 45670 86252 45722
rect 85956 45668 86012 45670
rect 86036 45668 86092 45670
rect 86116 45668 86172 45670
rect 86196 45668 86252 45670
rect 85956 44634 86012 44636
rect 86036 44634 86092 44636
rect 86116 44634 86172 44636
rect 86196 44634 86252 44636
rect 85956 44582 85982 44634
rect 85982 44582 86012 44634
rect 86036 44582 86046 44634
rect 86046 44582 86092 44634
rect 86116 44582 86162 44634
rect 86162 44582 86172 44634
rect 86196 44582 86226 44634
rect 86226 44582 86252 44634
rect 85956 44580 86012 44582
rect 86036 44580 86092 44582
rect 86116 44580 86172 44582
rect 86196 44580 86252 44582
rect 85956 43546 86012 43548
rect 86036 43546 86092 43548
rect 86116 43546 86172 43548
rect 86196 43546 86252 43548
rect 85956 43494 85982 43546
rect 85982 43494 86012 43546
rect 86036 43494 86046 43546
rect 86046 43494 86092 43546
rect 86116 43494 86162 43546
rect 86162 43494 86172 43546
rect 86196 43494 86226 43546
rect 86226 43494 86252 43546
rect 85956 43492 86012 43494
rect 86036 43492 86092 43494
rect 86116 43492 86172 43494
rect 86196 43492 86252 43494
rect 85956 42458 86012 42460
rect 86036 42458 86092 42460
rect 86116 42458 86172 42460
rect 86196 42458 86252 42460
rect 85956 42406 85982 42458
rect 85982 42406 86012 42458
rect 86036 42406 86046 42458
rect 86046 42406 86092 42458
rect 86116 42406 86162 42458
rect 86162 42406 86172 42458
rect 86196 42406 86226 42458
rect 86226 42406 86252 42458
rect 85956 42404 86012 42406
rect 86036 42404 86092 42406
rect 86116 42404 86172 42406
rect 86196 42404 86252 42406
rect 85956 41370 86012 41372
rect 86036 41370 86092 41372
rect 86116 41370 86172 41372
rect 86196 41370 86252 41372
rect 85956 41318 85982 41370
rect 85982 41318 86012 41370
rect 86036 41318 86046 41370
rect 86046 41318 86092 41370
rect 86116 41318 86162 41370
rect 86162 41318 86172 41370
rect 86196 41318 86226 41370
rect 86226 41318 86252 41370
rect 85956 41316 86012 41318
rect 86036 41316 86092 41318
rect 86116 41316 86172 41318
rect 86196 41316 86252 41318
rect 85956 40282 86012 40284
rect 86036 40282 86092 40284
rect 86116 40282 86172 40284
rect 86196 40282 86252 40284
rect 85956 40230 85982 40282
rect 85982 40230 86012 40282
rect 86036 40230 86046 40282
rect 86046 40230 86092 40282
rect 86116 40230 86162 40282
rect 86162 40230 86172 40282
rect 86196 40230 86226 40282
rect 86226 40230 86252 40282
rect 85956 40228 86012 40230
rect 86036 40228 86092 40230
rect 86116 40228 86172 40230
rect 86196 40228 86252 40230
rect 85956 39194 86012 39196
rect 86036 39194 86092 39196
rect 86116 39194 86172 39196
rect 86196 39194 86252 39196
rect 85956 39142 85982 39194
rect 85982 39142 86012 39194
rect 86036 39142 86046 39194
rect 86046 39142 86092 39194
rect 86116 39142 86162 39194
rect 86162 39142 86172 39194
rect 86196 39142 86226 39194
rect 86226 39142 86252 39194
rect 85956 39140 86012 39142
rect 86036 39140 86092 39142
rect 86116 39140 86172 39142
rect 86196 39140 86252 39142
rect 85956 38106 86012 38108
rect 86036 38106 86092 38108
rect 86116 38106 86172 38108
rect 86196 38106 86252 38108
rect 85956 38054 85982 38106
rect 85982 38054 86012 38106
rect 86036 38054 86046 38106
rect 86046 38054 86092 38106
rect 86116 38054 86162 38106
rect 86162 38054 86172 38106
rect 86196 38054 86226 38106
rect 86226 38054 86252 38106
rect 85956 38052 86012 38054
rect 86036 38052 86092 38054
rect 86116 38052 86172 38054
rect 86196 38052 86252 38054
rect 85956 37018 86012 37020
rect 86036 37018 86092 37020
rect 86116 37018 86172 37020
rect 86196 37018 86252 37020
rect 85956 36966 85982 37018
rect 85982 36966 86012 37018
rect 86036 36966 86046 37018
rect 86046 36966 86092 37018
rect 86116 36966 86162 37018
rect 86162 36966 86172 37018
rect 86196 36966 86226 37018
rect 86226 36966 86252 37018
rect 85956 36964 86012 36966
rect 86036 36964 86092 36966
rect 86116 36964 86172 36966
rect 86196 36964 86252 36966
rect 85956 35930 86012 35932
rect 86036 35930 86092 35932
rect 86116 35930 86172 35932
rect 86196 35930 86252 35932
rect 85956 35878 85982 35930
rect 85982 35878 86012 35930
rect 86036 35878 86046 35930
rect 86046 35878 86092 35930
rect 86116 35878 86162 35930
rect 86162 35878 86172 35930
rect 86196 35878 86226 35930
rect 86226 35878 86252 35930
rect 85956 35876 86012 35878
rect 86036 35876 86092 35878
rect 86116 35876 86172 35878
rect 86196 35876 86252 35878
rect 85956 34842 86012 34844
rect 86036 34842 86092 34844
rect 86116 34842 86172 34844
rect 86196 34842 86252 34844
rect 85956 34790 85982 34842
rect 85982 34790 86012 34842
rect 86036 34790 86046 34842
rect 86046 34790 86092 34842
rect 86116 34790 86162 34842
rect 86162 34790 86172 34842
rect 86196 34790 86226 34842
rect 86226 34790 86252 34842
rect 85956 34788 86012 34790
rect 86036 34788 86092 34790
rect 86116 34788 86172 34790
rect 86196 34788 86252 34790
rect 85956 33754 86012 33756
rect 86036 33754 86092 33756
rect 86116 33754 86172 33756
rect 86196 33754 86252 33756
rect 85956 33702 85982 33754
rect 85982 33702 86012 33754
rect 86036 33702 86046 33754
rect 86046 33702 86092 33754
rect 86116 33702 86162 33754
rect 86162 33702 86172 33754
rect 86196 33702 86226 33754
rect 86226 33702 86252 33754
rect 85956 33700 86012 33702
rect 86036 33700 86092 33702
rect 86116 33700 86172 33702
rect 86196 33700 86252 33702
rect 85956 32666 86012 32668
rect 86036 32666 86092 32668
rect 86116 32666 86172 32668
rect 86196 32666 86252 32668
rect 85956 32614 85982 32666
rect 85982 32614 86012 32666
rect 86036 32614 86046 32666
rect 86046 32614 86092 32666
rect 86116 32614 86162 32666
rect 86162 32614 86172 32666
rect 86196 32614 86226 32666
rect 86226 32614 86252 32666
rect 85956 32612 86012 32614
rect 86036 32612 86092 32614
rect 86116 32612 86172 32614
rect 86196 32612 86252 32614
rect 85956 31578 86012 31580
rect 86036 31578 86092 31580
rect 86116 31578 86172 31580
rect 86196 31578 86252 31580
rect 85956 31526 85982 31578
rect 85982 31526 86012 31578
rect 86036 31526 86046 31578
rect 86046 31526 86092 31578
rect 86116 31526 86162 31578
rect 86162 31526 86172 31578
rect 86196 31526 86226 31578
rect 86226 31526 86252 31578
rect 85956 31524 86012 31526
rect 86036 31524 86092 31526
rect 86116 31524 86172 31526
rect 86196 31524 86252 31526
rect 85956 30490 86012 30492
rect 86036 30490 86092 30492
rect 86116 30490 86172 30492
rect 86196 30490 86252 30492
rect 85956 30438 85982 30490
rect 85982 30438 86012 30490
rect 86036 30438 86046 30490
rect 86046 30438 86092 30490
rect 86116 30438 86162 30490
rect 86162 30438 86172 30490
rect 86196 30438 86226 30490
rect 86226 30438 86252 30490
rect 85956 30436 86012 30438
rect 86036 30436 86092 30438
rect 86116 30436 86172 30438
rect 86196 30436 86252 30438
rect 85956 29402 86012 29404
rect 86036 29402 86092 29404
rect 86116 29402 86172 29404
rect 86196 29402 86252 29404
rect 85956 29350 85982 29402
rect 85982 29350 86012 29402
rect 86036 29350 86046 29402
rect 86046 29350 86092 29402
rect 86116 29350 86162 29402
rect 86162 29350 86172 29402
rect 86196 29350 86226 29402
rect 86226 29350 86252 29402
rect 85956 29348 86012 29350
rect 86036 29348 86092 29350
rect 86116 29348 86172 29350
rect 86196 29348 86252 29350
rect 85956 28314 86012 28316
rect 86036 28314 86092 28316
rect 86116 28314 86172 28316
rect 86196 28314 86252 28316
rect 85956 28262 85982 28314
rect 85982 28262 86012 28314
rect 86036 28262 86046 28314
rect 86046 28262 86092 28314
rect 86116 28262 86162 28314
rect 86162 28262 86172 28314
rect 86196 28262 86226 28314
rect 86226 28262 86252 28314
rect 85956 28260 86012 28262
rect 86036 28260 86092 28262
rect 86116 28260 86172 28262
rect 86196 28260 86252 28262
rect 85956 27226 86012 27228
rect 86036 27226 86092 27228
rect 86116 27226 86172 27228
rect 86196 27226 86252 27228
rect 85956 27174 85982 27226
rect 85982 27174 86012 27226
rect 86036 27174 86046 27226
rect 86046 27174 86092 27226
rect 86116 27174 86162 27226
rect 86162 27174 86172 27226
rect 86196 27174 86226 27226
rect 86226 27174 86252 27226
rect 85956 27172 86012 27174
rect 86036 27172 86092 27174
rect 86116 27172 86172 27174
rect 86196 27172 86252 27174
rect 86682 99456 86738 99512
rect 86958 148824 87014 148880
rect 86866 134136 86922 134192
rect 86866 99728 86922 99784
rect 86774 95512 86830 95568
rect 87050 146512 87106 146568
rect 86958 97688 87014 97744
rect 86958 96600 87014 96656
rect 87234 149912 87290 149968
rect 87234 122304 87290 122360
rect 87234 118632 87290 118688
rect 87234 118496 87290 118552
rect 87234 109112 87290 109168
rect 87326 108704 87382 108760
rect 87234 108568 87290 108624
rect 87142 104216 87198 104272
rect 87326 104216 87382 104272
rect 87142 99332 87198 99388
rect 87234 97824 87290 97880
rect 87694 171672 87750 171728
rect 87326 96328 87382 96384
rect 86958 95376 87014 95432
rect 89956 177370 90012 177372
rect 90036 177370 90092 177372
rect 90116 177370 90172 177372
rect 90196 177370 90252 177372
rect 89956 177318 89982 177370
rect 89982 177318 90012 177370
rect 90036 177318 90046 177370
rect 90046 177318 90092 177370
rect 90116 177318 90162 177370
rect 90162 177318 90172 177370
rect 90196 177318 90226 177370
rect 90226 177318 90252 177370
rect 89956 177316 90012 177318
rect 90036 177316 90092 177318
rect 90116 177316 90172 177318
rect 90196 177316 90252 177318
rect 87956 176826 88012 176828
rect 88036 176826 88092 176828
rect 88116 176826 88172 176828
rect 88196 176826 88252 176828
rect 87956 176774 87982 176826
rect 87982 176774 88012 176826
rect 88036 176774 88046 176826
rect 88046 176774 88092 176826
rect 88116 176774 88162 176826
rect 88162 176774 88172 176826
rect 88196 176774 88226 176826
rect 88226 176774 88252 176826
rect 87956 176772 88012 176774
rect 88036 176772 88092 176774
rect 88116 176772 88172 176774
rect 88196 176772 88252 176774
rect 89956 176282 90012 176284
rect 90036 176282 90092 176284
rect 90116 176282 90172 176284
rect 90196 176282 90252 176284
rect 89956 176230 89982 176282
rect 89982 176230 90012 176282
rect 90036 176230 90046 176282
rect 90046 176230 90092 176282
rect 90116 176230 90162 176282
rect 90162 176230 90172 176282
rect 90196 176230 90226 176282
rect 90226 176230 90252 176282
rect 89956 176228 90012 176230
rect 90036 176228 90092 176230
rect 90116 176228 90172 176230
rect 90196 176228 90252 176230
rect 87956 175738 88012 175740
rect 88036 175738 88092 175740
rect 88116 175738 88172 175740
rect 88196 175738 88252 175740
rect 87956 175686 87982 175738
rect 87982 175686 88012 175738
rect 88036 175686 88046 175738
rect 88046 175686 88092 175738
rect 88116 175686 88162 175738
rect 88162 175686 88172 175738
rect 88196 175686 88226 175738
rect 88226 175686 88252 175738
rect 87956 175684 88012 175686
rect 88036 175684 88092 175686
rect 88116 175684 88172 175686
rect 88196 175684 88252 175686
rect 89956 175194 90012 175196
rect 90036 175194 90092 175196
rect 90116 175194 90172 175196
rect 90196 175194 90252 175196
rect 89956 175142 89982 175194
rect 89982 175142 90012 175194
rect 90036 175142 90046 175194
rect 90046 175142 90092 175194
rect 90116 175142 90162 175194
rect 90162 175142 90172 175194
rect 90196 175142 90226 175194
rect 90226 175142 90252 175194
rect 89956 175140 90012 175142
rect 90036 175140 90092 175142
rect 90116 175140 90172 175142
rect 90196 175140 90252 175142
rect 87956 174650 88012 174652
rect 88036 174650 88092 174652
rect 88116 174650 88172 174652
rect 88196 174650 88252 174652
rect 87956 174598 87982 174650
rect 87982 174598 88012 174650
rect 88036 174598 88046 174650
rect 88046 174598 88092 174650
rect 88116 174598 88162 174650
rect 88162 174598 88172 174650
rect 88196 174598 88226 174650
rect 88226 174598 88252 174650
rect 87956 174596 88012 174598
rect 88036 174596 88092 174598
rect 88116 174596 88172 174598
rect 88196 174596 88252 174598
rect 89956 174106 90012 174108
rect 90036 174106 90092 174108
rect 90116 174106 90172 174108
rect 90196 174106 90252 174108
rect 89956 174054 89982 174106
rect 89982 174054 90012 174106
rect 90036 174054 90046 174106
rect 90046 174054 90092 174106
rect 90116 174054 90162 174106
rect 90162 174054 90172 174106
rect 90196 174054 90226 174106
rect 90226 174054 90252 174106
rect 89956 174052 90012 174054
rect 90036 174052 90092 174054
rect 90116 174052 90172 174054
rect 90196 174052 90252 174054
rect 87956 173562 88012 173564
rect 88036 173562 88092 173564
rect 88116 173562 88172 173564
rect 88196 173562 88252 173564
rect 87956 173510 87982 173562
rect 87982 173510 88012 173562
rect 88036 173510 88046 173562
rect 88046 173510 88092 173562
rect 88116 173510 88162 173562
rect 88162 173510 88172 173562
rect 88196 173510 88226 173562
rect 88226 173510 88252 173562
rect 87956 173508 88012 173510
rect 88036 173508 88092 173510
rect 88116 173508 88172 173510
rect 88196 173508 88252 173510
rect 89956 173018 90012 173020
rect 90036 173018 90092 173020
rect 90116 173018 90172 173020
rect 90196 173018 90252 173020
rect 89956 172966 89982 173018
rect 89982 172966 90012 173018
rect 90036 172966 90046 173018
rect 90046 172966 90092 173018
rect 90116 172966 90162 173018
rect 90162 172966 90172 173018
rect 90196 172966 90226 173018
rect 90226 172966 90252 173018
rect 89956 172964 90012 172966
rect 90036 172964 90092 172966
rect 90116 172964 90172 172966
rect 90196 172964 90252 172966
rect 87956 172474 88012 172476
rect 88036 172474 88092 172476
rect 88116 172474 88172 172476
rect 88196 172474 88252 172476
rect 87956 172422 87982 172474
rect 87982 172422 88012 172474
rect 88036 172422 88046 172474
rect 88046 172422 88092 172474
rect 88116 172422 88162 172474
rect 88162 172422 88172 172474
rect 88196 172422 88226 172474
rect 88226 172422 88252 172474
rect 87956 172420 88012 172422
rect 88036 172420 88092 172422
rect 88116 172420 88172 172422
rect 88196 172420 88252 172422
rect 89956 171930 90012 171932
rect 90036 171930 90092 171932
rect 90116 171930 90172 171932
rect 90196 171930 90252 171932
rect 89956 171878 89982 171930
rect 89982 171878 90012 171930
rect 90036 171878 90046 171930
rect 90046 171878 90092 171930
rect 90116 171878 90162 171930
rect 90162 171878 90172 171930
rect 90196 171878 90226 171930
rect 90226 171878 90252 171930
rect 89956 171876 90012 171878
rect 90036 171876 90092 171878
rect 90116 171876 90172 171878
rect 90196 171876 90252 171878
rect 87956 171386 88012 171388
rect 88036 171386 88092 171388
rect 88116 171386 88172 171388
rect 88196 171386 88252 171388
rect 87956 171334 87982 171386
rect 87982 171334 88012 171386
rect 88036 171334 88046 171386
rect 88046 171334 88092 171386
rect 88116 171334 88162 171386
rect 88162 171334 88172 171386
rect 88196 171334 88226 171386
rect 88226 171334 88252 171386
rect 87956 171332 88012 171334
rect 88036 171332 88092 171334
rect 88116 171332 88172 171334
rect 88196 171332 88252 171334
rect 89956 170842 90012 170844
rect 90036 170842 90092 170844
rect 90116 170842 90172 170844
rect 90196 170842 90252 170844
rect 89956 170790 89982 170842
rect 89982 170790 90012 170842
rect 90036 170790 90046 170842
rect 90046 170790 90092 170842
rect 90116 170790 90162 170842
rect 90162 170790 90172 170842
rect 90196 170790 90226 170842
rect 90226 170790 90252 170842
rect 89956 170788 90012 170790
rect 90036 170788 90092 170790
rect 90116 170788 90172 170790
rect 90196 170788 90252 170790
rect 87956 170298 88012 170300
rect 88036 170298 88092 170300
rect 88116 170298 88172 170300
rect 88196 170298 88252 170300
rect 87956 170246 87982 170298
rect 87982 170246 88012 170298
rect 88036 170246 88046 170298
rect 88046 170246 88092 170298
rect 88116 170246 88162 170298
rect 88162 170246 88172 170298
rect 88196 170246 88226 170298
rect 88226 170246 88252 170298
rect 87956 170244 88012 170246
rect 88036 170244 88092 170246
rect 88116 170244 88172 170246
rect 88196 170244 88252 170246
rect 89956 169754 90012 169756
rect 90036 169754 90092 169756
rect 90116 169754 90172 169756
rect 90196 169754 90252 169756
rect 89956 169702 89982 169754
rect 89982 169702 90012 169754
rect 90036 169702 90046 169754
rect 90046 169702 90092 169754
rect 90116 169702 90162 169754
rect 90162 169702 90172 169754
rect 90196 169702 90226 169754
rect 90226 169702 90252 169754
rect 89956 169700 90012 169702
rect 90036 169700 90092 169702
rect 90116 169700 90172 169702
rect 90196 169700 90252 169702
rect 87878 169496 87934 169552
rect 87956 169210 88012 169212
rect 88036 169210 88092 169212
rect 88116 169210 88172 169212
rect 88196 169210 88252 169212
rect 87956 169158 87982 169210
rect 87982 169158 88012 169210
rect 88036 169158 88046 169210
rect 88046 169158 88092 169210
rect 88116 169158 88162 169210
rect 88162 169158 88172 169210
rect 88196 169158 88226 169210
rect 88226 169158 88252 169210
rect 87956 169156 88012 169158
rect 88036 169156 88092 169158
rect 88116 169156 88172 169158
rect 88196 169156 88252 169158
rect 89956 168666 90012 168668
rect 90036 168666 90092 168668
rect 90116 168666 90172 168668
rect 90196 168666 90252 168668
rect 89956 168614 89982 168666
rect 89982 168614 90012 168666
rect 90036 168614 90046 168666
rect 90046 168614 90092 168666
rect 90116 168614 90162 168666
rect 90162 168614 90172 168666
rect 90196 168614 90226 168666
rect 90226 168614 90252 168666
rect 89956 168612 90012 168614
rect 90036 168612 90092 168614
rect 90116 168612 90172 168614
rect 90196 168612 90252 168614
rect 87956 168122 88012 168124
rect 88036 168122 88092 168124
rect 88116 168122 88172 168124
rect 88196 168122 88252 168124
rect 87956 168070 87982 168122
rect 87982 168070 88012 168122
rect 88036 168070 88046 168122
rect 88046 168070 88092 168122
rect 88116 168070 88162 168122
rect 88162 168070 88172 168122
rect 88196 168070 88226 168122
rect 88226 168070 88252 168122
rect 87956 168068 88012 168070
rect 88036 168068 88092 168070
rect 88116 168068 88172 168070
rect 88196 168068 88252 168070
rect 89956 167578 90012 167580
rect 90036 167578 90092 167580
rect 90116 167578 90172 167580
rect 90196 167578 90252 167580
rect 89956 167526 89982 167578
rect 89982 167526 90012 167578
rect 90036 167526 90046 167578
rect 90046 167526 90092 167578
rect 90116 167526 90162 167578
rect 90162 167526 90172 167578
rect 90196 167526 90226 167578
rect 90226 167526 90252 167578
rect 89956 167524 90012 167526
rect 90036 167524 90092 167526
rect 90116 167524 90172 167526
rect 90196 167524 90252 167526
rect 87956 167034 88012 167036
rect 88036 167034 88092 167036
rect 88116 167034 88172 167036
rect 88196 167034 88252 167036
rect 87956 166982 87982 167034
rect 87982 166982 88012 167034
rect 88036 166982 88046 167034
rect 88046 166982 88092 167034
rect 88116 166982 88162 167034
rect 88162 166982 88172 167034
rect 88196 166982 88226 167034
rect 88226 166982 88252 167034
rect 87956 166980 88012 166982
rect 88036 166980 88092 166982
rect 88116 166980 88172 166982
rect 88196 166980 88252 166982
rect 89956 166490 90012 166492
rect 90036 166490 90092 166492
rect 90116 166490 90172 166492
rect 90196 166490 90252 166492
rect 89956 166438 89982 166490
rect 89982 166438 90012 166490
rect 90036 166438 90046 166490
rect 90046 166438 90092 166490
rect 90116 166438 90162 166490
rect 90162 166438 90172 166490
rect 90196 166438 90226 166490
rect 90226 166438 90252 166490
rect 89956 166436 90012 166438
rect 90036 166436 90092 166438
rect 90116 166436 90172 166438
rect 90196 166436 90252 166438
rect 87956 165946 88012 165948
rect 88036 165946 88092 165948
rect 88116 165946 88172 165948
rect 88196 165946 88252 165948
rect 87956 165894 87982 165946
rect 87982 165894 88012 165946
rect 88036 165894 88046 165946
rect 88046 165894 88092 165946
rect 88116 165894 88162 165946
rect 88162 165894 88172 165946
rect 88196 165894 88226 165946
rect 88226 165894 88252 165946
rect 87956 165892 88012 165894
rect 88036 165892 88092 165894
rect 88116 165892 88172 165894
rect 88196 165892 88252 165894
rect 89956 165402 90012 165404
rect 90036 165402 90092 165404
rect 90116 165402 90172 165404
rect 90196 165402 90252 165404
rect 89956 165350 89982 165402
rect 89982 165350 90012 165402
rect 90036 165350 90046 165402
rect 90046 165350 90092 165402
rect 90116 165350 90162 165402
rect 90162 165350 90172 165402
rect 90196 165350 90226 165402
rect 90226 165350 90252 165402
rect 89956 165348 90012 165350
rect 90036 165348 90092 165350
rect 90116 165348 90172 165350
rect 90196 165348 90252 165350
rect 87956 164858 88012 164860
rect 88036 164858 88092 164860
rect 88116 164858 88172 164860
rect 88196 164858 88252 164860
rect 87956 164806 87982 164858
rect 87982 164806 88012 164858
rect 88036 164806 88046 164858
rect 88046 164806 88092 164858
rect 88116 164806 88162 164858
rect 88162 164806 88172 164858
rect 88196 164806 88226 164858
rect 88226 164806 88252 164858
rect 87956 164804 88012 164806
rect 88036 164804 88092 164806
rect 88116 164804 88172 164806
rect 88196 164804 88252 164806
rect 87878 164600 87934 164656
rect 89956 164314 90012 164316
rect 90036 164314 90092 164316
rect 90116 164314 90172 164316
rect 90196 164314 90252 164316
rect 89956 164262 89982 164314
rect 89982 164262 90012 164314
rect 90036 164262 90046 164314
rect 90046 164262 90092 164314
rect 90116 164262 90162 164314
rect 90162 164262 90172 164314
rect 90196 164262 90226 164314
rect 90226 164262 90252 164314
rect 89956 164260 90012 164262
rect 90036 164260 90092 164262
rect 90116 164260 90172 164262
rect 90196 164260 90252 164262
rect 87956 163770 88012 163772
rect 88036 163770 88092 163772
rect 88116 163770 88172 163772
rect 88196 163770 88252 163772
rect 87956 163718 87982 163770
rect 87982 163718 88012 163770
rect 88036 163718 88046 163770
rect 88046 163718 88092 163770
rect 88116 163718 88162 163770
rect 88162 163718 88172 163770
rect 88196 163718 88226 163770
rect 88226 163718 88252 163770
rect 87956 163716 88012 163718
rect 88036 163716 88092 163718
rect 88116 163716 88172 163718
rect 88196 163716 88252 163718
rect 87878 163376 87934 163432
rect 89956 163226 90012 163228
rect 90036 163226 90092 163228
rect 90116 163226 90172 163228
rect 90196 163226 90252 163228
rect 89956 163174 89982 163226
rect 89982 163174 90012 163226
rect 90036 163174 90046 163226
rect 90046 163174 90092 163226
rect 90116 163174 90162 163226
rect 90162 163174 90172 163226
rect 90196 163174 90226 163226
rect 90226 163174 90252 163226
rect 89956 163172 90012 163174
rect 90036 163172 90092 163174
rect 90116 163172 90172 163174
rect 90196 163172 90252 163174
rect 87956 162682 88012 162684
rect 88036 162682 88092 162684
rect 88116 162682 88172 162684
rect 88196 162682 88252 162684
rect 87956 162630 87982 162682
rect 87982 162630 88012 162682
rect 88036 162630 88046 162682
rect 88046 162630 88092 162682
rect 88116 162630 88162 162682
rect 88162 162630 88172 162682
rect 88196 162630 88226 162682
rect 88226 162630 88252 162682
rect 87956 162628 88012 162630
rect 88036 162628 88092 162630
rect 88116 162628 88172 162630
rect 88196 162628 88252 162630
rect 89956 162138 90012 162140
rect 90036 162138 90092 162140
rect 90116 162138 90172 162140
rect 90196 162138 90252 162140
rect 89956 162086 89982 162138
rect 89982 162086 90012 162138
rect 90036 162086 90046 162138
rect 90046 162086 90092 162138
rect 90116 162086 90162 162138
rect 90162 162086 90172 162138
rect 90196 162086 90226 162138
rect 90226 162086 90252 162138
rect 89956 162084 90012 162086
rect 90036 162084 90092 162086
rect 90116 162084 90172 162086
rect 90196 162084 90252 162086
rect 87956 161594 88012 161596
rect 88036 161594 88092 161596
rect 88116 161594 88172 161596
rect 88196 161594 88252 161596
rect 87956 161542 87982 161594
rect 87982 161542 88012 161594
rect 88036 161542 88046 161594
rect 88046 161542 88092 161594
rect 88116 161542 88162 161594
rect 88162 161542 88172 161594
rect 88196 161542 88226 161594
rect 88226 161542 88252 161594
rect 87956 161540 88012 161542
rect 88036 161540 88092 161542
rect 88116 161540 88172 161542
rect 88196 161540 88252 161542
rect 89956 161050 90012 161052
rect 90036 161050 90092 161052
rect 90116 161050 90172 161052
rect 90196 161050 90252 161052
rect 89956 160998 89982 161050
rect 89982 160998 90012 161050
rect 90036 160998 90046 161050
rect 90046 160998 90092 161050
rect 90116 160998 90162 161050
rect 90162 160998 90172 161050
rect 90196 160998 90226 161050
rect 90226 160998 90252 161050
rect 89956 160996 90012 160998
rect 90036 160996 90092 160998
rect 90116 160996 90172 160998
rect 90196 160996 90252 160998
rect 87878 160792 87934 160848
rect 87956 160506 88012 160508
rect 88036 160506 88092 160508
rect 88116 160506 88172 160508
rect 88196 160506 88252 160508
rect 87956 160454 87982 160506
rect 87982 160454 88012 160506
rect 88036 160454 88046 160506
rect 88046 160454 88092 160506
rect 88116 160454 88162 160506
rect 88162 160454 88172 160506
rect 88196 160454 88226 160506
rect 88226 160454 88252 160506
rect 87956 160452 88012 160454
rect 88036 160452 88092 160454
rect 88116 160452 88172 160454
rect 88196 160452 88252 160454
rect 89956 159962 90012 159964
rect 90036 159962 90092 159964
rect 90116 159962 90172 159964
rect 90196 159962 90252 159964
rect 89956 159910 89982 159962
rect 89982 159910 90012 159962
rect 90036 159910 90046 159962
rect 90046 159910 90092 159962
rect 90116 159910 90162 159962
rect 90162 159910 90172 159962
rect 90196 159910 90226 159962
rect 90226 159910 90252 159962
rect 89956 159908 90012 159910
rect 90036 159908 90092 159910
rect 90116 159908 90172 159910
rect 90196 159908 90252 159910
rect 87956 159418 88012 159420
rect 88036 159418 88092 159420
rect 88116 159418 88172 159420
rect 88196 159418 88252 159420
rect 87956 159366 87982 159418
rect 87982 159366 88012 159418
rect 88036 159366 88046 159418
rect 88046 159366 88092 159418
rect 88116 159366 88162 159418
rect 88162 159366 88172 159418
rect 88196 159366 88226 159418
rect 88226 159366 88252 159418
rect 87956 159364 88012 159366
rect 88036 159364 88092 159366
rect 88116 159364 88172 159366
rect 88196 159364 88252 159366
rect 89956 158874 90012 158876
rect 90036 158874 90092 158876
rect 90116 158874 90172 158876
rect 90196 158874 90252 158876
rect 89956 158822 89982 158874
rect 89982 158822 90012 158874
rect 90036 158822 90046 158874
rect 90046 158822 90092 158874
rect 90116 158822 90162 158874
rect 90162 158822 90172 158874
rect 90196 158822 90226 158874
rect 90226 158822 90252 158874
rect 89956 158820 90012 158822
rect 90036 158820 90092 158822
rect 90116 158820 90172 158822
rect 90196 158820 90252 158822
rect 87956 158330 88012 158332
rect 88036 158330 88092 158332
rect 88116 158330 88172 158332
rect 88196 158330 88252 158332
rect 87956 158278 87982 158330
rect 87982 158278 88012 158330
rect 88036 158278 88046 158330
rect 88046 158278 88092 158330
rect 88116 158278 88162 158330
rect 88162 158278 88172 158330
rect 88196 158278 88226 158330
rect 88226 158278 88252 158330
rect 87956 158276 88012 158278
rect 88036 158276 88092 158278
rect 88116 158276 88172 158278
rect 88196 158276 88252 158278
rect 89956 157786 90012 157788
rect 90036 157786 90092 157788
rect 90116 157786 90172 157788
rect 90196 157786 90252 157788
rect 89956 157734 89982 157786
rect 89982 157734 90012 157786
rect 90036 157734 90046 157786
rect 90046 157734 90092 157786
rect 90116 157734 90162 157786
rect 90162 157734 90172 157786
rect 90196 157734 90226 157786
rect 90226 157734 90252 157786
rect 89956 157732 90012 157734
rect 90036 157732 90092 157734
rect 90116 157732 90172 157734
rect 90196 157732 90252 157734
rect 87956 157242 88012 157244
rect 88036 157242 88092 157244
rect 88116 157242 88172 157244
rect 88196 157242 88252 157244
rect 87956 157190 87982 157242
rect 87982 157190 88012 157242
rect 88036 157190 88046 157242
rect 88046 157190 88092 157242
rect 88116 157190 88162 157242
rect 88162 157190 88172 157242
rect 88196 157190 88226 157242
rect 88226 157190 88252 157242
rect 87956 157188 88012 157190
rect 88036 157188 88092 157190
rect 88116 157188 88172 157190
rect 88196 157188 88252 157190
rect 89956 156698 90012 156700
rect 90036 156698 90092 156700
rect 90116 156698 90172 156700
rect 90196 156698 90252 156700
rect 89956 156646 89982 156698
rect 89982 156646 90012 156698
rect 90036 156646 90046 156698
rect 90046 156646 90092 156698
rect 90116 156646 90162 156698
rect 90162 156646 90172 156698
rect 90196 156646 90226 156698
rect 90226 156646 90252 156698
rect 89956 156644 90012 156646
rect 90036 156644 90092 156646
rect 90116 156644 90172 156646
rect 90196 156644 90252 156646
rect 87956 156154 88012 156156
rect 88036 156154 88092 156156
rect 88116 156154 88172 156156
rect 88196 156154 88252 156156
rect 87956 156102 87982 156154
rect 87982 156102 88012 156154
rect 88036 156102 88046 156154
rect 88046 156102 88092 156154
rect 88116 156102 88162 156154
rect 88162 156102 88172 156154
rect 88196 156102 88226 156154
rect 88226 156102 88252 156154
rect 87956 156100 88012 156102
rect 88036 156100 88092 156102
rect 88116 156100 88172 156102
rect 88196 156100 88252 156102
rect 89956 155610 90012 155612
rect 90036 155610 90092 155612
rect 90116 155610 90172 155612
rect 90196 155610 90252 155612
rect 89956 155558 89982 155610
rect 89982 155558 90012 155610
rect 90036 155558 90046 155610
rect 90046 155558 90092 155610
rect 90116 155558 90162 155610
rect 90162 155558 90172 155610
rect 90196 155558 90226 155610
rect 90226 155558 90252 155610
rect 89956 155556 90012 155558
rect 90036 155556 90092 155558
rect 90116 155556 90172 155558
rect 90196 155556 90252 155558
rect 87956 155066 88012 155068
rect 88036 155066 88092 155068
rect 88116 155066 88172 155068
rect 88196 155066 88252 155068
rect 87956 155014 87982 155066
rect 87982 155014 88012 155066
rect 88036 155014 88046 155066
rect 88046 155014 88092 155066
rect 88116 155014 88162 155066
rect 88162 155014 88172 155066
rect 88196 155014 88226 155066
rect 88226 155014 88252 155066
rect 87956 155012 88012 155014
rect 88036 155012 88092 155014
rect 88116 155012 88172 155014
rect 88196 155012 88252 155014
rect 89956 154522 90012 154524
rect 90036 154522 90092 154524
rect 90116 154522 90172 154524
rect 90196 154522 90252 154524
rect 89956 154470 89982 154522
rect 89982 154470 90012 154522
rect 90036 154470 90046 154522
rect 90046 154470 90092 154522
rect 90116 154470 90162 154522
rect 90162 154470 90172 154522
rect 90196 154470 90226 154522
rect 90226 154470 90252 154522
rect 89956 154468 90012 154470
rect 90036 154468 90092 154470
rect 90116 154468 90172 154470
rect 90196 154468 90252 154470
rect 87956 153978 88012 153980
rect 88036 153978 88092 153980
rect 88116 153978 88172 153980
rect 88196 153978 88252 153980
rect 87956 153926 87982 153978
rect 87982 153926 88012 153978
rect 88036 153926 88046 153978
rect 88046 153926 88092 153978
rect 88116 153926 88162 153978
rect 88162 153926 88172 153978
rect 88196 153926 88226 153978
rect 88226 153926 88252 153978
rect 87956 153924 88012 153926
rect 88036 153924 88092 153926
rect 88116 153924 88172 153926
rect 88196 153924 88252 153926
rect 89956 153434 90012 153436
rect 90036 153434 90092 153436
rect 90116 153434 90172 153436
rect 90196 153434 90252 153436
rect 89956 153382 89982 153434
rect 89982 153382 90012 153434
rect 90036 153382 90046 153434
rect 90046 153382 90092 153434
rect 90116 153382 90162 153434
rect 90162 153382 90172 153434
rect 90196 153382 90226 153434
rect 90226 153382 90252 153434
rect 89956 153380 90012 153382
rect 90036 153380 90092 153382
rect 90116 153380 90172 153382
rect 90196 153380 90252 153382
rect 87956 152890 88012 152892
rect 88036 152890 88092 152892
rect 88116 152890 88172 152892
rect 88196 152890 88252 152892
rect 87956 152838 87982 152890
rect 87982 152838 88012 152890
rect 88036 152838 88046 152890
rect 88046 152838 88092 152890
rect 88116 152838 88162 152890
rect 88162 152838 88172 152890
rect 88196 152838 88226 152890
rect 88226 152838 88252 152890
rect 87956 152836 88012 152838
rect 88036 152836 88092 152838
rect 88116 152836 88172 152838
rect 88196 152836 88252 152838
rect 89956 152346 90012 152348
rect 90036 152346 90092 152348
rect 90116 152346 90172 152348
rect 90196 152346 90252 152348
rect 89956 152294 89982 152346
rect 89982 152294 90012 152346
rect 90036 152294 90046 152346
rect 90046 152294 90092 152346
rect 90116 152294 90162 152346
rect 90162 152294 90172 152346
rect 90196 152294 90226 152346
rect 90226 152294 90252 152346
rect 89956 152292 90012 152294
rect 90036 152292 90092 152294
rect 90116 152292 90172 152294
rect 90196 152292 90252 152294
rect 87956 151802 88012 151804
rect 88036 151802 88092 151804
rect 88116 151802 88172 151804
rect 88196 151802 88252 151804
rect 87956 151750 87982 151802
rect 87982 151750 88012 151802
rect 88036 151750 88046 151802
rect 88046 151750 88092 151802
rect 88116 151750 88162 151802
rect 88162 151750 88172 151802
rect 88196 151750 88226 151802
rect 88226 151750 88252 151802
rect 87956 151748 88012 151750
rect 88036 151748 88092 151750
rect 88116 151748 88172 151750
rect 88196 151748 88252 151750
rect 89956 151258 90012 151260
rect 90036 151258 90092 151260
rect 90116 151258 90172 151260
rect 90196 151258 90252 151260
rect 89956 151206 89982 151258
rect 89982 151206 90012 151258
rect 90036 151206 90046 151258
rect 90046 151206 90092 151258
rect 90116 151206 90162 151258
rect 90162 151206 90172 151258
rect 90196 151206 90226 151258
rect 90226 151206 90252 151258
rect 89956 151204 90012 151206
rect 90036 151204 90092 151206
rect 90116 151204 90172 151206
rect 90196 151204 90252 151206
rect 87956 150714 88012 150716
rect 88036 150714 88092 150716
rect 88116 150714 88172 150716
rect 88196 150714 88252 150716
rect 87956 150662 87982 150714
rect 87982 150662 88012 150714
rect 88036 150662 88046 150714
rect 88046 150662 88092 150714
rect 88116 150662 88162 150714
rect 88162 150662 88172 150714
rect 88196 150662 88226 150714
rect 88226 150662 88252 150714
rect 87956 150660 88012 150662
rect 88036 150660 88092 150662
rect 88116 150660 88172 150662
rect 88196 150660 88252 150662
rect 89956 150170 90012 150172
rect 90036 150170 90092 150172
rect 90116 150170 90172 150172
rect 90196 150170 90252 150172
rect 89956 150118 89982 150170
rect 89982 150118 90012 150170
rect 90036 150118 90046 150170
rect 90046 150118 90092 150170
rect 90116 150118 90162 150170
rect 90162 150118 90172 150170
rect 90196 150118 90226 150170
rect 90226 150118 90252 150170
rect 89956 150116 90012 150118
rect 90036 150116 90092 150118
rect 90116 150116 90172 150118
rect 90196 150116 90252 150118
rect 87956 149626 88012 149628
rect 88036 149626 88092 149628
rect 88116 149626 88172 149628
rect 88196 149626 88252 149628
rect 87956 149574 87982 149626
rect 87982 149574 88012 149626
rect 88036 149574 88046 149626
rect 88046 149574 88092 149626
rect 88116 149574 88162 149626
rect 88162 149574 88172 149626
rect 88196 149574 88226 149626
rect 88226 149574 88252 149626
rect 87956 149572 88012 149574
rect 88036 149572 88092 149574
rect 88116 149572 88172 149574
rect 88196 149572 88252 149574
rect 89956 149082 90012 149084
rect 90036 149082 90092 149084
rect 90116 149082 90172 149084
rect 90196 149082 90252 149084
rect 89956 149030 89982 149082
rect 89982 149030 90012 149082
rect 90036 149030 90046 149082
rect 90046 149030 90092 149082
rect 90116 149030 90162 149082
rect 90162 149030 90172 149082
rect 90196 149030 90226 149082
rect 90226 149030 90252 149082
rect 89956 149028 90012 149030
rect 90036 149028 90092 149030
rect 90116 149028 90172 149030
rect 90196 149028 90252 149030
rect 87956 148538 88012 148540
rect 88036 148538 88092 148540
rect 88116 148538 88172 148540
rect 88196 148538 88252 148540
rect 87956 148486 87982 148538
rect 87982 148486 88012 148538
rect 88036 148486 88046 148538
rect 88046 148486 88092 148538
rect 88116 148486 88162 148538
rect 88162 148486 88172 148538
rect 88196 148486 88226 148538
rect 88226 148486 88252 148538
rect 87956 148484 88012 148486
rect 88036 148484 88092 148486
rect 88116 148484 88172 148486
rect 88196 148484 88252 148486
rect 89956 147994 90012 147996
rect 90036 147994 90092 147996
rect 90116 147994 90172 147996
rect 90196 147994 90252 147996
rect 89956 147942 89982 147994
rect 89982 147942 90012 147994
rect 90036 147942 90046 147994
rect 90046 147942 90092 147994
rect 90116 147942 90162 147994
rect 90162 147942 90172 147994
rect 90196 147942 90226 147994
rect 90226 147942 90252 147994
rect 89956 147940 90012 147942
rect 90036 147940 90092 147942
rect 90116 147940 90172 147942
rect 90196 147940 90252 147942
rect 87956 147450 88012 147452
rect 88036 147450 88092 147452
rect 88116 147450 88172 147452
rect 88196 147450 88252 147452
rect 87956 147398 87982 147450
rect 87982 147398 88012 147450
rect 88036 147398 88046 147450
rect 88046 147398 88092 147450
rect 88116 147398 88162 147450
rect 88162 147398 88172 147450
rect 88196 147398 88226 147450
rect 88226 147398 88252 147450
rect 87956 147396 88012 147398
rect 88036 147396 88092 147398
rect 88116 147396 88172 147398
rect 88196 147396 88252 147398
rect 89956 146906 90012 146908
rect 90036 146906 90092 146908
rect 90116 146906 90172 146908
rect 90196 146906 90252 146908
rect 89956 146854 89982 146906
rect 89982 146854 90012 146906
rect 90036 146854 90046 146906
rect 90046 146854 90092 146906
rect 90116 146854 90162 146906
rect 90162 146854 90172 146906
rect 90196 146854 90226 146906
rect 90226 146854 90252 146906
rect 89956 146852 90012 146854
rect 90036 146852 90092 146854
rect 90116 146852 90172 146854
rect 90196 146852 90252 146854
rect 87956 146362 88012 146364
rect 88036 146362 88092 146364
rect 88116 146362 88172 146364
rect 88196 146362 88252 146364
rect 87956 146310 87982 146362
rect 87982 146310 88012 146362
rect 88036 146310 88046 146362
rect 88046 146310 88092 146362
rect 88116 146310 88162 146362
rect 88162 146310 88172 146362
rect 88196 146310 88226 146362
rect 88226 146310 88252 146362
rect 87956 146308 88012 146310
rect 88036 146308 88092 146310
rect 88116 146308 88172 146310
rect 88196 146308 88252 146310
rect 89956 145818 90012 145820
rect 90036 145818 90092 145820
rect 90116 145818 90172 145820
rect 90196 145818 90252 145820
rect 89956 145766 89982 145818
rect 89982 145766 90012 145818
rect 90036 145766 90046 145818
rect 90046 145766 90092 145818
rect 90116 145766 90162 145818
rect 90162 145766 90172 145818
rect 90196 145766 90226 145818
rect 90226 145766 90252 145818
rect 89956 145764 90012 145766
rect 90036 145764 90092 145766
rect 90116 145764 90172 145766
rect 90196 145764 90252 145766
rect 87956 145274 88012 145276
rect 88036 145274 88092 145276
rect 88116 145274 88172 145276
rect 88196 145274 88252 145276
rect 87956 145222 87982 145274
rect 87982 145222 88012 145274
rect 88036 145222 88046 145274
rect 88046 145222 88092 145274
rect 88116 145222 88162 145274
rect 88162 145222 88172 145274
rect 88196 145222 88226 145274
rect 88226 145222 88252 145274
rect 87956 145220 88012 145222
rect 88036 145220 88092 145222
rect 88116 145220 88172 145222
rect 88196 145220 88252 145222
rect 87970 145016 88026 145072
rect 89956 144730 90012 144732
rect 90036 144730 90092 144732
rect 90116 144730 90172 144732
rect 90196 144730 90252 144732
rect 89956 144678 89982 144730
rect 89982 144678 90012 144730
rect 90036 144678 90046 144730
rect 90046 144678 90092 144730
rect 90116 144678 90162 144730
rect 90162 144678 90172 144730
rect 90196 144678 90226 144730
rect 90226 144678 90252 144730
rect 89956 144676 90012 144678
rect 90036 144676 90092 144678
rect 90116 144676 90172 144678
rect 90196 144676 90252 144678
rect 87956 144186 88012 144188
rect 88036 144186 88092 144188
rect 88116 144186 88172 144188
rect 88196 144186 88252 144188
rect 87956 144134 87982 144186
rect 87982 144134 88012 144186
rect 88036 144134 88046 144186
rect 88046 144134 88092 144186
rect 88116 144134 88162 144186
rect 88162 144134 88172 144186
rect 88196 144134 88226 144186
rect 88226 144134 88252 144186
rect 87956 144132 88012 144134
rect 88036 144132 88092 144134
rect 88116 144132 88172 144134
rect 88196 144132 88252 144134
rect 88062 143928 88118 143984
rect 89956 143642 90012 143644
rect 90036 143642 90092 143644
rect 90116 143642 90172 143644
rect 90196 143642 90252 143644
rect 89956 143590 89982 143642
rect 89982 143590 90012 143642
rect 90036 143590 90046 143642
rect 90046 143590 90092 143642
rect 90116 143590 90162 143642
rect 90162 143590 90172 143642
rect 90196 143590 90226 143642
rect 90226 143590 90252 143642
rect 89956 143588 90012 143590
rect 90036 143588 90092 143590
rect 90116 143588 90172 143590
rect 90196 143588 90252 143590
rect 87956 143098 88012 143100
rect 88036 143098 88092 143100
rect 88116 143098 88172 143100
rect 88196 143098 88252 143100
rect 87956 143046 87982 143098
rect 87982 143046 88012 143098
rect 88036 143046 88046 143098
rect 88046 143046 88092 143098
rect 88116 143046 88162 143098
rect 88162 143046 88172 143098
rect 88196 143046 88226 143098
rect 88226 143046 88252 143098
rect 87956 143044 88012 143046
rect 88036 143044 88092 143046
rect 88116 143044 88172 143046
rect 88196 143044 88252 143046
rect 87970 142704 88026 142760
rect 89956 142554 90012 142556
rect 90036 142554 90092 142556
rect 90116 142554 90172 142556
rect 90196 142554 90252 142556
rect 89956 142502 89982 142554
rect 89982 142502 90012 142554
rect 90036 142502 90046 142554
rect 90046 142502 90092 142554
rect 90116 142502 90162 142554
rect 90162 142502 90172 142554
rect 90196 142502 90226 142554
rect 90226 142502 90252 142554
rect 89956 142500 90012 142502
rect 90036 142500 90092 142502
rect 90116 142500 90172 142502
rect 90196 142500 90252 142502
rect 87956 142010 88012 142012
rect 88036 142010 88092 142012
rect 88116 142010 88172 142012
rect 88196 142010 88252 142012
rect 87956 141958 87982 142010
rect 87982 141958 88012 142010
rect 88036 141958 88046 142010
rect 88046 141958 88092 142010
rect 88116 141958 88162 142010
rect 88162 141958 88172 142010
rect 88196 141958 88226 142010
rect 88226 141958 88252 142010
rect 87956 141956 88012 141958
rect 88036 141956 88092 141958
rect 88116 141956 88172 141958
rect 88196 141956 88252 141958
rect 89956 141466 90012 141468
rect 90036 141466 90092 141468
rect 90116 141466 90172 141468
rect 90196 141466 90252 141468
rect 89956 141414 89982 141466
rect 89982 141414 90012 141466
rect 90036 141414 90046 141466
rect 90046 141414 90092 141466
rect 90116 141414 90162 141466
rect 90162 141414 90172 141466
rect 90196 141414 90226 141466
rect 90226 141414 90252 141466
rect 89956 141412 90012 141414
rect 90036 141412 90092 141414
rect 90116 141412 90172 141414
rect 90196 141412 90252 141414
rect 87970 141228 88026 141264
rect 87970 141208 87972 141228
rect 87972 141208 88024 141228
rect 88024 141208 88026 141228
rect 87956 140922 88012 140924
rect 88036 140922 88092 140924
rect 88116 140922 88172 140924
rect 88196 140922 88252 140924
rect 87956 140870 87982 140922
rect 87982 140870 88012 140922
rect 88036 140870 88046 140922
rect 88046 140870 88092 140922
rect 88116 140870 88162 140922
rect 88162 140870 88172 140922
rect 88196 140870 88226 140922
rect 88226 140870 88252 140922
rect 87956 140868 88012 140870
rect 88036 140868 88092 140870
rect 88116 140868 88172 140870
rect 88196 140868 88252 140870
rect 89956 140378 90012 140380
rect 90036 140378 90092 140380
rect 90116 140378 90172 140380
rect 90196 140378 90252 140380
rect 89956 140326 89982 140378
rect 89982 140326 90012 140378
rect 90036 140326 90046 140378
rect 90046 140326 90092 140378
rect 90116 140326 90162 140378
rect 90162 140326 90172 140378
rect 90196 140326 90226 140378
rect 90226 140326 90252 140378
rect 89956 140324 90012 140326
rect 90036 140324 90092 140326
rect 90116 140324 90172 140326
rect 90196 140324 90252 140326
rect 88246 140120 88302 140176
rect 87956 139834 88012 139836
rect 88036 139834 88092 139836
rect 88116 139834 88172 139836
rect 88196 139834 88252 139836
rect 87956 139782 87982 139834
rect 87982 139782 88012 139834
rect 88036 139782 88046 139834
rect 88046 139782 88092 139834
rect 88116 139782 88162 139834
rect 88162 139782 88172 139834
rect 88196 139782 88226 139834
rect 88226 139782 88252 139834
rect 87956 139780 88012 139782
rect 88036 139780 88092 139782
rect 88116 139780 88172 139782
rect 88196 139780 88252 139782
rect 89956 139290 90012 139292
rect 90036 139290 90092 139292
rect 90116 139290 90172 139292
rect 90196 139290 90252 139292
rect 89956 139238 89982 139290
rect 89982 139238 90012 139290
rect 90036 139238 90046 139290
rect 90046 139238 90092 139290
rect 90116 139238 90162 139290
rect 90162 139238 90172 139290
rect 90196 139238 90226 139290
rect 90226 139238 90252 139290
rect 89956 139236 90012 139238
rect 90036 139236 90092 139238
rect 90116 139236 90172 139238
rect 90196 139236 90252 139238
rect 88062 139032 88118 139088
rect 87956 138746 88012 138748
rect 88036 138746 88092 138748
rect 88116 138746 88172 138748
rect 88196 138746 88252 138748
rect 87956 138694 87982 138746
rect 87982 138694 88012 138746
rect 88036 138694 88046 138746
rect 88046 138694 88092 138746
rect 88116 138694 88162 138746
rect 88162 138694 88172 138746
rect 88196 138694 88226 138746
rect 88226 138694 88252 138746
rect 87956 138692 88012 138694
rect 88036 138692 88092 138694
rect 88116 138692 88172 138694
rect 88196 138692 88252 138694
rect 89956 138202 90012 138204
rect 90036 138202 90092 138204
rect 90116 138202 90172 138204
rect 90196 138202 90252 138204
rect 89956 138150 89982 138202
rect 89982 138150 90012 138202
rect 90036 138150 90046 138202
rect 90046 138150 90092 138202
rect 90116 138150 90162 138202
rect 90162 138150 90172 138202
rect 90196 138150 90226 138202
rect 90226 138150 90252 138202
rect 89956 138148 90012 138150
rect 90036 138148 90092 138150
rect 90116 138148 90172 138150
rect 90196 138148 90252 138150
rect 87956 137658 88012 137660
rect 88036 137658 88092 137660
rect 88116 137658 88172 137660
rect 88196 137658 88252 137660
rect 87956 137606 87982 137658
rect 87982 137606 88012 137658
rect 88036 137606 88046 137658
rect 88046 137606 88092 137658
rect 88116 137606 88162 137658
rect 88162 137606 88172 137658
rect 88196 137606 88226 137658
rect 88226 137606 88252 137658
rect 87956 137604 88012 137606
rect 88036 137604 88092 137606
rect 88116 137604 88172 137606
rect 88196 137604 88252 137606
rect 89956 137114 90012 137116
rect 90036 137114 90092 137116
rect 90116 137114 90172 137116
rect 90196 137114 90252 137116
rect 89956 137062 89982 137114
rect 89982 137062 90012 137114
rect 90036 137062 90046 137114
rect 90046 137062 90092 137114
rect 90116 137062 90162 137114
rect 90162 137062 90172 137114
rect 90196 137062 90226 137114
rect 90226 137062 90252 137114
rect 89956 137060 90012 137062
rect 90036 137060 90092 137062
rect 90116 137060 90172 137062
rect 90196 137060 90252 137062
rect 87956 136570 88012 136572
rect 88036 136570 88092 136572
rect 88116 136570 88172 136572
rect 88196 136570 88252 136572
rect 87956 136518 87982 136570
rect 87982 136518 88012 136570
rect 88036 136518 88046 136570
rect 88046 136518 88092 136570
rect 88116 136518 88162 136570
rect 88162 136518 88172 136570
rect 88196 136518 88226 136570
rect 88226 136518 88252 136570
rect 87956 136516 88012 136518
rect 88036 136516 88092 136518
rect 88116 136516 88172 136518
rect 88196 136516 88252 136518
rect 89956 136026 90012 136028
rect 90036 136026 90092 136028
rect 90116 136026 90172 136028
rect 90196 136026 90252 136028
rect 89956 135974 89982 136026
rect 89982 135974 90012 136026
rect 90036 135974 90046 136026
rect 90046 135974 90092 136026
rect 90116 135974 90162 136026
rect 90162 135974 90172 136026
rect 90196 135974 90226 136026
rect 90226 135974 90252 136026
rect 89956 135972 90012 135974
rect 90036 135972 90092 135974
rect 90116 135972 90172 135974
rect 90196 135972 90252 135974
rect 87956 135482 88012 135484
rect 88036 135482 88092 135484
rect 88116 135482 88172 135484
rect 88196 135482 88252 135484
rect 87956 135430 87982 135482
rect 87982 135430 88012 135482
rect 88036 135430 88046 135482
rect 88046 135430 88092 135482
rect 88116 135430 88162 135482
rect 88162 135430 88172 135482
rect 88196 135430 88226 135482
rect 88226 135430 88252 135482
rect 87956 135428 88012 135430
rect 88036 135428 88092 135430
rect 88116 135428 88172 135430
rect 88196 135428 88252 135430
rect 89956 134938 90012 134940
rect 90036 134938 90092 134940
rect 90116 134938 90172 134940
rect 90196 134938 90252 134940
rect 89956 134886 89982 134938
rect 89982 134886 90012 134938
rect 90036 134886 90046 134938
rect 90046 134886 90092 134938
rect 90116 134886 90162 134938
rect 90162 134886 90172 134938
rect 90196 134886 90226 134938
rect 90226 134886 90252 134938
rect 89956 134884 90012 134886
rect 90036 134884 90092 134886
rect 90116 134884 90172 134886
rect 90196 134884 90252 134886
rect 87956 134394 88012 134396
rect 88036 134394 88092 134396
rect 88116 134394 88172 134396
rect 88196 134394 88252 134396
rect 87956 134342 87982 134394
rect 87982 134342 88012 134394
rect 88036 134342 88046 134394
rect 88046 134342 88092 134394
rect 88116 134342 88162 134394
rect 88162 134342 88172 134394
rect 88196 134342 88226 134394
rect 88226 134342 88252 134394
rect 87956 134340 88012 134342
rect 88036 134340 88092 134342
rect 88116 134340 88172 134342
rect 88196 134340 88252 134342
rect 89956 133850 90012 133852
rect 90036 133850 90092 133852
rect 90116 133850 90172 133852
rect 90196 133850 90252 133852
rect 89956 133798 89982 133850
rect 89982 133798 90012 133850
rect 90036 133798 90046 133850
rect 90046 133798 90092 133850
rect 90116 133798 90162 133850
rect 90162 133798 90172 133850
rect 90196 133798 90226 133850
rect 90226 133798 90252 133850
rect 89956 133796 90012 133798
rect 90036 133796 90092 133798
rect 90116 133796 90172 133798
rect 90196 133796 90252 133798
rect 87956 133306 88012 133308
rect 88036 133306 88092 133308
rect 88116 133306 88172 133308
rect 88196 133306 88252 133308
rect 87956 133254 87982 133306
rect 87982 133254 88012 133306
rect 88036 133254 88046 133306
rect 88046 133254 88092 133306
rect 88116 133254 88162 133306
rect 88162 133254 88172 133306
rect 88196 133254 88226 133306
rect 88226 133254 88252 133306
rect 87956 133252 88012 133254
rect 88036 133252 88092 133254
rect 88116 133252 88172 133254
rect 88196 133252 88252 133254
rect 89956 132762 90012 132764
rect 90036 132762 90092 132764
rect 90116 132762 90172 132764
rect 90196 132762 90252 132764
rect 89956 132710 89982 132762
rect 89982 132710 90012 132762
rect 90036 132710 90046 132762
rect 90046 132710 90092 132762
rect 90116 132710 90162 132762
rect 90162 132710 90172 132762
rect 90196 132710 90226 132762
rect 90226 132710 90252 132762
rect 89956 132708 90012 132710
rect 90036 132708 90092 132710
rect 90116 132708 90172 132710
rect 90196 132708 90252 132710
rect 87956 132218 88012 132220
rect 88036 132218 88092 132220
rect 88116 132218 88172 132220
rect 88196 132218 88252 132220
rect 87956 132166 87982 132218
rect 87982 132166 88012 132218
rect 88036 132166 88046 132218
rect 88046 132166 88092 132218
rect 88116 132166 88162 132218
rect 88162 132166 88172 132218
rect 88196 132166 88226 132218
rect 88226 132166 88252 132218
rect 87956 132164 88012 132166
rect 88036 132164 88092 132166
rect 88116 132164 88172 132166
rect 88196 132164 88252 132166
rect 88246 131824 88302 131880
rect 89956 131674 90012 131676
rect 90036 131674 90092 131676
rect 90116 131674 90172 131676
rect 90196 131674 90252 131676
rect 89956 131622 89982 131674
rect 89982 131622 90012 131674
rect 90036 131622 90046 131674
rect 90046 131622 90092 131674
rect 90116 131622 90162 131674
rect 90162 131622 90172 131674
rect 90196 131622 90226 131674
rect 90226 131622 90252 131674
rect 89956 131620 90012 131622
rect 90036 131620 90092 131622
rect 90116 131620 90172 131622
rect 90196 131620 90252 131622
rect 87956 131130 88012 131132
rect 88036 131130 88092 131132
rect 88116 131130 88172 131132
rect 88196 131130 88252 131132
rect 87956 131078 87982 131130
rect 87982 131078 88012 131130
rect 88036 131078 88046 131130
rect 88046 131078 88092 131130
rect 88116 131078 88162 131130
rect 88162 131078 88172 131130
rect 88196 131078 88226 131130
rect 88226 131078 88252 131130
rect 87956 131076 88012 131078
rect 88036 131076 88092 131078
rect 88116 131076 88172 131078
rect 88196 131076 88252 131078
rect 89956 130586 90012 130588
rect 90036 130586 90092 130588
rect 90116 130586 90172 130588
rect 90196 130586 90252 130588
rect 89956 130534 89982 130586
rect 89982 130534 90012 130586
rect 90036 130534 90046 130586
rect 90046 130534 90092 130586
rect 90116 130534 90162 130586
rect 90162 130534 90172 130586
rect 90196 130534 90226 130586
rect 90226 130534 90252 130586
rect 89956 130532 90012 130534
rect 90036 130532 90092 130534
rect 90116 130532 90172 130534
rect 90196 130532 90252 130534
rect 87956 130042 88012 130044
rect 88036 130042 88092 130044
rect 88116 130042 88172 130044
rect 88196 130042 88252 130044
rect 87956 129990 87982 130042
rect 87982 129990 88012 130042
rect 88036 129990 88046 130042
rect 88046 129990 88092 130042
rect 88116 129990 88162 130042
rect 88162 129990 88172 130042
rect 88196 129990 88226 130042
rect 88226 129990 88252 130042
rect 87956 129988 88012 129990
rect 88036 129988 88092 129990
rect 88116 129988 88172 129990
rect 88196 129988 88252 129990
rect 89956 129498 90012 129500
rect 90036 129498 90092 129500
rect 90116 129498 90172 129500
rect 90196 129498 90252 129500
rect 89956 129446 89982 129498
rect 89982 129446 90012 129498
rect 90036 129446 90046 129498
rect 90046 129446 90092 129498
rect 90116 129446 90162 129498
rect 90162 129446 90172 129498
rect 90196 129446 90226 129498
rect 90226 129446 90252 129498
rect 89956 129444 90012 129446
rect 90036 129444 90092 129446
rect 90116 129444 90172 129446
rect 90196 129444 90252 129446
rect 88246 129240 88302 129296
rect 87956 128954 88012 128956
rect 88036 128954 88092 128956
rect 88116 128954 88172 128956
rect 88196 128954 88252 128956
rect 87956 128902 87982 128954
rect 87982 128902 88012 128954
rect 88036 128902 88046 128954
rect 88046 128902 88092 128954
rect 88116 128902 88162 128954
rect 88162 128902 88172 128954
rect 88196 128902 88226 128954
rect 88226 128902 88252 128954
rect 87956 128900 88012 128902
rect 88036 128900 88092 128902
rect 88116 128900 88172 128902
rect 88196 128900 88252 128902
rect 89956 128410 90012 128412
rect 90036 128410 90092 128412
rect 90116 128410 90172 128412
rect 90196 128410 90252 128412
rect 89956 128358 89982 128410
rect 89982 128358 90012 128410
rect 90036 128358 90046 128410
rect 90046 128358 90092 128410
rect 90116 128358 90162 128410
rect 90162 128358 90172 128410
rect 90196 128358 90226 128410
rect 90226 128358 90252 128410
rect 89956 128356 90012 128358
rect 90036 128356 90092 128358
rect 90116 128356 90172 128358
rect 90196 128356 90252 128358
rect 88246 128152 88302 128208
rect 87956 127866 88012 127868
rect 88036 127866 88092 127868
rect 88116 127866 88172 127868
rect 88196 127866 88252 127868
rect 87956 127814 87982 127866
rect 87982 127814 88012 127866
rect 88036 127814 88046 127866
rect 88046 127814 88092 127866
rect 88116 127814 88162 127866
rect 88162 127814 88172 127866
rect 88196 127814 88226 127866
rect 88226 127814 88252 127866
rect 87956 127812 88012 127814
rect 88036 127812 88092 127814
rect 88116 127812 88172 127814
rect 88196 127812 88252 127814
rect 89956 127322 90012 127324
rect 90036 127322 90092 127324
rect 90116 127322 90172 127324
rect 90196 127322 90252 127324
rect 89956 127270 89982 127322
rect 89982 127270 90012 127322
rect 90036 127270 90046 127322
rect 90046 127270 90092 127322
rect 90116 127270 90162 127322
rect 90162 127270 90172 127322
rect 90196 127270 90226 127322
rect 90226 127270 90252 127322
rect 89956 127268 90012 127270
rect 90036 127268 90092 127270
rect 90116 127268 90172 127270
rect 90196 127268 90252 127270
rect 87956 126778 88012 126780
rect 88036 126778 88092 126780
rect 88116 126778 88172 126780
rect 88196 126778 88252 126780
rect 87956 126726 87982 126778
rect 87982 126726 88012 126778
rect 88036 126726 88046 126778
rect 88046 126726 88092 126778
rect 88116 126726 88162 126778
rect 88162 126726 88172 126778
rect 88196 126726 88226 126778
rect 88226 126726 88252 126778
rect 87956 126724 88012 126726
rect 88036 126724 88092 126726
rect 88116 126724 88172 126726
rect 88196 126724 88252 126726
rect 89956 126234 90012 126236
rect 90036 126234 90092 126236
rect 90116 126234 90172 126236
rect 90196 126234 90252 126236
rect 89956 126182 89982 126234
rect 89982 126182 90012 126234
rect 90036 126182 90046 126234
rect 90046 126182 90092 126234
rect 90116 126182 90162 126234
rect 90162 126182 90172 126234
rect 90196 126182 90226 126234
rect 90226 126182 90252 126234
rect 89956 126180 90012 126182
rect 90036 126180 90092 126182
rect 90116 126180 90172 126182
rect 90196 126180 90252 126182
rect 87970 125860 88026 125896
rect 87970 125840 87972 125860
rect 87972 125840 88024 125860
rect 88024 125840 88026 125860
rect 87956 125690 88012 125692
rect 88036 125690 88092 125692
rect 88116 125690 88172 125692
rect 88196 125690 88252 125692
rect 87956 125638 87982 125690
rect 87982 125638 88012 125690
rect 88036 125638 88046 125690
rect 88046 125638 88092 125690
rect 88116 125638 88162 125690
rect 88162 125638 88172 125690
rect 88196 125638 88226 125690
rect 88226 125638 88252 125690
rect 87956 125636 88012 125638
rect 88036 125636 88092 125638
rect 88116 125636 88172 125638
rect 88196 125636 88252 125638
rect 89956 125146 90012 125148
rect 90036 125146 90092 125148
rect 90116 125146 90172 125148
rect 90196 125146 90252 125148
rect 89956 125094 89982 125146
rect 89982 125094 90012 125146
rect 90036 125094 90046 125146
rect 90046 125094 90092 125146
rect 90116 125094 90162 125146
rect 90162 125094 90172 125146
rect 90196 125094 90226 125146
rect 90226 125094 90252 125146
rect 89956 125092 90012 125094
rect 90036 125092 90092 125094
rect 90116 125092 90172 125094
rect 90196 125092 90252 125094
rect 87956 124602 88012 124604
rect 88036 124602 88092 124604
rect 88116 124602 88172 124604
rect 88196 124602 88252 124604
rect 87956 124550 87982 124602
rect 87982 124550 88012 124602
rect 88036 124550 88046 124602
rect 88046 124550 88092 124602
rect 88116 124550 88162 124602
rect 88162 124550 88172 124602
rect 88196 124550 88226 124602
rect 88226 124550 88252 124602
rect 87956 124548 88012 124550
rect 88036 124548 88092 124550
rect 88116 124548 88172 124550
rect 88196 124548 88252 124550
rect 88246 124344 88302 124400
rect 89956 124058 90012 124060
rect 90036 124058 90092 124060
rect 90116 124058 90172 124060
rect 90196 124058 90252 124060
rect 89956 124006 89982 124058
rect 89982 124006 90012 124058
rect 90036 124006 90046 124058
rect 90046 124006 90092 124058
rect 90116 124006 90162 124058
rect 90162 124006 90172 124058
rect 90196 124006 90226 124058
rect 90226 124006 90252 124058
rect 89956 124004 90012 124006
rect 90036 124004 90092 124006
rect 90116 124004 90172 124006
rect 90196 124004 90252 124006
rect 87956 123514 88012 123516
rect 88036 123514 88092 123516
rect 88116 123514 88172 123516
rect 88196 123514 88252 123516
rect 87956 123462 87982 123514
rect 87982 123462 88012 123514
rect 88036 123462 88046 123514
rect 88046 123462 88092 123514
rect 88116 123462 88162 123514
rect 88162 123462 88172 123514
rect 88196 123462 88226 123514
rect 88226 123462 88252 123514
rect 87956 123460 88012 123462
rect 88036 123460 88092 123462
rect 88116 123460 88172 123462
rect 88196 123460 88252 123462
rect 87970 123256 88026 123312
rect 87956 122426 88012 122428
rect 88036 122426 88092 122428
rect 88116 122426 88172 122428
rect 88196 122426 88252 122428
rect 87956 122374 87982 122426
rect 87982 122374 88012 122426
rect 88036 122374 88046 122426
rect 88046 122374 88092 122426
rect 88116 122374 88162 122426
rect 88162 122374 88172 122426
rect 88196 122374 88226 122426
rect 88226 122374 88252 122426
rect 87956 122372 88012 122374
rect 88036 122372 88092 122374
rect 88116 122372 88172 122374
rect 88196 122372 88252 122374
rect 89956 122970 90012 122972
rect 90036 122970 90092 122972
rect 90116 122970 90172 122972
rect 90196 122970 90252 122972
rect 89956 122918 89982 122970
rect 89982 122918 90012 122970
rect 90036 122918 90046 122970
rect 90046 122918 90092 122970
rect 90116 122918 90162 122970
rect 90162 122918 90172 122970
rect 90196 122918 90226 122970
rect 90226 122918 90252 122970
rect 89956 122916 90012 122918
rect 90036 122916 90092 122918
rect 90116 122916 90172 122918
rect 90196 122916 90252 122918
rect 87878 122032 87934 122088
rect 89956 121882 90012 121884
rect 90036 121882 90092 121884
rect 90116 121882 90172 121884
rect 90196 121882 90252 121884
rect 89956 121830 89982 121882
rect 89982 121830 90012 121882
rect 90036 121830 90046 121882
rect 90046 121830 90092 121882
rect 90116 121830 90162 121882
rect 90162 121830 90172 121882
rect 90196 121830 90226 121882
rect 90226 121830 90252 121882
rect 89956 121828 90012 121830
rect 90036 121828 90092 121830
rect 90116 121828 90172 121830
rect 90196 121828 90252 121830
rect 87956 121338 88012 121340
rect 88036 121338 88092 121340
rect 88116 121338 88172 121340
rect 88196 121338 88252 121340
rect 87956 121286 87982 121338
rect 87982 121286 88012 121338
rect 88036 121286 88046 121338
rect 88046 121286 88092 121338
rect 88116 121286 88162 121338
rect 88162 121286 88172 121338
rect 88196 121286 88226 121338
rect 88226 121286 88252 121338
rect 87956 121284 88012 121286
rect 88036 121284 88092 121286
rect 88116 121284 88172 121286
rect 88196 121284 88252 121286
rect 87878 120536 87934 120592
rect 89956 120794 90012 120796
rect 90036 120794 90092 120796
rect 90116 120794 90172 120796
rect 90196 120794 90252 120796
rect 89956 120742 89982 120794
rect 89982 120742 90012 120794
rect 90036 120742 90046 120794
rect 90046 120742 90092 120794
rect 90116 120742 90162 120794
rect 90162 120742 90172 120794
rect 90196 120742 90226 120794
rect 90226 120742 90252 120794
rect 89956 120740 90012 120742
rect 90036 120740 90092 120742
rect 90116 120740 90172 120742
rect 90196 120740 90252 120742
rect 87956 120250 88012 120252
rect 88036 120250 88092 120252
rect 88116 120250 88172 120252
rect 88196 120250 88252 120252
rect 87956 120198 87982 120250
rect 87982 120198 88012 120250
rect 88036 120198 88046 120250
rect 88046 120198 88092 120250
rect 88116 120198 88162 120250
rect 88162 120198 88172 120250
rect 88196 120198 88226 120250
rect 88226 120198 88252 120250
rect 87956 120196 88012 120198
rect 88036 120196 88092 120198
rect 88116 120196 88172 120198
rect 88196 120196 88252 120198
rect 87878 119448 87934 119504
rect 89956 119706 90012 119708
rect 90036 119706 90092 119708
rect 90116 119706 90172 119708
rect 90196 119706 90252 119708
rect 89956 119654 89982 119706
rect 89982 119654 90012 119706
rect 90036 119654 90046 119706
rect 90046 119654 90092 119706
rect 90116 119654 90162 119706
rect 90162 119654 90172 119706
rect 90196 119654 90226 119706
rect 90226 119654 90252 119706
rect 89956 119652 90012 119654
rect 90036 119652 90092 119654
rect 90116 119652 90172 119654
rect 90196 119652 90252 119654
rect 87956 119162 88012 119164
rect 88036 119162 88092 119164
rect 88116 119162 88172 119164
rect 88196 119162 88252 119164
rect 87956 119110 87982 119162
rect 87982 119110 88012 119162
rect 88036 119110 88046 119162
rect 88046 119110 88092 119162
rect 88116 119110 88162 119162
rect 88162 119110 88172 119162
rect 88196 119110 88226 119162
rect 88226 119110 88252 119162
rect 87956 119108 88012 119110
rect 88036 119108 88092 119110
rect 88116 119108 88172 119110
rect 88196 119108 88252 119110
rect 89956 118618 90012 118620
rect 90036 118618 90092 118620
rect 90116 118618 90172 118620
rect 90196 118618 90252 118620
rect 89956 118566 89982 118618
rect 89982 118566 90012 118618
rect 90036 118566 90046 118618
rect 90046 118566 90092 118618
rect 90116 118566 90162 118618
rect 90162 118566 90172 118618
rect 90196 118566 90226 118618
rect 90226 118566 90252 118618
rect 89956 118564 90012 118566
rect 90036 118564 90092 118566
rect 90116 118564 90172 118566
rect 90196 118564 90252 118566
rect 88982 118360 89038 118416
rect 87956 118074 88012 118076
rect 88036 118074 88092 118076
rect 88116 118074 88172 118076
rect 88196 118074 88252 118076
rect 87956 118022 87982 118074
rect 87982 118022 88012 118074
rect 88036 118022 88046 118074
rect 88046 118022 88092 118074
rect 88116 118022 88162 118074
rect 88162 118022 88172 118074
rect 88196 118022 88226 118074
rect 88226 118022 88252 118074
rect 87956 118020 88012 118022
rect 88036 118020 88092 118022
rect 88116 118020 88172 118022
rect 88196 118020 88252 118022
rect 87956 116986 88012 116988
rect 88036 116986 88092 116988
rect 88116 116986 88172 116988
rect 88196 116986 88252 116988
rect 87956 116934 87982 116986
rect 87982 116934 88012 116986
rect 88036 116934 88046 116986
rect 88046 116934 88092 116986
rect 88116 116934 88162 116986
rect 88162 116934 88172 116986
rect 88196 116934 88226 116986
rect 88226 116934 88252 116986
rect 87956 116932 88012 116934
rect 88036 116932 88092 116934
rect 88116 116932 88172 116934
rect 88196 116932 88252 116934
rect 88246 116728 88302 116784
rect 87956 115898 88012 115900
rect 88036 115898 88092 115900
rect 88116 115898 88172 115900
rect 88196 115898 88252 115900
rect 87956 115846 87982 115898
rect 87982 115846 88012 115898
rect 88036 115846 88046 115898
rect 88046 115846 88092 115898
rect 88116 115846 88162 115898
rect 88162 115846 88172 115898
rect 88196 115846 88226 115898
rect 88226 115846 88252 115898
rect 87956 115844 88012 115846
rect 88036 115844 88092 115846
rect 88116 115844 88172 115846
rect 88196 115844 88252 115846
rect 87956 114810 88012 114812
rect 88036 114810 88092 114812
rect 88116 114810 88172 114812
rect 88196 114810 88252 114812
rect 87956 114758 87982 114810
rect 87982 114758 88012 114810
rect 88036 114758 88046 114810
rect 88046 114758 88092 114810
rect 88116 114758 88162 114810
rect 88162 114758 88172 114810
rect 88196 114758 88226 114810
rect 88226 114758 88252 114810
rect 87956 114756 88012 114758
rect 88036 114756 88092 114758
rect 88116 114756 88172 114758
rect 88196 114756 88252 114758
rect 87970 114572 88026 114608
rect 87970 114552 87972 114572
rect 87972 114552 88024 114572
rect 88024 114552 88026 114572
rect 87956 113722 88012 113724
rect 88036 113722 88092 113724
rect 88116 113722 88172 113724
rect 88196 113722 88252 113724
rect 87956 113670 87982 113722
rect 87982 113670 88012 113722
rect 88036 113670 88046 113722
rect 88046 113670 88092 113722
rect 88116 113670 88162 113722
rect 88162 113670 88172 113722
rect 88196 113670 88226 113722
rect 88226 113670 88252 113722
rect 87956 113668 88012 113670
rect 88036 113668 88092 113670
rect 88116 113668 88172 113670
rect 88196 113668 88252 113670
rect 87956 112634 88012 112636
rect 88036 112634 88092 112636
rect 88116 112634 88172 112636
rect 88196 112634 88252 112636
rect 87956 112582 87982 112634
rect 87982 112582 88012 112634
rect 88036 112582 88046 112634
rect 88046 112582 88092 112634
rect 88116 112582 88162 112634
rect 88162 112582 88172 112634
rect 88196 112582 88226 112634
rect 88226 112582 88252 112634
rect 87956 112580 88012 112582
rect 88036 112580 88092 112582
rect 88116 112580 88172 112582
rect 88196 112580 88252 112582
rect 87970 112376 88026 112432
rect 87956 111546 88012 111548
rect 88036 111546 88092 111548
rect 88116 111546 88172 111548
rect 88196 111546 88252 111548
rect 87956 111494 87982 111546
rect 87982 111494 88012 111546
rect 88036 111494 88046 111546
rect 88046 111494 88092 111546
rect 88116 111494 88162 111546
rect 88162 111494 88172 111546
rect 88196 111494 88226 111546
rect 88226 111494 88252 111546
rect 87956 111492 88012 111494
rect 88036 111492 88092 111494
rect 88116 111492 88172 111494
rect 88196 111492 88252 111494
rect 88246 111152 88302 111208
rect 87956 110458 88012 110460
rect 88036 110458 88092 110460
rect 88116 110458 88172 110460
rect 88196 110458 88252 110460
rect 87956 110406 87982 110458
rect 87982 110406 88012 110458
rect 88036 110406 88046 110458
rect 88046 110406 88092 110458
rect 88116 110406 88162 110458
rect 88162 110406 88172 110458
rect 88196 110406 88226 110458
rect 88226 110406 88252 110458
rect 87956 110404 88012 110406
rect 88036 110404 88092 110406
rect 88116 110404 88172 110406
rect 88196 110404 88252 110406
rect 87956 109370 88012 109372
rect 88036 109370 88092 109372
rect 88116 109370 88172 109372
rect 88196 109370 88252 109372
rect 87956 109318 87982 109370
rect 87982 109318 88012 109370
rect 88036 109318 88046 109370
rect 88046 109318 88092 109370
rect 88116 109318 88162 109370
rect 88162 109318 88172 109370
rect 88196 109318 88226 109370
rect 88226 109318 88252 109370
rect 87956 109316 88012 109318
rect 88036 109316 88092 109318
rect 88116 109316 88172 109318
rect 88196 109316 88252 109318
rect 88246 109112 88302 109168
rect 87970 108604 87972 108624
rect 87972 108604 88024 108624
rect 88024 108604 88026 108624
rect 87970 108568 88026 108604
rect 87956 108282 88012 108284
rect 88036 108282 88092 108284
rect 88116 108282 88172 108284
rect 88196 108282 88252 108284
rect 87956 108230 87982 108282
rect 87982 108230 88012 108282
rect 88036 108230 88046 108282
rect 88046 108230 88092 108282
rect 88116 108230 88162 108282
rect 88162 108230 88172 108282
rect 88196 108230 88226 108282
rect 88226 108230 88252 108282
rect 87956 108228 88012 108230
rect 88036 108228 88092 108230
rect 88116 108228 88172 108230
rect 88196 108228 88252 108230
rect 87970 107480 88026 107536
rect 87956 107194 88012 107196
rect 88036 107194 88092 107196
rect 88116 107194 88172 107196
rect 88196 107194 88252 107196
rect 87956 107142 87982 107194
rect 87982 107142 88012 107194
rect 88036 107142 88046 107194
rect 88046 107142 88092 107194
rect 88116 107142 88162 107194
rect 88162 107142 88172 107194
rect 88196 107142 88226 107194
rect 88226 107142 88252 107194
rect 87956 107140 88012 107142
rect 88036 107140 88092 107142
rect 88116 107140 88172 107142
rect 88196 107140 88252 107142
rect 87956 106106 88012 106108
rect 88036 106106 88092 106108
rect 88116 106106 88172 106108
rect 88196 106106 88252 106108
rect 87956 106054 87982 106106
rect 87982 106054 88012 106106
rect 88036 106054 88046 106106
rect 88046 106054 88092 106106
rect 88116 106054 88162 106106
rect 88162 106054 88172 106106
rect 88196 106054 88226 106106
rect 88226 106054 88252 106106
rect 87956 106052 88012 106054
rect 88036 106052 88092 106054
rect 88116 106052 88172 106054
rect 88196 106052 88252 106054
rect 87956 105018 88012 105020
rect 88036 105018 88092 105020
rect 88116 105018 88172 105020
rect 88196 105018 88252 105020
rect 87956 104966 87982 105018
rect 87982 104966 88012 105018
rect 88036 104966 88046 105018
rect 88046 104966 88092 105018
rect 88116 104966 88162 105018
rect 88162 104966 88172 105018
rect 88196 104966 88226 105018
rect 88226 104966 88252 105018
rect 87956 104964 88012 104966
rect 88036 104964 88092 104966
rect 88116 104964 88172 104966
rect 88196 104964 88252 104966
rect 87602 98776 87658 98832
rect 87956 103930 88012 103932
rect 88036 103930 88092 103932
rect 88116 103930 88172 103932
rect 88196 103930 88252 103932
rect 87956 103878 87982 103930
rect 87982 103878 88012 103930
rect 88036 103878 88046 103930
rect 88046 103878 88092 103930
rect 88116 103878 88162 103930
rect 88162 103878 88172 103930
rect 88196 103878 88226 103930
rect 88226 103878 88252 103930
rect 87956 103876 88012 103878
rect 88036 103876 88092 103878
rect 88116 103876 88172 103878
rect 88196 103876 88252 103878
rect 87956 102842 88012 102844
rect 88036 102842 88092 102844
rect 88116 102842 88172 102844
rect 88196 102842 88252 102844
rect 87956 102790 87982 102842
rect 87982 102790 88012 102842
rect 88036 102790 88046 102842
rect 88046 102790 88092 102842
rect 88116 102790 88162 102842
rect 88162 102790 88172 102842
rect 88196 102790 88226 102842
rect 88226 102790 88252 102842
rect 87956 102788 88012 102790
rect 88036 102788 88092 102790
rect 88116 102788 88172 102790
rect 88196 102788 88252 102790
rect 87956 101754 88012 101756
rect 88036 101754 88092 101756
rect 88116 101754 88172 101756
rect 88196 101754 88252 101756
rect 87956 101702 87982 101754
rect 87982 101702 88012 101754
rect 88036 101702 88046 101754
rect 88046 101702 88092 101754
rect 88116 101702 88162 101754
rect 88162 101702 88172 101754
rect 88196 101702 88226 101754
rect 88226 101702 88252 101754
rect 87956 101700 88012 101702
rect 88036 101700 88092 101702
rect 88116 101700 88172 101702
rect 88196 101700 88252 101702
rect 87956 100666 88012 100668
rect 88036 100666 88092 100668
rect 88116 100666 88172 100668
rect 88196 100666 88252 100668
rect 87956 100614 87982 100666
rect 87982 100614 88012 100666
rect 88036 100614 88046 100666
rect 88046 100614 88092 100666
rect 88116 100614 88162 100666
rect 88162 100614 88172 100666
rect 88196 100614 88226 100666
rect 88226 100614 88252 100666
rect 87956 100612 88012 100614
rect 88036 100612 88092 100614
rect 88116 100612 88172 100614
rect 88196 100612 88252 100614
rect 87956 99578 88012 99580
rect 88036 99578 88092 99580
rect 88116 99578 88172 99580
rect 88196 99578 88252 99580
rect 87956 99526 87982 99578
rect 87982 99526 88012 99578
rect 88036 99526 88046 99578
rect 88046 99526 88092 99578
rect 88116 99526 88162 99578
rect 88162 99526 88172 99578
rect 88196 99526 88226 99578
rect 88226 99526 88252 99578
rect 87956 99524 88012 99526
rect 88036 99524 88092 99526
rect 88116 99524 88172 99526
rect 88196 99524 88252 99526
rect 86682 89528 86738 89584
rect 86682 86808 86738 86864
rect 86958 94288 87014 94344
rect 88522 105032 88578 105088
rect 87956 98490 88012 98492
rect 88036 98490 88092 98492
rect 88116 98490 88172 98492
rect 88196 98490 88252 98492
rect 87956 98438 87982 98490
rect 87982 98438 88012 98490
rect 88036 98438 88046 98490
rect 88046 98438 88092 98490
rect 88116 98438 88162 98490
rect 88162 98438 88172 98490
rect 88196 98438 88226 98490
rect 88226 98438 88252 98490
rect 87956 98436 88012 98438
rect 88036 98436 88092 98438
rect 88116 98436 88172 98438
rect 88196 98436 88252 98438
rect 87786 95920 87842 95976
rect 86866 89528 86922 89584
rect 87050 89528 87106 89584
rect 87050 85040 87106 85096
rect 86866 80144 86922 80200
rect 86958 80008 87014 80064
rect 87050 78512 87106 78568
rect 87510 89800 87566 89856
rect 87418 85040 87474 85096
rect 87234 84632 87290 84688
rect 87142 77016 87198 77072
rect 87050 75928 87106 75984
rect 86958 74704 87014 74760
rect 86958 73616 87014 73672
rect 87326 84496 87382 84552
rect 87326 80012 87382 80068
rect 87234 72528 87290 72584
rect 87142 71032 87198 71088
rect 86682 38256 86738 38312
rect 86590 30776 86646 30832
rect 85956 26138 86012 26140
rect 86036 26138 86092 26140
rect 86116 26138 86172 26140
rect 86196 26138 86252 26140
rect 85956 26086 85982 26138
rect 85982 26086 86012 26138
rect 86036 26086 86046 26138
rect 86046 26086 86092 26138
rect 86116 26086 86162 26138
rect 86162 26086 86172 26138
rect 86196 26086 86226 26138
rect 86226 26086 86252 26138
rect 85956 26084 86012 26086
rect 86036 26084 86092 26086
rect 86116 26084 86172 26086
rect 86196 26084 86252 26086
rect 85956 25050 86012 25052
rect 86036 25050 86092 25052
rect 86116 25050 86172 25052
rect 86196 25050 86252 25052
rect 85956 24998 85982 25050
rect 85982 24998 86012 25050
rect 86036 24998 86046 25050
rect 86046 24998 86092 25050
rect 86116 24998 86162 25050
rect 86162 24998 86172 25050
rect 86196 24998 86226 25050
rect 86226 24998 86252 25050
rect 85956 24996 86012 24998
rect 86036 24996 86092 24998
rect 86116 24996 86172 24998
rect 86196 24996 86252 24998
rect 85956 23962 86012 23964
rect 86036 23962 86092 23964
rect 86116 23962 86172 23964
rect 86196 23962 86252 23964
rect 85956 23910 85982 23962
rect 85982 23910 86012 23962
rect 86036 23910 86046 23962
rect 86046 23910 86092 23962
rect 86116 23910 86162 23962
rect 86162 23910 86172 23962
rect 86196 23910 86226 23962
rect 86226 23910 86252 23962
rect 85956 23908 86012 23910
rect 86036 23908 86092 23910
rect 86116 23908 86172 23910
rect 86196 23908 86252 23910
rect 85956 22874 86012 22876
rect 86036 22874 86092 22876
rect 86116 22874 86172 22876
rect 86196 22874 86252 22876
rect 85956 22822 85982 22874
rect 85982 22822 86012 22874
rect 86036 22822 86046 22874
rect 86046 22822 86092 22874
rect 86116 22822 86162 22874
rect 86162 22822 86172 22874
rect 86196 22822 86226 22874
rect 86226 22822 86252 22874
rect 85956 22820 86012 22822
rect 86036 22820 86092 22822
rect 86116 22820 86172 22822
rect 86196 22820 86252 22822
rect 85956 21786 86012 21788
rect 86036 21786 86092 21788
rect 86116 21786 86172 21788
rect 86196 21786 86252 21788
rect 85956 21734 85982 21786
rect 85982 21734 86012 21786
rect 86036 21734 86046 21786
rect 86046 21734 86092 21786
rect 86116 21734 86162 21786
rect 86162 21734 86172 21786
rect 86196 21734 86226 21786
rect 86226 21734 86252 21786
rect 85956 21732 86012 21734
rect 86036 21732 86092 21734
rect 86116 21732 86172 21734
rect 86196 21732 86252 21734
rect 85956 20698 86012 20700
rect 86036 20698 86092 20700
rect 86116 20698 86172 20700
rect 86196 20698 86252 20700
rect 85956 20646 85982 20698
rect 85982 20646 86012 20698
rect 86036 20646 86046 20698
rect 86046 20646 86092 20698
rect 86116 20646 86162 20698
rect 86162 20646 86172 20698
rect 86196 20646 86226 20698
rect 86226 20646 86252 20698
rect 85956 20644 86012 20646
rect 86036 20644 86092 20646
rect 86116 20644 86172 20646
rect 86196 20644 86252 20646
rect 86314 19896 86370 19952
rect 85956 19610 86012 19612
rect 86036 19610 86092 19612
rect 86116 19610 86172 19612
rect 86196 19610 86252 19612
rect 85956 19558 85982 19610
rect 85982 19558 86012 19610
rect 86036 19558 86046 19610
rect 86046 19558 86092 19610
rect 86116 19558 86162 19610
rect 86162 19558 86172 19610
rect 86196 19558 86226 19610
rect 86226 19558 86252 19610
rect 85956 19556 86012 19558
rect 86036 19556 86092 19558
rect 86116 19556 86172 19558
rect 86196 19556 86252 19558
rect 85956 18522 86012 18524
rect 86036 18522 86092 18524
rect 86116 18522 86172 18524
rect 86196 18522 86252 18524
rect 85956 18470 85982 18522
rect 85982 18470 86012 18522
rect 86036 18470 86046 18522
rect 86046 18470 86092 18522
rect 86116 18470 86162 18522
rect 86162 18470 86172 18522
rect 86196 18470 86226 18522
rect 86226 18470 86252 18522
rect 85956 18468 86012 18470
rect 86036 18468 86092 18470
rect 86116 18468 86172 18470
rect 86196 18468 86252 18470
rect 85956 17434 86012 17436
rect 86036 17434 86092 17436
rect 86116 17434 86172 17436
rect 86196 17434 86252 17436
rect 85956 17382 85982 17434
rect 85982 17382 86012 17434
rect 86036 17382 86046 17434
rect 86046 17382 86092 17434
rect 86116 17382 86162 17434
rect 86162 17382 86172 17434
rect 86196 17382 86226 17434
rect 86226 17382 86252 17434
rect 85956 17380 86012 17382
rect 86036 17380 86092 17382
rect 86116 17380 86172 17382
rect 86196 17380 86252 17382
rect 85956 16346 86012 16348
rect 86036 16346 86092 16348
rect 86116 16346 86172 16348
rect 86196 16346 86252 16348
rect 85956 16294 85982 16346
rect 85982 16294 86012 16346
rect 86036 16294 86046 16346
rect 86046 16294 86092 16346
rect 86116 16294 86162 16346
rect 86162 16294 86172 16346
rect 86196 16294 86226 16346
rect 86226 16294 86252 16346
rect 85956 16292 86012 16294
rect 86036 16292 86092 16294
rect 86116 16292 86172 16294
rect 86196 16292 86252 16294
rect 85956 15258 86012 15260
rect 86036 15258 86092 15260
rect 86116 15258 86172 15260
rect 86196 15258 86252 15260
rect 85956 15206 85982 15258
rect 85982 15206 86012 15258
rect 86036 15206 86046 15258
rect 86046 15206 86092 15258
rect 86116 15206 86162 15258
rect 86162 15206 86172 15258
rect 86196 15206 86226 15258
rect 86226 15206 86252 15258
rect 85956 15204 86012 15206
rect 86036 15204 86092 15206
rect 86116 15204 86172 15206
rect 86196 15204 86252 15206
rect 85956 14170 86012 14172
rect 86036 14170 86092 14172
rect 86116 14170 86172 14172
rect 86196 14170 86252 14172
rect 85956 14118 85982 14170
rect 85982 14118 86012 14170
rect 86036 14118 86046 14170
rect 86046 14118 86092 14170
rect 86116 14118 86162 14170
rect 86162 14118 86172 14170
rect 86196 14118 86226 14170
rect 86226 14118 86252 14170
rect 85956 14116 86012 14118
rect 86036 14116 86092 14118
rect 86116 14116 86172 14118
rect 86196 14116 86252 14118
rect 85956 13082 86012 13084
rect 86036 13082 86092 13084
rect 86116 13082 86172 13084
rect 86196 13082 86252 13084
rect 85956 13030 85982 13082
rect 85982 13030 86012 13082
rect 86036 13030 86046 13082
rect 86046 13030 86092 13082
rect 86116 13030 86162 13082
rect 86162 13030 86172 13082
rect 86196 13030 86226 13082
rect 86226 13030 86252 13082
rect 85956 13028 86012 13030
rect 86036 13028 86092 13030
rect 86116 13028 86172 13030
rect 86196 13028 86252 13030
rect 85956 11994 86012 11996
rect 86036 11994 86092 11996
rect 86116 11994 86172 11996
rect 86196 11994 86252 11996
rect 85956 11942 85982 11994
rect 85982 11942 86012 11994
rect 86036 11942 86046 11994
rect 86046 11942 86092 11994
rect 86116 11942 86162 11994
rect 86162 11942 86172 11994
rect 86196 11942 86226 11994
rect 86226 11942 86252 11994
rect 85956 11940 86012 11942
rect 86036 11940 86092 11942
rect 86116 11940 86172 11942
rect 86196 11940 86252 11942
rect 85956 10906 86012 10908
rect 86036 10906 86092 10908
rect 86116 10906 86172 10908
rect 86196 10906 86252 10908
rect 85956 10854 85982 10906
rect 85982 10854 86012 10906
rect 86036 10854 86046 10906
rect 86046 10854 86092 10906
rect 86116 10854 86162 10906
rect 86162 10854 86172 10906
rect 86196 10854 86226 10906
rect 86226 10854 86252 10906
rect 85956 10852 86012 10854
rect 86036 10852 86092 10854
rect 86116 10852 86172 10854
rect 86196 10852 86252 10854
rect 85956 9818 86012 9820
rect 86036 9818 86092 9820
rect 86116 9818 86172 9820
rect 86196 9818 86252 9820
rect 85956 9766 85982 9818
rect 85982 9766 86012 9818
rect 86036 9766 86046 9818
rect 86046 9766 86092 9818
rect 86116 9766 86162 9818
rect 86162 9766 86172 9818
rect 86196 9766 86226 9818
rect 86226 9766 86252 9818
rect 85956 9764 86012 9766
rect 86036 9764 86092 9766
rect 86116 9764 86172 9766
rect 86196 9764 86252 9766
rect 85956 8730 86012 8732
rect 86036 8730 86092 8732
rect 86116 8730 86172 8732
rect 86196 8730 86252 8732
rect 85956 8678 85982 8730
rect 85982 8678 86012 8730
rect 86036 8678 86046 8730
rect 86046 8678 86092 8730
rect 86116 8678 86162 8730
rect 86162 8678 86172 8730
rect 86196 8678 86226 8730
rect 86226 8678 86252 8730
rect 85956 8676 86012 8678
rect 86036 8676 86092 8678
rect 86116 8676 86172 8678
rect 86196 8676 86252 8678
rect 85956 7642 86012 7644
rect 86036 7642 86092 7644
rect 86116 7642 86172 7644
rect 86196 7642 86252 7644
rect 85956 7590 85982 7642
rect 85982 7590 86012 7642
rect 86036 7590 86046 7642
rect 86046 7590 86092 7642
rect 86116 7590 86162 7642
rect 86162 7590 86172 7642
rect 86196 7590 86226 7642
rect 86226 7590 86252 7642
rect 85956 7588 86012 7590
rect 86036 7588 86092 7590
rect 86116 7588 86172 7590
rect 86196 7588 86252 7590
rect 85956 6554 86012 6556
rect 86036 6554 86092 6556
rect 86116 6554 86172 6556
rect 86196 6554 86252 6556
rect 85956 6502 85982 6554
rect 85982 6502 86012 6554
rect 86036 6502 86046 6554
rect 86046 6502 86092 6554
rect 86116 6502 86162 6554
rect 86162 6502 86172 6554
rect 86196 6502 86226 6554
rect 86226 6502 86252 6554
rect 85956 6500 86012 6502
rect 86036 6500 86092 6502
rect 86116 6500 86172 6502
rect 86196 6500 86252 6502
rect 85956 5466 86012 5468
rect 86036 5466 86092 5468
rect 86116 5466 86172 5468
rect 86196 5466 86252 5468
rect 85956 5414 85982 5466
rect 85982 5414 86012 5466
rect 86036 5414 86046 5466
rect 86046 5414 86092 5466
rect 86116 5414 86162 5466
rect 86162 5414 86172 5466
rect 86196 5414 86226 5466
rect 86226 5414 86252 5466
rect 85956 5412 86012 5414
rect 86036 5412 86092 5414
rect 86116 5412 86172 5414
rect 86196 5412 86252 5414
rect 85956 4378 86012 4380
rect 86036 4378 86092 4380
rect 86116 4378 86172 4380
rect 86196 4378 86252 4380
rect 85956 4326 85982 4378
rect 85982 4326 86012 4378
rect 86036 4326 86046 4378
rect 86046 4326 86092 4378
rect 86116 4326 86162 4378
rect 86162 4326 86172 4378
rect 86196 4326 86226 4378
rect 86226 4326 86252 4378
rect 85956 4324 86012 4326
rect 86036 4324 86092 4326
rect 86116 4324 86172 4326
rect 86196 4324 86252 4326
rect 85956 3290 86012 3292
rect 86036 3290 86092 3292
rect 86116 3290 86172 3292
rect 86196 3290 86252 3292
rect 85956 3238 85982 3290
rect 85982 3238 86012 3290
rect 86036 3238 86046 3290
rect 86046 3238 86092 3290
rect 86116 3238 86162 3290
rect 86162 3238 86172 3290
rect 86196 3238 86226 3290
rect 86226 3238 86252 3290
rect 85956 3236 86012 3238
rect 86036 3236 86092 3238
rect 86116 3236 86172 3238
rect 86196 3236 86252 3238
rect 85956 2202 86012 2204
rect 86036 2202 86092 2204
rect 86116 2202 86172 2204
rect 86196 2202 86252 2204
rect 85956 2150 85982 2202
rect 85982 2150 86012 2202
rect 86036 2150 86046 2202
rect 86046 2150 86092 2202
rect 86116 2150 86162 2202
rect 86162 2150 86172 2202
rect 86196 2150 86226 2202
rect 86226 2150 86252 2202
rect 85956 2148 86012 2150
rect 86036 2148 86092 2150
rect 86116 2148 86172 2150
rect 86196 2148 86252 2150
rect 86406 13912 86462 13968
rect 86498 10104 86554 10160
rect 86774 33360 86830 33416
rect 87142 68720 87198 68776
rect 87418 79872 87474 79928
rect 87326 67224 87382 67280
rect 87326 64912 87382 64968
rect 87510 63824 87566 63880
rect 87418 58928 87474 58984
rect 86958 57876 86960 57896
rect 86960 57876 87012 57896
rect 87012 57876 87014 57896
rect 86958 57840 87014 57876
rect 87050 56380 87052 56400
rect 87052 56380 87104 56400
rect 87104 56380 87106 56400
rect 87050 56344 87106 56380
rect 86958 55256 87014 55312
rect 86958 54032 87014 54088
rect 86958 52944 87014 53000
rect 87694 85176 87750 85232
rect 87786 84768 87842 84824
rect 87786 69808 87842 69864
rect 87786 66172 87788 66192
rect 87788 66172 87840 66192
rect 87840 66172 87842 66192
rect 87786 66136 87842 66172
rect 87786 62736 87842 62792
rect 87786 61240 87842 61296
rect 87694 60016 87750 60072
rect 87694 49136 87750 49192
rect 87602 48048 87658 48104
rect 87694 46552 87750 46608
rect 87602 45464 87658 45520
rect 86958 36760 87014 36816
rect 87510 39344 87566 39400
rect 86958 34584 87014 34640
rect 86958 31864 87014 31920
rect 87326 35672 87382 35728
rect 86958 29688 87014 29744
rect 86958 28464 87014 28520
rect 86958 26968 87014 27024
rect 87234 25880 87290 25936
rect 86958 24792 87014 24848
rect 87050 23588 87106 23624
rect 87050 23568 87052 23588
rect 87052 23568 87104 23588
rect 87104 23568 87106 23588
rect 87142 22480 87198 22536
rect 87142 18808 87198 18864
rect 87234 17584 87290 17640
rect 87142 16088 87198 16144
rect 87142 15000 87198 15056
rect 86958 12688 87014 12744
rect 86958 11192 87014 11248
rect 86958 9016 87014 9072
rect 87050 5208 87106 5264
rect 87050 2896 87106 2952
rect 86866 1672 86922 1728
rect 87326 6296 87382 6352
rect 87694 44240 87750 44296
rect 87694 43152 87750 43208
rect 87786 41656 87842 41712
rect 88706 97552 88762 97608
rect 87956 97402 88012 97404
rect 88036 97402 88092 97404
rect 88116 97402 88172 97404
rect 88196 97402 88252 97404
rect 87956 97350 87982 97402
rect 87982 97350 88012 97402
rect 88036 97350 88046 97402
rect 88046 97350 88092 97402
rect 88116 97350 88162 97402
rect 88162 97350 88172 97402
rect 88196 97350 88226 97402
rect 88226 97350 88252 97402
rect 87956 97348 88012 97350
rect 88036 97348 88092 97350
rect 88116 97348 88172 97350
rect 88196 97348 88252 97350
rect 89956 117530 90012 117532
rect 90036 117530 90092 117532
rect 90116 117530 90172 117532
rect 90196 117530 90252 117532
rect 89956 117478 89982 117530
rect 89982 117478 90012 117530
rect 90036 117478 90046 117530
rect 90046 117478 90092 117530
rect 90116 117478 90162 117530
rect 90162 117478 90172 117530
rect 90196 117478 90226 117530
rect 90226 117478 90252 117530
rect 89956 117476 90012 117478
rect 90036 117476 90092 117478
rect 90116 117476 90172 117478
rect 90196 117476 90252 117478
rect 89956 116442 90012 116444
rect 90036 116442 90092 116444
rect 90116 116442 90172 116444
rect 90196 116442 90252 116444
rect 89956 116390 89982 116442
rect 89982 116390 90012 116442
rect 90036 116390 90046 116442
rect 90046 116390 90092 116442
rect 90116 116390 90162 116442
rect 90162 116390 90172 116442
rect 90196 116390 90226 116442
rect 90226 116390 90252 116442
rect 89956 116388 90012 116390
rect 90036 116388 90092 116390
rect 90116 116388 90172 116390
rect 90196 116388 90252 116390
rect 89956 115354 90012 115356
rect 90036 115354 90092 115356
rect 90116 115354 90172 115356
rect 90196 115354 90252 115356
rect 89956 115302 89982 115354
rect 89982 115302 90012 115354
rect 90036 115302 90046 115354
rect 90046 115302 90092 115354
rect 90116 115302 90162 115354
rect 90162 115302 90172 115354
rect 90196 115302 90226 115354
rect 90226 115302 90252 115354
rect 89956 115300 90012 115302
rect 90036 115300 90092 115302
rect 90116 115300 90172 115302
rect 90196 115300 90252 115302
rect 89956 114266 90012 114268
rect 90036 114266 90092 114268
rect 90116 114266 90172 114268
rect 90196 114266 90252 114268
rect 89956 114214 89982 114266
rect 89982 114214 90012 114266
rect 90036 114214 90046 114266
rect 90046 114214 90092 114266
rect 90116 114214 90162 114266
rect 90162 114214 90172 114266
rect 90196 114214 90226 114266
rect 90226 114214 90252 114266
rect 89956 114212 90012 114214
rect 90036 114212 90092 114214
rect 90116 114212 90172 114214
rect 90196 114212 90252 114214
rect 89956 113178 90012 113180
rect 90036 113178 90092 113180
rect 90116 113178 90172 113180
rect 90196 113178 90252 113180
rect 89956 113126 89982 113178
rect 89982 113126 90012 113178
rect 90036 113126 90046 113178
rect 90046 113126 90092 113178
rect 90116 113126 90162 113178
rect 90162 113126 90172 113178
rect 90196 113126 90226 113178
rect 90226 113126 90252 113178
rect 89956 113124 90012 113126
rect 90036 113124 90092 113126
rect 90116 113124 90172 113126
rect 90196 113124 90252 113126
rect 89956 112090 90012 112092
rect 90036 112090 90092 112092
rect 90116 112090 90172 112092
rect 90196 112090 90252 112092
rect 89956 112038 89982 112090
rect 89982 112038 90012 112090
rect 90036 112038 90046 112090
rect 90046 112038 90092 112090
rect 90116 112038 90162 112090
rect 90162 112038 90172 112090
rect 90196 112038 90226 112090
rect 90226 112038 90252 112090
rect 89956 112036 90012 112038
rect 90036 112036 90092 112038
rect 90116 112036 90172 112038
rect 90196 112036 90252 112038
rect 89956 111002 90012 111004
rect 90036 111002 90092 111004
rect 90116 111002 90172 111004
rect 90196 111002 90252 111004
rect 89956 110950 89982 111002
rect 89982 110950 90012 111002
rect 90036 110950 90046 111002
rect 90046 110950 90092 111002
rect 90116 110950 90162 111002
rect 90162 110950 90172 111002
rect 90196 110950 90226 111002
rect 90226 110950 90252 111002
rect 89956 110948 90012 110950
rect 90036 110948 90092 110950
rect 90116 110948 90172 110950
rect 90196 110948 90252 110950
rect 89956 109914 90012 109916
rect 90036 109914 90092 109916
rect 90116 109914 90172 109916
rect 90196 109914 90252 109916
rect 89956 109862 89982 109914
rect 89982 109862 90012 109914
rect 90036 109862 90046 109914
rect 90046 109862 90092 109914
rect 90116 109862 90162 109914
rect 90162 109862 90172 109914
rect 90196 109862 90226 109914
rect 90226 109862 90252 109914
rect 89956 109860 90012 109862
rect 90036 109860 90092 109862
rect 90116 109860 90172 109862
rect 90196 109860 90252 109862
rect 89956 108826 90012 108828
rect 90036 108826 90092 108828
rect 90116 108826 90172 108828
rect 90196 108826 90252 108828
rect 89956 108774 89982 108826
rect 89982 108774 90012 108826
rect 90036 108774 90046 108826
rect 90046 108774 90092 108826
rect 90116 108774 90162 108826
rect 90162 108774 90172 108826
rect 90196 108774 90226 108826
rect 90226 108774 90252 108826
rect 89956 108772 90012 108774
rect 90036 108772 90092 108774
rect 90116 108772 90172 108774
rect 90196 108772 90252 108774
rect 89956 107738 90012 107740
rect 90036 107738 90092 107740
rect 90116 107738 90172 107740
rect 90196 107738 90252 107740
rect 89956 107686 89982 107738
rect 89982 107686 90012 107738
rect 90036 107686 90046 107738
rect 90046 107686 90092 107738
rect 90116 107686 90162 107738
rect 90162 107686 90172 107738
rect 90196 107686 90226 107738
rect 90226 107686 90252 107738
rect 89956 107684 90012 107686
rect 90036 107684 90092 107686
rect 90116 107684 90172 107686
rect 90196 107684 90252 107686
rect 89956 106650 90012 106652
rect 90036 106650 90092 106652
rect 90116 106650 90172 106652
rect 90196 106650 90252 106652
rect 89956 106598 89982 106650
rect 89982 106598 90012 106650
rect 90036 106598 90046 106650
rect 90046 106598 90092 106650
rect 90116 106598 90162 106650
rect 90162 106598 90172 106650
rect 90196 106598 90226 106650
rect 90226 106598 90252 106650
rect 89956 106596 90012 106598
rect 90036 106596 90092 106598
rect 90116 106596 90172 106598
rect 90196 106596 90252 106598
rect 89956 105562 90012 105564
rect 90036 105562 90092 105564
rect 90116 105562 90172 105564
rect 90196 105562 90252 105564
rect 89956 105510 89982 105562
rect 89982 105510 90012 105562
rect 90036 105510 90046 105562
rect 90046 105510 90092 105562
rect 90116 105510 90162 105562
rect 90162 105510 90172 105562
rect 90196 105510 90226 105562
rect 90226 105510 90252 105562
rect 89956 105508 90012 105510
rect 90036 105508 90092 105510
rect 90116 105508 90172 105510
rect 90196 105508 90252 105510
rect 89956 104474 90012 104476
rect 90036 104474 90092 104476
rect 90116 104474 90172 104476
rect 90196 104474 90252 104476
rect 89956 104422 89982 104474
rect 89982 104422 90012 104474
rect 90036 104422 90046 104474
rect 90046 104422 90092 104474
rect 90116 104422 90162 104474
rect 90162 104422 90172 104474
rect 90196 104422 90226 104474
rect 90226 104422 90252 104474
rect 89956 104420 90012 104422
rect 90036 104420 90092 104422
rect 90116 104420 90172 104422
rect 90196 104420 90252 104422
rect 89956 103386 90012 103388
rect 90036 103386 90092 103388
rect 90116 103386 90172 103388
rect 90196 103386 90252 103388
rect 89956 103334 89982 103386
rect 89982 103334 90012 103386
rect 90036 103334 90046 103386
rect 90046 103334 90092 103386
rect 90116 103334 90162 103386
rect 90162 103334 90172 103386
rect 90196 103334 90226 103386
rect 90226 103334 90252 103386
rect 89956 103332 90012 103334
rect 90036 103332 90092 103334
rect 90116 103332 90172 103334
rect 90196 103332 90252 103334
rect 89956 102298 90012 102300
rect 90036 102298 90092 102300
rect 90116 102298 90172 102300
rect 90196 102298 90252 102300
rect 89956 102246 89982 102298
rect 89982 102246 90012 102298
rect 90036 102246 90046 102298
rect 90046 102246 90092 102298
rect 90116 102246 90162 102298
rect 90162 102246 90172 102298
rect 90196 102246 90226 102298
rect 90226 102246 90252 102298
rect 89956 102244 90012 102246
rect 90036 102244 90092 102246
rect 90116 102244 90172 102246
rect 90196 102244 90252 102246
rect 89956 101210 90012 101212
rect 90036 101210 90092 101212
rect 90116 101210 90172 101212
rect 90196 101210 90252 101212
rect 89956 101158 89982 101210
rect 89982 101158 90012 101210
rect 90036 101158 90046 101210
rect 90046 101158 90092 101210
rect 90116 101158 90162 101210
rect 90162 101158 90172 101210
rect 90196 101158 90226 101210
rect 90226 101158 90252 101210
rect 89956 101156 90012 101158
rect 90036 101156 90092 101158
rect 90116 101156 90172 101158
rect 90196 101156 90252 101158
rect 90362 100136 90418 100192
rect 89956 100122 90012 100124
rect 90036 100122 90092 100124
rect 90116 100122 90172 100124
rect 90196 100122 90252 100124
rect 89956 100070 89982 100122
rect 89982 100070 90012 100122
rect 90036 100070 90046 100122
rect 90046 100070 90092 100122
rect 90116 100070 90162 100122
rect 90162 100070 90172 100122
rect 90196 100070 90226 100122
rect 90226 100070 90252 100122
rect 89956 100068 90012 100070
rect 90036 100068 90092 100070
rect 90116 100068 90172 100070
rect 90196 100068 90252 100070
rect 89956 99034 90012 99036
rect 90036 99034 90092 99036
rect 90116 99034 90172 99036
rect 90196 99034 90252 99036
rect 89956 98982 89982 99034
rect 89982 98982 90012 99034
rect 90036 98982 90046 99034
rect 90046 98982 90092 99034
rect 90116 98982 90162 99034
rect 90162 98982 90172 99034
rect 90196 98982 90226 99034
rect 90226 98982 90252 99034
rect 89956 98980 90012 98982
rect 90036 98980 90092 98982
rect 90116 98980 90172 98982
rect 90196 98980 90252 98982
rect 89956 97946 90012 97948
rect 90036 97946 90092 97948
rect 90116 97946 90172 97948
rect 90196 97946 90252 97948
rect 89956 97894 89982 97946
rect 89982 97894 90012 97946
rect 90036 97894 90046 97946
rect 90046 97894 90092 97946
rect 90116 97894 90162 97946
rect 90162 97894 90172 97946
rect 90196 97894 90226 97946
rect 90226 97894 90252 97946
rect 89956 97892 90012 97894
rect 90036 97892 90092 97894
rect 90116 97892 90172 97894
rect 90196 97892 90252 97894
rect 89956 96858 90012 96860
rect 90036 96858 90092 96860
rect 90116 96858 90172 96860
rect 90196 96858 90252 96860
rect 89956 96806 89982 96858
rect 89982 96806 90012 96858
rect 90036 96806 90046 96858
rect 90046 96806 90092 96858
rect 90116 96806 90162 96858
rect 90162 96806 90172 96858
rect 90196 96806 90226 96858
rect 90226 96806 90252 96858
rect 89956 96804 90012 96806
rect 90036 96804 90092 96806
rect 90116 96804 90172 96806
rect 90196 96804 90252 96806
rect 87956 96314 88012 96316
rect 88036 96314 88092 96316
rect 88116 96314 88172 96316
rect 88196 96314 88252 96316
rect 87956 96262 87982 96314
rect 87982 96262 88012 96314
rect 88036 96262 88046 96314
rect 88046 96262 88092 96314
rect 88116 96262 88162 96314
rect 88162 96262 88172 96314
rect 88196 96262 88226 96314
rect 88226 96262 88252 96314
rect 87956 96260 88012 96262
rect 88036 96260 88092 96262
rect 88116 96260 88172 96262
rect 88196 96260 88252 96262
rect 89956 95770 90012 95772
rect 90036 95770 90092 95772
rect 90116 95770 90172 95772
rect 90196 95770 90252 95772
rect 89956 95718 89982 95770
rect 89982 95718 90012 95770
rect 90036 95718 90046 95770
rect 90046 95718 90092 95770
rect 90116 95718 90162 95770
rect 90162 95718 90172 95770
rect 90196 95718 90226 95770
rect 90226 95718 90252 95770
rect 89956 95716 90012 95718
rect 90036 95716 90092 95718
rect 90116 95716 90172 95718
rect 90196 95716 90252 95718
rect 87956 95226 88012 95228
rect 88036 95226 88092 95228
rect 88116 95226 88172 95228
rect 88196 95226 88252 95228
rect 87956 95174 87982 95226
rect 87982 95174 88012 95226
rect 88036 95174 88046 95226
rect 88046 95174 88092 95226
rect 88116 95174 88162 95226
rect 88162 95174 88172 95226
rect 88196 95174 88226 95226
rect 88226 95174 88252 95226
rect 87956 95172 88012 95174
rect 88036 95172 88092 95174
rect 88116 95172 88172 95174
rect 88196 95172 88252 95174
rect 89956 94682 90012 94684
rect 90036 94682 90092 94684
rect 90116 94682 90172 94684
rect 90196 94682 90252 94684
rect 89956 94630 89982 94682
rect 89982 94630 90012 94682
rect 90036 94630 90046 94682
rect 90046 94630 90092 94682
rect 90116 94630 90162 94682
rect 90162 94630 90172 94682
rect 90196 94630 90226 94682
rect 90226 94630 90252 94682
rect 89956 94628 90012 94630
rect 90036 94628 90092 94630
rect 90116 94628 90172 94630
rect 90196 94628 90252 94630
rect 87956 94138 88012 94140
rect 88036 94138 88092 94140
rect 88116 94138 88172 94140
rect 88196 94138 88252 94140
rect 87956 94086 87982 94138
rect 87982 94086 88012 94138
rect 88036 94086 88046 94138
rect 88046 94086 88092 94138
rect 88116 94086 88162 94138
rect 88162 94086 88172 94138
rect 88196 94086 88226 94138
rect 88226 94086 88252 94138
rect 87956 94084 88012 94086
rect 88036 94084 88092 94086
rect 88116 94084 88172 94086
rect 88196 94084 88252 94086
rect 89956 93594 90012 93596
rect 90036 93594 90092 93596
rect 90116 93594 90172 93596
rect 90196 93594 90252 93596
rect 89956 93542 89982 93594
rect 89982 93542 90012 93594
rect 90036 93542 90046 93594
rect 90046 93542 90092 93594
rect 90116 93542 90162 93594
rect 90162 93542 90172 93594
rect 90196 93542 90226 93594
rect 90226 93542 90252 93594
rect 89956 93540 90012 93542
rect 90036 93540 90092 93542
rect 90116 93540 90172 93542
rect 90196 93540 90252 93542
rect 87956 93050 88012 93052
rect 88036 93050 88092 93052
rect 88116 93050 88172 93052
rect 88196 93050 88252 93052
rect 87956 92998 87982 93050
rect 87982 92998 88012 93050
rect 88036 92998 88046 93050
rect 88046 92998 88092 93050
rect 88116 92998 88162 93050
rect 88162 92998 88172 93050
rect 88196 92998 88226 93050
rect 88226 92998 88252 93050
rect 87956 92996 88012 92998
rect 88036 92996 88092 92998
rect 88116 92996 88172 92998
rect 88196 92996 88252 92998
rect 89956 92506 90012 92508
rect 90036 92506 90092 92508
rect 90116 92506 90172 92508
rect 90196 92506 90252 92508
rect 89956 92454 89982 92506
rect 89982 92454 90012 92506
rect 90036 92454 90046 92506
rect 90046 92454 90092 92506
rect 90116 92454 90162 92506
rect 90162 92454 90172 92506
rect 90196 92454 90226 92506
rect 90226 92454 90252 92506
rect 89956 92452 90012 92454
rect 90036 92452 90092 92454
rect 90116 92452 90172 92454
rect 90196 92452 90252 92454
rect 87956 91962 88012 91964
rect 88036 91962 88092 91964
rect 88116 91962 88172 91964
rect 88196 91962 88252 91964
rect 87956 91910 87982 91962
rect 87982 91910 88012 91962
rect 88036 91910 88046 91962
rect 88046 91910 88092 91962
rect 88116 91910 88162 91962
rect 88162 91910 88172 91962
rect 88196 91910 88226 91962
rect 88226 91910 88252 91962
rect 87956 91908 88012 91910
rect 88036 91908 88092 91910
rect 88116 91908 88172 91910
rect 88196 91908 88252 91910
rect 87956 90874 88012 90876
rect 88036 90874 88092 90876
rect 88116 90874 88172 90876
rect 88196 90874 88252 90876
rect 87956 90822 87982 90874
rect 87982 90822 88012 90874
rect 88036 90822 88046 90874
rect 88046 90822 88092 90874
rect 88116 90822 88162 90874
rect 88162 90822 88172 90874
rect 88196 90822 88226 90874
rect 88226 90822 88252 90874
rect 87956 90820 88012 90822
rect 88036 90820 88092 90822
rect 88116 90820 88172 90822
rect 88196 90820 88252 90822
rect 87956 89786 88012 89788
rect 88036 89786 88092 89788
rect 88116 89786 88172 89788
rect 88196 89786 88252 89788
rect 87956 89734 87982 89786
rect 87982 89734 88012 89786
rect 88036 89734 88046 89786
rect 88046 89734 88092 89786
rect 88116 89734 88162 89786
rect 88162 89734 88172 89786
rect 88196 89734 88226 89786
rect 88226 89734 88252 89786
rect 87956 89732 88012 89734
rect 88036 89732 88092 89734
rect 88116 89732 88172 89734
rect 88196 89732 88252 89734
rect 89956 91418 90012 91420
rect 90036 91418 90092 91420
rect 90116 91418 90172 91420
rect 90196 91418 90252 91420
rect 89956 91366 89982 91418
rect 89982 91366 90012 91418
rect 90036 91366 90046 91418
rect 90046 91366 90092 91418
rect 90116 91366 90162 91418
rect 90162 91366 90172 91418
rect 90196 91366 90226 91418
rect 90226 91366 90252 91418
rect 89956 91364 90012 91366
rect 90036 91364 90092 91366
rect 90116 91364 90172 91366
rect 90196 91364 90252 91366
rect 89956 90330 90012 90332
rect 90036 90330 90092 90332
rect 90116 90330 90172 90332
rect 90196 90330 90252 90332
rect 89956 90278 89982 90330
rect 89982 90278 90012 90330
rect 90036 90278 90046 90330
rect 90046 90278 90092 90330
rect 90116 90278 90162 90330
rect 90162 90278 90172 90330
rect 90196 90278 90226 90330
rect 90226 90278 90252 90330
rect 89956 90276 90012 90278
rect 90036 90276 90092 90278
rect 90116 90276 90172 90278
rect 90196 90276 90252 90278
rect 89956 89242 90012 89244
rect 90036 89242 90092 89244
rect 90116 89242 90172 89244
rect 90196 89242 90252 89244
rect 89956 89190 89982 89242
rect 89982 89190 90012 89242
rect 90036 89190 90046 89242
rect 90046 89190 90092 89242
rect 90116 89190 90162 89242
rect 90162 89190 90172 89242
rect 90196 89190 90226 89242
rect 90226 89190 90252 89242
rect 89956 89188 90012 89190
rect 90036 89188 90092 89190
rect 90116 89188 90172 89190
rect 90196 89188 90252 89190
rect 87956 88698 88012 88700
rect 88036 88698 88092 88700
rect 88116 88698 88172 88700
rect 88196 88698 88252 88700
rect 87956 88646 87982 88698
rect 87982 88646 88012 88698
rect 88036 88646 88046 88698
rect 88046 88646 88092 88698
rect 88116 88646 88162 88698
rect 88162 88646 88172 88698
rect 88196 88646 88226 88698
rect 88226 88646 88252 88698
rect 87956 88644 88012 88646
rect 88036 88644 88092 88646
rect 88116 88644 88172 88646
rect 88196 88644 88252 88646
rect 89956 88154 90012 88156
rect 90036 88154 90092 88156
rect 90116 88154 90172 88156
rect 90196 88154 90252 88156
rect 89956 88102 89982 88154
rect 89982 88102 90012 88154
rect 90036 88102 90046 88154
rect 90046 88102 90092 88154
rect 90116 88102 90162 88154
rect 90162 88102 90172 88154
rect 90196 88102 90226 88154
rect 90226 88102 90252 88154
rect 89956 88100 90012 88102
rect 90036 88100 90092 88102
rect 90116 88100 90172 88102
rect 90196 88100 90252 88102
rect 87970 87896 88026 87952
rect 87956 87610 88012 87612
rect 88036 87610 88092 87612
rect 88116 87610 88172 87612
rect 88196 87610 88252 87612
rect 87956 87558 87982 87610
rect 87982 87558 88012 87610
rect 88036 87558 88046 87610
rect 88046 87558 88092 87610
rect 88116 87558 88162 87610
rect 88162 87558 88172 87610
rect 88196 87558 88226 87610
rect 88226 87558 88252 87610
rect 87956 87556 88012 87558
rect 88036 87556 88092 87558
rect 88116 87556 88172 87558
rect 88196 87556 88252 87558
rect 89956 87066 90012 87068
rect 90036 87066 90092 87068
rect 90116 87066 90172 87068
rect 90196 87066 90252 87068
rect 89956 87014 89982 87066
rect 89982 87014 90012 87066
rect 90036 87014 90046 87066
rect 90046 87014 90092 87066
rect 90116 87014 90162 87066
rect 90162 87014 90172 87066
rect 90196 87014 90226 87066
rect 90226 87014 90252 87066
rect 89956 87012 90012 87014
rect 90036 87012 90092 87014
rect 90116 87012 90172 87014
rect 90196 87012 90252 87014
rect 87956 86522 88012 86524
rect 88036 86522 88092 86524
rect 88116 86522 88172 86524
rect 88196 86522 88252 86524
rect 87956 86470 87982 86522
rect 87982 86470 88012 86522
rect 88036 86470 88046 86522
rect 88046 86470 88092 86522
rect 88116 86470 88162 86522
rect 88162 86470 88172 86522
rect 88196 86470 88226 86522
rect 88226 86470 88252 86522
rect 87956 86468 88012 86470
rect 88036 86468 88092 86470
rect 88116 86468 88172 86470
rect 88196 86468 88252 86470
rect 89956 85978 90012 85980
rect 90036 85978 90092 85980
rect 90116 85978 90172 85980
rect 90196 85978 90252 85980
rect 89956 85926 89982 85978
rect 89982 85926 90012 85978
rect 90036 85926 90046 85978
rect 90046 85926 90092 85978
rect 90116 85926 90162 85978
rect 90162 85926 90172 85978
rect 90196 85926 90226 85978
rect 90226 85926 90252 85978
rect 89956 85924 90012 85926
rect 90036 85924 90092 85926
rect 90116 85924 90172 85926
rect 90196 85924 90252 85926
rect 87970 85584 88026 85640
rect 87956 85434 88012 85436
rect 88036 85434 88092 85436
rect 88116 85434 88172 85436
rect 88196 85434 88252 85436
rect 87956 85382 87982 85434
rect 87982 85382 88012 85434
rect 88036 85382 88046 85434
rect 88046 85382 88092 85434
rect 88116 85382 88162 85434
rect 88162 85382 88172 85434
rect 88196 85382 88226 85434
rect 88226 85382 88252 85434
rect 87956 85380 88012 85382
rect 88036 85380 88092 85382
rect 88116 85380 88172 85382
rect 88196 85380 88252 85382
rect 89956 84890 90012 84892
rect 90036 84890 90092 84892
rect 90116 84890 90172 84892
rect 90196 84890 90252 84892
rect 89956 84838 89982 84890
rect 89982 84838 90012 84890
rect 90036 84838 90046 84890
rect 90046 84838 90092 84890
rect 90116 84838 90162 84890
rect 90162 84838 90172 84890
rect 90196 84838 90226 84890
rect 90226 84838 90252 84890
rect 89956 84836 90012 84838
rect 90036 84836 90092 84838
rect 90116 84836 90172 84838
rect 90196 84836 90252 84838
rect 87970 84496 88026 84552
rect 87956 84346 88012 84348
rect 88036 84346 88092 84348
rect 88116 84346 88172 84348
rect 88196 84346 88252 84348
rect 87956 84294 87982 84346
rect 87982 84294 88012 84346
rect 88036 84294 88046 84346
rect 88046 84294 88092 84346
rect 88116 84294 88162 84346
rect 88162 84294 88172 84346
rect 88196 84294 88226 84346
rect 88226 84294 88252 84346
rect 87956 84292 88012 84294
rect 88036 84292 88092 84294
rect 88116 84292 88172 84294
rect 88196 84292 88252 84294
rect 89956 83802 90012 83804
rect 90036 83802 90092 83804
rect 90116 83802 90172 83804
rect 90196 83802 90252 83804
rect 89956 83750 89982 83802
rect 89982 83750 90012 83802
rect 90036 83750 90046 83802
rect 90046 83750 90092 83802
rect 90116 83750 90162 83802
rect 90162 83750 90172 83802
rect 90196 83750 90226 83802
rect 90226 83750 90252 83802
rect 89956 83748 90012 83750
rect 90036 83748 90092 83750
rect 90116 83748 90172 83750
rect 90196 83748 90252 83750
rect 87970 83408 88026 83464
rect 87956 83258 88012 83260
rect 88036 83258 88092 83260
rect 88116 83258 88172 83260
rect 88196 83258 88252 83260
rect 87956 83206 87982 83258
rect 87982 83206 88012 83258
rect 88036 83206 88046 83258
rect 88046 83206 88092 83258
rect 88116 83206 88162 83258
rect 88162 83206 88172 83258
rect 88196 83206 88226 83258
rect 88226 83206 88252 83258
rect 87956 83204 88012 83206
rect 88036 83204 88092 83206
rect 88116 83204 88172 83206
rect 88196 83204 88252 83206
rect 89956 82714 90012 82716
rect 90036 82714 90092 82716
rect 90116 82714 90172 82716
rect 90196 82714 90252 82716
rect 89956 82662 89982 82714
rect 89982 82662 90012 82714
rect 90036 82662 90046 82714
rect 90046 82662 90092 82714
rect 90116 82662 90162 82714
rect 90162 82662 90172 82714
rect 90196 82662 90226 82714
rect 90226 82662 90252 82714
rect 89956 82660 90012 82662
rect 90036 82660 90092 82662
rect 90116 82660 90172 82662
rect 90196 82660 90252 82662
rect 87956 82170 88012 82172
rect 88036 82170 88092 82172
rect 88116 82170 88172 82172
rect 88196 82170 88252 82172
rect 87956 82118 87982 82170
rect 87982 82118 88012 82170
rect 88036 82118 88046 82170
rect 88046 82118 88092 82170
rect 88116 82118 88162 82170
rect 88162 82118 88172 82170
rect 88196 82118 88226 82170
rect 88226 82118 88252 82170
rect 87956 82116 88012 82118
rect 88036 82116 88092 82118
rect 88116 82116 88172 82118
rect 88196 82116 88252 82118
rect 87970 81948 87972 81968
rect 87972 81948 88024 81968
rect 88024 81948 88026 81968
rect 87970 81912 88026 81948
rect 89956 81626 90012 81628
rect 90036 81626 90092 81628
rect 90116 81626 90172 81628
rect 90196 81626 90252 81628
rect 89956 81574 89982 81626
rect 89982 81574 90012 81626
rect 90036 81574 90046 81626
rect 90046 81574 90092 81626
rect 90116 81574 90162 81626
rect 90162 81574 90172 81626
rect 90196 81574 90226 81626
rect 90226 81574 90252 81626
rect 89956 81572 90012 81574
rect 90036 81572 90092 81574
rect 90116 81572 90172 81574
rect 90196 81572 90252 81574
rect 87956 81082 88012 81084
rect 88036 81082 88092 81084
rect 88116 81082 88172 81084
rect 88196 81082 88252 81084
rect 87956 81030 87982 81082
rect 87982 81030 88012 81082
rect 88036 81030 88046 81082
rect 88046 81030 88092 81082
rect 88116 81030 88162 81082
rect 88162 81030 88172 81082
rect 88196 81030 88226 81082
rect 88226 81030 88252 81082
rect 87956 81028 88012 81030
rect 88036 81028 88092 81030
rect 88116 81028 88172 81030
rect 88196 81028 88252 81030
rect 87970 80688 88026 80744
rect 89956 80538 90012 80540
rect 90036 80538 90092 80540
rect 90116 80538 90172 80540
rect 90196 80538 90252 80540
rect 89956 80486 89982 80538
rect 89982 80486 90012 80538
rect 90036 80486 90046 80538
rect 90046 80486 90092 80538
rect 90116 80486 90162 80538
rect 90162 80486 90172 80538
rect 90196 80486 90226 80538
rect 90226 80486 90252 80538
rect 89956 80484 90012 80486
rect 90036 80484 90092 80486
rect 90116 80484 90172 80486
rect 90196 80484 90252 80486
rect 87956 79994 88012 79996
rect 88036 79994 88092 79996
rect 88116 79994 88172 79996
rect 88196 79994 88252 79996
rect 87956 79942 87982 79994
rect 87982 79942 88012 79994
rect 88036 79942 88046 79994
rect 88046 79942 88092 79994
rect 88116 79942 88162 79994
rect 88162 79942 88172 79994
rect 88196 79942 88226 79994
rect 88226 79942 88252 79994
rect 87956 79940 88012 79942
rect 88036 79940 88092 79942
rect 88116 79940 88172 79942
rect 88196 79940 88252 79942
rect 88246 79600 88302 79656
rect 89956 79450 90012 79452
rect 90036 79450 90092 79452
rect 90116 79450 90172 79452
rect 90196 79450 90252 79452
rect 89956 79398 89982 79450
rect 89982 79398 90012 79450
rect 90036 79398 90046 79450
rect 90046 79398 90092 79450
rect 90116 79398 90162 79450
rect 90162 79398 90172 79450
rect 90196 79398 90226 79450
rect 90226 79398 90252 79450
rect 89956 79396 90012 79398
rect 90036 79396 90092 79398
rect 90116 79396 90172 79398
rect 90196 79396 90252 79398
rect 87956 78906 88012 78908
rect 88036 78906 88092 78908
rect 88116 78906 88172 78908
rect 88196 78906 88252 78908
rect 87956 78854 87982 78906
rect 87982 78854 88012 78906
rect 88036 78854 88046 78906
rect 88046 78854 88092 78906
rect 88116 78854 88162 78906
rect 88162 78854 88172 78906
rect 88196 78854 88226 78906
rect 88226 78854 88252 78906
rect 87956 78852 88012 78854
rect 88036 78852 88092 78854
rect 88116 78852 88172 78854
rect 88196 78852 88252 78854
rect 89956 78362 90012 78364
rect 90036 78362 90092 78364
rect 90116 78362 90172 78364
rect 90196 78362 90252 78364
rect 89956 78310 89982 78362
rect 89982 78310 90012 78362
rect 90036 78310 90046 78362
rect 90046 78310 90092 78362
rect 90116 78310 90162 78362
rect 90162 78310 90172 78362
rect 90196 78310 90226 78362
rect 90226 78310 90252 78362
rect 89956 78308 90012 78310
rect 90036 78308 90092 78310
rect 90116 78308 90172 78310
rect 90196 78308 90252 78310
rect 87956 77818 88012 77820
rect 88036 77818 88092 77820
rect 88116 77818 88172 77820
rect 88196 77818 88252 77820
rect 87956 77766 87982 77818
rect 87982 77766 88012 77818
rect 88036 77766 88046 77818
rect 88046 77766 88092 77818
rect 88116 77766 88162 77818
rect 88162 77766 88172 77818
rect 88196 77766 88226 77818
rect 88226 77766 88252 77818
rect 87956 77764 88012 77766
rect 88036 77764 88092 77766
rect 88116 77764 88172 77766
rect 88196 77764 88252 77766
rect 89956 77274 90012 77276
rect 90036 77274 90092 77276
rect 90116 77274 90172 77276
rect 90196 77274 90252 77276
rect 89956 77222 89982 77274
rect 89982 77222 90012 77274
rect 90036 77222 90046 77274
rect 90046 77222 90092 77274
rect 90116 77222 90162 77274
rect 90162 77222 90172 77274
rect 90196 77222 90226 77274
rect 90226 77222 90252 77274
rect 89956 77220 90012 77222
rect 90036 77220 90092 77222
rect 90116 77220 90172 77222
rect 90196 77220 90252 77222
rect 87956 76730 88012 76732
rect 88036 76730 88092 76732
rect 88116 76730 88172 76732
rect 88196 76730 88252 76732
rect 87956 76678 87982 76730
rect 87982 76678 88012 76730
rect 88036 76678 88046 76730
rect 88046 76678 88092 76730
rect 88116 76678 88162 76730
rect 88162 76678 88172 76730
rect 88196 76678 88226 76730
rect 88226 76678 88252 76730
rect 87956 76676 88012 76678
rect 88036 76676 88092 76678
rect 88116 76676 88172 76678
rect 88196 76676 88252 76678
rect 89956 76186 90012 76188
rect 90036 76186 90092 76188
rect 90116 76186 90172 76188
rect 90196 76186 90252 76188
rect 89956 76134 89982 76186
rect 89982 76134 90012 76186
rect 90036 76134 90046 76186
rect 90046 76134 90092 76186
rect 90116 76134 90162 76186
rect 90162 76134 90172 76186
rect 90196 76134 90226 76186
rect 90226 76134 90252 76186
rect 89956 76132 90012 76134
rect 90036 76132 90092 76134
rect 90116 76132 90172 76134
rect 90196 76132 90252 76134
rect 87956 75642 88012 75644
rect 88036 75642 88092 75644
rect 88116 75642 88172 75644
rect 88196 75642 88252 75644
rect 87956 75590 87982 75642
rect 87982 75590 88012 75642
rect 88036 75590 88046 75642
rect 88046 75590 88092 75642
rect 88116 75590 88162 75642
rect 88162 75590 88172 75642
rect 88196 75590 88226 75642
rect 88226 75590 88252 75642
rect 87956 75588 88012 75590
rect 88036 75588 88092 75590
rect 88116 75588 88172 75590
rect 88196 75588 88252 75590
rect 89956 75098 90012 75100
rect 90036 75098 90092 75100
rect 90116 75098 90172 75100
rect 90196 75098 90252 75100
rect 89956 75046 89982 75098
rect 89982 75046 90012 75098
rect 90036 75046 90046 75098
rect 90046 75046 90092 75098
rect 90116 75046 90162 75098
rect 90162 75046 90172 75098
rect 90196 75046 90226 75098
rect 90226 75046 90252 75098
rect 89956 75044 90012 75046
rect 90036 75044 90092 75046
rect 90116 75044 90172 75046
rect 90196 75044 90252 75046
rect 87956 74554 88012 74556
rect 88036 74554 88092 74556
rect 88116 74554 88172 74556
rect 88196 74554 88252 74556
rect 87956 74502 87982 74554
rect 87982 74502 88012 74554
rect 88036 74502 88046 74554
rect 88046 74502 88092 74554
rect 88116 74502 88162 74554
rect 88162 74502 88172 74554
rect 88196 74502 88226 74554
rect 88226 74502 88252 74554
rect 87956 74500 88012 74502
rect 88036 74500 88092 74502
rect 88116 74500 88172 74502
rect 88196 74500 88252 74502
rect 89956 74010 90012 74012
rect 90036 74010 90092 74012
rect 90116 74010 90172 74012
rect 90196 74010 90252 74012
rect 89956 73958 89982 74010
rect 89982 73958 90012 74010
rect 90036 73958 90046 74010
rect 90046 73958 90092 74010
rect 90116 73958 90162 74010
rect 90162 73958 90172 74010
rect 90196 73958 90226 74010
rect 90226 73958 90252 74010
rect 89956 73956 90012 73958
rect 90036 73956 90092 73958
rect 90116 73956 90172 73958
rect 90196 73956 90252 73958
rect 87956 73466 88012 73468
rect 88036 73466 88092 73468
rect 88116 73466 88172 73468
rect 88196 73466 88252 73468
rect 87956 73414 87982 73466
rect 87982 73414 88012 73466
rect 88036 73414 88046 73466
rect 88046 73414 88092 73466
rect 88116 73414 88162 73466
rect 88162 73414 88172 73466
rect 88196 73414 88226 73466
rect 88226 73414 88252 73466
rect 87956 73412 88012 73414
rect 88036 73412 88092 73414
rect 88116 73412 88172 73414
rect 88196 73412 88252 73414
rect 89956 72922 90012 72924
rect 90036 72922 90092 72924
rect 90116 72922 90172 72924
rect 90196 72922 90252 72924
rect 89956 72870 89982 72922
rect 89982 72870 90012 72922
rect 90036 72870 90046 72922
rect 90046 72870 90092 72922
rect 90116 72870 90162 72922
rect 90162 72870 90172 72922
rect 90196 72870 90226 72922
rect 90226 72870 90252 72922
rect 89956 72868 90012 72870
rect 90036 72868 90092 72870
rect 90116 72868 90172 72870
rect 90196 72868 90252 72870
rect 87956 72378 88012 72380
rect 88036 72378 88092 72380
rect 88116 72378 88172 72380
rect 88196 72378 88252 72380
rect 87956 72326 87982 72378
rect 87982 72326 88012 72378
rect 88036 72326 88046 72378
rect 88046 72326 88092 72378
rect 88116 72326 88162 72378
rect 88162 72326 88172 72378
rect 88196 72326 88226 72378
rect 88226 72326 88252 72378
rect 87956 72324 88012 72326
rect 88036 72324 88092 72326
rect 88116 72324 88172 72326
rect 88196 72324 88252 72326
rect 89956 71834 90012 71836
rect 90036 71834 90092 71836
rect 90116 71834 90172 71836
rect 90196 71834 90252 71836
rect 89956 71782 89982 71834
rect 89982 71782 90012 71834
rect 90036 71782 90046 71834
rect 90046 71782 90092 71834
rect 90116 71782 90162 71834
rect 90162 71782 90172 71834
rect 90196 71782 90226 71834
rect 90226 71782 90252 71834
rect 89956 71780 90012 71782
rect 90036 71780 90092 71782
rect 90116 71780 90172 71782
rect 90196 71780 90252 71782
rect 87956 71290 88012 71292
rect 88036 71290 88092 71292
rect 88116 71290 88172 71292
rect 88196 71290 88252 71292
rect 87956 71238 87982 71290
rect 87982 71238 88012 71290
rect 88036 71238 88046 71290
rect 88046 71238 88092 71290
rect 88116 71238 88162 71290
rect 88162 71238 88172 71290
rect 88196 71238 88226 71290
rect 88226 71238 88252 71290
rect 87956 71236 88012 71238
rect 88036 71236 88092 71238
rect 88116 71236 88172 71238
rect 88196 71236 88252 71238
rect 89956 70746 90012 70748
rect 90036 70746 90092 70748
rect 90116 70746 90172 70748
rect 90196 70746 90252 70748
rect 89956 70694 89982 70746
rect 89982 70694 90012 70746
rect 90036 70694 90046 70746
rect 90046 70694 90092 70746
rect 90116 70694 90162 70746
rect 90162 70694 90172 70746
rect 90196 70694 90226 70746
rect 90226 70694 90252 70746
rect 89956 70692 90012 70694
rect 90036 70692 90092 70694
rect 90116 70692 90172 70694
rect 90196 70692 90252 70694
rect 87956 70202 88012 70204
rect 88036 70202 88092 70204
rect 88116 70202 88172 70204
rect 88196 70202 88252 70204
rect 87956 70150 87982 70202
rect 87982 70150 88012 70202
rect 88036 70150 88046 70202
rect 88046 70150 88092 70202
rect 88116 70150 88162 70202
rect 88162 70150 88172 70202
rect 88196 70150 88226 70202
rect 88226 70150 88252 70202
rect 87956 70148 88012 70150
rect 88036 70148 88092 70150
rect 88116 70148 88172 70150
rect 88196 70148 88252 70150
rect 89956 69658 90012 69660
rect 90036 69658 90092 69660
rect 90116 69658 90172 69660
rect 90196 69658 90252 69660
rect 89956 69606 89982 69658
rect 89982 69606 90012 69658
rect 90036 69606 90046 69658
rect 90046 69606 90092 69658
rect 90116 69606 90162 69658
rect 90162 69606 90172 69658
rect 90196 69606 90226 69658
rect 90226 69606 90252 69658
rect 89956 69604 90012 69606
rect 90036 69604 90092 69606
rect 90116 69604 90172 69606
rect 90196 69604 90252 69606
rect 87956 69114 88012 69116
rect 88036 69114 88092 69116
rect 88116 69114 88172 69116
rect 88196 69114 88252 69116
rect 87956 69062 87982 69114
rect 87982 69062 88012 69114
rect 88036 69062 88046 69114
rect 88046 69062 88092 69114
rect 88116 69062 88162 69114
rect 88162 69062 88172 69114
rect 88196 69062 88226 69114
rect 88226 69062 88252 69114
rect 87956 69060 88012 69062
rect 88036 69060 88092 69062
rect 88116 69060 88172 69062
rect 88196 69060 88252 69062
rect 89956 68570 90012 68572
rect 90036 68570 90092 68572
rect 90116 68570 90172 68572
rect 90196 68570 90252 68572
rect 89956 68518 89982 68570
rect 89982 68518 90012 68570
rect 90036 68518 90046 68570
rect 90046 68518 90092 68570
rect 90116 68518 90162 68570
rect 90162 68518 90172 68570
rect 90196 68518 90226 68570
rect 90226 68518 90252 68570
rect 89956 68516 90012 68518
rect 90036 68516 90092 68518
rect 90116 68516 90172 68518
rect 90196 68516 90252 68518
rect 87956 68026 88012 68028
rect 88036 68026 88092 68028
rect 88116 68026 88172 68028
rect 88196 68026 88252 68028
rect 87956 67974 87982 68026
rect 87982 67974 88012 68026
rect 88036 67974 88046 68026
rect 88046 67974 88092 68026
rect 88116 67974 88162 68026
rect 88162 67974 88172 68026
rect 88196 67974 88226 68026
rect 88226 67974 88252 68026
rect 87956 67972 88012 67974
rect 88036 67972 88092 67974
rect 88116 67972 88172 67974
rect 88196 67972 88252 67974
rect 89956 67482 90012 67484
rect 90036 67482 90092 67484
rect 90116 67482 90172 67484
rect 90196 67482 90252 67484
rect 89956 67430 89982 67482
rect 89982 67430 90012 67482
rect 90036 67430 90046 67482
rect 90046 67430 90092 67482
rect 90116 67430 90162 67482
rect 90162 67430 90172 67482
rect 90196 67430 90226 67482
rect 90226 67430 90252 67482
rect 89956 67428 90012 67430
rect 90036 67428 90092 67430
rect 90116 67428 90172 67430
rect 90196 67428 90252 67430
rect 87956 66938 88012 66940
rect 88036 66938 88092 66940
rect 88116 66938 88172 66940
rect 88196 66938 88252 66940
rect 87956 66886 87982 66938
rect 87982 66886 88012 66938
rect 88036 66886 88046 66938
rect 88046 66886 88092 66938
rect 88116 66886 88162 66938
rect 88162 66886 88172 66938
rect 88196 66886 88226 66938
rect 88226 66886 88252 66938
rect 87956 66884 88012 66886
rect 88036 66884 88092 66886
rect 88116 66884 88172 66886
rect 88196 66884 88252 66886
rect 89956 66394 90012 66396
rect 90036 66394 90092 66396
rect 90116 66394 90172 66396
rect 90196 66394 90252 66396
rect 89956 66342 89982 66394
rect 89982 66342 90012 66394
rect 90036 66342 90046 66394
rect 90046 66342 90092 66394
rect 90116 66342 90162 66394
rect 90162 66342 90172 66394
rect 90196 66342 90226 66394
rect 90226 66342 90252 66394
rect 89956 66340 90012 66342
rect 90036 66340 90092 66342
rect 90116 66340 90172 66342
rect 90196 66340 90252 66342
rect 87956 65850 88012 65852
rect 88036 65850 88092 65852
rect 88116 65850 88172 65852
rect 88196 65850 88252 65852
rect 87956 65798 87982 65850
rect 87982 65798 88012 65850
rect 88036 65798 88046 65850
rect 88046 65798 88092 65850
rect 88116 65798 88162 65850
rect 88162 65798 88172 65850
rect 88196 65798 88226 65850
rect 88226 65798 88252 65850
rect 87956 65796 88012 65798
rect 88036 65796 88092 65798
rect 88116 65796 88172 65798
rect 88196 65796 88252 65798
rect 89956 65306 90012 65308
rect 90036 65306 90092 65308
rect 90116 65306 90172 65308
rect 90196 65306 90252 65308
rect 89956 65254 89982 65306
rect 89982 65254 90012 65306
rect 90036 65254 90046 65306
rect 90046 65254 90092 65306
rect 90116 65254 90162 65306
rect 90162 65254 90172 65306
rect 90196 65254 90226 65306
rect 90226 65254 90252 65306
rect 89956 65252 90012 65254
rect 90036 65252 90092 65254
rect 90116 65252 90172 65254
rect 90196 65252 90252 65254
rect 87956 64762 88012 64764
rect 88036 64762 88092 64764
rect 88116 64762 88172 64764
rect 88196 64762 88252 64764
rect 87956 64710 87982 64762
rect 87982 64710 88012 64762
rect 88036 64710 88046 64762
rect 88046 64710 88092 64762
rect 88116 64710 88162 64762
rect 88162 64710 88172 64762
rect 88196 64710 88226 64762
rect 88226 64710 88252 64762
rect 87956 64708 88012 64710
rect 88036 64708 88092 64710
rect 88116 64708 88172 64710
rect 88196 64708 88252 64710
rect 89956 64218 90012 64220
rect 90036 64218 90092 64220
rect 90116 64218 90172 64220
rect 90196 64218 90252 64220
rect 89956 64166 89982 64218
rect 89982 64166 90012 64218
rect 90036 64166 90046 64218
rect 90046 64166 90092 64218
rect 90116 64166 90162 64218
rect 90162 64166 90172 64218
rect 90196 64166 90226 64218
rect 90226 64166 90252 64218
rect 89956 64164 90012 64166
rect 90036 64164 90092 64166
rect 90116 64164 90172 64166
rect 90196 64164 90252 64166
rect 87956 63674 88012 63676
rect 88036 63674 88092 63676
rect 88116 63674 88172 63676
rect 88196 63674 88252 63676
rect 87956 63622 87982 63674
rect 87982 63622 88012 63674
rect 88036 63622 88046 63674
rect 88046 63622 88092 63674
rect 88116 63622 88162 63674
rect 88162 63622 88172 63674
rect 88196 63622 88226 63674
rect 88226 63622 88252 63674
rect 87956 63620 88012 63622
rect 88036 63620 88092 63622
rect 88116 63620 88172 63622
rect 88196 63620 88252 63622
rect 89956 63130 90012 63132
rect 90036 63130 90092 63132
rect 90116 63130 90172 63132
rect 90196 63130 90252 63132
rect 89956 63078 89982 63130
rect 89982 63078 90012 63130
rect 90036 63078 90046 63130
rect 90046 63078 90092 63130
rect 90116 63078 90162 63130
rect 90162 63078 90172 63130
rect 90196 63078 90226 63130
rect 90226 63078 90252 63130
rect 89956 63076 90012 63078
rect 90036 63076 90092 63078
rect 90116 63076 90172 63078
rect 90196 63076 90252 63078
rect 87956 62586 88012 62588
rect 88036 62586 88092 62588
rect 88116 62586 88172 62588
rect 88196 62586 88252 62588
rect 87956 62534 87982 62586
rect 87982 62534 88012 62586
rect 88036 62534 88046 62586
rect 88046 62534 88092 62586
rect 88116 62534 88162 62586
rect 88162 62534 88172 62586
rect 88196 62534 88226 62586
rect 88226 62534 88252 62586
rect 87956 62532 88012 62534
rect 88036 62532 88092 62534
rect 88116 62532 88172 62534
rect 88196 62532 88252 62534
rect 89956 62042 90012 62044
rect 90036 62042 90092 62044
rect 90116 62042 90172 62044
rect 90196 62042 90252 62044
rect 89956 61990 89982 62042
rect 89982 61990 90012 62042
rect 90036 61990 90046 62042
rect 90046 61990 90092 62042
rect 90116 61990 90162 62042
rect 90162 61990 90172 62042
rect 90196 61990 90226 62042
rect 90226 61990 90252 62042
rect 89956 61988 90012 61990
rect 90036 61988 90092 61990
rect 90116 61988 90172 61990
rect 90196 61988 90252 61990
rect 87956 61498 88012 61500
rect 88036 61498 88092 61500
rect 88116 61498 88172 61500
rect 88196 61498 88252 61500
rect 87956 61446 87982 61498
rect 87982 61446 88012 61498
rect 88036 61446 88046 61498
rect 88046 61446 88092 61498
rect 88116 61446 88162 61498
rect 88162 61446 88172 61498
rect 88196 61446 88226 61498
rect 88226 61446 88252 61498
rect 87956 61444 88012 61446
rect 88036 61444 88092 61446
rect 88116 61444 88172 61446
rect 88196 61444 88252 61446
rect 89956 60954 90012 60956
rect 90036 60954 90092 60956
rect 90116 60954 90172 60956
rect 90196 60954 90252 60956
rect 89956 60902 89982 60954
rect 89982 60902 90012 60954
rect 90036 60902 90046 60954
rect 90046 60902 90092 60954
rect 90116 60902 90162 60954
rect 90162 60902 90172 60954
rect 90196 60902 90226 60954
rect 90226 60902 90252 60954
rect 89956 60900 90012 60902
rect 90036 60900 90092 60902
rect 90116 60900 90172 60902
rect 90196 60900 90252 60902
rect 87956 60410 88012 60412
rect 88036 60410 88092 60412
rect 88116 60410 88172 60412
rect 88196 60410 88252 60412
rect 87956 60358 87982 60410
rect 87982 60358 88012 60410
rect 88036 60358 88046 60410
rect 88046 60358 88092 60410
rect 88116 60358 88162 60410
rect 88162 60358 88172 60410
rect 88196 60358 88226 60410
rect 88226 60358 88252 60410
rect 87956 60356 88012 60358
rect 88036 60356 88092 60358
rect 88116 60356 88172 60358
rect 88196 60356 88252 60358
rect 89956 59866 90012 59868
rect 90036 59866 90092 59868
rect 90116 59866 90172 59868
rect 90196 59866 90252 59868
rect 89956 59814 89982 59866
rect 89982 59814 90012 59866
rect 90036 59814 90046 59866
rect 90046 59814 90092 59866
rect 90116 59814 90162 59866
rect 90162 59814 90172 59866
rect 90196 59814 90226 59866
rect 90226 59814 90252 59866
rect 89956 59812 90012 59814
rect 90036 59812 90092 59814
rect 90116 59812 90172 59814
rect 90196 59812 90252 59814
rect 87956 59322 88012 59324
rect 88036 59322 88092 59324
rect 88116 59322 88172 59324
rect 88196 59322 88252 59324
rect 87956 59270 87982 59322
rect 87982 59270 88012 59322
rect 88036 59270 88046 59322
rect 88046 59270 88092 59322
rect 88116 59270 88162 59322
rect 88162 59270 88172 59322
rect 88196 59270 88226 59322
rect 88226 59270 88252 59322
rect 87956 59268 88012 59270
rect 88036 59268 88092 59270
rect 88116 59268 88172 59270
rect 88196 59268 88252 59270
rect 89956 58778 90012 58780
rect 90036 58778 90092 58780
rect 90116 58778 90172 58780
rect 90196 58778 90252 58780
rect 89956 58726 89982 58778
rect 89982 58726 90012 58778
rect 90036 58726 90046 58778
rect 90046 58726 90092 58778
rect 90116 58726 90162 58778
rect 90162 58726 90172 58778
rect 90196 58726 90226 58778
rect 90226 58726 90252 58778
rect 89956 58724 90012 58726
rect 90036 58724 90092 58726
rect 90116 58724 90172 58726
rect 90196 58724 90252 58726
rect 87956 58234 88012 58236
rect 88036 58234 88092 58236
rect 88116 58234 88172 58236
rect 88196 58234 88252 58236
rect 87956 58182 87982 58234
rect 87982 58182 88012 58234
rect 88036 58182 88046 58234
rect 88046 58182 88092 58234
rect 88116 58182 88162 58234
rect 88162 58182 88172 58234
rect 88196 58182 88226 58234
rect 88226 58182 88252 58234
rect 87956 58180 88012 58182
rect 88036 58180 88092 58182
rect 88116 58180 88172 58182
rect 88196 58180 88252 58182
rect 89956 57690 90012 57692
rect 90036 57690 90092 57692
rect 90116 57690 90172 57692
rect 90196 57690 90252 57692
rect 89956 57638 89982 57690
rect 89982 57638 90012 57690
rect 90036 57638 90046 57690
rect 90046 57638 90092 57690
rect 90116 57638 90162 57690
rect 90162 57638 90172 57690
rect 90196 57638 90226 57690
rect 90226 57638 90252 57690
rect 89956 57636 90012 57638
rect 90036 57636 90092 57638
rect 90116 57636 90172 57638
rect 90196 57636 90252 57638
rect 87956 57146 88012 57148
rect 88036 57146 88092 57148
rect 88116 57146 88172 57148
rect 88196 57146 88252 57148
rect 87956 57094 87982 57146
rect 87982 57094 88012 57146
rect 88036 57094 88046 57146
rect 88046 57094 88092 57146
rect 88116 57094 88162 57146
rect 88162 57094 88172 57146
rect 88196 57094 88226 57146
rect 88226 57094 88252 57146
rect 87956 57092 88012 57094
rect 88036 57092 88092 57094
rect 88116 57092 88172 57094
rect 88196 57092 88252 57094
rect 89956 56602 90012 56604
rect 90036 56602 90092 56604
rect 90116 56602 90172 56604
rect 90196 56602 90252 56604
rect 89956 56550 89982 56602
rect 89982 56550 90012 56602
rect 90036 56550 90046 56602
rect 90046 56550 90092 56602
rect 90116 56550 90162 56602
rect 90162 56550 90172 56602
rect 90196 56550 90226 56602
rect 90226 56550 90252 56602
rect 89956 56548 90012 56550
rect 90036 56548 90092 56550
rect 90116 56548 90172 56550
rect 90196 56548 90252 56550
rect 87956 56058 88012 56060
rect 88036 56058 88092 56060
rect 88116 56058 88172 56060
rect 88196 56058 88252 56060
rect 87956 56006 87982 56058
rect 87982 56006 88012 56058
rect 88036 56006 88046 56058
rect 88046 56006 88092 56058
rect 88116 56006 88162 56058
rect 88162 56006 88172 56058
rect 88196 56006 88226 56058
rect 88226 56006 88252 56058
rect 87956 56004 88012 56006
rect 88036 56004 88092 56006
rect 88116 56004 88172 56006
rect 88196 56004 88252 56006
rect 89956 55514 90012 55516
rect 90036 55514 90092 55516
rect 90116 55514 90172 55516
rect 90196 55514 90252 55516
rect 89956 55462 89982 55514
rect 89982 55462 90012 55514
rect 90036 55462 90046 55514
rect 90046 55462 90092 55514
rect 90116 55462 90162 55514
rect 90162 55462 90172 55514
rect 90196 55462 90226 55514
rect 90226 55462 90252 55514
rect 89956 55460 90012 55462
rect 90036 55460 90092 55462
rect 90116 55460 90172 55462
rect 90196 55460 90252 55462
rect 87956 54970 88012 54972
rect 88036 54970 88092 54972
rect 88116 54970 88172 54972
rect 88196 54970 88252 54972
rect 87956 54918 87982 54970
rect 87982 54918 88012 54970
rect 88036 54918 88046 54970
rect 88046 54918 88092 54970
rect 88116 54918 88162 54970
rect 88162 54918 88172 54970
rect 88196 54918 88226 54970
rect 88226 54918 88252 54970
rect 87956 54916 88012 54918
rect 88036 54916 88092 54918
rect 88116 54916 88172 54918
rect 88196 54916 88252 54918
rect 89956 54426 90012 54428
rect 90036 54426 90092 54428
rect 90116 54426 90172 54428
rect 90196 54426 90252 54428
rect 89956 54374 89982 54426
rect 89982 54374 90012 54426
rect 90036 54374 90046 54426
rect 90046 54374 90092 54426
rect 90116 54374 90162 54426
rect 90162 54374 90172 54426
rect 90196 54374 90226 54426
rect 90226 54374 90252 54426
rect 89956 54372 90012 54374
rect 90036 54372 90092 54374
rect 90116 54372 90172 54374
rect 90196 54372 90252 54374
rect 87956 53882 88012 53884
rect 88036 53882 88092 53884
rect 88116 53882 88172 53884
rect 88196 53882 88252 53884
rect 87956 53830 87982 53882
rect 87982 53830 88012 53882
rect 88036 53830 88046 53882
rect 88046 53830 88092 53882
rect 88116 53830 88162 53882
rect 88162 53830 88172 53882
rect 88196 53830 88226 53882
rect 88226 53830 88252 53882
rect 87956 53828 88012 53830
rect 88036 53828 88092 53830
rect 88116 53828 88172 53830
rect 88196 53828 88252 53830
rect 89956 53338 90012 53340
rect 90036 53338 90092 53340
rect 90116 53338 90172 53340
rect 90196 53338 90252 53340
rect 89956 53286 89982 53338
rect 89982 53286 90012 53338
rect 90036 53286 90046 53338
rect 90046 53286 90092 53338
rect 90116 53286 90162 53338
rect 90162 53286 90172 53338
rect 90196 53286 90226 53338
rect 90226 53286 90252 53338
rect 89956 53284 90012 53286
rect 90036 53284 90092 53286
rect 90116 53284 90172 53286
rect 90196 53284 90252 53286
rect 87956 52794 88012 52796
rect 88036 52794 88092 52796
rect 88116 52794 88172 52796
rect 88196 52794 88252 52796
rect 87956 52742 87982 52794
rect 87982 52742 88012 52794
rect 88036 52742 88046 52794
rect 88046 52742 88092 52794
rect 88116 52742 88162 52794
rect 88162 52742 88172 52794
rect 88196 52742 88226 52794
rect 88226 52742 88252 52794
rect 87956 52740 88012 52742
rect 88036 52740 88092 52742
rect 88116 52740 88172 52742
rect 88196 52740 88252 52742
rect 89956 52250 90012 52252
rect 90036 52250 90092 52252
rect 90116 52250 90172 52252
rect 90196 52250 90252 52252
rect 89956 52198 89982 52250
rect 89982 52198 90012 52250
rect 90036 52198 90046 52250
rect 90046 52198 90092 52250
rect 90116 52198 90162 52250
rect 90162 52198 90172 52250
rect 90196 52198 90226 52250
rect 90226 52198 90252 52250
rect 89956 52196 90012 52198
rect 90036 52196 90092 52198
rect 90116 52196 90172 52198
rect 90196 52196 90252 52198
rect 87956 51706 88012 51708
rect 88036 51706 88092 51708
rect 88116 51706 88172 51708
rect 88196 51706 88252 51708
rect 87956 51654 87982 51706
rect 87982 51654 88012 51706
rect 88036 51654 88046 51706
rect 88046 51654 88092 51706
rect 88116 51654 88162 51706
rect 88162 51654 88172 51706
rect 88196 51654 88226 51706
rect 88226 51654 88252 51706
rect 87956 51652 88012 51654
rect 88036 51652 88092 51654
rect 88116 51652 88172 51654
rect 88196 51652 88252 51654
rect 89956 51162 90012 51164
rect 90036 51162 90092 51164
rect 90116 51162 90172 51164
rect 90196 51162 90252 51164
rect 89956 51110 89982 51162
rect 89982 51110 90012 51162
rect 90036 51110 90046 51162
rect 90046 51110 90092 51162
rect 90116 51110 90162 51162
rect 90162 51110 90172 51162
rect 90196 51110 90226 51162
rect 90226 51110 90252 51162
rect 89956 51108 90012 51110
rect 90036 51108 90092 51110
rect 90116 51108 90172 51110
rect 90196 51108 90252 51110
rect 87956 50618 88012 50620
rect 88036 50618 88092 50620
rect 88116 50618 88172 50620
rect 88196 50618 88252 50620
rect 87956 50566 87982 50618
rect 87982 50566 88012 50618
rect 88036 50566 88046 50618
rect 88046 50566 88092 50618
rect 88116 50566 88162 50618
rect 88162 50566 88172 50618
rect 88196 50566 88226 50618
rect 88226 50566 88252 50618
rect 87956 50564 88012 50566
rect 88036 50564 88092 50566
rect 88116 50564 88172 50566
rect 88196 50564 88252 50566
rect 89956 50074 90012 50076
rect 90036 50074 90092 50076
rect 90116 50074 90172 50076
rect 90196 50074 90252 50076
rect 89956 50022 89982 50074
rect 89982 50022 90012 50074
rect 90036 50022 90046 50074
rect 90046 50022 90092 50074
rect 90116 50022 90162 50074
rect 90162 50022 90172 50074
rect 90196 50022 90226 50074
rect 90226 50022 90252 50074
rect 89956 50020 90012 50022
rect 90036 50020 90092 50022
rect 90116 50020 90172 50022
rect 90196 50020 90252 50022
rect 87956 49530 88012 49532
rect 88036 49530 88092 49532
rect 88116 49530 88172 49532
rect 88196 49530 88252 49532
rect 87956 49478 87982 49530
rect 87982 49478 88012 49530
rect 88036 49478 88046 49530
rect 88046 49478 88092 49530
rect 88116 49478 88162 49530
rect 88162 49478 88172 49530
rect 88196 49478 88226 49530
rect 88226 49478 88252 49530
rect 87956 49476 88012 49478
rect 88036 49476 88092 49478
rect 88116 49476 88172 49478
rect 88196 49476 88252 49478
rect 89956 48986 90012 48988
rect 90036 48986 90092 48988
rect 90116 48986 90172 48988
rect 90196 48986 90252 48988
rect 89956 48934 89982 48986
rect 89982 48934 90012 48986
rect 90036 48934 90046 48986
rect 90046 48934 90092 48986
rect 90116 48934 90162 48986
rect 90162 48934 90172 48986
rect 90196 48934 90226 48986
rect 90226 48934 90252 48986
rect 89956 48932 90012 48934
rect 90036 48932 90092 48934
rect 90116 48932 90172 48934
rect 90196 48932 90252 48934
rect 87956 48442 88012 48444
rect 88036 48442 88092 48444
rect 88116 48442 88172 48444
rect 88196 48442 88252 48444
rect 87956 48390 87982 48442
rect 87982 48390 88012 48442
rect 88036 48390 88046 48442
rect 88046 48390 88092 48442
rect 88116 48390 88162 48442
rect 88162 48390 88172 48442
rect 88196 48390 88226 48442
rect 88226 48390 88252 48442
rect 87956 48388 88012 48390
rect 88036 48388 88092 48390
rect 88116 48388 88172 48390
rect 88196 48388 88252 48390
rect 89956 47898 90012 47900
rect 90036 47898 90092 47900
rect 90116 47898 90172 47900
rect 90196 47898 90252 47900
rect 89956 47846 89982 47898
rect 89982 47846 90012 47898
rect 90036 47846 90046 47898
rect 90046 47846 90092 47898
rect 90116 47846 90162 47898
rect 90162 47846 90172 47898
rect 90196 47846 90226 47898
rect 90226 47846 90252 47898
rect 89956 47844 90012 47846
rect 90036 47844 90092 47846
rect 90116 47844 90172 47846
rect 90196 47844 90252 47846
rect 87956 47354 88012 47356
rect 88036 47354 88092 47356
rect 88116 47354 88172 47356
rect 88196 47354 88252 47356
rect 87956 47302 87982 47354
rect 87982 47302 88012 47354
rect 88036 47302 88046 47354
rect 88046 47302 88092 47354
rect 88116 47302 88162 47354
rect 88162 47302 88172 47354
rect 88196 47302 88226 47354
rect 88226 47302 88252 47354
rect 87956 47300 88012 47302
rect 88036 47300 88092 47302
rect 88116 47300 88172 47302
rect 88196 47300 88252 47302
rect 89956 46810 90012 46812
rect 90036 46810 90092 46812
rect 90116 46810 90172 46812
rect 90196 46810 90252 46812
rect 89956 46758 89982 46810
rect 89982 46758 90012 46810
rect 90036 46758 90046 46810
rect 90046 46758 90092 46810
rect 90116 46758 90162 46810
rect 90162 46758 90172 46810
rect 90196 46758 90226 46810
rect 90226 46758 90252 46810
rect 89956 46756 90012 46758
rect 90036 46756 90092 46758
rect 90116 46756 90172 46758
rect 90196 46756 90252 46758
rect 87956 46266 88012 46268
rect 88036 46266 88092 46268
rect 88116 46266 88172 46268
rect 88196 46266 88252 46268
rect 87956 46214 87982 46266
rect 87982 46214 88012 46266
rect 88036 46214 88046 46266
rect 88046 46214 88092 46266
rect 88116 46214 88162 46266
rect 88162 46214 88172 46266
rect 88196 46214 88226 46266
rect 88226 46214 88252 46266
rect 87956 46212 88012 46214
rect 88036 46212 88092 46214
rect 88116 46212 88172 46214
rect 88196 46212 88252 46214
rect 89956 45722 90012 45724
rect 90036 45722 90092 45724
rect 90116 45722 90172 45724
rect 90196 45722 90252 45724
rect 89956 45670 89982 45722
rect 89982 45670 90012 45722
rect 90036 45670 90046 45722
rect 90046 45670 90092 45722
rect 90116 45670 90162 45722
rect 90162 45670 90172 45722
rect 90196 45670 90226 45722
rect 90226 45670 90252 45722
rect 89956 45668 90012 45670
rect 90036 45668 90092 45670
rect 90116 45668 90172 45670
rect 90196 45668 90252 45670
rect 87956 45178 88012 45180
rect 88036 45178 88092 45180
rect 88116 45178 88172 45180
rect 88196 45178 88252 45180
rect 87956 45126 87982 45178
rect 87982 45126 88012 45178
rect 88036 45126 88046 45178
rect 88046 45126 88092 45178
rect 88116 45126 88162 45178
rect 88162 45126 88172 45178
rect 88196 45126 88226 45178
rect 88226 45126 88252 45178
rect 87956 45124 88012 45126
rect 88036 45124 88092 45126
rect 88116 45124 88172 45126
rect 88196 45124 88252 45126
rect 89956 44634 90012 44636
rect 90036 44634 90092 44636
rect 90116 44634 90172 44636
rect 90196 44634 90252 44636
rect 89956 44582 89982 44634
rect 89982 44582 90012 44634
rect 90036 44582 90046 44634
rect 90046 44582 90092 44634
rect 90116 44582 90162 44634
rect 90162 44582 90172 44634
rect 90196 44582 90226 44634
rect 90226 44582 90252 44634
rect 89956 44580 90012 44582
rect 90036 44580 90092 44582
rect 90116 44580 90172 44582
rect 90196 44580 90252 44582
rect 87956 44090 88012 44092
rect 88036 44090 88092 44092
rect 88116 44090 88172 44092
rect 88196 44090 88252 44092
rect 87956 44038 87982 44090
rect 87982 44038 88012 44090
rect 88036 44038 88046 44090
rect 88046 44038 88092 44090
rect 88116 44038 88162 44090
rect 88162 44038 88172 44090
rect 88196 44038 88226 44090
rect 88226 44038 88252 44090
rect 87956 44036 88012 44038
rect 88036 44036 88092 44038
rect 88116 44036 88172 44038
rect 88196 44036 88252 44038
rect 89956 43546 90012 43548
rect 90036 43546 90092 43548
rect 90116 43546 90172 43548
rect 90196 43546 90252 43548
rect 89956 43494 89982 43546
rect 89982 43494 90012 43546
rect 90036 43494 90046 43546
rect 90046 43494 90092 43546
rect 90116 43494 90162 43546
rect 90162 43494 90172 43546
rect 90196 43494 90226 43546
rect 90226 43494 90252 43546
rect 89956 43492 90012 43494
rect 90036 43492 90092 43494
rect 90116 43492 90172 43494
rect 90196 43492 90252 43494
rect 87956 43002 88012 43004
rect 88036 43002 88092 43004
rect 88116 43002 88172 43004
rect 88196 43002 88252 43004
rect 87956 42950 87982 43002
rect 87982 42950 88012 43002
rect 88036 42950 88046 43002
rect 88046 42950 88092 43002
rect 88116 42950 88162 43002
rect 88162 42950 88172 43002
rect 88196 42950 88226 43002
rect 88226 42950 88252 43002
rect 87956 42948 88012 42950
rect 88036 42948 88092 42950
rect 88116 42948 88172 42950
rect 88196 42948 88252 42950
rect 89956 42458 90012 42460
rect 90036 42458 90092 42460
rect 90116 42458 90172 42460
rect 90196 42458 90252 42460
rect 89956 42406 89982 42458
rect 89982 42406 90012 42458
rect 90036 42406 90046 42458
rect 90046 42406 90092 42458
rect 90116 42406 90162 42458
rect 90162 42406 90172 42458
rect 90196 42406 90226 42458
rect 90226 42406 90252 42458
rect 89956 42404 90012 42406
rect 90036 42404 90092 42406
rect 90116 42404 90172 42406
rect 90196 42404 90252 42406
rect 87956 41914 88012 41916
rect 88036 41914 88092 41916
rect 88116 41914 88172 41916
rect 88196 41914 88252 41916
rect 87956 41862 87982 41914
rect 87982 41862 88012 41914
rect 88036 41862 88046 41914
rect 88046 41862 88092 41914
rect 88116 41862 88162 41914
rect 88162 41862 88172 41914
rect 88196 41862 88226 41914
rect 88226 41862 88252 41914
rect 87956 41860 88012 41862
rect 88036 41860 88092 41862
rect 88116 41860 88172 41862
rect 88196 41860 88252 41862
rect 89956 41370 90012 41372
rect 90036 41370 90092 41372
rect 90116 41370 90172 41372
rect 90196 41370 90252 41372
rect 89956 41318 89982 41370
rect 89982 41318 90012 41370
rect 90036 41318 90046 41370
rect 90046 41318 90092 41370
rect 90116 41318 90162 41370
rect 90162 41318 90172 41370
rect 90196 41318 90226 41370
rect 90226 41318 90252 41370
rect 89956 41316 90012 41318
rect 90036 41316 90092 41318
rect 90116 41316 90172 41318
rect 90196 41316 90252 41318
rect 87956 40826 88012 40828
rect 88036 40826 88092 40828
rect 88116 40826 88172 40828
rect 88196 40826 88252 40828
rect 87956 40774 87982 40826
rect 87982 40774 88012 40826
rect 88036 40774 88046 40826
rect 88046 40774 88092 40826
rect 88116 40774 88162 40826
rect 88162 40774 88172 40826
rect 88196 40774 88226 40826
rect 88226 40774 88252 40826
rect 87956 40772 88012 40774
rect 88036 40772 88092 40774
rect 88116 40772 88172 40774
rect 88196 40772 88252 40774
rect 87878 40568 87934 40624
rect 89956 40282 90012 40284
rect 90036 40282 90092 40284
rect 90116 40282 90172 40284
rect 90196 40282 90252 40284
rect 89956 40230 89982 40282
rect 89982 40230 90012 40282
rect 90036 40230 90046 40282
rect 90046 40230 90092 40282
rect 90116 40230 90162 40282
rect 90162 40230 90172 40282
rect 90196 40230 90226 40282
rect 90226 40230 90252 40282
rect 89956 40228 90012 40230
rect 90036 40228 90092 40230
rect 90116 40228 90172 40230
rect 90196 40228 90252 40230
rect 87956 39738 88012 39740
rect 88036 39738 88092 39740
rect 88116 39738 88172 39740
rect 88196 39738 88252 39740
rect 87956 39686 87982 39738
rect 87982 39686 88012 39738
rect 88036 39686 88046 39738
rect 88046 39686 88092 39738
rect 88116 39686 88162 39738
rect 88162 39686 88172 39738
rect 88196 39686 88226 39738
rect 88226 39686 88252 39738
rect 87956 39684 88012 39686
rect 88036 39684 88092 39686
rect 88116 39684 88172 39686
rect 88196 39684 88252 39686
rect 89956 39194 90012 39196
rect 90036 39194 90092 39196
rect 90116 39194 90172 39196
rect 90196 39194 90252 39196
rect 89956 39142 89982 39194
rect 89982 39142 90012 39194
rect 90036 39142 90046 39194
rect 90046 39142 90092 39194
rect 90116 39142 90162 39194
rect 90162 39142 90172 39194
rect 90196 39142 90226 39194
rect 90226 39142 90252 39194
rect 89956 39140 90012 39142
rect 90036 39140 90092 39142
rect 90116 39140 90172 39142
rect 90196 39140 90252 39142
rect 87956 38650 88012 38652
rect 88036 38650 88092 38652
rect 88116 38650 88172 38652
rect 88196 38650 88252 38652
rect 87956 38598 87982 38650
rect 87982 38598 88012 38650
rect 88036 38598 88046 38650
rect 88046 38598 88092 38650
rect 88116 38598 88162 38650
rect 88162 38598 88172 38650
rect 88196 38598 88226 38650
rect 88226 38598 88252 38650
rect 87956 38596 88012 38598
rect 88036 38596 88092 38598
rect 88116 38596 88172 38598
rect 88196 38596 88252 38598
rect 89956 38106 90012 38108
rect 90036 38106 90092 38108
rect 90116 38106 90172 38108
rect 90196 38106 90252 38108
rect 89956 38054 89982 38106
rect 89982 38054 90012 38106
rect 90036 38054 90046 38106
rect 90046 38054 90092 38106
rect 90116 38054 90162 38106
rect 90162 38054 90172 38106
rect 90196 38054 90226 38106
rect 90226 38054 90252 38106
rect 89956 38052 90012 38054
rect 90036 38052 90092 38054
rect 90116 38052 90172 38054
rect 90196 38052 90252 38054
rect 87956 37562 88012 37564
rect 88036 37562 88092 37564
rect 88116 37562 88172 37564
rect 88196 37562 88252 37564
rect 87956 37510 87982 37562
rect 87982 37510 88012 37562
rect 88036 37510 88046 37562
rect 88046 37510 88092 37562
rect 88116 37510 88162 37562
rect 88162 37510 88172 37562
rect 88196 37510 88226 37562
rect 88226 37510 88252 37562
rect 87956 37508 88012 37510
rect 88036 37508 88092 37510
rect 88116 37508 88172 37510
rect 88196 37508 88252 37510
rect 89956 37018 90012 37020
rect 90036 37018 90092 37020
rect 90116 37018 90172 37020
rect 90196 37018 90252 37020
rect 89956 36966 89982 37018
rect 89982 36966 90012 37018
rect 90036 36966 90046 37018
rect 90046 36966 90092 37018
rect 90116 36966 90162 37018
rect 90162 36966 90172 37018
rect 90196 36966 90226 37018
rect 90226 36966 90252 37018
rect 89956 36964 90012 36966
rect 90036 36964 90092 36966
rect 90116 36964 90172 36966
rect 90196 36964 90252 36966
rect 87956 36474 88012 36476
rect 88036 36474 88092 36476
rect 88116 36474 88172 36476
rect 88196 36474 88252 36476
rect 87956 36422 87982 36474
rect 87982 36422 88012 36474
rect 88036 36422 88046 36474
rect 88046 36422 88092 36474
rect 88116 36422 88162 36474
rect 88162 36422 88172 36474
rect 88196 36422 88226 36474
rect 88226 36422 88252 36474
rect 87956 36420 88012 36422
rect 88036 36420 88092 36422
rect 88116 36420 88172 36422
rect 88196 36420 88252 36422
rect 89956 35930 90012 35932
rect 90036 35930 90092 35932
rect 90116 35930 90172 35932
rect 90196 35930 90252 35932
rect 89956 35878 89982 35930
rect 89982 35878 90012 35930
rect 90036 35878 90046 35930
rect 90046 35878 90092 35930
rect 90116 35878 90162 35930
rect 90162 35878 90172 35930
rect 90196 35878 90226 35930
rect 90226 35878 90252 35930
rect 89956 35876 90012 35878
rect 90036 35876 90092 35878
rect 90116 35876 90172 35878
rect 90196 35876 90252 35878
rect 87956 35386 88012 35388
rect 88036 35386 88092 35388
rect 88116 35386 88172 35388
rect 88196 35386 88252 35388
rect 87956 35334 87982 35386
rect 87982 35334 88012 35386
rect 88036 35334 88046 35386
rect 88046 35334 88092 35386
rect 88116 35334 88162 35386
rect 88162 35334 88172 35386
rect 88196 35334 88226 35386
rect 88226 35334 88252 35386
rect 87956 35332 88012 35334
rect 88036 35332 88092 35334
rect 88116 35332 88172 35334
rect 88196 35332 88252 35334
rect 89956 34842 90012 34844
rect 90036 34842 90092 34844
rect 90116 34842 90172 34844
rect 90196 34842 90252 34844
rect 89956 34790 89982 34842
rect 89982 34790 90012 34842
rect 90036 34790 90046 34842
rect 90046 34790 90092 34842
rect 90116 34790 90162 34842
rect 90162 34790 90172 34842
rect 90196 34790 90226 34842
rect 90226 34790 90252 34842
rect 89956 34788 90012 34790
rect 90036 34788 90092 34790
rect 90116 34788 90172 34790
rect 90196 34788 90252 34790
rect 87956 34298 88012 34300
rect 88036 34298 88092 34300
rect 88116 34298 88172 34300
rect 88196 34298 88252 34300
rect 87956 34246 87982 34298
rect 87982 34246 88012 34298
rect 88036 34246 88046 34298
rect 88046 34246 88092 34298
rect 88116 34246 88162 34298
rect 88162 34246 88172 34298
rect 88196 34246 88226 34298
rect 88226 34246 88252 34298
rect 87956 34244 88012 34246
rect 88036 34244 88092 34246
rect 88116 34244 88172 34246
rect 88196 34244 88252 34246
rect 89956 33754 90012 33756
rect 90036 33754 90092 33756
rect 90116 33754 90172 33756
rect 90196 33754 90252 33756
rect 89956 33702 89982 33754
rect 89982 33702 90012 33754
rect 90036 33702 90046 33754
rect 90046 33702 90092 33754
rect 90116 33702 90162 33754
rect 90162 33702 90172 33754
rect 90196 33702 90226 33754
rect 90226 33702 90252 33754
rect 89956 33700 90012 33702
rect 90036 33700 90092 33702
rect 90116 33700 90172 33702
rect 90196 33700 90252 33702
rect 87956 33210 88012 33212
rect 88036 33210 88092 33212
rect 88116 33210 88172 33212
rect 88196 33210 88252 33212
rect 87956 33158 87982 33210
rect 87982 33158 88012 33210
rect 88036 33158 88046 33210
rect 88046 33158 88092 33210
rect 88116 33158 88162 33210
rect 88162 33158 88172 33210
rect 88196 33158 88226 33210
rect 88226 33158 88252 33210
rect 87956 33156 88012 33158
rect 88036 33156 88092 33158
rect 88116 33156 88172 33158
rect 88196 33156 88252 33158
rect 89956 32666 90012 32668
rect 90036 32666 90092 32668
rect 90116 32666 90172 32668
rect 90196 32666 90252 32668
rect 89956 32614 89982 32666
rect 89982 32614 90012 32666
rect 90036 32614 90046 32666
rect 90046 32614 90092 32666
rect 90116 32614 90162 32666
rect 90162 32614 90172 32666
rect 90196 32614 90226 32666
rect 90226 32614 90252 32666
rect 89956 32612 90012 32614
rect 90036 32612 90092 32614
rect 90116 32612 90172 32614
rect 90196 32612 90252 32614
rect 87956 32122 88012 32124
rect 88036 32122 88092 32124
rect 88116 32122 88172 32124
rect 88196 32122 88252 32124
rect 87956 32070 87982 32122
rect 87982 32070 88012 32122
rect 88036 32070 88046 32122
rect 88046 32070 88092 32122
rect 88116 32070 88162 32122
rect 88162 32070 88172 32122
rect 88196 32070 88226 32122
rect 88226 32070 88252 32122
rect 87956 32068 88012 32070
rect 88036 32068 88092 32070
rect 88116 32068 88172 32070
rect 88196 32068 88252 32070
rect 89956 31578 90012 31580
rect 90036 31578 90092 31580
rect 90116 31578 90172 31580
rect 90196 31578 90252 31580
rect 89956 31526 89982 31578
rect 89982 31526 90012 31578
rect 90036 31526 90046 31578
rect 90046 31526 90092 31578
rect 90116 31526 90162 31578
rect 90162 31526 90172 31578
rect 90196 31526 90226 31578
rect 90226 31526 90252 31578
rect 89956 31524 90012 31526
rect 90036 31524 90092 31526
rect 90116 31524 90172 31526
rect 90196 31524 90252 31526
rect 87956 31034 88012 31036
rect 88036 31034 88092 31036
rect 88116 31034 88172 31036
rect 88196 31034 88252 31036
rect 87956 30982 87982 31034
rect 87982 30982 88012 31034
rect 88036 30982 88046 31034
rect 88046 30982 88092 31034
rect 88116 30982 88162 31034
rect 88162 30982 88172 31034
rect 88196 30982 88226 31034
rect 88226 30982 88252 31034
rect 87956 30980 88012 30982
rect 88036 30980 88092 30982
rect 88116 30980 88172 30982
rect 88196 30980 88252 30982
rect 89956 30490 90012 30492
rect 90036 30490 90092 30492
rect 90116 30490 90172 30492
rect 90196 30490 90252 30492
rect 89956 30438 89982 30490
rect 89982 30438 90012 30490
rect 90036 30438 90046 30490
rect 90046 30438 90092 30490
rect 90116 30438 90162 30490
rect 90162 30438 90172 30490
rect 90196 30438 90226 30490
rect 90226 30438 90252 30490
rect 89956 30436 90012 30438
rect 90036 30436 90092 30438
rect 90116 30436 90172 30438
rect 90196 30436 90252 30438
rect 87956 29946 88012 29948
rect 88036 29946 88092 29948
rect 88116 29946 88172 29948
rect 88196 29946 88252 29948
rect 87956 29894 87982 29946
rect 87982 29894 88012 29946
rect 88036 29894 88046 29946
rect 88046 29894 88092 29946
rect 88116 29894 88162 29946
rect 88162 29894 88172 29946
rect 88196 29894 88226 29946
rect 88226 29894 88252 29946
rect 87956 29892 88012 29894
rect 88036 29892 88092 29894
rect 88116 29892 88172 29894
rect 88196 29892 88252 29894
rect 89956 29402 90012 29404
rect 90036 29402 90092 29404
rect 90116 29402 90172 29404
rect 90196 29402 90252 29404
rect 89956 29350 89982 29402
rect 89982 29350 90012 29402
rect 90036 29350 90046 29402
rect 90046 29350 90092 29402
rect 90116 29350 90162 29402
rect 90162 29350 90172 29402
rect 90196 29350 90226 29402
rect 90226 29350 90252 29402
rect 89956 29348 90012 29350
rect 90036 29348 90092 29350
rect 90116 29348 90172 29350
rect 90196 29348 90252 29350
rect 87956 28858 88012 28860
rect 88036 28858 88092 28860
rect 88116 28858 88172 28860
rect 88196 28858 88252 28860
rect 87956 28806 87982 28858
rect 87982 28806 88012 28858
rect 88036 28806 88046 28858
rect 88046 28806 88092 28858
rect 88116 28806 88162 28858
rect 88162 28806 88172 28858
rect 88196 28806 88226 28858
rect 88226 28806 88252 28858
rect 87956 28804 88012 28806
rect 88036 28804 88092 28806
rect 88116 28804 88172 28806
rect 88196 28804 88252 28806
rect 89956 28314 90012 28316
rect 90036 28314 90092 28316
rect 90116 28314 90172 28316
rect 90196 28314 90252 28316
rect 89956 28262 89982 28314
rect 89982 28262 90012 28314
rect 90036 28262 90046 28314
rect 90046 28262 90092 28314
rect 90116 28262 90162 28314
rect 90162 28262 90172 28314
rect 90196 28262 90226 28314
rect 90226 28262 90252 28314
rect 89956 28260 90012 28262
rect 90036 28260 90092 28262
rect 90116 28260 90172 28262
rect 90196 28260 90252 28262
rect 87956 27770 88012 27772
rect 88036 27770 88092 27772
rect 88116 27770 88172 27772
rect 88196 27770 88252 27772
rect 87956 27718 87982 27770
rect 87982 27718 88012 27770
rect 88036 27718 88046 27770
rect 88046 27718 88092 27770
rect 88116 27718 88162 27770
rect 88162 27718 88172 27770
rect 88196 27718 88226 27770
rect 88226 27718 88252 27770
rect 87956 27716 88012 27718
rect 88036 27716 88092 27718
rect 88116 27716 88172 27718
rect 88196 27716 88252 27718
rect 89956 27226 90012 27228
rect 90036 27226 90092 27228
rect 90116 27226 90172 27228
rect 90196 27226 90252 27228
rect 89956 27174 89982 27226
rect 89982 27174 90012 27226
rect 90036 27174 90046 27226
rect 90046 27174 90092 27226
rect 90116 27174 90162 27226
rect 90162 27174 90172 27226
rect 90196 27174 90226 27226
rect 90226 27174 90252 27226
rect 89956 27172 90012 27174
rect 90036 27172 90092 27174
rect 90116 27172 90172 27174
rect 90196 27172 90252 27174
rect 87956 26682 88012 26684
rect 88036 26682 88092 26684
rect 88116 26682 88172 26684
rect 88196 26682 88252 26684
rect 87956 26630 87982 26682
rect 87982 26630 88012 26682
rect 88036 26630 88046 26682
rect 88046 26630 88092 26682
rect 88116 26630 88162 26682
rect 88162 26630 88172 26682
rect 88196 26630 88226 26682
rect 88226 26630 88252 26682
rect 87956 26628 88012 26630
rect 88036 26628 88092 26630
rect 88116 26628 88172 26630
rect 88196 26628 88252 26630
rect 89956 26138 90012 26140
rect 90036 26138 90092 26140
rect 90116 26138 90172 26140
rect 90196 26138 90252 26140
rect 89956 26086 89982 26138
rect 89982 26086 90012 26138
rect 90036 26086 90046 26138
rect 90046 26086 90092 26138
rect 90116 26086 90162 26138
rect 90162 26086 90172 26138
rect 90196 26086 90226 26138
rect 90226 26086 90252 26138
rect 89956 26084 90012 26086
rect 90036 26084 90092 26086
rect 90116 26084 90172 26086
rect 90196 26084 90252 26086
rect 87956 25594 88012 25596
rect 88036 25594 88092 25596
rect 88116 25594 88172 25596
rect 88196 25594 88252 25596
rect 87956 25542 87982 25594
rect 87982 25542 88012 25594
rect 88036 25542 88046 25594
rect 88046 25542 88092 25594
rect 88116 25542 88162 25594
rect 88162 25542 88172 25594
rect 88196 25542 88226 25594
rect 88226 25542 88252 25594
rect 87956 25540 88012 25542
rect 88036 25540 88092 25542
rect 88116 25540 88172 25542
rect 88196 25540 88252 25542
rect 89956 25050 90012 25052
rect 90036 25050 90092 25052
rect 90116 25050 90172 25052
rect 90196 25050 90252 25052
rect 89956 24998 89982 25050
rect 89982 24998 90012 25050
rect 90036 24998 90046 25050
rect 90046 24998 90092 25050
rect 90116 24998 90162 25050
rect 90162 24998 90172 25050
rect 90196 24998 90226 25050
rect 90226 24998 90252 25050
rect 89956 24996 90012 24998
rect 90036 24996 90092 24998
rect 90116 24996 90172 24998
rect 90196 24996 90252 24998
rect 87956 24506 88012 24508
rect 88036 24506 88092 24508
rect 88116 24506 88172 24508
rect 88196 24506 88252 24508
rect 87956 24454 87982 24506
rect 87982 24454 88012 24506
rect 88036 24454 88046 24506
rect 88046 24454 88092 24506
rect 88116 24454 88162 24506
rect 88162 24454 88172 24506
rect 88196 24454 88226 24506
rect 88226 24454 88252 24506
rect 87956 24452 88012 24454
rect 88036 24452 88092 24454
rect 88116 24452 88172 24454
rect 88196 24452 88252 24454
rect 89956 23962 90012 23964
rect 90036 23962 90092 23964
rect 90116 23962 90172 23964
rect 90196 23962 90252 23964
rect 89956 23910 89982 23962
rect 89982 23910 90012 23962
rect 90036 23910 90046 23962
rect 90046 23910 90092 23962
rect 90116 23910 90162 23962
rect 90162 23910 90172 23962
rect 90196 23910 90226 23962
rect 90226 23910 90252 23962
rect 89956 23908 90012 23910
rect 90036 23908 90092 23910
rect 90116 23908 90172 23910
rect 90196 23908 90252 23910
rect 87956 23418 88012 23420
rect 88036 23418 88092 23420
rect 88116 23418 88172 23420
rect 88196 23418 88252 23420
rect 87956 23366 87982 23418
rect 87982 23366 88012 23418
rect 88036 23366 88046 23418
rect 88046 23366 88092 23418
rect 88116 23366 88162 23418
rect 88162 23366 88172 23418
rect 88196 23366 88226 23418
rect 88226 23366 88252 23418
rect 87956 23364 88012 23366
rect 88036 23364 88092 23366
rect 88116 23364 88172 23366
rect 88196 23364 88252 23366
rect 89956 22874 90012 22876
rect 90036 22874 90092 22876
rect 90116 22874 90172 22876
rect 90196 22874 90252 22876
rect 89956 22822 89982 22874
rect 89982 22822 90012 22874
rect 90036 22822 90046 22874
rect 90046 22822 90092 22874
rect 90116 22822 90162 22874
rect 90162 22822 90172 22874
rect 90196 22822 90226 22874
rect 90226 22822 90252 22874
rect 89956 22820 90012 22822
rect 90036 22820 90092 22822
rect 90116 22820 90172 22822
rect 90196 22820 90252 22822
rect 87956 22330 88012 22332
rect 88036 22330 88092 22332
rect 88116 22330 88172 22332
rect 88196 22330 88252 22332
rect 87956 22278 87982 22330
rect 87982 22278 88012 22330
rect 88036 22278 88046 22330
rect 88046 22278 88092 22330
rect 88116 22278 88162 22330
rect 88162 22278 88172 22330
rect 88196 22278 88226 22330
rect 88226 22278 88252 22330
rect 87956 22276 88012 22278
rect 88036 22276 88092 22278
rect 88116 22276 88172 22278
rect 88196 22276 88252 22278
rect 89956 21786 90012 21788
rect 90036 21786 90092 21788
rect 90116 21786 90172 21788
rect 90196 21786 90252 21788
rect 89956 21734 89982 21786
rect 89982 21734 90012 21786
rect 90036 21734 90046 21786
rect 90046 21734 90092 21786
rect 90116 21734 90162 21786
rect 90162 21734 90172 21786
rect 90196 21734 90226 21786
rect 90226 21734 90252 21786
rect 89956 21732 90012 21734
rect 90036 21732 90092 21734
rect 90116 21732 90172 21734
rect 90196 21732 90252 21734
rect 87956 21242 88012 21244
rect 88036 21242 88092 21244
rect 88116 21242 88172 21244
rect 88196 21242 88252 21244
rect 87956 21190 87982 21242
rect 87982 21190 88012 21242
rect 88036 21190 88046 21242
rect 88046 21190 88092 21242
rect 88116 21190 88162 21242
rect 88162 21190 88172 21242
rect 88196 21190 88226 21242
rect 88226 21190 88252 21242
rect 87956 21188 88012 21190
rect 88036 21188 88092 21190
rect 88116 21188 88172 21190
rect 88196 21188 88252 21190
rect 87878 20984 87934 21040
rect 89956 20698 90012 20700
rect 90036 20698 90092 20700
rect 90116 20698 90172 20700
rect 90196 20698 90252 20700
rect 89956 20646 89982 20698
rect 89982 20646 90012 20698
rect 90036 20646 90046 20698
rect 90046 20646 90092 20698
rect 90116 20646 90162 20698
rect 90162 20646 90172 20698
rect 90196 20646 90226 20698
rect 90226 20646 90252 20698
rect 89956 20644 90012 20646
rect 90036 20644 90092 20646
rect 90116 20644 90172 20646
rect 90196 20644 90252 20646
rect 87956 20154 88012 20156
rect 88036 20154 88092 20156
rect 88116 20154 88172 20156
rect 88196 20154 88252 20156
rect 87956 20102 87982 20154
rect 87982 20102 88012 20154
rect 88036 20102 88046 20154
rect 88046 20102 88092 20154
rect 88116 20102 88162 20154
rect 88162 20102 88172 20154
rect 88196 20102 88226 20154
rect 88226 20102 88252 20154
rect 87956 20100 88012 20102
rect 88036 20100 88092 20102
rect 88116 20100 88172 20102
rect 88196 20100 88252 20102
rect 89956 19610 90012 19612
rect 90036 19610 90092 19612
rect 90116 19610 90172 19612
rect 90196 19610 90252 19612
rect 89956 19558 89982 19610
rect 89982 19558 90012 19610
rect 90036 19558 90046 19610
rect 90046 19558 90092 19610
rect 90116 19558 90162 19610
rect 90162 19558 90172 19610
rect 90196 19558 90226 19610
rect 90226 19558 90252 19610
rect 89956 19556 90012 19558
rect 90036 19556 90092 19558
rect 90116 19556 90172 19558
rect 90196 19556 90252 19558
rect 87956 19066 88012 19068
rect 88036 19066 88092 19068
rect 88116 19066 88172 19068
rect 88196 19066 88252 19068
rect 87956 19014 87982 19066
rect 87982 19014 88012 19066
rect 88036 19014 88046 19066
rect 88046 19014 88092 19066
rect 88116 19014 88162 19066
rect 88162 19014 88172 19066
rect 88196 19014 88226 19066
rect 88226 19014 88252 19066
rect 87956 19012 88012 19014
rect 88036 19012 88092 19014
rect 88116 19012 88172 19014
rect 88196 19012 88252 19014
rect 89956 18522 90012 18524
rect 90036 18522 90092 18524
rect 90116 18522 90172 18524
rect 90196 18522 90252 18524
rect 89956 18470 89982 18522
rect 89982 18470 90012 18522
rect 90036 18470 90046 18522
rect 90046 18470 90092 18522
rect 90116 18470 90162 18522
rect 90162 18470 90172 18522
rect 90196 18470 90226 18522
rect 90226 18470 90252 18522
rect 89956 18468 90012 18470
rect 90036 18468 90092 18470
rect 90116 18468 90172 18470
rect 90196 18468 90252 18470
rect 87956 17978 88012 17980
rect 88036 17978 88092 17980
rect 88116 17978 88172 17980
rect 88196 17978 88252 17980
rect 87956 17926 87982 17978
rect 87982 17926 88012 17978
rect 88036 17926 88046 17978
rect 88046 17926 88092 17978
rect 88116 17926 88162 17978
rect 88162 17926 88172 17978
rect 88196 17926 88226 17978
rect 88226 17926 88252 17978
rect 87956 17924 88012 17926
rect 88036 17924 88092 17926
rect 88116 17924 88172 17926
rect 88196 17924 88252 17926
rect 89956 17434 90012 17436
rect 90036 17434 90092 17436
rect 90116 17434 90172 17436
rect 90196 17434 90252 17436
rect 89956 17382 89982 17434
rect 89982 17382 90012 17434
rect 90036 17382 90046 17434
rect 90046 17382 90092 17434
rect 90116 17382 90162 17434
rect 90162 17382 90172 17434
rect 90196 17382 90226 17434
rect 90226 17382 90252 17434
rect 89956 17380 90012 17382
rect 90036 17380 90092 17382
rect 90116 17380 90172 17382
rect 90196 17380 90252 17382
rect 87956 16890 88012 16892
rect 88036 16890 88092 16892
rect 88116 16890 88172 16892
rect 88196 16890 88252 16892
rect 87956 16838 87982 16890
rect 87982 16838 88012 16890
rect 88036 16838 88046 16890
rect 88046 16838 88092 16890
rect 88116 16838 88162 16890
rect 88162 16838 88172 16890
rect 88196 16838 88226 16890
rect 88226 16838 88252 16890
rect 87956 16836 88012 16838
rect 88036 16836 88092 16838
rect 88116 16836 88172 16838
rect 88196 16836 88252 16838
rect 89956 16346 90012 16348
rect 90036 16346 90092 16348
rect 90116 16346 90172 16348
rect 90196 16346 90252 16348
rect 89956 16294 89982 16346
rect 89982 16294 90012 16346
rect 90036 16294 90046 16346
rect 90046 16294 90092 16346
rect 90116 16294 90162 16346
rect 90162 16294 90172 16346
rect 90196 16294 90226 16346
rect 90226 16294 90252 16346
rect 89956 16292 90012 16294
rect 90036 16292 90092 16294
rect 90116 16292 90172 16294
rect 90196 16292 90252 16294
rect 87956 15802 88012 15804
rect 88036 15802 88092 15804
rect 88116 15802 88172 15804
rect 88196 15802 88252 15804
rect 87956 15750 87982 15802
rect 87982 15750 88012 15802
rect 88036 15750 88046 15802
rect 88046 15750 88092 15802
rect 88116 15750 88162 15802
rect 88162 15750 88172 15802
rect 88196 15750 88226 15802
rect 88226 15750 88252 15802
rect 87956 15748 88012 15750
rect 88036 15748 88092 15750
rect 88116 15748 88172 15750
rect 88196 15748 88252 15750
rect 89956 15258 90012 15260
rect 90036 15258 90092 15260
rect 90116 15258 90172 15260
rect 90196 15258 90252 15260
rect 89956 15206 89982 15258
rect 89982 15206 90012 15258
rect 90036 15206 90046 15258
rect 90046 15206 90092 15258
rect 90116 15206 90162 15258
rect 90162 15206 90172 15258
rect 90196 15206 90226 15258
rect 90226 15206 90252 15258
rect 89956 15204 90012 15206
rect 90036 15204 90092 15206
rect 90116 15204 90172 15206
rect 90196 15204 90252 15206
rect 87956 14714 88012 14716
rect 88036 14714 88092 14716
rect 88116 14714 88172 14716
rect 88196 14714 88252 14716
rect 87956 14662 87982 14714
rect 87982 14662 88012 14714
rect 88036 14662 88046 14714
rect 88046 14662 88092 14714
rect 88116 14662 88162 14714
rect 88162 14662 88172 14714
rect 88196 14662 88226 14714
rect 88226 14662 88252 14714
rect 87956 14660 88012 14662
rect 88036 14660 88092 14662
rect 88116 14660 88172 14662
rect 88196 14660 88252 14662
rect 89956 14170 90012 14172
rect 90036 14170 90092 14172
rect 90116 14170 90172 14172
rect 90196 14170 90252 14172
rect 89956 14118 89982 14170
rect 89982 14118 90012 14170
rect 90036 14118 90046 14170
rect 90046 14118 90092 14170
rect 90116 14118 90162 14170
rect 90162 14118 90172 14170
rect 90196 14118 90226 14170
rect 90226 14118 90252 14170
rect 89956 14116 90012 14118
rect 90036 14116 90092 14118
rect 90116 14116 90172 14118
rect 90196 14116 90252 14118
rect 87956 13626 88012 13628
rect 88036 13626 88092 13628
rect 88116 13626 88172 13628
rect 88196 13626 88252 13628
rect 87956 13574 87982 13626
rect 87982 13574 88012 13626
rect 88036 13574 88046 13626
rect 88046 13574 88092 13626
rect 88116 13574 88162 13626
rect 88162 13574 88172 13626
rect 88196 13574 88226 13626
rect 88226 13574 88252 13626
rect 87956 13572 88012 13574
rect 88036 13572 88092 13574
rect 88116 13572 88172 13574
rect 88196 13572 88252 13574
rect 89956 13082 90012 13084
rect 90036 13082 90092 13084
rect 90116 13082 90172 13084
rect 90196 13082 90252 13084
rect 89956 13030 89982 13082
rect 89982 13030 90012 13082
rect 90036 13030 90046 13082
rect 90046 13030 90092 13082
rect 90116 13030 90162 13082
rect 90162 13030 90172 13082
rect 90196 13030 90226 13082
rect 90226 13030 90252 13082
rect 89956 13028 90012 13030
rect 90036 13028 90092 13030
rect 90116 13028 90172 13030
rect 90196 13028 90252 13030
rect 87956 12538 88012 12540
rect 88036 12538 88092 12540
rect 88116 12538 88172 12540
rect 88196 12538 88252 12540
rect 87956 12486 87982 12538
rect 87982 12486 88012 12538
rect 88036 12486 88046 12538
rect 88046 12486 88092 12538
rect 88116 12486 88162 12538
rect 88162 12486 88172 12538
rect 88196 12486 88226 12538
rect 88226 12486 88252 12538
rect 87956 12484 88012 12486
rect 88036 12484 88092 12486
rect 88116 12484 88172 12486
rect 88196 12484 88252 12486
rect 89956 11994 90012 11996
rect 90036 11994 90092 11996
rect 90116 11994 90172 11996
rect 90196 11994 90252 11996
rect 89956 11942 89982 11994
rect 89982 11942 90012 11994
rect 90036 11942 90046 11994
rect 90046 11942 90092 11994
rect 90116 11942 90162 11994
rect 90162 11942 90172 11994
rect 90196 11942 90226 11994
rect 90226 11942 90252 11994
rect 89956 11940 90012 11942
rect 90036 11940 90092 11942
rect 90116 11940 90172 11942
rect 90196 11940 90252 11942
rect 87956 11450 88012 11452
rect 88036 11450 88092 11452
rect 88116 11450 88172 11452
rect 88196 11450 88252 11452
rect 87956 11398 87982 11450
rect 87982 11398 88012 11450
rect 88036 11398 88046 11450
rect 88046 11398 88092 11450
rect 88116 11398 88162 11450
rect 88162 11398 88172 11450
rect 88196 11398 88226 11450
rect 88226 11398 88252 11450
rect 87956 11396 88012 11398
rect 88036 11396 88092 11398
rect 88116 11396 88172 11398
rect 88196 11396 88252 11398
rect 89956 10906 90012 10908
rect 90036 10906 90092 10908
rect 90116 10906 90172 10908
rect 90196 10906 90252 10908
rect 89956 10854 89982 10906
rect 89982 10854 90012 10906
rect 90036 10854 90046 10906
rect 90046 10854 90092 10906
rect 90116 10854 90162 10906
rect 90162 10854 90172 10906
rect 90196 10854 90226 10906
rect 90226 10854 90252 10906
rect 89956 10852 90012 10854
rect 90036 10852 90092 10854
rect 90116 10852 90172 10854
rect 90196 10852 90252 10854
rect 87956 10362 88012 10364
rect 88036 10362 88092 10364
rect 88116 10362 88172 10364
rect 88196 10362 88252 10364
rect 87956 10310 87982 10362
rect 87982 10310 88012 10362
rect 88036 10310 88046 10362
rect 88046 10310 88092 10362
rect 88116 10310 88162 10362
rect 88162 10310 88172 10362
rect 88196 10310 88226 10362
rect 88226 10310 88252 10362
rect 87956 10308 88012 10310
rect 88036 10308 88092 10310
rect 88116 10308 88172 10310
rect 88196 10308 88252 10310
rect 89956 9818 90012 9820
rect 90036 9818 90092 9820
rect 90116 9818 90172 9820
rect 90196 9818 90252 9820
rect 89956 9766 89982 9818
rect 89982 9766 90012 9818
rect 90036 9766 90046 9818
rect 90046 9766 90092 9818
rect 90116 9766 90162 9818
rect 90162 9766 90172 9818
rect 90196 9766 90226 9818
rect 90226 9766 90252 9818
rect 89956 9764 90012 9766
rect 90036 9764 90092 9766
rect 90116 9764 90172 9766
rect 90196 9764 90252 9766
rect 87956 9274 88012 9276
rect 88036 9274 88092 9276
rect 88116 9274 88172 9276
rect 88196 9274 88252 9276
rect 87956 9222 87982 9274
rect 87982 9222 88012 9274
rect 88036 9222 88046 9274
rect 88046 9222 88092 9274
rect 88116 9222 88162 9274
rect 88162 9222 88172 9274
rect 88196 9222 88226 9274
rect 88226 9222 88252 9274
rect 87956 9220 88012 9222
rect 88036 9220 88092 9222
rect 88116 9220 88172 9222
rect 88196 9220 88252 9222
rect 89956 8730 90012 8732
rect 90036 8730 90092 8732
rect 90116 8730 90172 8732
rect 90196 8730 90252 8732
rect 89956 8678 89982 8730
rect 89982 8678 90012 8730
rect 90036 8678 90046 8730
rect 90046 8678 90092 8730
rect 90116 8678 90162 8730
rect 90162 8678 90172 8730
rect 90196 8678 90226 8730
rect 90226 8678 90252 8730
rect 89956 8676 90012 8678
rect 90036 8676 90092 8678
rect 90116 8676 90172 8678
rect 90196 8676 90252 8678
rect 87956 8186 88012 8188
rect 88036 8186 88092 8188
rect 88116 8186 88172 8188
rect 88196 8186 88252 8188
rect 87956 8134 87982 8186
rect 87982 8134 88012 8186
rect 88036 8134 88046 8186
rect 88046 8134 88092 8186
rect 88116 8134 88162 8186
rect 88162 8134 88172 8186
rect 88196 8134 88226 8186
rect 88226 8134 88252 8186
rect 87956 8132 88012 8134
rect 88036 8132 88092 8134
rect 88116 8132 88172 8134
rect 88196 8132 88252 8134
rect 87878 7792 87934 7848
rect 87602 4120 87658 4176
rect 89956 7642 90012 7644
rect 90036 7642 90092 7644
rect 90116 7642 90172 7644
rect 90196 7642 90252 7644
rect 89956 7590 89982 7642
rect 89982 7590 90012 7642
rect 90036 7590 90046 7642
rect 90046 7590 90092 7642
rect 90116 7590 90162 7642
rect 90162 7590 90172 7642
rect 90196 7590 90226 7642
rect 90226 7590 90252 7642
rect 89956 7588 90012 7590
rect 90036 7588 90092 7590
rect 90116 7588 90172 7590
rect 90196 7588 90252 7590
rect 87956 7098 88012 7100
rect 88036 7098 88092 7100
rect 88116 7098 88172 7100
rect 88196 7098 88252 7100
rect 87956 7046 87982 7098
rect 87982 7046 88012 7098
rect 88036 7046 88046 7098
rect 88046 7046 88092 7098
rect 88116 7046 88162 7098
rect 88162 7046 88172 7098
rect 88196 7046 88226 7098
rect 88226 7046 88252 7098
rect 87956 7044 88012 7046
rect 88036 7044 88092 7046
rect 88116 7044 88172 7046
rect 88196 7044 88252 7046
rect 89956 6554 90012 6556
rect 90036 6554 90092 6556
rect 90116 6554 90172 6556
rect 90196 6554 90252 6556
rect 89956 6502 89982 6554
rect 89982 6502 90012 6554
rect 90036 6502 90046 6554
rect 90046 6502 90092 6554
rect 90116 6502 90162 6554
rect 90162 6502 90172 6554
rect 90196 6502 90226 6554
rect 90226 6502 90252 6554
rect 89956 6500 90012 6502
rect 90036 6500 90092 6502
rect 90116 6500 90172 6502
rect 90196 6500 90252 6502
rect 87956 6010 88012 6012
rect 88036 6010 88092 6012
rect 88116 6010 88172 6012
rect 88196 6010 88252 6012
rect 87956 5958 87982 6010
rect 87982 5958 88012 6010
rect 88036 5958 88046 6010
rect 88046 5958 88092 6010
rect 88116 5958 88162 6010
rect 88162 5958 88172 6010
rect 88196 5958 88226 6010
rect 88226 5958 88252 6010
rect 87956 5956 88012 5958
rect 88036 5956 88092 5958
rect 88116 5956 88172 5958
rect 88196 5956 88252 5958
rect 89956 5466 90012 5468
rect 90036 5466 90092 5468
rect 90116 5466 90172 5468
rect 90196 5466 90252 5468
rect 89956 5414 89982 5466
rect 89982 5414 90012 5466
rect 90036 5414 90046 5466
rect 90046 5414 90092 5466
rect 90116 5414 90162 5466
rect 90162 5414 90172 5466
rect 90196 5414 90226 5466
rect 90226 5414 90252 5466
rect 89956 5412 90012 5414
rect 90036 5412 90092 5414
rect 90116 5412 90172 5414
rect 90196 5412 90252 5414
rect 87956 4922 88012 4924
rect 88036 4922 88092 4924
rect 88116 4922 88172 4924
rect 88196 4922 88252 4924
rect 87956 4870 87982 4922
rect 87982 4870 88012 4922
rect 88036 4870 88046 4922
rect 88046 4870 88092 4922
rect 88116 4870 88162 4922
rect 88162 4870 88172 4922
rect 88196 4870 88226 4922
rect 88226 4870 88252 4922
rect 87956 4868 88012 4870
rect 88036 4868 88092 4870
rect 88116 4868 88172 4870
rect 88196 4868 88252 4870
rect 89956 4378 90012 4380
rect 90036 4378 90092 4380
rect 90116 4378 90172 4380
rect 90196 4378 90252 4380
rect 89956 4326 89982 4378
rect 89982 4326 90012 4378
rect 90036 4326 90046 4378
rect 90046 4326 90092 4378
rect 90116 4326 90162 4378
rect 90162 4326 90172 4378
rect 90196 4326 90226 4378
rect 90226 4326 90252 4378
rect 89956 4324 90012 4326
rect 90036 4324 90092 4326
rect 90116 4324 90172 4326
rect 90196 4324 90252 4326
rect 87956 3834 88012 3836
rect 88036 3834 88092 3836
rect 88116 3834 88172 3836
rect 88196 3834 88252 3836
rect 87956 3782 87982 3834
rect 87982 3782 88012 3834
rect 88036 3782 88046 3834
rect 88046 3782 88092 3834
rect 88116 3782 88162 3834
rect 88162 3782 88172 3834
rect 88196 3782 88226 3834
rect 88226 3782 88252 3834
rect 87956 3780 88012 3782
rect 88036 3780 88092 3782
rect 88116 3780 88172 3782
rect 88196 3780 88252 3782
rect 89956 3290 90012 3292
rect 90036 3290 90092 3292
rect 90116 3290 90172 3292
rect 90196 3290 90252 3292
rect 89956 3238 89982 3290
rect 89982 3238 90012 3290
rect 90036 3238 90046 3290
rect 90046 3238 90092 3290
rect 90116 3238 90162 3290
rect 90162 3238 90172 3290
rect 90196 3238 90226 3290
rect 90226 3238 90252 3290
rect 89956 3236 90012 3238
rect 90036 3236 90092 3238
rect 90116 3236 90172 3238
rect 90196 3236 90252 3238
rect 87956 2746 88012 2748
rect 88036 2746 88092 2748
rect 88116 2746 88172 2748
rect 88196 2746 88252 2748
rect 87956 2694 87982 2746
rect 87982 2694 88012 2746
rect 88036 2694 88046 2746
rect 88046 2694 88092 2746
rect 88116 2694 88162 2746
rect 88162 2694 88172 2746
rect 88196 2694 88226 2746
rect 88226 2694 88252 2746
rect 87956 2692 88012 2694
rect 88036 2692 88092 2694
rect 88116 2692 88172 2694
rect 88196 2692 88252 2694
rect 89956 2202 90012 2204
rect 90036 2202 90092 2204
rect 90116 2202 90172 2204
rect 90196 2202 90252 2204
rect 89956 2150 89982 2202
rect 89982 2150 90012 2202
rect 90036 2150 90046 2202
rect 90046 2150 90092 2202
rect 90116 2150 90162 2202
rect 90162 2150 90172 2202
rect 90196 2150 90226 2202
rect 90226 2150 90252 2202
rect 89956 2148 90012 2150
rect 90036 2148 90092 2150
rect 90116 2148 90172 2150
rect 90196 2148 90252 2150
rect 86958 584 87014 640
<< metal3 >>
rect 89294 191388 89300 191452
rect 89364 191450 89370 191452
rect 91200 191450 92000 191480
rect 89364 191390 92000 191450
rect 89364 191388 89370 191390
rect 91200 191360 92000 191390
rect 88926 190164 88932 190228
rect 88996 190226 89002 190228
rect 91200 190226 92000 190256
rect 88996 190166 92000 190226
rect 88996 190164 89002 190166
rect 91200 190136 92000 190166
rect 1944 189344 2264 189345
rect 1944 189280 1952 189344
rect 2016 189280 2032 189344
rect 2096 189280 2112 189344
rect 2176 189280 2192 189344
rect 2256 189280 2264 189344
rect 1944 189279 2264 189280
rect 85944 189344 86264 189345
rect 85944 189280 85952 189344
rect 86016 189280 86032 189344
rect 86096 189280 86112 189344
rect 86176 189280 86192 189344
rect 86256 189280 86264 189344
rect 85944 189279 86264 189280
rect 89944 189344 90264 189345
rect 89944 189280 89952 189344
rect 90016 189280 90032 189344
rect 90096 189280 90112 189344
rect 90176 189280 90192 189344
rect 90256 189280 90264 189344
rect 89944 189279 90264 189280
rect 75126 189076 75132 189140
rect 75196 189138 75202 189140
rect 75821 189138 75887 189141
rect 75196 189136 75887 189138
rect 75196 189080 75826 189136
rect 75882 189080 75887 189136
rect 75196 189078 75887 189080
rect 75196 189076 75202 189078
rect 75821 189075 75887 189078
rect 89110 188940 89116 189004
rect 89180 189002 89186 189004
rect 91200 189002 92000 189032
rect 89180 188942 92000 189002
rect 89180 188940 89186 188942
rect 91200 188912 92000 188942
rect 3944 188800 4264 188801
rect 3944 188736 3952 188800
rect 4016 188736 4032 188800
rect 4096 188736 4112 188800
rect 4176 188736 4192 188800
rect 4256 188736 4264 188800
rect 3944 188735 4264 188736
rect 87944 188800 88264 188801
rect 87944 188736 87952 188800
rect 88016 188736 88032 188800
rect 88096 188736 88112 188800
rect 88176 188736 88192 188800
rect 88256 188736 88264 188800
rect 87944 188735 88264 188736
rect 1944 188256 2264 188257
rect 1944 188192 1952 188256
rect 2016 188192 2032 188256
rect 2096 188192 2112 188256
rect 2176 188192 2192 188256
rect 2256 188192 2264 188256
rect 1944 188191 2264 188192
rect 85944 188256 86264 188257
rect 85944 188192 85952 188256
rect 86016 188192 86032 188256
rect 86096 188192 86112 188256
rect 86176 188192 86192 188256
rect 86256 188192 86264 188256
rect 85944 188191 86264 188192
rect 89944 188256 90264 188257
rect 89944 188192 89952 188256
rect 90016 188192 90032 188256
rect 90096 188192 90112 188256
rect 90176 188192 90192 188256
rect 90256 188192 90264 188256
rect 89944 188191 90264 188192
rect 89478 187716 89484 187780
rect 89548 187778 89554 187780
rect 91200 187778 92000 187808
rect 89548 187718 92000 187778
rect 89548 187716 89554 187718
rect 3944 187712 4264 187713
rect 3944 187648 3952 187712
rect 4016 187648 4032 187712
rect 4096 187648 4112 187712
rect 4176 187648 4192 187712
rect 4256 187648 4264 187712
rect 3944 187647 4264 187648
rect 87944 187712 88264 187713
rect 87944 187648 87952 187712
rect 88016 187648 88032 187712
rect 88096 187648 88112 187712
rect 88176 187648 88192 187712
rect 88256 187648 88264 187712
rect 91200 187688 92000 187718
rect 87944 187647 88264 187648
rect 1944 187168 2264 187169
rect 1944 187104 1952 187168
rect 2016 187104 2032 187168
rect 2096 187104 2112 187168
rect 2176 187104 2192 187168
rect 2256 187104 2264 187168
rect 1944 187103 2264 187104
rect 85944 187168 86264 187169
rect 85944 187104 85952 187168
rect 86016 187104 86032 187168
rect 86096 187104 86112 187168
rect 86176 187104 86192 187168
rect 86256 187104 86264 187168
rect 85944 187103 86264 187104
rect 89944 187168 90264 187169
rect 89944 187104 89952 187168
rect 90016 187104 90032 187168
rect 90096 187104 90112 187168
rect 90176 187104 90192 187168
rect 90256 187104 90264 187168
rect 89944 187103 90264 187104
rect 79317 187100 79383 187101
rect 79317 187096 79364 187100
rect 79428 187098 79434 187100
rect 79317 187040 79322 187096
rect 79317 187036 79364 187040
rect 79428 187038 79474 187098
rect 79428 187036 79434 187038
rect 79317 187035 79383 187036
rect 3944 186624 4264 186625
rect 3944 186560 3952 186624
rect 4016 186560 4032 186624
rect 4096 186560 4112 186624
rect 4176 186560 4192 186624
rect 4256 186560 4264 186624
rect 3944 186559 4264 186560
rect 87944 186624 88264 186625
rect 87944 186560 87952 186624
rect 88016 186560 88032 186624
rect 88096 186560 88112 186624
rect 88176 186560 88192 186624
rect 88256 186560 88264 186624
rect 87944 186559 88264 186560
rect 88742 186492 88748 186556
rect 88812 186554 88818 186556
rect 91200 186554 92000 186584
rect 88812 186494 92000 186554
rect 88812 186492 88818 186494
rect 91200 186464 92000 186494
rect 84377 186282 84443 186285
rect 83230 186280 84443 186282
rect 83230 186224 84382 186280
rect 84438 186224 84443 186280
rect 83230 186222 84443 186224
rect 83230 186091 83290 186222
rect 84377 186219 84443 186222
rect 1944 186080 2264 186081
rect 1944 186016 1952 186080
rect 2016 186016 2032 186080
rect 2096 186016 2112 186080
rect 2176 186016 2192 186080
rect 2256 186016 2264 186080
rect 1944 186015 2264 186016
rect 85944 186080 86264 186081
rect 85944 186016 85952 186080
rect 86016 186016 86032 186080
rect 86096 186016 86112 186080
rect 86176 186016 86192 186080
rect 86256 186016 86264 186080
rect 85944 186015 86264 186016
rect 89944 186080 90264 186081
rect 89944 186016 89952 186080
rect 90016 186016 90032 186080
rect 90096 186016 90112 186080
rect 90176 186016 90192 186080
rect 90256 186016 90264 186080
rect 89944 186015 90264 186016
rect 3944 185536 4264 185537
rect 3944 185472 3952 185536
rect 4016 185472 4032 185536
rect 4096 185472 4112 185536
rect 4176 185472 4192 185536
rect 4256 185472 4264 185536
rect 3944 185471 4264 185472
rect 87944 185536 88264 185537
rect 87944 185472 87952 185536
rect 88016 185472 88032 185536
rect 88096 185472 88112 185536
rect 88176 185472 88192 185536
rect 88256 185472 88264 185536
rect 87944 185471 88264 185472
rect 88374 185268 88380 185332
rect 88444 185330 88450 185332
rect 91200 185330 92000 185360
rect 88444 185270 92000 185330
rect 88444 185268 88450 185270
rect 91200 185240 92000 185270
rect 1944 184992 2264 184993
rect 1944 184928 1952 184992
rect 2016 184928 2032 184992
rect 2096 184928 2112 184992
rect 2176 184928 2192 184992
rect 2256 184928 2264 184992
rect 1944 184927 2264 184928
rect 85944 184992 86264 184993
rect 85944 184928 85952 184992
rect 86016 184928 86032 184992
rect 86096 184928 86112 184992
rect 86176 184928 86192 184992
rect 86256 184928 86264 184992
rect 85944 184927 86264 184928
rect 89944 184992 90264 184993
rect 89944 184928 89952 184992
rect 90016 184928 90032 184992
rect 90096 184928 90112 184992
rect 90176 184928 90192 184992
rect 90256 184928 90264 184992
rect 89944 184927 90264 184928
rect 3944 184448 4264 184449
rect 3944 184384 3952 184448
rect 4016 184384 4032 184448
rect 4096 184384 4112 184448
rect 4176 184384 4192 184448
rect 4256 184384 4264 184448
rect 3944 184383 4264 184384
rect 87944 184448 88264 184449
rect 87944 184384 87952 184448
rect 88016 184384 88032 184448
rect 88096 184384 88112 184448
rect 88176 184384 88192 184448
rect 88256 184384 88264 184448
rect 87944 184383 88264 184384
rect 87454 184044 87460 184108
rect 87524 184106 87530 184108
rect 91200 184106 92000 184136
rect 87524 184046 92000 184106
rect 87524 184044 87530 184046
rect 91200 184016 92000 184046
rect 1944 183904 2264 183905
rect 1944 183840 1952 183904
rect 2016 183840 2032 183904
rect 2096 183840 2112 183904
rect 2176 183840 2192 183904
rect 2256 183840 2264 183904
rect 1944 183839 2264 183840
rect 85944 183904 86264 183905
rect 85944 183840 85952 183904
rect 86016 183840 86032 183904
rect 86096 183840 86112 183904
rect 86176 183840 86192 183904
rect 86256 183840 86264 183904
rect 85944 183839 86264 183840
rect 89944 183904 90264 183905
rect 89944 183840 89952 183904
rect 90016 183840 90032 183904
rect 90096 183840 90112 183904
rect 90176 183840 90192 183904
rect 90256 183840 90264 183904
rect 89944 183839 90264 183840
rect 3944 183360 4264 183361
rect 3944 183296 3952 183360
rect 4016 183296 4032 183360
rect 4096 183296 4112 183360
rect 4176 183296 4192 183360
rect 4256 183296 4264 183360
rect 3944 183295 4264 183296
rect 87944 183360 88264 183361
rect 87944 183296 87952 183360
rect 88016 183296 88032 183360
rect 88096 183296 88112 183360
rect 88176 183296 88192 183360
rect 88256 183296 88264 183360
rect 87944 183295 88264 183296
rect 4797 183018 4863 183021
rect 5165 183018 5231 183021
rect 4797 183016 6194 183018
rect 4797 182960 4802 183016
rect 4858 182960 5170 183016
rect 5226 182960 6194 183016
rect 4797 182958 6194 182960
rect 4797 182955 4863 182958
rect 5165 182955 5231 182958
rect 91200 182882 92000 182912
rect 90406 182822 92000 182882
rect 1944 182816 2264 182817
rect 1944 182752 1952 182816
rect 2016 182752 2032 182816
rect 2096 182752 2112 182816
rect 2176 182752 2192 182816
rect 2256 182752 2264 182816
rect 1944 182751 2264 182752
rect 85944 182816 86264 182817
rect 85944 182752 85952 182816
rect 86016 182752 86032 182816
rect 86096 182752 86112 182816
rect 86176 182752 86192 182816
rect 86256 182752 86264 182816
rect 85944 182751 86264 182752
rect 89944 182816 90264 182817
rect 89944 182752 89952 182816
rect 90016 182752 90032 182816
rect 90096 182752 90112 182816
rect 90176 182752 90192 182816
rect 90256 182752 90264 182816
rect 89944 182751 90264 182752
rect 87086 182548 87092 182612
rect 87156 182610 87162 182612
rect 90406 182610 90466 182822
rect 91200 182792 92000 182822
rect 87156 182550 90466 182610
rect 87156 182548 87162 182550
rect 3944 182272 4264 182273
rect 3944 182208 3952 182272
rect 4016 182208 4032 182272
rect 4096 182208 4112 182272
rect 4176 182208 4192 182272
rect 4256 182208 4264 182272
rect 3944 182207 4264 182208
rect 87944 182272 88264 182273
rect 87944 182208 87952 182272
rect 88016 182208 88032 182272
rect 88096 182208 88112 182272
rect 88176 182208 88192 182272
rect 88256 182208 88264 182272
rect 87944 182207 88264 182208
rect 4797 181930 4863 181933
rect 4797 181928 6194 181930
rect 4797 181872 4802 181928
rect 4858 181872 6194 181928
rect 4797 181870 6194 181872
rect 4797 181867 4863 181870
rect 6134 181867 6194 181870
rect 1944 181728 2264 181729
rect 1944 181664 1952 181728
rect 2016 181664 2032 181728
rect 2096 181664 2112 181728
rect 2176 181664 2192 181728
rect 2256 181664 2264 181728
rect 1944 181663 2264 181664
rect 85944 181728 86264 181729
rect 85944 181664 85952 181728
rect 86016 181664 86032 181728
rect 86096 181664 86112 181728
rect 86176 181664 86192 181728
rect 86256 181664 86264 181728
rect 85944 181663 86264 181664
rect 89944 181728 90264 181729
rect 89944 181664 89952 181728
rect 90016 181664 90032 181728
rect 90096 181664 90112 181728
rect 90176 181664 90192 181728
rect 90256 181664 90264 181728
rect 89944 181663 90264 181664
rect 91200 181658 92000 181688
rect 90406 181598 92000 181658
rect 87689 181522 87755 181525
rect 90406 181522 90466 181598
rect 91200 181568 92000 181598
rect 87689 181520 90466 181522
rect 87689 181464 87694 181520
rect 87750 181464 90466 181520
rect 87689 181462 90466 181464
rect 87689 181459 87755 181462
rect 3944 181184 4264 181185
rect 3944 181120 3952 181184
rect 4016 181120 4032 181184
rect 4096 181120 4112 181184
rect 4176 181120 4192 181184
rect 4256 181120 4264 181184
rect 3944 181119 4264 181120
rect 87944 181184 88264 181185
rect 87944 181120 87952 181184
rect 88016 181120 88032 181184
rect 88096 181120 88112 181184
rect 88176 181120 88192 181184
rect 88256 181120 88264 181184
rect 87944 181119 88264 181120
rect 1944 180640 2264 180641
rect 1944 180576 1952 180640
rect 2016 180576 2032 180640
rect 2096 180576 2112 180640
rect 2176 180576 2192 180640
rect 2256 180576 2264 180640
rect 1944 180575 2264 180576
rect 85944 180640 86264 180641
rect 85944 180576 85952 180640
rect 86016 180576 86032 180640
rect 86096 180576 86112 180640
rect 86176 180576 86192 180640
rect 86256 180576 86264 180640
rect 85944 180575 86264 180576
rect 89944 180640 90264 180641
rect 89944 180576 89952 180640
rect 90016 180576 90032 180640
rect 90096 180576 90112 180640
rect 90176 180576 90192 180640
rect 90256 180576 90264 180640
rect 89944 180575 90264 180576
rect 87638 180372 87644 180436
rect 87708 180434 87714 180436
rect 91200 180434 92000 180464
rect 87708 180374 92000 180434
rect 87708 180372 87714 180374
rect 91200 180344 92000 180374
rect 4613 180162 4679 180165
rect 6134 180162 6194 180167
rect 4613 180160 6194 180162
rect 4613 180104 4618 180160
rect 4674 180104 6194 180160
rect 4613 180102 6194 180104
rect 4613 180099 4679 180102
rect 3944 180096 4264 180097
rect 3944 180032 3952 180096
rect 4016 180032 4032 180096
rect 4096 180032 4112 180096
rect 4176 180032 4192 180096
rect 4256 180032 4264 180096
rect 3944 180031 4264 180032
rect 87944 180096 88264 180097
rect 87944 180032 87952 180096
rect 88016 180032 88032 180096
rect 88096 180032 88112 180096
rect 88176 180032 88192 180096
rect 88256 180032 88264 180096
rect 87944 180031 88264 180032
rect 1944 179552 2264 179553
rect 1944 179488 1952 179552
rect 2016 179488 2032 179552
rect 2096 179488 2112 179552
rect 2176 179488 2192 179552
rect 2256 179488 2264 179552
rect 1944 179487 2264 179488
rect 85944 179552 86264 179553
rect 85944 179488 85952 179552
rect 86016 179488 86032 179552
rect 86096 179488 86112 179552
rect 86176 179488 86192 179552
rect 86256 179488 86264 179552
rect 85944 179487 86264 179488
rect 89944 179552 90264 179553
rect 89944 179488 89952 179552
rect 90016 179488 90032 179552
rect 90096 179488 90112 179552
rect 90176 179488 90192 179552
rect 90256 179488 90264 179552
rect 89944 179487 90264 179488
rect 87270 179148 87276 179212
rect 87340 179210 87346 179212
rect 91200 179210 92000 179240
rect 87340 179150 92000 179210
rect 87340 179148 87346 179150
rect 91200 179120 92000 179150
rect 4521 179074 4587 179077
rect 4521 179072 6194 179074
rect 4521 179016 4526 179072
rect 4582 179016 6194 179072
rect 4521 179014 6194 179016
rect 4521 179011 4587 179014
rect 3944 179008 4264 179009
rect 3944 178944 3952 179008
rect 4016 178944 4032 179008
rect 4096 178944 4112 179008
rect 4176 178944 4192 179008
rect 4256 178944 4264 179008
rect 3944 178943 4264 178944
rect 87944 179008 88264 179009
rect 87944 178944 87952 179008
rect 88016 178944 88032 179008
rect 88096 178944 88112 179008
rect 88176 178944 88192 179008
rect 88256 178944 88264 179008
rect 87944 178943 88264 178944
rect 1944 178464 2264 178465
rect 1944 178400 1952 178464
rect 2016 178400 2032 178464
rect 2096 178400 2112 178464
rect 2176 178400 2192 178464
rect 2256 178400 2264 178464
rect 1944 178399 2264 178400
rect 85944 178464 86264 178465
rect 85944 178400 85952 178464
rect 86016 178400 86032 178464
rect 86096 178400 86112 178464
rect 86176 178400 86192 178464
rect 86256 178400 86264 178464
rect 85944 178399 86264 178400
rect 89944 178464 90264 178465
rect 89944 178400 89952 178464
rect 90016 178400 90032 178464
rect 90096 178400 90112 178464
rect 90176 178400 90192 178464
rect 90256 178400 90264 178464
rect 89944 178399 90264 178400
rect 91200 177986 92000 178016
rect 88382 177926 92000 177986
rect 3944 177920 4264 177921
rect 3944 177856 3952 177920
rect 4016 177856 4032 177920
rect 4096 177856 4112 177920
rect 4176 177856 4192 177920
rect 4256 177856 4264 177920
rect 3944 177855 4264 177856
rect 87944 177920 88264 177921
rect 87944 177856 87952 177920
rect 88016 177856 88032 177920
rect 88096 177856 88112 177920
rect 88176 177856 88192 177920
rect 88256 177856 88264 177920
rect 87944 177855 88264 177856
rect 87781 177714 87847 177717
rect 88382 177714 88442 177926
rect 91200 177896 92000 177926
rect 87781 177712 88442 177714
rect 87781 177656 87786 177712
rect 87842 177656 88442 177712
rect 87781 177654 88442 177656
rect 87781 177651 87847 177654
rect 1944 177376 2264 177377
rect 1944 177312 1952 177376
rect 2016 177312 2032 177376
rect 2096 177312 2112 177376
rect 2176 177312 2192 177376
rect 2256 177312 2264 177376
rect 85944 177376 86264 177377
rect 1944 177311 2264 177312
rect 4705 177034 4771 177037
rect 6134 177034 6194 177339
rect 85944 177312 85952 177376
rect 86016 177312 86032 177376
rect 86096 177312 86112 177376
rect 86176 177312 86192 177376
rect 86256 177312 86264 177376
rect 85944 177311 86264 177312
rect 89944 177376 90264 177377
rect 89944 177312 89952 177376
rect 90016 177312 90032 177376
rect 90096 177312 90112 177376
rect 90176 177312 90192 177376
rect 90256 177312 90264 177376
rect 89944 177311 90264 177312
rect 4705 177032 6194 177034
rect 4705 176976 4710 177032
rect 4766 176976 6194 177032
rect 4705 176974 6194 176976
rect 4705 176971 4771 176974
rect 83406 176972 83412 177036
rect 83476 177034 83482 177036
rect 83476 176974 88442 177034
rect 83476 176972 83482 176974
rect 3944 176832 4264 176833
rect 3944 176768 3952 176832
rect 4016 176768 4032 176832
rect 4096 176768 4112 176832
rect 4176 176768 4192 176832
rect 4256 176768 4264 176832
rect 3944 176767 4264 176768
rect 87944 176832 88264 176833
rect 87944 176768 87952 176832
rect 88016 176768 88032 176832
rect 88096 176768 88112 176832
rect 88176 176768 88192 176832
rect 88256 176768 88264 176832
rect 87944 176767 88264 176768
rect 88382 176762 88442 176974
rect 91200 176762 92000 176792
rect 88382 176702 92000 176762
rect 91200 176672 92000 176702
rect 1944 176288 2264 176289
rect 1944 176224 1952 176288
rect 2016 176224 2032 176288
rect 2096 176224 2112 176288
rect 2176 176224 2192 176288
rect 2256 176224 2264 176288
rect 1944 176223 2264 176224
rect 85944 176288 86264 176289
rect 85944 176224 85952 176288
rect 86016 176224 86032 176288
rect 86096 176224 86112 176288
rect 86176 176224 86192 176288
rect 86256 176224 86264 176288
rect 85944 176223 86264 176224
rect 89944 176288 90264 176289
rect 89944 176224 89952 176288
rect 90016 176224 90032 176288
rect 90096 176224 90112 176288
rect 90176 176224 90192 176288
rect 90256 176224 90264 176288
rect 89944 176223 90264 176224
rect 4797 176218 4863 176221
rect 5257 176218 5323 176221
rect 4797 176216 6194 176218
rect 4797 176160 4802 176216
rect 4858 176160 5262 176216
rect 5318 176160 6194 176216
rect 4797 176158 6194 176160
rect 4797 176155 4863 176158
rect 5257 176155 5323 176158
rect 3944 175744 4264 175745
rect 3944 175680 3952 175744
rect 4016 175680 4032 175744
rect 4096 175680 4112 175744
rect 4176 175680 4192 175744
rect 4256 175680 4264 175744
rect 3944 175679 4264 175680
rect 87944 175744 88264 175745
rect 87944 175680 87952 175744
rect 88016 175680 88032 175744
rect 88096 175680 88112 175744
rect 88176 175680 88192 175744
rect 88256 175680 88264 175744
rect 87944 175679 88264 175680
rect 91200 175538 92000 175568
rect 84150 175478 92000 175538
rect 83590 175340 83596 175404
rect 83660 175402 83666 175404
rect 84150 175402 84210 175478
rect 91200 175448 92000 175478
rect 83660 175342 84210 175402
rect 83660 175340 83666 175342
rect 1944 175200 2264 175201
rect 1944 175136 1952 175200
rect 2016 175136 2032 175200
rect 2096 175136 2112 175200
rect 2176 175136 2192 175200
rect 2256 175136 2264 175200
rect 1944 175135 2264 175136
rect 85944 175200 86264 175201
rect 85944 175136 85952 175200
rect 86016 175136 86032 175200
rect 86096 175136 86112 175200
rect 86176 175136 86192 175200
rect 86256 175136 86264 175200
rect 85944 175135 86264 175136
rect 89944 175200 90264 175201
rect 89944 175136 89952 175200
rect 90016 175136 90032 175200
rect 90096 175136 90112 175200
rect 90176 175136 90192 175200
rect 90256 175136 90264 175200
rect 89944 175135 90264 175136
rect 3944 174656 4264 174657
rect 3944 174592 3952 174656
rect 4016 174592 4032 174656
rect 4096 174592 4112 174656
rect 4176 174592 4192 174656
rect 4256 174592 4264 174656
rect 3944 174591 4264 174592
rect 87944 174656 88264 174657
rect 87944 174592 87952 174656
rect 88016 174592 88032 174656
rect 88096 174592 88112 174656
rect 88176 174592 88192 174656
rect 88256 174592 88264 174656
rect 87944 174591 88264 174592
rect 4797 174586 4863 174589
rect 5257 174586 5323 174589
rect 4797 174584 6194 174586
rect 4797 174528 4802 174584
rect 4858 174528 5262 174584
rect 5318 174528 6194 174584
rect 4797 174526 6194 174528
rect 4797 174523 4863 174526
rect 5257 174523 5323 174526
rect 6134 174511 6194 174526
rect 87413 174314 87479 174317
rect 91200 174314 92000 174344
rect 87413 174312 92000 174314
rect 87413 174256 87418 174312
rect 87474 174256 92000 174312
rect 87413 174254 92000 174256
rect 87413 174251 87479 174254
rect 91200 174224 92000 174254
rect 1944 174112 2264 174113
rect 1944 174048 1952 174112
rect 2016 174048 2032 174112
rect 2096 174048 2112 174112
rect 2176 174048 2192 174112
rect 2256 174048 2264 174112
rect 1944 174047 2264 174048
rect 85944 174112 86264 174113
rect 85944 174048 85952 174112
rect 86016 174048 86032 174112
rect 86096 174048 86112 174112
rect 86176 174048 86192 174112
rect 86256 174048 86264 174112
rect 85944 174047 86264 174048
rect 89944 174112 90264 174113
rect 89944 174048 89952 174112
rect 90016 174048 90032 174112
rect 90096 174048 90112 174112
rect 90176 174048 90192 174112
rect 90256 174048 90264 174112
rect 89944 174047 90264 174048
rect 3944 173568 4264 173569
rect 3944 173504 3952 173568
rect 4016 173504 4032 173568
rect 4096 173504 4112 173568
rect 4176 173504 4192 173568
rect 4256 173504 4264 173568
rect 3944 173503 4264 173504
rect 87944 173568 88264 173569
rect 87944 173504 87952 173568
rect 88016 173504 88032 173568
rect 88096 173504 88112 173568
rect 88176 173504 88192 173568
rect 88256 173504 88264 173568
rect 87944 173503 88264 173504
rect 87597 173226 87663 173229
rect 91200 173226 92000 173256
rect 87597 173224 92000 173226
rect 87597 173168 87602 173224
rect 87658 173168 92000 173224
rect 87597 173166 92000 173168
rect 87597 173163 87663 173166
rect 91200 173136 92000 173166
rect 1944 173024 2264 173025
rect 1944 172960 1952 173024
rect 2016 172960 2032 173024
rect 2096 172960 2112 173024
rect 2176 172960 2192 173024
rect 2256 172960 2264 173024
rect 1944 172959 2264 172960
rect 85944 173024 86264 173025
rect 85944 172960 85952 173024
rect 86016 172960 86032 173024
rect 86096 172960 86112 173024
rect 86176 172960 86192 173024
rect 86256 172960 86264 173024
rect 85944 172959 86264 172960
rect 89944 173024 90264 173025
rect 89944 172960 89952 173024
rect 90016 172960 90032 173024
rect 90096 172960 90112 173024
rect 90176 172960 90192 173024
rect 90256 172960 90264 173024
rect 89944 172959 90264 172960
rect 3944 172480 4264 172481
rect 3944 172416 3952 172480
rect 4016 172416 4032 172480
rect 4096 172416 4112 172480
rect 4176 172416 4192 172480
rect 4256 172416 4264 172480
rect 3944 172415 4264 172416
rect 87944 172480 88264 172481
rect 87944 172416 87952 172480
rect 88016 172416 88032 172480
rect 88096 172416 88112 172480
rect 88176 172416 88192 172480
rect 88256 172416 88264 172480
rect 87944 172415 88264 172416
rect 91200 172002 92000 172032
rect 90406 171942 92000 172002
rect 1944 171936 2264 171937
rect 1944 171872 1952 171936
rect 2016 171872 2032 171936
rect 2096 171872 2112 171936
rect 2176 171872 2192 171936
rect 2256 171872 2264 171936
rect 1944 171871 2264 171872
rect 85944 171936 86264 171937
rect 85944 171872 85952 171936
rect 86016 171872 86032 171936
rect 86096 171872 86112 171936
rect 86176 171872 86192 171936
rect 86256 171872 86264 171936
rect 85944 171871 86264 171872
rect 89944 171936 90264 171937
rect 89944 171872 89952 171936
rect 90016 171872 90032 171936
rect 90096 171872 90112 171936
rect 90176 171872 90192 171936
rect 90256 171872 90264 171936
rect 89944 171871 90264 171872
rect 87689 171730 87755 171733
rect 90406 171730 90466 171942
rect 91200 171912 92000 171942
rect 87689 171728 90466 171730
rect 87689 171672 87694 171728
rect 87750 171672 90466 171728
rect 87689 171670 90466 171672
rect 87689 171667 87755 171670
rect 3944 171392 4264 171393
rect 3944 171328 3952 171392
rect 4016 171328 4032 171392
rect 4096 171328 4112 171392
rect 4176 171328 4192 171392
rect 4256 171328 4264 171392
rect 3944 171327 4264 171328
rect 87944 171392 88264 171393
rect 87944 171328 87952 171392
rect 88016 171328 88032 171392
rect 88096 171328 88112 171392
rect 88176 171328 88192 171392
rect 88256 171328 88264 171392
rect 87944 171327 88264 171328
rect 1944 170848 2264 170849
rect 1944 170784 1952 170848
rect 2016 170784 2032 170848
rect 2096 170784 2112 170848
rect 2176 170784 2192 170848
rect 2256 170784 2264 170848
rect 1944 170783 2264 170784
rect 85944 170848 86264 170849
rect 85944 170784 85952 170848
rect 86016 170784 86032 170848
rect 86096 170784 86112 170848
rect 86176 170784 86192 170848
rect 86256 170784 86264 170848
rect 85944 170783 86264 170784
rect 89944 170848 90264 170849
rect 89944 170784 89952 170848
rect 90016 170784 90032 170848
rect 90096 170784 90112 170848
rect 90176 170784 90192 170848
rect 90256 170784 90264 170848
rect 89944 170783 90264 170784
rect 91200 170778 92000 170808
rect 90406 170718 92000 170778
rect 3944 170304 4264 170305
rect 3944 170240 3952 170304
rect 4016 170240 4032 170304
rect 4096 170240 4112 170304
rect 4176 170240 4192 170304
rect 4256 170240 4264 170304
rect 3944 170239 4264 170240
rect 87944 170304 88264 170305
rect 87944 170240 87952 170304
rect 88016 170240 88032 170304
rect 88096 170240 88112 170304
rect 88176 170240 88192 170304
rect 88256 170240 88264 170304
rect 87944 170239 88264 170240
rect 90406 170098 90466 170718
rect 91200 170688 92000 170718
rect 84150 170038 90466 170098
rect 84150 169965 84210 170038
rect 84101 169960 84210 169965
rect 84101 169904 84106 169960
rect 84162 169904 84210 169960
rect 84101 169902 84210 169904
rect 84101 169899 84167 169902
rect 1944 169760 2264 169761
rect 1944 169696 1952 169760
rect 2016 169696 2032 169760
rect 2096 169696 2112 169760
rect 2176 169696 2192 169760
rect 2256 169696 2264 169760
rect 1944 169695 2264 169696
rect 85944 169760 86264 169761
rect 85944 169696 85952 169760
rect 86016 169696 86032 169760
rect 86096 169696 86112 169760
rect 86176 169696 86192 169760
rect 86256 169696 86264 169760
rect 85944 169695 86264 169696
rect 89944 169760 90264 169761
rect 89944 169696 89952 169760
rect 90016 169696 90032 169760
rect 90096 169696 90112 169760
rect 90176 169696 90192 169760
rect 90256 169696 90264 169760
rect 89944 169695 90264 169696
rect 87873 169554 87939 169557
rect 91200 169554 92000 169584
rect 87873 169552 92000 169554
rect 87873 169496 87878 169552
rect 87934 169496 92000 169552
rect 87873 169494 92000 169496
rect 87873 169491 87939 169494
rect 91200 169464 92000 169494
rect 3944 169216 4264 169217
rect 3944 169152 3952 169216
rect 4016 169152 4032 169216
rect 4096 169152 4112 169216
rect 4176 169152 4192 169216
rect 4256 169152 4264 169216
rect 3944 169151 4264 169152
rect 87944 169216 88264 169217
rect 87944 169152 87952 169216
rect 88016 169152 88032 169216
rect 88096 169152 88112 169216
rect 88176 169152 88192 169216
rect 88256 169152 88264 169216
rect 87944 169151 88264 169152
rect 1944 168672 2264 168673
rect 1944 168608 1952 168672
rect 2016 168608 2032 168672
rect 2096 168608 2112 168672
rect 2176 168608 2192 168672
rect 2256 168608 2264 168672
rect 1944 168607 2264 168608
rect 85944 168672 86264 168673
rect 85944 168608 85952 168672
rect 86016 168608 86032 168672
rect 86096 168608 86112 168672
rect 86176 168608 86192 168672
rect 86256 168608 86264 168672
rect 85944 168607 86264 168608
rect 89944 168672 90264 168673
rect 89944 168608 89952 168672
rect 90016 168608 90032 168672
rect 90096 168608 90112 168672
rect 90176 168608 90192 168672
rect 90256 168608 90264 168672
rect 89944 168607 90264 168608
rect 87045 168330 87111 168333
rect 91200 168330 92000 168360
rect 87045 168328 92000 168330
rect 87045 168272 87050 168328
rect 87106 168272 92000 168328
rect 87045 168270 92000 168272
rect 87045 168267 87111 168270
rect 91200 168240 92000 168270
rect 3944 168128 4264 168129
rect 3944 168064 3952 168128
rect 4016 168064 4032 168128
rect 4096 168064 4112 168128
rect 4176 168064 4192 168128
rect 4256 168064 4264 168128
rect 3944 168063 4264 168064
rect 87944 168128 88264 168129
rect 87944 168064 87952 168128
rect 88016 168064 88032 168128
rect 88096 168064 88112 168128
rect 88176 168064 88192 168128
rect 88256 168064 88264 168128
rect 87944 168063 88264 168064
rect 1944 167584 2264 167585
rect 1944 167520 1952 167584
rect 2016 167520 2032 167584
rect 2096 167520 2112 167584
rect 2176 167520 2192 167584
rect 2256 167520 2264 167584
rect 1944 167519 2264 167520
rect 85944 167584 86264 167585
rect 85944 167520 85952 167584
rect 86016 167520 86032 167584
rect 86096 167520 86112 167584
rect 86176 167520 86192 167584
rect 86256 167520 86264 167584
rect 85944 167519 86264 167520
rect 89944 167584 90264 167585
rect 89944 167520 89952 167584
rect 90016 167520 90032 167584
rect 90096 167520 90112 167584
rect 90176 167520 90192 167584
rect 90256 167520 90264 167584
rect 89944 167519 90264 167520
rect 83774 167316 83780 167380
rect 83844 167378 83850 167380
rect 83844 167318 88442 167378
rect 83844 167316 83850 167318
rect 88382 167106 88442 167318
rect 91200 167106 92000 167136
rect 88382 167046 92000 167106
rect 3944 167040 4264 167041
rect 3944 166976 3952 167040
rect 4016 166976 4032 167040
rect 4096 166976 4112 167040
rect 4176 166976 4192 167040
rect 4256 166976 4264 167040
rect 3944 166975 4264 166976
rect 87944 167040 88264 167041
rect 87944 166976 87952 167040
rect 88016 166976 88032 167040
rect 88096 166976 88112 167040
rect 88176 166976 88192 167040
rect 88256 166976 88264 167040
rect 91200 167016 92000 167046
rect 87944 166975 88264 166976
rect 1944 166496 2264 166497
rect 1944 166432 1952 166496
rect 2016 166432 2032 166496
rect 2096 166432 2112 166496
rect 2176 166432 2192 166496
rect 2256 166432 2264 166496
rect 1944 166431 2264 166432
rect 85944 166496 86264 166497
rect 85944 166432 85952 166496
rect 86016 166432 86032 166496
rect 86096 166432 86112 166496
rect 86176 166432 86192 166496
rect 86256 166432 86264 166496
rect 85944 166431 86264 166432
rect 89944 166496 90264 166497
rect 89944 166432 89952 166496
rect 90016 166432 90032 166496
rect 90096 166432 90112 166496
rect 90176 166432 90192 166496
rect 90256 166432 90264 166496
rect 89944 166431 90264 166432
rect 3944 165952 4264 165953
rect 3944 165888 3952 165952
rect 4016 165888 4032 165952
rect 4096 165888 4112 165952
rect 4176 165888 4192 165952
rect 4256 165888 4264 165952
rect 3944 165887 4264 165888
rect 87944 165952 88264 165953
rect 87944 165888 87952 165952
rect 88016 165888 88032 165952
rect 88096 165888 88112 165952
rect 88176 165888 88192 165952
rect 88256 165888 88264 165952
rect 87944 165887 88264 165888
rect 91200 165882 92000 165912
rect 88382 165822 92000 165882
rect 87505 165746 87571 165749
rect 88382 165746 88442 165822
rect 91200 165792 92000 165822
rect 87505 165744 88442 165746
rect 87505 165688 87510 165744
rect 87566 165688 88442 165744
rect 87505 165686 88442 165688
rect 87505 165683 87571 165686
rect 1944 165408 2264 165409
rect 1944 165344 1952 165408
rect 2016 165344 2032 165408
rect 2096 165344 2112 165408
rect 2176 165344 2192 165408
rect 2256 165344 2264 165408
rect 1944 165343 2264 165344
rect 85944 165408 86264 165409
rect 85944 165344 85952 165408
rect 86016 165344 86032 165408
rect 86096 165344 86112 165408
rect 86176 165344 86192 165408
rect 86256 165344 86264 165408
rect 85944 165343 86264 165344
rect 89944 165408 90264 165409
rect 89944 165344 89952 165408
rect 90016 165344 90032 165408
rect 90096 165344 90112 165408
rect 90176 165344 90192 165408
rect 90256 165344 90264 165408
rect 89944 165343 90264 165344
rect 3944 164864 4264 164865
rect 3944 164800 3952 164864
rect 4016 164800 4032 164864
rect 4096 164800 4112 164864
rect 4176 164800 4192 164864
rect 4256 164800 4264 164864
rect 3944 164799 4264 164800
rect 87944 164864 88264 164865
rect 87944 164800 87952 164864
rect 88016 164800 88032 164864
rect 88096 164800 88112 164864
rect 88176 164800 88192 164864
rect 88256 164800 88264 164864
rect 87944 164799 88264 164800
rect 87873 164658 87939 164661
rect 91200 164658 92000 164688
rect 87873 164656 92000 164658
rect 87873 164600 87878 164656
rect 87934 164600 92000 164656
rect 87873 164598 92000 164600
rect 87873 164595 87939 164598
rect 91200 164568 92000 164598
rect 1944 164320 2264 164321
rect 1944 164256 1952 164320
rect 2016 164256 2032 164320
rect 2096 164256 2112 164320
rect 2176 164256 2192 164320
rect 2256 164256 2264 164320
rect 1944 164255 2264 164256
rect 85944 164320 86264 164321
rect 85944 164256 85952 164320
rect 86016 164256 86032 164320
rect 86096 164256 86112 164320
rect 86176 164256 86192 164320
rect 86256 164256 86264 164320
rect 85944 164255 86264 164256
rect 89944 164320 90264 164321
rect 89944 164256 89952 164320
rect 90016 164256 90032 164320
rect 90096 164256 90112 164320
rect 90176 164256 90192 164320
rect 90256 164256 90264 164320
rect 89944 164255 90264 164256
rect 84101 164114 84167 164117
rect 84326 164114 84332 164116
rect 84101 164112 84332 164114
rect 84101 164056 84106 164112
rect 84162 164056 84332 164112
rect 84101 164054 84332 164056
rect 84101 164051 84167 164054
rect 84326 164052 84332 164054
rect 84396 164052 84402 164116
rect 3944 163776 4264 163777
rect 3944 163712 3952 163776
rect 4016 163712 4032 163776
rect 4096 163712 4112 163776
rect 4176 163712 4192 163776
rect 4256 163712 4264 163776
rect 3944 163711 4264 163712
rect 87944 163776 88264 163777
rect 87944 163712 87952 163776
rect 88016 163712 88032 163776
rect 88096 163712 88112 163776
rect 88176 163712 88192 163776
rect 88256 163712 88264 163776
rect 87944 163711 88264 163712
rect 87873 163434 87939 163437
rect 91200 163434 92000 163464
rect 87873 163432 92000 163434
rect 87873 163376 87878 163432
rect 87934 163376 92000 163432
rect 87873 163374 92000 163376
rect 87873 163371 87939 163374
rect 91200 163344 92000 163374
rect 1944 163232 2264 163233
rect 1944 163168 1952 163232
rect 2016 163168 2032 163232
rect 2096 163168 2112 163232
rect 2176 163168 2192 163232
rect 2256 163168 2264 163232
rect 1944 163167 2264 163168
rect 85944 163232 86264 163233
rect 85944 163168 85952 163232
rect 86016 163168 86032 163232
rect 86096 163168 86112 163232
rect 86176 163168 86192 163232
rect 86256 163168 86264 163232
rect 85944 163167 86264 163168
rect 89944 163232 90264 163233
rect 89944 163168 89952 163232
rect 90016 163168 90032 163232
rect 90096 163168 90112 163232
rect 90176 163168 90192 163232
rect 90256 163168 90264 163232
rect 89944 163167 90264 163168
rect 3944 162688 4264 162689
rect 3944 162624 3952 162688
rect 4016 162624 4032 162688
rect 4096 162624 4112 162688
rect 4176 162624 4192 162688
rect 4256 162624 4264 162688
rect 3944 162623 4264 162624
rect 87944 162688 88264 162689
rect 87944 162624 87952 162688
rect 88016 162624 88032 162688
rect 88096 162624 88112 162688
rect 88176 162624 88192 162688
rect 88256 162624 88264 162688
rect 87944 162623 88264 162624
rect 91200 162210 92000 162240
rect 90406 162150 92000 162210
rect 1944 162144 2264 162145
rect 1944 162080 1952 162144
rect 2016 162080 2032 162144
rect 2096 162080 2112 162144
rect 2176 162080 2192 162144
rect 2256 162080 2264 162144
rect 1944 162079 2264 162080
rect 85944 162144 86264 162145
rect 85944 162080 85952 162144
rect 86016 162080 86032 162144
rect 86096 162080 86112 162144
rect 86176 162080 86192 162144
rect 86256 162080 86264 162144
rect 85944 162079 86264 162080
rect 89944 162144 90264 162145
rect 89944 162080 89952 162144
rect 90016 162080 90032 162144
rect 90096 162080 90112 162144
rect 90176 162080 90192 162144
rect 90256 162080 90264 162144
rect 89944 162079 90264 162080
rect 86350 161876 86356 161940
rect 86420 161938 86426 161940
rect 90406 161938 90466 162150
rect 91200 162120 92000 162150
rect 86420 161878 90466 161938
rect 86420 161876 86426 161878
rect 85113 161804 85179 161805
rect 85062 161802 85068 161804
rect 85022 161742 85068 161802
rect 85132 161800 85179 161804
rect 85174 161744 85179 161800
rect 85062 161740 85068 161742
rect 85132 161740 85179 161744
rect 85113 161739 85179 161740
rect 3944 161600 4264 161601
rect 3944 161536 3952 161600
rect 4016 161536 4032 161600
rect 4096 161536 4112 161600
rect 4176 161536 4192 161600
rect 4256 161536 4264 161600
rect 3944 161535 4264 161536
rect 87944 161600 88264 161601
rect 87944 161536 87952 161600
rect 88016 161536 88032 161600
rect 88096 161536 88112 161600
rect 88176 161536 88192 161600
rect 88256 161536 88264 161600
rect 87944 161535 88264 161536
rect 1944 161056 2264 161057
rect 1944 160992 1952 161056
rect 2016 160992 2032 161056
rect 2096 160992 2112 161056
rect 2176 160992 2192 161056
rect 2256 160992 2264 161056
rect 1944 160991 2264 160992
rect 85944 161056 86264 161057
rect 85944 160992 85952 161056
rect 86016 160992 86032 161056
rect 86096 160992 86112 161056
rect 86176 160992 86192 161056
rect 86256 160992 86264 161056
rect 85944 160991 86264 160992
rect 89944 161056 90264 161057
rect 89944 160992 89952 161056
rect 90016 160992 90032 161056
rect 90096 160992 90112 161056
rect 90176 160992 90192 161056
rect 90256 160992 90264 161056
rect 89944 160991 90264 160992
rect 91200 160986 92000 161016
rect 90406 160926 92000 160986
rect 87873 160850 87939 160853
rect 90406 160850 90466 160926
rect 91200 160896 92000 160926
rect 87873 160848 90466 160850
rect 87873 160792 87878 160848
rect 87934 160792 90466 160848
rect 87873 160790 90466 160792
rect 87873 160787 87939 160790
rect 3944 160512 4264 160513
rect 3944 160448 3952 160512
rect 4016 160448 4032 160512
rect 4096 160448 4112 160512
rect 4176 160448 4192 160512
rect 4256 160448 4264 160512
rect 3944 160447 4264 160448
rect 87944 160512 88264 160513
rect 87944 160448 87952 160512
rect 88016 160448 88032 160512
rect 88096 160448 88112 160512
rect 88176 160448 88192 160512
rect 88256 160448 88264 160512
rect 87944 160447 88264 160448
rect 1944 159968 2264 159969
rect 1944 159904 1952 159968
rect 2016 159904 2032 159968
rect 2096 159904 2112 159968
rect 2176 159904 2192 159968
rect 2256 159904 2264 159968
rect 1944 159903 2264 159904
rect 85944 159968 86264 159969
rect 85944 159904 85952 159968
rect 86016 159904 86032 159968
rect 86096 159904 86112 159968
rect 86176 159904 86192 159968
rect 86256 159904 86264 159968
rect 85944 159903 86264 159904
rect 89944 159968 90264 159969
rect 89944 159904 89952 159968
rect 90016 159904 90032 159968
rect 90096 159904 90112 159968
rect 90176 159904 90192 159968
rect 90256 159904 90264 159968
rect 89944 159903 90264 159904
rect 87413 159762 87479 159765
rect 91200 159762 92000 159792
rect 87413 159760 92000 159762
rect 87413 159704 87418 159760
rect 87474 159704 92000 159760
rect 87413 159702 92000 159704
rect 87413 159699 87479 159702
rect 91200 159672 92000 159702
rect 3944 159424 4264 159425
rect 3944 159360 3952 159424
rect 4016 159360 4032 159424
rect 4096 159360 4112 159424
rect 4176 159360 4192 159424
rect 4256 159360 4264 159424
rect 3944 159359 4264 159360
rect 87944 159424 88264 159425
rect 87944 159360 87952 159424
rect 88016 159360 88032 159424
rect 88096 159360 88112 159424
rect 88176 159360 88192 159424
rect 88256 159360 88264 159424
rect 87944 159359 88264 159360
rect 1944 158880 2264 158881
rect 1944 158816 1952 158880
rect 2016 158816 2032 158880
rect 2096 158816 2112 158880
rect 2176 158816 2192 158880
rect 2256 158816 2264 158880
rect 1944 158815 2264 158816
rect 85944 158880 86264 158881
rect 85944 158816 85952 158880
rect 86016 158816 86032 158880
rect 86096 158816 86112 158880
rect 86176 158816 86192 158880
rect 86256 158816 86264 158880
rect 85944 158815 86264 158816
rect 89944 158880 90264 158881
rect 89944 158816 89952 158880
rect 90016 158816 90032 158880
rect 90096 158816 90112 158880
rect 90176 158816 90192 158880
rect 90256 158816 90264 158880
rect 89944 158815 90264 158816
rect 86585 158538 86651 158541
rect 91200 158538 92000 158568
rect 86585 158536 92000 158538
rect 86585 158480 86590 158536
rect 86646 158480 92000 158536
rect 86585 158478 92000 158480
rect 86585 158475 86651 158478
rect 91200 158448 92000 158478
rect 3944 158336 4264 158337
rect 3944 158272 3952 158336
rect 4016 158272 4032 158336
rect 4096 158272 4112 158336
rect 4176 158272 4192 158336
rect 4256 158272 4264 158336
rect 3944 158271 4264 158272
rect 87944 158336 88264 158337
rect 87944 158272 87952 158336
rect 88016 158272 88032 158336
rect 88096 158272 88112 158336
rect 88176 158272 88192 158336
rect 88256 158272 88264 158336
rect 87944 158271 88264 158272
rect 1944 157792 2264 157793
rect 1944 157728 1952 157792
rect 2016 157728 2032 157792
rect 2096 157728 2112 157792
rect 2176 157728 2192 157792
rect 2256 157728 2264 157792
rect 1944 157727 2264 157728
rect 85944 157792 86264 157793
rect 85944 157728 85952 157792
rect 86016 157728 86032 157792
rect 86096 157728 86112 157792
rect 86176 157728 86192 157792
rect 86256 157728 86264 157792
rect 85944 157727 86264 157728
rect 89944 157792 90264 157793
rect 89944 157728 89952 157792
rect 90016 157728 90032 157792
rect 90096 157728 90112 157792
rect 90176 157728 90192 157792
rect 90256 157728 90264 157792
rect 89944 157727 90264 157728
rect 91200 157314 92000 157344
rect 88382 157254 92000 157314
rect 3944 157248 4264 157249
rect 3944 157184 3952 157248
rect 4016 157184 4032 157248
rect 4096 157184 4112 157248
rect 4176 157184 4192 157248
rect 4256 157184 4264 157248
rect 3944 157183 4264 157184
rect 87944 157248 88264 157249
rect 87944 157184 87952 157248
rect 88016 157184 88032 157248
rect 88096 157184 88112 157248
rect 88176 157184 88192 157248
rect 88256 157184 88264 157248
rect 87944 157183 88264 157184
rect 87321 157042 87387 157045
rect 88382 157042 88442 157254
rect 91200 157224 92000 157254
rect 87321 157040 88442 157042
rect 87321 156984 87326 157040
rect 87382 156984 88442 157040
rect 87321 156982 88442 156984
rect 87321 156979 87387 156982
rect 1944 156704 2264 156705
rect 1944 156640 1952 156704
rect 2016 156640 2032 156704
rect 2096 156640 2112 156704
rect 2176 156640 2192 156704
rect 2256 156640 2264 156704
rect 1944 156639 2264 156640
rect 85944 156704 86264 156705
rect 85944 156640 85952 156704
rect 86016 156640 86032 156704
rect 86096 156640 86112 156704
rect 86176 156640 86192 156704
rect 86256 156640 86264 156704
rect 85944 156639 86264 156640
rect 89944 156704 90264 156705
rect 89944 156640 89952 156704
rect 90016 156640 90032 156704
rect 90096 156640 90112 156704
rect 90176 156640 90192 156704
rect 90256 156640 90264 156704
rect 89944 156639 90264 156640
rect 85798 156300 85804 156364
rect 85868 156362 85874 156364
rect 85868 156302 88442 156362
rect 85868 156300 85874 156302
rect 3944 156160 4264 156161
rect 3944 156096 3952 156160
rect 4016 156096 4032 156160
rect 4096 156096 4112 156160
rect 4176 156096 4192 156160
rect 4256 156096 4264 156160
rect 3944 156095 4264 156096
rect 87944 156160 88264 156161
rect 87944 156096 87952 156160
rect 88016 156096 88032 156160
rect 88096 156096 88112 156160
rect 88176 156096 88192 156160
rect 88256 156096 88264 156160
rect 87944 156095 88264 156096
rect 88382 156090 88442 156302
rect 91200 156090 92000 156120
rect 88382 156030 92000 156090
rect 91200 156000 92000 156030
rect 1944 155616 2264 155617
rect 1944 155552 1952 155616
rect 2016 155552 2032 155616
rect 2096 155552 2112 155616
rect 2176 155552 2192 155616
rect 2256 155552 2264 155616
rect 1944 155551 2264 155552
rect 85944 155616 86264 155617
rect 85944 155552 85952 155616
rect 86016 155552 86032 155616
rect 86096 155552 86112 155616
rect 86176 155552 86192 155616
rect 86256 155552 86264 155616
rect 85944 155551 86264 155552
rect 89944 155616 90264 155617
rect 89944 155552 89952 155616
rect 90016 155552 90032 155616
rect 90096 155552 90112 155616
rect 90176 155552 90192 155616
rect 90256 155552 90264 155616
rect 89944 155551 90264 155552
rect 3944 155072 4264 155073
rect 3944 155008 3952 155072
rect 4016 155008 4032 155072
rect 4096 155008 4112 155072
rect 4176 155008 4192 155072
rect 4256 155008 4264 155072
rect 3944 155007 4264 155008
rect 87944 155072 88264 155073
rect 87944 155008 87952 155072
rect 88016 155008 88032 155072
rect 88096 155008 88112 155072
rect 88176 155008 88192 155072
rect 88256 155008 88264 155072
rect 87944 155007 88264 155008
rect 87137 154866 87203 154869
rect 91200 154866 92000 154896
rect 87137 154864 92000 154866
rect 87137 154808 87142 154864
rect 87198 154808 92000 154864
rect 87137 154806 92000 154808
rect 87137 154803 87203 154806
rect 91200 154776 92000 154806
rect 1944 154528 2264 154529
rect 1944 154464 1952 154528
rect 2016 154464 2032 154528
rect 2096 154464 2112 154528
rect 2176 154464 2192 154528
rect 2256 154464 2264 154528
rect 1944 154463 2264 154464
rect 85944 154528 86264 154529
rect 85944 154464 85952 154528
rect 86016 154464 86032 154528
rect 86096 154464 86112 154528
rect 86176 154464 86192 154528
rect 86256 154464 86264 154528
rect 85944 154463 86264 154464
rect 89944 154528 90264 154529
rect 89944 154464 89952 154528
rect 90016 154464 90032 154528
rect 90096 154464 90112 154528
rect 90176 154464 90192 154528
rect 90256 154464 90264 154528
rect 89944 154463 90264 154464
rect 82537 154050 82603 154053
rect 84326 154050 84332 154052
rect 82537 154048 84332 154050
rect 82537 153992 82542 154048
rect 82598 153992 84332 154048
rect 82537 153990 84332 153992
rect 82537 153987 82603 153990
rect 84326 153988 84332 153990
rect 84396 153988 84402 154052
rect 3944 153984 4264 153985
rect 3944 153920 3952 153984
rect 4016 153920 4032 153984
rect 4096 153920 4112 153984
rect 4176 153920 4192 153984
rect 4256 153920 4264 153984
rect 3944 153919 4264 153920
rect 87944 153984 88264 153985
rect 87944 153920 87952 153984
rect 88016 153920 88032 153984
rect 88096 153920 88112 153984
rect 88176 153920 88192 153984
rect 88256 153920 88264 153984
rect 87944 153919 88264 153920
rect 86534 153716 86540 153780
rect 86604 153778 86610 153780
rect 91200 153778 92000 153808
rect 86604 153718 92000 153778
rect 86604 153716 86610 153718
rect 91200 153688 92000 153718
rect 1944 153440 2264 153441
rect 1944 153376 1952 153440
rect 2016 153376 2032 153440
rect 2096 153376 2112 153440
rect 2176 153376 2192 153440
rect 2256 153376 2264 153440
rect 1944 153375 2264 153376
rect 85944 153440 86264 153441
rect 85944 153376 85952 153440
rect 86016 153376 86032 153440
rect 86096 153376 86112 153440
rect 86176 153376 86192 153440
rect 86256 153376 86264 153440
rect 85944 153375 86264 153376
rect 89944 153440 90264 153441
rect 89944 153376 89952 153440
rect 90016 153376 90032 153440
rect 90096 153376 90112 153440
rect 90176 153376 90192 153440
rect 90256 153376 90264 153440
rect 89944 153375 90264 153376
rect 3944 152896 4264 152897
rect 3944 152832 3952 152896
rect 4016 152832 4032 152896
rect 4096 152832 4112 152896
rect 4176 152832 4192 152896
rect 4256 152832 4264 152896
rect 3944 152831 4264 152832
rect 87944 152896 88264 152897
rect 87944 152832 87952 152896
rect 88016 152832 88032 152896
rect 88096 152832 88112 152896
rect 88176 152832 88192 152896
rect 88256 152832 88264 152896
rect 87944 152831 88264 152832
rect 86769 152554 86835 152557
rect 91200 152554 92000 152584
rect 86769 152552 92000 152554
rect 86769 152496 86774 152552
rect 86830 152496 92000 152552
rect 86769 152494 92000 152496
rect 86769 152491 86835 152494
rect 91200 152464 92000 152494
rect 1944 152352 2264 152353
rect 1944 152288 1952 152352
rect 2016 152288 2032 152352
rect 2096 152288 2112 152352
rect 2176 152288 2192 152352
rect 2256 152288 2264 152352
rect 1944 152287 2264 152288
rect 85944 152352 86264 152353
rect 85944 152288 85952 152352
rect 86016 152288 86032 152352
rect 86096 152288 86112 152352
rect 86176 152288 86192 152352
rect 86256 152288 86264 152352
rect 85944 152287 86264 152288
rect 89944 152352 90264 152353
rect 89944 152288 89952 152352
rect 90016 152288 90032 152352
rect 90096 152288 90112 152352
rect 90176 152288 90192 152352
rect 90256 152288 90264 152352
rect 89944 152287 90264 152288
rect 3944 151808 4264 151809
rect 3944 151744 3952 151808
rect 4016 151744 4032 151808
rect 4096 151744 4112 151808
rect 4176 151744 4192 151808
rect 4256 151744 4264 151808
rect 3944 151743 4264 151744
rect 87944 151808 88264 151809
rect 87944 151744 87952 151808
rect 88016 151744 88032 151808
rect 88096 151744 88112 151808
rect 88176 151744 88192 151808
rect 88256 151744 88264 151808
rect 87944 151743 88264 151744
rect 91200 151330 92000 151360
rect 90406 151270 92000 151330
rect 1944 151264 2264 151265
rect 1944 151200 1952 151264
rect 2016 151200 2032 151264
rect 2096 151200 2112 151264
rect 2176 151200 2192 151264
rect 2256 151200 2264 151264
rect 1944 151199 2264 151200
rect 85944 151264 86264 151265
rect 85944 151200 85952 151264
rect 86016 151200 86032 151264
rect 86096 151200 86112 151264
rect 86176 151200 86192 151264
rect 86256 151200 86264 151264
rect 85944 151199 86264 151200
rect 89944 151264 90264 151265
rect 89944 151200 89952 151264
rect 90016 151200 90032 151264
rect 90096 151200 90112 151264
rect 90176 151200 90192 151264
rect 90256 151200 90264 151264
rect 89944 151199 90264 151200
rect 86677 151058 86743 151061
rect 90406 151058 90466 151270
rect 91200 151240 92000 151270
rect 86677 151056 90466 151058
rect 86677 151000 86682 151056
rect 86738 151000 90466 151056
rect 86677 150998 90466 151000
rect 86677 150995 86743 150998
rect 3944 150720 4264 150721
rect 3944 150656 3952 150720
rect 4016 150656 4032 150720
rect 4096 150656 4112 150720
rect 4176 150656 4192 150720
rect 4256 150656 4264 150720
rect 3944 150655 4264 150656
rect 87944 150720 88264 150721
rect 87944 150656 87952 150720
rect 88016 150656 88032 150720
rect 88096 150656 88112 150720
rect 88176 150656 88192 150720
rect 88256 150656 88264 150720
rect 87944 150655 88264 150656
rect 1944 150176 2264 150177
rect 1944 150112 1952 150176
rect 2016 150112 2032 150176
rect 2096 150112 2112 150176
rect 2176 150112 2192 150176
rect 2256 150112 2264 150176
rect 1944 150111 2264 150112
rect 85944 150176 86264 150177
rect 85944 150112 85952 150176
rect 86016 150112 86032 150176
rect 86096 150112 86112 150176
rect 86176 150112 86192 150176
rect 86256 150112 86264 150176
rect 85944 150111 86264 150112
rect 89944 150176 90264 150177
rect 89944 150112 89952 150176
rect 90016 150112 90032 150176
rect 90096 150112 90112 150176
rect 90176 150112 90192 150176
rect 90256 150112 90264 150176
rect 89944 150111 90264 150112
rect 91200 150106 92000 150136
rect 90406 150046 92000 150106
rect 87229 149970 87295 149973
rect 90406 149970 90466 150046
rect 91200 150016 92000 150046
rect 87229 149968 90466 149970
rect 87229 149912 87234 149968
rect 87290 149912 90466 149968
rect 87229 149910 90466 149912
rect 87229 149907 87295 149910
rect 3944 149632 4264 149633
rect 3944 149568 3952 149632
rect 4016 149568 4032 149632
rect 4096 149568 4112 149632
rect 4176 149568 4192 149632
rect 4256 149568 4264 149632
rect 3944 149567 4264 149568
rect 87944 149632 88264 149633
rect 87944 149568 87952 149632
rect 88016 149568 88032 149632
rect 88096 149568 88112 149632
rect 88176 149568 88192 149632
rect 88256 149568 88264 149632
rect 87944 149567 88264 149568
rect 1944 149088 2264 149089
rect 1944 149024 1952 149088
rect 2016 149024 2032 149088
rect 2096 149024 2112 149088
rect 2176 149024 2192 149088
rect 2256 149024 2264 149088
rect 1944 149023 2264 149024
rect 85944 149088 86264 149089
rect 85944 149024 85952 149088
rect 86016 149024 86032 149088
rect 86096 149024 86112 149088
rect 86176 149024 86192 149088
rect 86256 149024 86264 149088
rect 85944 149023 86264 149024
rect 89944 149088 90264 149089
rect 89944 149024 89952 149088
rect 90016 149024 90032 149088
rect 90096 149024 90112 149088
rect 90176 149024 90192 149088
rect 90256 149024 90264 149088
rect 89944 149023 90264 149024
rect 86953 148882 87019 148885
rect 91200 148882 92000 148912
rect 86953 148880 92000 148882
rect 86953 148824 86958 148880
rect 87014 148824 92000 148880
rect 86953 148822 92000 148824
rect 86953 148819 87019 148822
rect 91200 148792 92000 148822
rect 3944 148544 4264 148545
rect 3944 148480 3952 148544
rect 4016 148480 4032 148544
rect 4096 148480 4112 148544
rect 4176 148480 4192 148544
rect 4256 148480 4264 148544
rect 3944 148479 4264 148480
rect 87944 148544 88264 148545
rect 87944 148480 87952 148544
rect 88016 148480 88032 148544
rect 88096 148480 88112 148544
rect 88176 148480 88192 148544
rect 88256 148480 88264 148544
rect 87944 148479 88264 148480
rect 1944 148000 2264 148001
rect 1944 147936 1952 148000
rect 2016 147936 2032 148000
rect 2096 147936 2112 148000
rect 2176 147936 2192 148000
rect 2256 147936 2264 148000
rect 1944 147935 2264 147936
rect 85944 148000 86264 148001
rect 85944 147936 85952 148000
rect 86016 147936 86032 148000
rect 86096 147936 86112 148000
rect 86176 147936 86192 148000
rect 86256 147936 86264 148000
rect 85944 147935 86264 147936
rect 89944 148000 90264 148001
rect 89944 147936 89952 148000
rect 90016 147936 90032 148000
rect 90096 147936 90112 148000
rect 90176 147936 90192 148000
rect 90256 147936 90264 148000
rect 89944 147935 90264 147936
rect 86902 147596 86908 147660
rect 86972 147658 86978 147660
rect 91200 147658 92000 147688
rect 86972 147598 92000 147658
rect 86972 147596 86978 147598
rect 91200 147568 92000 147598
rect 3944 147456 4264 147457
rect 3944 147392 3952 147456
rect 4016 147392 4032 147456
rect 4096 147392 4112 147456
rect 4176 147392 4192 147456
rect 4256 147392 4264 147456
rect 3944 147391 4264 147392
rect 87944 147456 88264 147457
rect 87944 147392 87952 147456
rect 88016 147392 88032 147456
rect 88096 147392 88112 147456
rect 88176 147392 88192 147456
rect 88256 147392 88264 147456
rect 87944 147391 88264 147392
rect 1944 146912 2264 146913
rect 1944 146848 1952 146912
rect 2016 146848 2032 146912
rect 2096 146848 2112 146912
rect 2176 146848 2192 146912
rect 2256 146848 2264 146912
rect 1944 146847 2264 146848
rect 85944 146912 86264 146913
rect 85944 146848 85952 146912
rect 86016 146848 86032 146912
rect 86096 146848 86112 146912
rect 86176 146848 86192 146912
rect 86256 146848 86264 146912
rect 85944 146847 86264 146848
rect 89944 146912 90264 146913
rect 89944 146848 89952 146912
rect 90016 146848 90032 146912
rect 90096 146848 90112 146912
rect 90176 146848 90192 146912
rect 90256 146848 90264 146912
rect 89944 146847 90264 146848
rect 87045 146570 87111 146573
rect 87045 146568 88442 146570
rect 87045 146512 87050 146568
rect 87106 146512 88442 146568
rect 87045 146510 88442 146512
rect 87045 146507 87111 146510
rect 88382 146434 88442 146510
rect 91200 146434 92000 146464
rect 88382 146374 92000 146434
rect 3944 146368 4264 146369
rect 3944 146304 3952 146368
rect 4016 146304 4032 146368
rect 4096 146304 4112 146368
rect 4176 146304 4192 146368
rect 4256 146304 4264 146368
rect 3944 146303 4264 146304
rect 87944 146368 88264 146369
rect 87944 146304 87952 146368
rect 88016 146304 88032 146368
rect 88096 146304 88112 146368
rect 88176 146304 88192 146368
rect 88256 146304 88264 146368
rect 91200 146344 92000 146374
rect 87944 146303 88264 146304
rect 1944 145824 2264 145825
rect 1944 145760 1952 145824
rect 2016 145760 2032 145824
rect 2096 145760 2112 145824
rect 2176 145760 2192 145824
rect 2256 145760 2264 145824
rect 1944 145759 2264 145760
rect 85944 145824 86264 145825
rect 85944 145760 85952 145824
rect 86016 145760 86032 145824
rect 86096 145760 86112 145824
rect 86176 145760 86192 145824
rect 86256 145760 86264 145824
rect 85944 145759 86264 145760
rect 89944 145824 90264 145825
rect 89944 145760 89952 145824
rect 90016 145760 90032 145824
rect 90096 145760 90112 145824
rect 90176 145760 90192 145824
rect 90256 145760 90264 145824
rect 89944 145759 90264 145760
rect 3944 145280 4264 145281
rect 3944 145216 3952 145280
rect 4016 145216 4032 145280
rect 4096 145216 4112 145280
rect 4176 145216 4192 145280
rect 4256 145216 4264 145280
rect 3944 145215 4264 145216
rect 87944 145280 88264 145281
rect 87944 145216 87952 145280
rect 88016 145216 88032 145280
rect 88096 145216 88112 145280
rect 88176 145216 88192 145280
rect 88256 145216 88264 145280
rect 87944 145215 88264 145216
rect 91200 145210 92000 145240
rect 88382 145150 92000 145210
rect 87965 145074 88031 145077
rect 88382 145074 88442 145150
rect 91200 145120 92000 145150
rect 87965 145072 88442 145074
rect 87965 145016 87970 145072
rect 88026 145016 88442 145072
rect 87965 145014 88442 145016
rect 87965 145011 88031 145014
rect 1944 144736 2264 144737
rect 1944 144672 1952 144736
rect 2016 144672 2032 144736
rect 2096 144672 2112 144736
rect 2176 144672 2192 144736
rect 2256 144672 2264 144736
rect 1944 144671 2264 144672
rect 85944 144736 86264 144737
rect 85944 144672 85952 144736
rect 86016 144672 86032 144736
rect 86096 144672 86112 144736
rect 86176 144672 86192 144736
rect 86256 144672 86264 144736
rect 85944 144671 86264 144672
rect 89944 144736 90264 144737
rect 89944 144672 89952 144736
rect 90016 144672 90032 144736
rect 90096 144672 90112 144736
rect 90176 144672 90192 144736
rect 90256 144672 90264 144736
rect 89944 144671 90264 144672
rect 3944 144192 4264 144193
rect 3944 144128 3952 144192
rect 4016 144128 4032 144192
rect 4096 144128 4112 144192
rect 4176 144128 4192 144192
rect 4256 144128 4264 144192
rect 3944 144127 4264 144128
rect 87944 144192 88264 144193
rect 87944 144128 87952 144192
rect 88016 144128 88032 144192
rect 88096 144128 88112 144192
rect 88176 144128 88192 144192
rect 88256 144128 88264 144192
rect 87944 144127 88264 144128
rect 88057 143986 88123 143989
rect 91200 143986 92000 144016
rect 88057 143984 92000 143986
rect 88057 143928 88062 143984
rect 88118 143928 92000 143984
rect 88057 143926 92000 143928
rect 88057 143923 88123 143926
rect 91200 143896 92000 143926
rect 1944 143648 2264 143649
rect 1944 143584 1952 143648
rect 2016 143584 2032 143648
rect 2096 143584 2112 143648
rect 2176 143584 2192 143648
rect 2256 143584 2264 143648
rect 1944 143583 2264 143584
rect 85944 143648 86264 143649
rect 85944 143584 85952 143648
rect 86016 143584 86032 143648
rect 86096 143584 86112 143648
rect 86176 143584 86192 143648
rect 86256 143584 86264 143648
rect 85944 143583 86264 143584
rect 89944 143648 90264 143649
rect 89944 143584 89952 143648
rect 90016 143584 90032 143648
rect 90096 143584 90112 143648
rect 90176 143584 90192 143648
rect 90256 143584 90264 143648
rect 89944 143583 90264 143584
rect 3944 143104 4264 143105
rect 3944 143040 3952 143104
rect 4016 143040 4032 143104
rect 4096 143040 4112 143104
rect 4176 143040 4192 143104
rect 4256 143040 4264 143104
rect 3944 143039 4264 143040
rect 87944 143104 88264 143105
rect 87944 143040 87952 143104
rect 88016 143040 88032 143104
rect 88096 143040 88112 143104
rect 88176 143040 88192 143104
rect 88256 143040 88264 143104
rect 87944 143039 88264 143040
rect 87965 142762 88031 142765
rect 91200 142762 92000 142792
rect 87965 142760 92000 142762
rect 87965 142704 87970 142760
rect 88026 142704 92000 142760
rect 87965 142702 92000 142704
rect 87965 142699 88031 142702
rect 91200 142672 92000 142702
rect 1944 142560 2264 142561
rect 1944 142496 1952 142560
rect 2016 142496 2032 142560
rect 2096 142496 2112 142560
rect 2176 142496 2192 142560
rect 2256 142496 2264 142560
rect 1944 142495 2264 142496
rect 85944 142560 86264 142561
rect 85944 142496 85952 142560
rect 86016 142496 86032 142560
rect 86096 142496 86112 142560
rect 86176 142496 86192 142560
rect 86256 142496 86264 142560
rect 85944 142495 86264 142496
rect 89944 142560 90264 142561
rect 89944 142496 89952 142560
rect 90016 142496 90032 142560
rect 90096 142496 90112 142560
rect 90176 142496 90192 142560
rect 90256 142496 90264 142560
rect 89944 142495 90264 142496
rect 3944 142016 4264 142017
rect 3944 141952 3952 142016
rect 4016 141952 4032 142016
rect 4096 141952 4112 142016
rect 4176 141952 4192 142016
rect 4256 141952 4264 142016
rect 3944 141951 4264 141952
rect 87944 142016 88264 142017
rect 87944 141952 87952 142016
rect 88016 141952 88032 142016
rect 88096 141952 88112 142016
rect 88176 141952 88192 142016
rect 88256 141952 88264 142016
rect 87944 141951 88264 141952
rect 91200 141538 92000 141568
rect 90406 141478 92000 141538
rect 1944 141472 2264 141473
rect 1944 141408 1952 141472
rect 2016 141408 2032 141472
rect 2096 141408 2112 141472
rect 2176 141408 2192 141472
rect 2256 141408 2264 141472
rect 1944 141407 2264 141408
rect 85944 141472 86264 141473
rect 85944 141408 85952 141472
rect 86016 141408 86032 141472
rect 86096 141408 86112 141472
rect 86176 141408 86192 141472
rect 86256 141408 86264 141472
rect 85944 141407 86264 141408
rect 89944 141472 90264 141473
rect 89944 141408 89952 141472
rect 90016 141408 90032 141472
rect 90096 141408 90112 141472
rect 90176 141408 90192 141472
rect 90256 141408 90264 141472
rect 89944 141407 90264 141408
rect 87965 141266 88031 141269
rect 90406 141266 90466 141478
rect 91200 141448 92000 141478
rect 87965 141264 90466 141266
rect 87965 141208 87970 141264
rect 88026 141208 90466 141264
rect 87965 141206 90466 141208
rect 87965 141203 88031 141206
rect 3944 140928 4264 140929
rect 3944 140864 3952 140928
rect 4016 140864 4032 140928
rect 4096 140864 4112 140928
rect 4176 140864 4192 140928
rect 4256 140864 4264 140928
rect 3944 140863 4264 140864
rect 87944 140928 88264 140929
rect 87944 140864 87952 140928
rect 88016 140864 88032 140928
rect 88096 140864 88112 140928
rect 88176 140864 88192 140928
rect 88256 140864 88264 140928
rect 87944 140863 88264 140864
rect 1944 140384 2264 140385
rect 1944 140320 1952 140384
rect 2016 140320 2032 140384
rect 2096 140320 2112 140384
rect 2176 140320 2192 140384
rect 2256 140320 2264 140384
rect 1944 140319 2264 140320
rect 85944 140384 86264 140385
rect 85944 140320 85952 140384
rect 86016 140320 86032 140384
rect 86096 140320 86112 140384
rect 86176 140320 86192 140384
rect 86256 140320 86264 140384
rect 85944 140319 86264 140320
rect 89944 140384 90264 140385
rect 89944 140320 89952 140384
rect 90016 140320 90032 140384
rect 90096 140320 90112 140384
rect 90176 140320 90192 140384
rect 90256 140320 90264 140384
rect 89944 140319 90264 140320
rect 91200 140314 92000 140344
rect 90406 140254 92000 140314
rect 88241 140178 88307 140181
rect 90406 140178 90466 140254
rect 91200 140224 92000 140254
rect 88241 140176 90466 140178
rect 88241 140120 88246 140176
rect 88302 140120 90466 140176
rect 88241 140118 90466 140120
rect 88241 140115 88307 140118
rect 3944 139840 4264 139841
rect 3944 139776 3952 139840
rect 4016 139776 4032 139840
rect 4096 139776 4112 139840
rect 4176 139776 4192 139840
rect 4256 139776 4264 139840
rect 3944 139775 4264 139776
rect 87944 139840 88264 139841
rect 87944 139776 87952 139840
rect 88016 139776 88032 139840
rect 88096 139776 88112 139840
rect 88176 139776 88192 139840
rect 88256 139776 88264 139840
rect 87944 139775 88264 139776
rect 1944 139296 2264 139297
rect 1944 139232 1952 139296
rect 2016 139232 2032 139296
rect 2096 139232 2112 139296
rect 2176 139232 2192 139296
rect 2256 139232 2264 139296
rect 1944 139231 2264 139232
rect 85944 139296 86264 139297
rect 85944 139232 85952 139296
rect 86016 139232 86032 139296
rect 86096 139232 86112 139296
rect 86176 139232 86192 139296
rect 86256 139232 86264 139296
rect 85944 139231 86264 139232
rect 89944 139296 90264 139297
rect 89944 139232 89952 139296
rect 90016 139232 90032 139296
rect 90096 139232 90112 139296
rect 90176 139232 90192 139296
rect 90256 139232 90264 139296
rect 89944 139231 90264 139232
rect 88057 139090 88123 139093
rect 91200 139090 92000 139120
rect 88057 139088 92000 139090
rect 88057 139032 88062 139088
rect 88118 139032 92000 139088
rect 88057 139030 92000 139032
rect 88057 139027 88123 139030
rect 91200 139000 92000 139030
rect 3944 138752 4264 138753
rect 3944 138688 3952 138752
rect 4016 138688 4032 138752
rect 4096 138688 4112 138752
rect 4176 138688 4192 138752
rect 4256 138688 4264 138752
rect 3944 138687 4264 138688
rect 87944 138752 88264 138753
rect 87944 138688 87952 138752
rect 88016 138688 88032 138752
rect 88096 138688 88112 138752
rect 88176 138688 88192 138752
rect 88256 138688 88264 138752
rect 87944 138687 88264 138688
rect 1944 138208 2264 138209
rect 1944 138144 1952 138208
rect 2016 138144 2032 138208
rect 2096 138144 2112 138208
rect 2176 138144 2192 138208
rect 2256 138144 2264 138208
rect 1944 138143 2264 138144
rect 85944 138208 86264 138209
rect 85944 138144 85952 138208
rect 86016 138144 86032 138208
rect 86096 138144 86112 138208
rect 86176 138144 86192 138208
rect 86256 138144 86264 138208
rect 85944 138143 86264 138144
rect 89944 138208 90264 138209
rect 89944 138144 89952 138208
rect 90016 138144 90032 138208
rect 90096 138144 90112 138208
rect 90176 138144 90192 138208
rect 90256 138144 90264 138208
rect 89944 138143 90264 138144
rect 86493 137866 86559 137869
rect 91200 137866 92000 137896
rect 86493 137864 92000 137866
rect 86493 137808 86498 137864
rect 86554 137808 92000 137864
rect 86493 137806 92000 137808
rect 86493 137803 86559 137806
rect 91200 137776 92000 137806
rect 3944 137664 4264 137665
rect 3944 137600 3952 137664
rect 4016 137600 4032 137664
rect 4096 137600 4112 137664
rect 4176 137600 4192 137664
rect 4256 137600 4264 137664
rect 3944 137599 4264 137600
rect 87944 137664 88264 137665
rect 87944 137600 87952 137664
rect 88016 137600 88032 137664
rect 88096 137600 88112 137664
rect 88176 137600 88192 137664
rect 88256 137600 88264 137664
rect 87944 137599 88264 137600
rect 1944 137120 2264 137121
rect 1944 137056 1952 137120
rect 2016 137056 2032 137120
rect 2096 137056 2112 137120
rect 2176 137056 2192 137120
rect 2256 137056 2264 137120
rect 1944 137055 2264 137056
rect 85944 137120 86264 137121
rect 85944 137056 85952 137120
rect 86016 137056 86032 137120
rect 86096 137056 86112 137120
rect 86176 137056 86192 137120
rect 86256 137056 86264 137120
rect 85944 137055 86264 137056
rect 89944 137120 90264 137121
rect 89944 137056 89952 137120
rect 90016 137056 90032 137120
rect 90096 137056 90112 137120
rect 90176 137056 90192 137120
rect 90256 137056 90264 137120
rect 89944 137055 90264 137056
rect 91200 136642 92000 136672
rect 88382 136582 92000 136642
rect 3944 136576 4264 136577
rect 3944 136512 3952 136576
rect 4016 136512 4032 136576
rect 4096 136512 4112 136576
rect 4176 136512 4192 136576
rect 4256 136512 4264 136576
rect 3944 136511 4264 136512
rect 87944 136576 88264 136577
rect 87944 136512 87952 136576
rect 88016 136512 88032 136576
rect 88096 136512 88112 136576
rect 88176 136512 88192 136576
rect 88256 136512 88264 136576
rect 87944 136511 88264 136512
rect 86309 136370 86375 136373
rect 88382 136370 88442 136582
rect 91200 136552 92000 136582
rect 86309 136368 88442 136370
rect 86309 136312 86314 136368
rect 86370 136312 88442 136368
rect 86309 136310 88442 136312
rect 86309 136307 86375 136310
rect 1944 136032 2264 136033
rect 1944 135968 1952 136032
rect 2016 135968 2032 136032
rect 2096 135968 2112 136032
rect 2176 135968 2192 136032
rect 2256 135968 2264 136032
rect 1944 135967 2264 135968
rect 85944 136032 86264 136033
rect 85944 135968 85952 136032
rect 86016 135968 86032 136032
rect 86096 135968 86112 136032
rect 86176 135968 86192 136032
rect 86256 135968 86264 136032
rect 85944 135967 86264 135968
rect 89944 136032 90264 136033
rect 89944 135968 89952 136032
rect 90016 135968 90032 136032
rect 90096 135968 90112 136032
rect 90176 135968 90192 136032
rect 90256 135968 90264 136032
rect 89944 135967 90264 135968
rect 3944 135488 4264 135489
rect 3944 135424 3952 135488
rect 4016 135424 4032 135488
rect 4096 135424 4112 135488
rect 4176 135424 4192 135488
rect 4256 135424 4264 135488
rect 3944 135423 4264 135424
rect 87944 135488 88264 135489
rect 87944 135424 87952 135488
rect 88016 135424 88032 135488
rect 88096 135424 88112 135488
rect 88176 135424 88192 135488
rect 88256 135424 88264 135488
rect 87944 135423 88264 135424
rect 91200 135418 92000 135448
rect 88382 135358 92000 135418
rect 86401 135282 86467 135285
rect 88382 135282 88442 135358
rect 91200 135328 92000 135358
rect 86401 135280 88442 135282
rect 86401 135224 86406 135280
rect 86462 135224 88442 135280
rect 86401 135222 88442 135224
rect 86401 135219 86467 135222
rect 1944 134944 2264 134945
rect 1944 134880 1952 134944
rect 2016 134880 2032 134944
rect 2096 134880 2112 134944
rect 2176 134880 2192 134944
rect 2256 134880 2264 134944
rect 1944 134879 2264 134880
rect 85944 134944 86264 134945
rect 85944 134880 85952 134944
rect 86016 134880 86032 134944
rect 86096 134880 86112 134944
rect 86176 134880 86192 134944
rect 86256 134880 86264 134944
rect 85944 134879 86264 134880
rect 89944 134944 90264 134945
rect 89944 134880 89952 134944
rect 90016 134880 90032 134944
rect 90096 134880 90112 134944
rect 90176 134880 90192 134944
rect 90256 134880 90264 134944
rect 89944 134879 90264 134880
rect 3944 134400 4264 134401
rect 3944 134336 3952 134400
rect 4016 134336 4032 134400
rect 4096 134336 4112 134400
rect 4176 134336 4192 134400
rect 4256 134336 4264 134400
rect 3944 134335 4264 134336
rect 87944 134400 88264 134401
rect 87944 134336 87952 134400
rect 88016 134336 88032 134400
rect 88096 134336 88112 134400
rect 88176 134336 88192 134400
rect 88256 134336 88264 134400
rect 87944 134335 88264 134336
rect 91200 134330 92000 134360
rect 88382 134270 92000 134330
rect 86861 134194 86927 134197
rect 88382 134194 88442 134270
rect 91200 134240 92000 134270
rect 86861 134192 88442 134194
rect 86861 134136 86866 134192
rect 86922 134136 88442 134192
rect 86861 134134 88442 134136
rect 86861 134131 86927 134134
rect 1944 133856 2264 133857
rect 1944 133792 1952 133856
rect 2016 133792 2032 133856
rect 2096 133792 2112 133856
rect 2176 133792 2192 133856
rect 2256 133792 2264 133856
rect 1944 133791 2264 133792
rect 85944 133856 86264 133857
rect 85944 133792 85952 133856
rect 86016 133792 86032 133856
rect 86096 133792 86112 133856
rect 86176 133792 86192 133856
rect 86256 133792 86264 133856
rect 85944 133791 86264 133792
rect 89944 133856 90264 133857
rect 89944 133792 89952 133856
rect 90016 133792 90032 133856
rect 90096 133792 90112 133856
rect 90176 133792 90192 133856
rect 90256 133792 90264 133856
rect 89944 133791 90264 133792
rect 3944 133312 4264 133313
rect 3944 133248 3952 133312
rect 4016 133248 4032 133312
rect 4096 133248 4112 133312
rect 4176 133248 4192 133312
rect 4256 133248 4264 133312
rect 3944 133247 4264 133248
rect 87944 133312 88264 133313
rect 87944 133248 87952 133312
rect 88016 133248 88032 133312
rect 88096 133248 88112 133312
rect 88176 133248 88192 133312
rect 88256 133248 88264 133312
rect 87944 133247 88264 133248
rect 84878 133044 84884 133108
rect 84948 133106 84954 133108
rect 91200 133106 92000 133136
rect 84948 133046 92000 133106
rect 84948 133044 84954 133046
rect 91200 133016 92000 133046
rect 1944 132768 2264 132769
rect 1944 132704 1952 132768
rect 2016 132704 2032 132768
rect 2096 132704 2112 132768
rect 2176 132704 2192 132768
rect 2256 132704 2264 132768
rect 1944 132703 2264 132704
rect 85944 132768 86264 132769
rect 85944 132704 85952 132768
rect 86016 132704 86032 132768
rect 86096 132704 86112 132768
rect 86176 132704 86192 132768
rect 86256 132704 86264 132768
rect 85944 132703 86264 132704
rect 89944 132768 90264 132769
rect 89944 132704 89952 132768
rect 90016 132704 90032 132768
rect 90096 132704 90112 132768
rect 90176 132704 90192 132768
rect 90256 132704 90264 132768
rect 89944 132703 90264 132704
rect 83406 132364 83412 132428
rect 83476 132426 83482 132428
rect 83958 132426 83964 132428
rect 83476 132366 83964 132426
rect 83476 132364 83482 132366
rect 83958 132364 83964 132366
rect 84028 132364 84034 132428
rect 82537 132290 82603 132293
rect 83406 132290 83412 132292
rect 82537 132288 83412 132290
rect 82537 132232 82542 132288
rect 82598 132232 83412 132288
rect 82537 132230 83412 132232
rect 82537 132227 82603 132230
rect 83406 132228 83412 132230
rect 83476 132228 83482 132292
rect 3944 132224 4264 132225
rect 3944 132160 3952 132224
rect 4016 132160 4032 132224
rect 4096 132160 4112 132224
rect 4176 132160 4192 132224
rect 4256 132160 4264 132224
rect 3944 132159 4264 132160
rect 87944 132224 88264 132225
rect 87944 132160 87952 132224
rect 88016 132160 88032 132224
rect 88096 132160 88112 132224
rect 88176 132160 88192 132224
rect 88256 132160 88264 132224
rect 87944 132159 88264 132160
rect 88241 131882 88307 131885
rect 91200 131882 92000 131912
rect 88241 131880 92000 131882
rect 88241 131824 88246 131880
rect 88302 131824 92000 131880
rect 88241 131822 92000 131824
rect 88241 131819 88307 131822
rect 91200 131792 92000 131822
rect 1944 131680 2264 131681
rect 1944 131616 1952 131680
rect 2016 131616 2032 131680
rect 2096 131616 2112 131680
rect 2176 131616 2192 131680
rect 2256 131616 2264 131680
rect 1944 131615 2264 131616
rect 85944 131680 86264 131681
rect 85944 131616 85952 131680
rect 86016 131616 86032 131680
rect 86096 131616 86112 131680
rect 86176 131616 86192 131680
rect 86256 131616 86264 131680
rect 85944 131615 86264 131616
rect 89944 131680 90264 131681
rect 89944 131616 89952 131680
rect 90016 131616 90032 131680
rect 90096 131616 90112 131680
rect 90176 131616 90192 131680
rect 90256 131616 90264 131680
rect 89944 131615 90264 131616
rect 3944 131136 4264 131137
rect 3944 131072 3952 131136
rect 4016 131072 4032 131136
rect 4096 131072 4112 131136
rect 4176 131072 4192 131136
rect 4256 131072 4264 131136
rect 3944 131071 4264 131072
rect 87944 131136 88264 131137
rect 87944 131072 87952 131136
rect 88016 131072 88032 131136
rect 88096 131072 88112 131136
rect 88176 131072 88192 131136
rect 88256 131072 88264 131136
rect 87944 131071 88264 131072
rect 91200 130658 92000 130688
rect 90406 130598 92000 130658
rect 1944 130592 2264 130593
rect 1944 130528 1952 130592
rect 2016 130528 2032 130592
rect 2096 130528 2112 130592
rect 2176 130528 2192 130592
rect 2256 130528 2264 130592
rect 1944 130527 2264 130528
rect 85944 130592 86264 130593
rect 85944 130528 85952 130592
rect 86016 130528 86032 130592
rect 86096 130528 86112 130592
rect 86176 130528 86192 130592
rect 86256 130528 86264 130592
rect 85944 130527 86264 130528
rect 89944 130592 90264 130593
rect 89944 130528 89952 130592
rect 90016 130528 90032 130592
rect 90096 130528 90112 130592
rect 90176 130528 90192 130592
rect 90256 130528 90264 130592
rect 89944 130527 90264 130528
rect 85246 130324 85252 130388
rect 85316 130386 85322 130388
rect 90406 130386 90466 130598
rect 91200 130568 92000 130598
rect 85316 130326 90466 130386
rect 85316 130324 85322 130326
rect 3944 130048 4264 130049
rect 3944 129984 3952 130048
rect 4016 129984 4032 130048
rect 4096 129984 4112 130048
rect 4176 129984 4192 130048
rect 4256 129984 4264 130048
rect 3944 129983 4264 129984
rect 87944 130048 88264 130049
rect 87944 129984 87952 130048
rect 88016 129984 88032 130048
rect 88096 129984 88112 130048
rect 88176 129984 88192 130048
rect 88256 129984 88264 130048
rect 87944 129983 88264 129984
rect 1944 129504 2264 129505
rect 1944 129440 1952 129504
rect 2016 129440 2032 129504
rect 2096 129440 2112 129504
rect 2176 129440 2192 129504
rect 2256 129440 2264 129504
rect 1944 129439 2264 129440
rect 85944 129504 86264 129505
rect 85944 129440 85952 129504
rect 86016 129440 86032 129504
rect 86096 129440 86112 129504
rect 86176 129440 86192 129504
rect 86256 129440 86264 129504
rect 85944 129439 86264 129440
rect 89944 129504 90264 129505
rect 89944 129440 89952 129504
rect 90016 129440 90032 129504
rect 90096 129440 90112 129504
rect 90176 129440 90192 129504
rect 90256 129440 90264 129504
rect 89944 129439 90264 129440
rect 91200 129434 92000 129464
rect 90406 129374 92000 129434
rect 88241 129298 88307 129301
rect 90406 129298 90466 129374
rect 91200 129344 92000 129374
rect 88241 129296 90466 129298
rect 88241 129240 88246 129296
rect 88302 129240 90466 129296
rect 88241 129238 90466 129240
rect 88241 129235 88307 129238
rect 3944 128960 4264 128961
rect 3944 128896 3952 128960
rect 4016 128896 4032 128960
rect 4096 128896 4112 128960
rect 4176 128896 4192 128960
rect 4256 128896 4264 128960
rect 3944 128895 4264 128896
rect 87944 128960 88264 128961
rect 87944 128896 87952 128960
rect 88016 128896 88032 128960
rect 88096 128896 88112 128960
rect 88176 128896 88192 128960
rect 88256 128896 88264 128960
rect 87944 128895 88264 128896
rect 1944 128416 2264 128417
rect 1944 128352 1952 128416
rect 2016 128352 2032 128416
rect 2096 128352 2112 128416
rect 2176 128352 2192 128416
rect 2256 128352 2264 128416
rect 1944 128351 2264 128352
rect 85944 128416 86264 128417
rect 85944 128352 85952 128416
rect 86016 128352 86032 128416
rect 86096 128352 86112 128416
rect 86176 128352 86192 128416
rect 86256 128352 86264 128416
rect 85944 128351 86264 128352
rect 89944 128416 90264 128417
rect 89944 128352 89952 128416
rect 90016 128352 90032 128416
rect 90096 128352 90112 128416
rect 90176 128352 90192 128416
rect 90256 128352 90264 128416
rect 89944 128351 90264 128352
rect 88241 128210 88307 128213
rect 91200 128210 92000 128240
rect 88241 128208 92000 128210
rect 88241 128152 88246 128208
rect 88302 128152 92000 128208
rect 88241 128150 92000 128152
rect 88241 128147 88307 128150
rect 91200 128120 92000 128150
rect 3944 127872 4264 127873
rect 3944 127808 3952 127872
rect 4016 127808 4032 127872
rect 4096 127808 4112 127872
rect 4176 127808 4192 127872
rect 4256 127808 4264 127872
rect 3944 127807 4264 127808
rect 87944 127872 88264 127873
rect 87944 127808 87952 127872
rect 88016 127808 88032 127872
rect 88096 127808 88112 127872
rect 88176 127808 88192 127872
rect 88256 127808 88264 127872
rect 87944 127807 88264 127808
rect 1944 127328 2264 127329
rect 1944 127264 1952 127328
rect 2016 127264 2032 127328
rect 2096 127264 2112 127328
rect 2176 127264 2192 127328
rect 2256 127264 2264 127328
rect 1944 127263 2264 127264
rect 85944 127328 86264 127329
rect 85944 127264 85952 127328
rect 86016 127264 86032 127328
rect 86096 127264 86112 127328
rect 86176 127264 86192 127328
rect 86256 127264 86264 127328
rect 85944 127263 86264 127264
rect 89944 127328 90264 127329
rect 89944 127264 89952 127328
rect 90016 127264 90032 127328
rect 90096 127264 90112 127328
rect 90176 127264 90192 127328
rect 90256 127264 90264 127328
rect 89944 127263 90264 127264
rect 84510 126924 84516 126988
rect 84580 126986 84586 126988
rect 91200 126986 92000 127016
rect 84580 126926 92000 126986
rect 84580 126924 84586 126926
rect 91200 126896 92000 126926
rect 3944 126784 4264 126785
rect 3944 126720 3952 126784
rect 4016 126720 4032 126784
rect 4096 126720 4112 126784
rect 4176 126720 4192 126784
rect 4256 126720 4264 126784
rect 3944 126719 4264 126720
rect 87944 126784 88264 126785
rect 87944 126720 87952 126784
rect 88016 126720 88032 126784
rect 88096 126720 88112 126784
rect 88176 126720 88192 126784
rect 88256 126720 88264 126784
rect 87944 126719 88264 126720
rect 1944 126240 2264 126241
rect 1944 126176 1952 126240
rect 2016 126176 2032 126240
rect 2096 126176 2112 126240
rect 2176 126176 2192 126240
rect 2256 126176 2264 126240
rect 1944 126175 2264 126176
rect 85944 126240 86264 126241
rect 85944 126176 85952 126240
rect 86016 126176 86032 126240
rect 86096 126176 86112 126240
rect 86176 126176 86192 126240
rect 86256 126176 86264 126240
rect 85944 126175 86264 126176
rect 89944 126240 90264 126241
rect 89944 126176 89952 126240
rect 90016 126176 90032 126240
rect 90096 126176 90112 126240
rect 90176 126176 90192 126240
rect 90256 126176 90264 126240
rect 89944 126175 90264 126176
rect 87965 125898 88031 125901
rect 87965 125896 88442 125898
rect 83260 125790 83474 125850
rect 87965 125840 87970 125896
rect 88026 125840 88442 125896
rect 87965 125838 88442 125840
rect 87965 125835 88031 125838
rect 83414 125762 83474 125790
rect 84561 125762 84627 125765
rect 84694 125762 84700 125764
rect 83414 125760 84700 125762
rect 83414 125704 84566 125760
rect 84622 125704 84700 125760
rect 83414 125702 84700 125704
rect 84561 125699 84627 125702
rect 84694 125700 84700 125702
rect 84764 125700 84770 125764
rect 88382 125762 88442 125838
rect 91200 125762 92000 125792
rect 88382 125702 92000 125762
rect 3944 125696 4264 125697
rect 3944 125632 3952 125696
rect 4016 125632 4032 125696
rect 4096 125632 4112 125696
rect 4176 125632 4192 125696
rect 4256 125632 4264 125696
rect 3944 125631 4264 125632
rect 87944 125696 88264 125697
rect 87944 125632 87952 125696
rect 88016 125632 88032 125696
rect 88096 125632 88112 125696
rect 88176 125632 88192 125696
rect 88256 125632 88264 125696
rect 91200 125672 92000 125702
rect 87944 125631 88264 125632
rect 1944 125152 2264 125153
rect 1944 125088 1952 125152
rect 2016 125088 2032 125152
rect 2096 125088 2112 125152
rect 2176 125088 2192 125152
rect 2256 125088 2264 125152
rect 1944 125087 2264 125088
rect 85944 125152 86264 125153
rect 85944 125088 85952 125152
rect 86016 125088 86032 125152
rect 86096 125088 86112 125152
rect 86176 125088 86192 125152
rect 86256 125088 86264 125152
rect 85944 125087 86264 125088
rect 89944 125152 90264 125153
rect 89944 125088 89952 125152
rect 90016 125088 90032 125152
rect 90096 125088 90112 125152
rect 90176 125088 90192 125152
rect 90256 125088 90264 125152
rect 89944 125087 90264 125088
rect 3944 124608 4264 124609
rect 3944 124544 3952 124608
rect 4016 124544 4032 124608
rect 4096 124544 4112 124608
rect 4176 124544 4192 124608
rect 4256 124544 4264 124608
rect 3944 124543 4264 124544
rect 87944 124608 88264 124609
rect 87944 124544 87952 124608
rect 88016 124544 88032 124608
rect 88096 124544 88112 124608
rect 88176 124544 88192 124608
rect 88256 124544 88264 124608
rect 87944 124543 88264 124544
rect 91200 124538 92000 124568
rect 88382 124478 92000 124538
rect 88241 124402 88307 124405
rect 88382 124402 88442 124478
rect 91200 124448 92000 124478
rect 88241 124400 88442 124402
rect 88241 124344 88246 124400
rect 88302 124344 88442 124400
rect 88241 124342 88442 124344
rect 88241 124339 88307 124342
rect 84469 124130 84535 124133
rect 83230 124128 84535 124130
rect 83230 124072 84474 124128
rect 84530 124072 84535 124128
rect 83230 124070 84535 124072
rect 84469 124067 84535 124070
rect 1944 124064 2264 124065
rect 1944 124000 1952 124064
rect 2016 124000 2032 124064
rect 2096 124000 2112 124064
rect 2176 124000 2192 124064
rect 2256 124000 2264 124064
rect 1944 123999 2264 124000
rect 85944 124064 86264 124065
rect 85944 124000 85952 124064
rect 86016 124000 86032 124064
rect 86096 124000 86112 124064
rect 86176 124000 86192 124064
rect 86256 124000 86264 124064
rect 85944 123999 86264 124000
rect 89944 124064 90264 124065
rect 89944 124000 89952 124064
rect 90016 124000 90032 124064
rect 90096 124000 90112 124064
rect 90176 124000 90192 124064
rect 90256 124000 90264 124064
rect 89944 123999 90264 124000
rect 3944 123520 4264 123521
rect 3944 123456 3952 123520
rect 4016 123456 4032 123520
rect 4096 123456 4112 123520
rect 4176 123456 4192 123520
rect 4256 123456 4264 123520
rect 3944 123455 4264 123456
rect 87944 123520 88264 123521
rect 87944 123456 87952 123520
rect 88016 123456 88032 123520
rect 88096 123456 88112 123520
rect 88176 123456 88192 123520
rect 88256 123456 88264 123520
rect 87944 123455 88264 123456
rect 87965 123314 88031 123317
rect 91200 123314 92000 123344
rect 87965 123312 92000 123314
rect 87965 123256 87970 123312
rect 88026 123256 92000 123312
rect 87965 123254 92000 123256
rect 87965 123251 88031 123254
rect 91200 123224 92000 123254
rect 84377 123042 84443 123045
rect 83230 123040 84443 123042
rect 83230 122984 84382 123040
rect 84438 122984 84443 123040
rect 83230 122982 84443 122984
rect 84377 122979 84443 122982
rect 1944 122976 2264 122977
rect 1944 122912 1952 122976
rect 2016 122912 2032 122976
rect 2096 122912 2112 122976
rect 2176 122912 2192 122976
rect 2256 122912 2264 122976
rect 1944 122911 2264 122912
rect 85944 122976 86264 122977
rect 85944 122912 85952 122976
rect 86016 122912 86032 122976
rect 86096 122912 86112 122976
rect 86176 122912 86192 122976
rect 86256 122912 86264 122976
rect 85944 122911 86264 122912
rect 89944 122976 90264 122977
rect 89944 122912 89952 122976
rect 90016 122912 90032 122976
rect 90096 122912 90112 122976
rect 90176 122912 90192 122976
rect 90256 122912 90264 122976
rect 89944 122911 90264 122912
rect 86902 122572 86908 122636
rect 86972 122634 86978 122636
rect 90582 122634 90588 122636
rect 86972 122574 90588 122634
rect 86972 122572 86978 122574
rect 90582 122572 90588 122574
rect 90652 122572 90658 122636
rect 3944 122432 4264 122433
rect 3944 122368 3952 122432
rect 4016 122368 4032 122432
rect 4096 122368 4112 122432
rect 4176 122368 4192 122432
rect 4256 122368 4264 122432
rect 3944 122367 4264 122368
rect 87944 122432 88264 122433
rect 87944 122368 87952 122432
rect 88016 122368 88032 122432
rect 88096 122368 88112 122432
rect 88176 122368 88192 122432
rect 88256 122368 88264 122432
rect 87944 122367 88264 122368
rect 86902 122300 86908 122364
rect 86972 122362 86978 122364
rect 87229 122362 87295 122365
rect 86972 122360 87295 122362
rect 86972 122304 87234 122360
rect 87290 122304 87295 122360
rect 86972 122302 87295 122304
rect 86972 122300 86978 122302
rect 87229 122299 87295 122302
rect 87873 122090 87939 122093
rect 91200 122090 92000 122120
rect 87873 122088 92000 122090
rect 87873 122032 87878 122088
rect 87934 122032 92000 122088
rect 87873 122030 92000 122032
rect 87873 122027 87939 122030
rect 91200 122000 92000 122030
rect 1944 121888 2264 121889
rect 1944 121824 1952 121888
rect 2016 121824 2032 121888
rect 2096 121824 2112 121888
rect 2176 121824 2192 121888
rect 2256 121824 2264 121888
rect 1944 121823 2264 121824
rect 85944 121888 86264 121889
rect 85944 121824 85952 121888
rect 86016 121824 86032 121888
rect 86096 121824 86112 121888
rect 86176 121824 86192 121888
rect 86256 121824 86264 121888
rect 85944 121823 86264 121824
rect 89944 121888 90264 121889
rect 89944 121824 89952 121888
rect 90016 121824 90032 121888
rect 90096 121824 90112 121888
rect 90176 121824 90192 121888
rect 90256 121824 90264 121888
rect 89944 121823 90264 121824
rect 5441 121546 5507 121549
rect 6126 121546 6132 121548
rect 5441 121544 6132 121546
rect 5441 121488 5446 121544
rect 5502 121488 6132 121544
rect 5441 121486 6132 121488
rect 5441 121483 5507 121486
rect 6126 121484 6132 121486
rect 6196 121484 6202 121548
rect 3944 121344 4264 121345
rect 3944 121280 3952 121344
rect 4016 121280 4032 121344
rect 4096 121280 4112 121344
rect 4176 121280 4192 121344
rect 4256 121280 4264 121344
rect 87944 121344 88264 121345
rect 3944 121279 4264 121280
rect 83230 121002 83290 121292
rect 87944 121280 87952 121344
rect 88016 121280 88032 121344
rect 88096 121280 88112 121344
rect 88176 121280 88192 121344
rect 88256 121280 88264 121344
rect 87944 121279 88264 121280
rect 84469 121002 84535 121005
rect 83230 121000 84535 121002
rect 83230 120944 84474 121000
rect 84530 120944 84535 121000
rect 83230 120942 84535 120944
rect 84469 120939 84535 120942
rect 91200 120866 92000 120896
rect 90406 120806 92000 120866
rect 1944 120800 2264 120801
rect 1944 120736 1952 120800
rect 2016 120736 2032 120800
rect 2096 120736 2112 120800
rect 2176 120736 2192 120800
rect 2256 120736 2264 120800
rect 1944 120735 2264 120736
rect 85944 120800 86264 120801
rect 85944 120736 85952 120800
rect 86016 120736 86032 120800
rect 86096 120736 86112 120800
rect 86176 120736 86192 120800
rect 86256 120736 86264 120800
rect 85944 120735 86264 120736
rect 89944 120800 90264 120801
rect 89944 120736 89952 120800
rect 90016 120736 90032 120800
rect 90096 120736 90112 120800
rect 90176 120736 90192 120800
rect 90256 120736 90264 120800
rect 89944 120735 90264 120736
rect 87873 120594 87939 120597
rect 90406 120594 90466 120806
rect 91200 120776 92000 120806
rect 87873 120592 90466 120594
rect 87873 120536 87878 120592
rect 87934 120536 90466 120592
rect 87873 120534 90466 120536
rect 87873 120531 87939 120534
rect 3944 120256 4264 120257
rect 3944 120192 3952 120256
rect 4016 120192 4032 120256
rect 4096 120192 4112 120256
rect 4176 120192 4192 120256
rect 4256 120192 4264 120256
rect 3944 120191 4264 120192
rect 87944 120256 88264 120257
rect 87944 120192 87952 120256
rect 88016 120192 88032 120256
rect 88096 120192 88112 120256
rect 88176 120192 88192 120256
rect 88256 120192 88264 120256
rect 87944 120191 88264 120192
rect 84326 120186 84332 120188
rect 83230 120126 84332 120186
rect 84326 120124 84332 120126
rect 84396 120186 84402 120188
rect 84561 120186 84627 120189
rect 84396 120184 84627 120186
rect 84396 120128 84566 120184
rect 84622 120128 84627 120184
rect 84396 120126 84627 120128
rect 84396 120124 84402 120126
rect 84561 120123 84627 120126
rect 1944 119712 2264 119713
rect 1944 119648 1952 119712
rect 2016 119648 2032 119712
rect 2096 119648 2112 119712
rect 2176 119648 2192 119712
rect 2256 119648 2264 119712
rect 1944 119647 2264 119648
rect 85944 119712 86264 119713
rect 85944 119648 85952 119712
rect 86016 119648 86032 119712
rect 86096 119648 86112 119712
rect 86176 119648 86192 119712
rect 86256 119648 86264 119712
rect 85944 119647 86264 119648
rect 89944 119712 90264 119713
rect 89944 119648 89952 119712
rect 90016 119648 90032 119712
rect 90096 119648 90112 119712
rect 90176 119648 90192 119712
rect 90256 119648 90264 119712
rect 89944 119647 90264 119648
rect 91200 119642 92000 119672
rect 90406 119582 92000 119642
rect 87873 119506 87939 119509
rect 90406 119506 90466 119582
rect 91200 119552 92000 119582
rect 87873 119504 90466 119506
rect 87873 119448 87878 119504
rect 87934 119448 90466 119504
rect 87873 119446 90466 119448
rect 87873 119443 87939 119446
rect 3944 119168 4264 119169
rect 3944 119104 3952 119168
rect 4016 119104 4032 119168
rect 4096 119104 4112 119168
rect 4176 119104 4192 119168
rect 4256 119104 4264 119168
rect 3944 119103 4264 119104
rect 87944 119168 88264 119169
rect 87944 119104 87952 119168
rect 88016 119104 88032 119168
rect 88096 119104 88112 119168
rect 88176 119104 88192 119168
rect 88256 119104 88264 119168
rect 87944 119103 88264 119104
rect 87229 118690 87295 118693
rect 86358 118688 87295 118690
rect 86358 118632 87234 118688
rect 87290 118632 87295 118688
rect 86358 118630 87295 118632
rect 1944 118624 2264 118625
rect 1944 118560 1952 118624
rect 2016 118560 2032 118624
rect 2096 118560 2112 118624
rect 2176 118560 2192 118624
rect 2256 118560 2264 118624
rect 1944 118559 2264 118560
rect 85944 118624 86264 118625
rect 85944 118560 85952 118624
rect 86016 118560 86032 118624
rect 86096 118560 86112 118624
rect 86176 118560 86192 118624
rect 86256 118560 86264 118624
rect 85944 118559 86264 118560
rect 83230 118282 83290 118464
rect 85481 118418 85547 118421
rect 86358 118418 86418 118630
rect 87229 118627 87295 118630
rect 89944 118624 90264 118625
rect 89944 118560 89952 118624
rect 90016 118560 90032 118624
rect 90096 118560 90112 118624
rect 90176 118560 90192 118624
rect 90256 118560 90264 118624
rect 89944 118559 90264 118560
rect 86902 118492 86908 118556
rect 86972 118554 86978 118556
rect 87229 118554 87295 118557
rect 86972 118552 87295 118554
rect 86972 118496 87234 118552
rect 87290 118496 87295 118552
rect 86972 118494 87295 118496
rect 86972 118492 86978 118494
rect 87229 118491 87295 118494
rect 85481 118416 86418 118418
rect 85481 118360 85486 118416
rect 85542 118360 86418 118416
rect 85481 118358 86418 118360
rect 88977 118418 89043 118421
rect 91200 118418 92000 118448
rect 88977 118416 92000 118418
rect 88977 118360 88982 118416
rect 89038 118360 92000 118416
rect 88977 118358 92000 118360
rect 85481 118355 85547 118358
rect 88977 118355 89043 118358
rect 91200 118328 92000 118358
rect 84377 118282 84443 118285
rect 83230 118280 84443 118282
rect 83230 118224 84382 118280
rect 84438 118224 84443 118280
rect 83230 118222 84443 118224
rect 84377 118219 84443 118222
rect 3944 118080 4264 118081
rect 3944 118016 3952 118080
rect 4016 118016 4032 118080
rect 4096 118016 4112 118080
rect 4176 118016 4192 118080
rect 4256 118016 4264 118080
rect 3944 118015 4264 118016
rect 87944 118080 88264 118081
rect 87944 118016 87952 118080
rect 88016 118016 88032 118080
rect 88096 118016 88112 118080
rect 88176 118016 88192 118080
rect 88256 118016 88264 118080
rect 87944 118015 88264 118016
rect 1944 117536 2264 117537
rect 1944 117472 1952 117536
rect 2016 117472 2032 117536
rect 2096 117472 2112 117536
rect 2176 117472 2192 117536
rect 2256 117472 2264 117536
rect 1944 117471 2264 117472
rect 85944 117536 86264 117537
rect 85944 117472 85952 117536
rect 86016 117472 86032 117536
rect 86096 117472 86112 117536
rect 86176 117472 86192 117536
rect 86256 117472 86264 117536
rect 85944 117471 86264 117472
rect 89944 117536 90264 117537
rect 89944 117472 89952 117536
rect 90016 117472 90032 117536
rect 90096 117472 90112 117536
rect 90176 117472 90192 117536
rect 90256 117472 90264 117536
rect 89944 117471 90264 117472
rect 83230 117330 83290 117336
rect 84561 117330 84627 117333
rect 83230 117328 84627 117330
rect 83230 117272 84566 117328
rect 84622 117272 84627 117328
rect 83230 117270 84627 117272
rect 84561 117267 84627 117270
rect 91200 117194 92000 117224
rect 89670 117134 92000 117194
rect 3944 116992 4264 116993
rect 3944 116928 3952 116992
rect 4016 116928 4032 116992
rect 4096 116928 4112 116992
rect 4176 116928 4192 116992
rect 4256 116928 4264 116992
rect 3944 116927 4264 116928
rect 87944 116992 88264 116993
rect 87944 116928 87952 116992
rect 88016 116928 88032 116992
rect 88096 116928 88112 116992
rect 88176 116928 88192 116992
rect 88256 116928 88264 116992
rect 87944 116927 88264 116928
rect 88241 116786 88307 116789
rect 89670 116786 89730 117134
rect 91200 117104 92000 117134
rect 88241 116784 89730 116786
rect 88241 116728 88246 116784
rect 88302 116728 89730 116784
rect 88241 116726 89730 116728
rect 88241 116723 88307 116726
rect 5349 116652 5415 116653
rect 5349 116650 5396 116652
rect 5268 116648 5396 116650
rect 5460 116650 5466 116652
rect 6134 116650 6194 116663
rect 5268 116592 5354 116648
rect 5268 116590 5396 116592
rect 5349 116588 5396 116590
rect 5460 116590 6194 116650
rect 5460 116588 5466 116590
rect 5349 116587 5415 116588
rect 1944 116448 2264 116449
rect 1944 116384 1952 116448
rect 2016 116384 2032 116448
rect 2096 116384 2112 116448
rect 2176 116384 2192 116448
rect 2256 116384 2264 116448
rect 1944 116383 2264 116384
rect 85944 116448 86264 116449
rect 85944 116384 85952 116448
rect 86016 116384 86032 116448
rect 86096 116384 86112 116448
rect 86176 116384 86192 116448
rect 86256 116384 86264 116448
rect 85944 116383 86264 116384
rect 89944 116448 90264 116449
rect 89944 116384 89952 116448
rect 90016 116384 90032 116448
rect 90096 116384 90112 116448
rect 90176 116384 90192 116448
rect 90256 116384 90264 116448
rect 89944 116383 90264 116384
rect 86309 116106 86375 116109
rect 86309 116104 89730 116106
rect 86309 116048 86314 116104
rect 86370 116048 89730 116104
rect 86309 116046 89730 116048
rect 86309 116043 86375 116046
rect 89670 115970 89730 116046
rect 91200 115970 92000 116000
rect 89670 115910 92000 115970
rect 3944 115904 4264 115905
rect 3944 115840 3952 115904
rect 4016 115840 4032 115904
rect 4096 115840 4112 115904
rect 4176 115840 4192 115904
rect 4256 115840 4264 115904
rect 3944 115839 4264 115840
rect 87944 115904 88264 115905
rect 87944 115840 87952 115904
rect 88016 115840 88032 115904
rect 88096 115840 88112 115904
rect 88176 115840 88192 115904
rect 88256 115840 88264 115904
rect 91200 115880 92000 115910
rect 87944 115839 88264 115840
rect 1944 115360 2264 115361
rect 1944 115296 1952 115360
rect 2016 115296 2032 115360
rect 2096 115296 2112 115360
rect 2176 115296 2192 115360
rect 2256 115296 2264 115360
rect 1944 115295 2264 115296
rect 85944 115360 86264 115361
rect 85944 115296 85952 115360
rect 86016 115296 86032 115360
rect 86096 115296 86112 115360
rect 86176 115296 86192 115360
rect 86256 115296 86264 115360
rect 85944 115295 86264 115296
rect 89944 115360 90264 115361
rect 89944 115296 89952 115360
rect 90016 115296 90032 115360
rect 90096 115296 90112 115360
rect 90176 115296 90192 115360
rect 90256 115296 90264 115360
rect 89944 115295 90264 115296
rect 5441 115018 5507 115021
rect 5441 115016 6194 115018
rect 5441 114960 5446 115016
rect 5502 114960 6194 115016
rect 5441 114958 6194 114960
rect 5441 114955 5507 114958
rect 91200 114882 92000 114912
rect 89670 114822 92000 114882
rect 3944 114816 4264 114817
rect 3944 114752 3952 114816
rect 4016 114752 4032 114816
rect 4096 114752 4112 114816
rect 4176 114752 4192 114816
rect 4256 114752 4264 114816
rect 3944 114751 4264 114752
rect 87944 114816 88264 114817
rect 87944 114752 87952 114816
rect 88016 114752 88032 114816
rect 88096 114752 88112 114816
rect 88176 114752 88192 114816
rect 88256 114752 88264 114816
rect 87944 114751 88264 114752
rect 87965 114610 88031 114613
rect 89670 114610 89730 114822
rect 91200 114792 92000 114822
rect 87965 114608 89730 114610
rect 87965 114552 87970 114608
rect 88026 114552 89730 114608
rect 87965 114550 89730 114552
rect 87965 114547 88031 114550
rect 82629 114338 82695 114341
rect 83406 114338 83412 114340
rect 82629 114336 83412 114338
rect 82629 114280 82634 114336
rect 82690 114280 83412 114336
rect 82629 114278 83412 114280
rect 82629 114275 82695 114278
rect 83406 114276 83412 114278
rect 83476 114276 83482 114340
rect 1944 114272 2264 114273
rect 1944 114208 1952 114272
rect 2016 114208 2032 114272
rect 2096 114208 2112 114272
rect 2176 114208 2192 114272
rect 2256 114208 2264 114272
rect 1944 114207 2264 114208
rect 85944 114272 86264 114273
rect 85944 114208 85952 114272
rect 86016 114208 86032 114272
rect 86096 114208 86112 114272
rect 86176 114208 86192 114272
rect 86256 114208 86264 114272
rect 85944 114207 86264 114208
rect 89944 114272 90264 114273
rect 89944 114208 89952 114272
rect 90016 114208 90032 114272
rect 90096 114208 90112 114272
rect 90176 114208 90192 114272
rect 90256 114208 90264 114272
rect 89944 114207 90264 114208
rect 83406 113868 83412 113932
rect 83476 113930 83482 113932
rect 83958 113930 83964 113932
rect 83476 113870 83964 113930
rect 83476 113868 83482 113870
rect 83958 113868 83964 113870
rect 84028 113868 84034 113932
rect 3944 113728 4264 113729
rect 3944 113664 3952 113728
rect 4016 113664 4032 113728
rect 4096 113664 4112 113728
rect 4176 113664 4192 113728
rect 4256 113664 4264 113728
rect 3944 113663 4264 113664
rect 87944 113728 88264 113729
rect 87944 113664 87952 113728
rect 88016 113664 88032 113728
rect 88096 113664 88112 113728
rect 88176 113664 88192 113728
rect 88256 113664 88264 113728
rect 87944 113663 88264 113664
rect 91200 113658 92000 113688
rect 89670 113598 92000 113658
rect 86493 113522 86559 113525
rect 89670 113522 89730 113598
rect 91200 113568 92000 113598
rect 86493 113520 89730 113522
rect 86493 113464 86498 113520
rect 86554 113464 89730 113520
rect 86493 113462 89730 113464
rect 86493 113459 86559 113462
rect 1944 113184 2264 113185
rect 1944 113120 1952 113184
rect 2016 113120 2032 113184
rect 2096 113120 2112 113184
rect 2176 113120 2192 113184
rect 2256 113120 2264 113184
rect 1944 113119 2264 113120
rect 85944 113184 86264 113185
rect 85944 113120 85952 113184
rect 86016 113120 86032 113184
rect 86096 113120 86112 113184
rect 86176 113120 86192 113184
rect 86256 113120 86264 113184
rect 85944 113119 86264 113120
rect 89944 113184 90264 113185
rect 89944 113120 89952 113184
rect 90016 113120 90032 113184
rect 90096 113120 90112 113184
rect 90176 113120 90192 113184
rect 90256 113120 90264 113184
rect 89944 113119 90264 113120
rect 3944 112640 4264 112641
rect 3944 112576 3952 112640
rect 4016 112576 4032 112640
rect 4096 112576 4112 112640
rect 4176 112576 4192 112640
rect 4256 112576 4264 112640
rect 3944 112575 4264 112576
rect 87944 112640 88264 112641
rect 87944 112576 87952 112640
rect 88016 112576 88032 112640
rect 88096 112576 88112 112640
rect 88176 112576 88192 112640
rect 88256 112576 88264 112640
rect 87944 112575 88264 112576
rect 87965 112434 88031 112437
rect 91200 112434 92000 112464
rect 87965 112432 92000 112434
rect 87965 112376 87970 112432
rect 88026 112376 92000 112432
rect 87965 112374 92000 112376
rect 87965 112371 88031 112374
rect 91200 112344 92000 112374
rect 1944 112096 2264 112097
rect 1944 112032 1952 112096
rect 2016 112032 2032 112096
rect 2096 112032 2112 112096
rect 2176 112032 2192 112096
rect 2256 112032 2264 112096
rect 1944 112031 2264 112032
rect 85944 112096 86264 112097
rect 85944 112032 85952 112096
rect 86016 112032 86032 112096
rect 86096 112032 86112 112096
rect 86176 112032 86192 112096
rect 86256 112032 86264 112096
rect 85944 112031 86264 112032
rect 89944 112096 90264 112097
rect 89944 112032 89952 112096
rect 90016 112032 90032 112096
rect 90096 112032 90112 112096
rect 90176 112032 90192 112096
rect 90256 112032 90264 112096
rect 89944 112031 90264 112032
rect 3944 111552 4264 111553
rect 3944 111488 3952 111552
rect 4016 111488 4032 111552
rect 4096 111488 4112 111552
rect 4176 111488 4192 111552
rect 4256 111488 4264 111552
rect 3944 111487 4264 111488
rect 87944 111552 88264 111553
rect 87944 111488 87952 111552
rect 88016 111488 88032 111552
rect 88096 111488 88112 111552
rect 88176 111488 88192 111552
rect 88256 111488 88264 111552
rect 87944 111487 88264 111488
rect 88241 111210 88307 111213
rect 91200 111210 92000 111240
rect 88241 111208 92000 111210
rect 88241 111152 88246 111208
rect 88302 111152 92000 111208
rect 88241 111150 92000 111152
rect 88241 111147 88307 111150
rect 91200 111120 92000 111150
rect 1944 111008 2264 111009
rect 1944 110944 1952 111008
rect 2016 110944 2032 111008
rect 2096 110944 2112 111008
rect 2176 110944 2192 111008
rect 2256 110944 2264 111008
rect 1944 110943 2264 110944
rect 85944 111008 86264 111009
rect 85944 110944 85952 111008
rect 86016 110944 86032 111008
rect 86096 110944 86112 111008
rect 86176 110944 86192 111008
rect 86256 110944 86264 111008
rect 85944 110943 86264 110944
rect 89944 111008 90264 111009
rect 89944 110944 89952 111008
rect 90016 110944 90032 111008
rect 90096 110944 90112 111008
rect 90176 110944 90192 111008
rect 90256 110944 90264 111008
rect 89944 110943 90264 110944
rect 3944 110464 4264 110465
rect 3944 110400 3952 110464
rect 4016 110400 4032 110464
rect 4096 110400 4112 110464
rect 4176 110400 4192 110464
rect 4256 110400 4264 110464
rect 3944 110399 4264 110400
rect 87944 110464 88264 110465
rect 87944 110400 87952 110464
rect 88016 110400 88032 110464
rect 88096 110400 88112 110464
rect 88176 110400 88192 110464
rect 88256 110400 88264 110464
rect 87944 110399 88264 110400
rect 91200 109986 92000 110016
rect 90406 109926 92000 109986
rect 1944 109920 2264 109921
rect 1944 109856 1952 109920
rect 2016 109856 2032 109920
rect 2096 109856 2112 109920
rect 2176 109856 2192 109920
rect 2256 109856 2264 109920
rect 1944 109855 2264 109856
rect 85944 109920 86264 109921
rect 85944 109856 85952 109920
rect 86016 109856 86032 109920
rect 86096 109856 86112 109920
rect 86176 109856 86192 109920
rect 86256 109856 86264 109920
rect 85944 109855 86264 109856
rect 89944 109920 90264 109921
rect 89944 109856 89952 109920
rect 90016 109856 90032 109920
rect 90096 109856 90112 109920
rect 90176 109856 90192 109920
rect 90256 109856 90264 109920
rect 89944 109855 90264 109856
rect 90406 109714 90466 109926
rect 91200 109896 92000 109926
rect 89670 109654 90466 109714
rect 3944 109376 4264 109377
rect 3944 109312 3952 109376
rect 4016 109312 4032 109376
rect 4096 109312 4112 109376
rect 4176 109312 4192 109376
rect 4256 109312 4264 109376
rect 3944 109311 4264 109312
rect 87944 109376 88264 109377
rect 87944 109312 87952 109376
rect 88016 109312 88032 109376
rect 88096 109312 88112 109376
rect 88176 109312 88192 109376
rect 88256 109312 88264 109376
rect 87944 109311 88264 109312
rect 86902 109108 86908 109172
rect 86972 109170 86978 109172
rect 87229 109170 87295 109173
rect 86972 109168 87295 109170
rect 86972 109112 87234 109168
rect 87290 109112 87295 109168
rect 86972 109110 87295 109112
rect 86972 109108 86978 109110
rect 87229 109107 87295 109110
rect 88241 109170 88307 109173
rect 89670 109170 89730 109654
rect 88241 109168 89730 109170
rect 88241 109112 88246 109168
rect 88302 109112 89730 109168
rect 88241 109110 89730 109112
rect 88241 109107 88307 109110
rect 1944 108832 2264 108833
rect 1944 108768 1952 108832
rect 2016 108768 2032 108832
rect 2096 108768 2112 108832
rect 2176 108768 2192 108832
rect 2256 108768 2264 108832
rect 1944 108767 2264 108768
rect 85944 108832 86264 108833
rect 85944 108768 85952 108832
rect 86016 108768 86032 108832
rect 86096 108768 86112 108832
rect 86176 108768 86192 108832
rect 86256 108768 86264 108832
rect 85944 108767 86264 108768
rect 89944 108832 90264 108833
rect 89944 108768 89952 108832
rect 90016 108768 90032 108832
rect 90096 108768 90112 108832
rect 90176 108768 90192 108832
rect 90256 108768 90264 108832
rect 89944 108767 90264 108768
rect 86902 108700 86908 108764
rect 86972 108762 86978 108764
rect 87321 108762 87387 108765
rect 91200 108762 92000 108792
rect 86972 108760 87387 108762
rect 86972 108704 87326 108760
rect 87382 108704 87387 108760
rect 86972 108702 87387 108704
rect 86972 108700 86978 108702
rect 87321 108699 87387 108702
rect 90406 108702 92000 108762
rect 85614 108564 85620 108628
rect 85684 108626 85690 108628
rect 87229 108626 87295 108629
rect 85684 108624 87295 108626
rect 85684 108568 87234 108624
rect 87290 108568 87295 108624
rect 85684 108566 87295 108568
rect 85684 108564 85690 108566
rect 87229 108563 87295 108566
rect 87965 108626 88031 108629
rect 90406 108626 90466 108702
rect 91200 108672 92000 108702
rect 87965 108624 90466 108626
rect 87965 108568 87970 108624
rect 88026 108568 90466 108624
rect 87965 108566 90466 108568
rect 87965 108563 88031 108566
rect 3944 108288 4264 108289
rect 3944 108224 3952 108288
rect 4016 108224 4032 108288
rect 4096 108224 4112 108288
rect 4176 108224 4192 108288
rect 4256 108224 4264 108288
rect 3944 108223 4264 108224
rect 87944 108288 88264 108289
rect 87944 108224 87952 108288
rect 88016 108224 88032 108288
rect 88096 108224 88112 108288
rect 88176 108224 88192 108288
rect 88256 108224 88264 108288
rect 87944 108223 88264 108224
rect 1944 107744 2264 107745
rect 1944 107680 1952 107744
rect 2016 107680 2032 107744
rect 2096 107680 2112 107744
rect 2176 107680 2192 107744
rect 2256 107680 2264 107744
rect 1944 107679 2264 107680
rect 85944 107744 86264 107745
rect 85944 107680 85952 107744
rect 86016 107680 86032 107744
rect 86096 107680 86112 107744
rect 86176 107680 86192 107744
rect 86256 107680 86264 107744
rect 85944 107679 86264 107680
rect 89944 107744 90264 107745
rect 89944 107680 89952 107744
rect 90016 107680 90032 107744
rect 90096 107680 90112 107744
rect 90176 107680 90192 107744
rect 90256 107680 90264 107744
rect 89944 107679 90264 107680
rect 87965 107538 88031 107541
rect 91200 107538 92000 107568
rect 87965 107536 92000 107538
rect 87965 107480 87970 107536
rect 88026 107480 92000 107536
rect 87965 107478 92000 107480
rect 87965 107475 88031 107478
rect 91200 107448 92000 107478
rect 3944 107200 4264 107201
rect 3944 107136 3952 107200
rect 4016 107136 4032 107200
rect 4096 107136 4112 107200
rect 4176 107136 4192 107200
rect 4256 107136 4264 107200
rect 3944 107135 4264 107136
rect 87944 107200 88264 107201
rect 87944 107136 87952 107200
rect 88016 107136 88032 107200
rect 88096 107136 88112 107200
rect 88176 107136 88192 107200
rect 88256 107136 88264 107200
rect 87944 107135 88264 107136
rect 1944 106656 2264 106657
rect 1944 106592 1952 106656
rect 2016 106592 2032 106656
rect 2096 106592 2112 106656
rect 2176 106592 2192 106656
rect 2256 106592 2264 106656
rect 1944 106591 2264 106592
rect 85944 106656 86264 106657
rect 85944 106592 85952 106656
rect 86016 106592 86032 106656
rect 86096 106592 86112 106656
rect 86176 106592 86192 106656
rect 86256 106592 86264 106656
rect 85944 106591 86264 106592
rect 89944 106656 90264 106657
rect 89944 106592 89952 106656
rect 90016 106592 90032 106656
rect 90096 106592 90112 106656
rect 90176 106592 90192 106656
rect 90256 106592 90264 106656
rect 89944 106591 90264 106592
rect 86401 106314 86467 106317
rect 91200 106314 92000 106344
rect 86401 106312 92000 106314
rect 86401 106256 86406 106312
rect 86462 106256 92000 106312
rect 86401 106254 92000 106256
rect 86401 106251 86467 106254
rect 91200 106224 92000 106254
rect 3944 106112 4264 106113
rect 3944 106048 3952 106112
rect 4016 106048 4032 106112
rect 4096 106048 4112 106112
rect 4176 106048 4192 106112
rect 4256 106048 4264 106112
rect 3944 106047 4264 106048
rect 87944 106112 88264 106113
rect 87944 106048 87952 106112
rect 88016 106048 88032 106112
rect 88096 106048 88112 106112
rect 88176 106048 88192 106112
rect 88256 106048 88264 106112
rect 87944 106047 88264 106048
rect 1944 105568 2264 105569
rect 1944 105504 1952 105568
rect 2016 105504 2032 105568
rect 2096 105504 2112 105568
rect 2176 105504 2192 105568
rect 2256 105504 2264 105568
rect 1944 105503 2264 105504
rect 85944 105568 86264 105569
rect 85944 105504 85952 105568
rect 86016 105504 86032 105568
rect 86096 105504 86112 105568
rect 86176 105504 86192 105568
rect 86256 105504 86264 105568
rect 85944 105503 86264 105504
rect 89944 105568 90264 105569
rect 89944 105504 89952 105568
rect 90016 105504 90032 105568
rect 90096 105504 90112 105568
rect 90176 105504 90192 105568
rect 90256 105504 90264 105568
rect 89944 105503 90264 105504
rect 88517 105090 88583 105093
rect 91200 105090 92000 105120
rect 88517 105088 92000 105090
rect 88517 105032 88522 105088
rect 88578 105032 92000 105088
rect 88517 105030 92000 105032
rect 88517 105027 88583 105030
rect 3944 105024 4264 105025
rect 3944 104960 3952 105024
rect 4016 104960 4032 105024
rect 4096 104960 4112 105024
rect 4176 104960 4192 105024
rect 4256 104960 4264 105024
rect 3944 104959 4264 104960
rect 87944 105024 88264 105025
rect 87944 104960 87952 105024
rect 88016 104960 88032 105024
rect 88096 104960 88112 105024
rect 88176 104960 88192 105024
rect 88256 104960 88264 105024
rect 91200 105000 92000 105030
rect 87944 104959 88264 104960
rect 86677 104682 86743 104685
rect 86358 104680 86743 104682
rect 86358 104624 86682 104680
rect 86738 104624 86743 104680
rect 86358 104622 86743 104624
rect 1944 104480 2264 104481
rect 1944 104416 1952 104480
rect 2016 104416 2032 104480
rect 2096 104416 2112 104480
rect 2176 104416 2192 104480
rect 2256 104416 2264 104480
rect 1944 104415 2264 104416
rect 85944 104480 86264 104481
rect 85944 104416 85952 104480
rect 86016 104416 86032 104480
rect 86096 104416 86112 104480
rect 86176 104416 86192 104480
rect 86256 104416 86264 104480
rect 85944 104415 86264 104416
rect 85665 104138 85731 104141
rect 86358 104138 86418 104622
rect 86677 104619 86743 104622
rect 89944 104480 90264 104481
rect 89944 104416 89952 104480
rect 90016 104416 90032 104480
rect 90096 104416 90112 104480
rect 90176 104416 90192 104480
rect 90256 104416 90264 104480
rect 89944 104415 90264 104416
rect 87137 104274 87203 104277
rect 87321 104274 87387 104277
rect 87137 104272 87387 104274
rect 87137 104216 87142 104272
rect 87198 104216 87326 104272
rect 87382 104216 87387 104272
rect 87137 104214 87387 104216
rect 87137 104211 87203 104214
rect 87321 104211 87387 104214
rect 85665 104136 86418 104138
rect 85665 104080 85670 104136
rect 85726 104080 86418 104136
rect 85665 104078 86418 104080
rect 85665 104075 85731 104078
rect 3944 103936 4264 103937
rect 3944 103872 3952 103936
rect 4016 103872 4032 103936
rect 4096 103872 4112 103936
rect 4176 103872 4192 103936
rect 4256 103872 4264 103936
rect 3944 103871 4264 103872
rect 87944 103936 88264 103937
rect 87944 103872 87952 103936
rect 88016 103872 88032 103936
rect 88096 103872 88112 103936
rect 88176 103872 88192 103936
rect 88256 103872 88264 103936
rect 87944 103871 88264 103872
rect 91200 103866 92000 103896
rect 89670 103806 92000 103866
rect 86718 103668 86724 103732
rect 86788 103730 86794 103732
rect 89670 103730 89730 103806
rect 91200 103776 92000 103806
rect 86788 103670 89730 103730
rect 86788 103668 86794 103670
rect 1944 103392 2264 103393
rect 1944 103328 1952 103392
rect 2016 103328 2032 103392
rect 2096 103328 2112 103392
rect 2176 103328 2192 103392
rect 2256 103328 2264 103392
rect 1944 103327 2264 103328
rect 85944 103392 86264 103393
rect 85944 103328 85952 103392
rect 86016 103328 86032 103392
rect 86096 103328 86112 103392
rect 86176 103328 86192 103392
rect 86256 103328 86264 103392
rect 85944 103327 86264 103328
rect 89944 103392 90264 103393
rect 89944 103328 89952 103392
rect 90016 103328 90032 103392
rect 90096 103328 90112 103392
rect 90176 103328 90192 103392
rect 90256 103328 90264 103392
rect 89944 103327 90264 103328
rect 3944 102848 4264 102849
rect 3944 102784 3952 102848
rect 4016 102784 4032 102848
rect 4096 102784 4112 102848
rect 4176 102784 4192 102848
rect 4256 102784 4264 102848
rect 3944 102783 4264 102784
rect 87944 102848 88264 102849
rect 87944 102784 87952 102848
rect 88016 102784 88032 102848
rect 88096 102784 88112 102848
rect 88176 102784 88192 102848
rect 88256 102784 88264 102848
rect 87944 102783 88264 102784
rect 86902 102580 86908 102644
rect 86972 102642 86978 102644
rect 91200 102642 92000 102672
rect 86972 102582 92000 102642
rect 86972 102580 86978 102582
rect 91200 102552 92000 102582
rect 1944 102304 2264 102305
rect 1944 102240 1952 102304
rect 2016 102240 2032 102304
rect 2096 102240 2112 102304
rect 2176 102240 2192 102304
rect 2256 102240 2264 102304
rect 1944 102239 2264 102240
rect 85944 102304 86264 102305
rect 85944 102240 85952 102304
rect 86016 102240 86032 102304
rect 86096 102240 86112 102304
rect 86176 102240 86192 102304
rect 86256 102240 86264 102304
rect 85944 102239 86264 102240
rect 89944 102304 90264 102305
rect 89944 102240 89952 102304
rect 90016 102240 90032 102304
rect 90096 102240 90112 102304
rect 90176 102240 90192 102304
rect 90256 102240 90264 102304
rect 89944 102239 90264 102240
rect 3944 101760 4264 101761
rect 3944 101696 3952 101760
rect 4016 101696 4032 101760
rect 4096 101696 4112 101760
rect 4176 101696 4192 101760
rect 4256 101696 4264 101760
rect 3944 101695 4264 101696
rect 87944 101760 88264 101761
rect 87944 101696 87952 101760
rect 88016 101696 88032 101760
rect 88096 101696 88112 101760
rect 88176 101696 88192 101760
rect 88256 101696 88264 101760
rect 87944 101695 88264 101696
rect 86585 101418 86651 101421
rect 91200 101418 92000 101448
rect 86585 101416 92000 101418
rect 86585 101360 86590 101416
rect 86646 101360 92000 101416
rect 86585 101358 92000 101360
rect 86585 101355 86651 101358
rect 91200 101328 92000 101358
rect 1944 101216 2264 101217
rect 1944 101152 1952 101216
rect 2016 101152 2032 101216
rect 2096 101152 2112 101216
rect 2176 101152 2192 101216
rect 2256 101152 2264 101216
rect 1944 101151 2264 101152
rect 85944 101216 86264 101217
rect 85944 101152 85952 101216
rect 86016 101152 86032 101216
rect 86096 101152 86112 101216
rect 86176 101152 86192 101216
rect 86256 101152 86264 101216
rect 85944 101151 86264 101152
rect 89944 101216 90264 101217
rect 89944 101152 89952 101216
rect 90016 101152 90032 101216
rect 90096 101152 90112 101216
rect 90176 101152 90192 101216
rect 90256 101152 90264 101216
rect 89944 101151 90264 101152
rect 3944 100672 4264 100673
rect 3944 100608 3952 100672
rect 4016 100608 4032 100672
rect 4096 100608 4112 100672
rect 4176 100608 4192 100672
rect 4256 100608 4264 100672
rect 3944 100607 4264 100608
rect 87944 100672 88264 100673
rect 87944 100608 87952 100672
rect 88016 100608 88032 100672
rect 88096 100608 88112 100672
rect 88176 100608 88192 100672
rect 88256 100608 88264 100672
rect 87944 100607 88264 100608
rect 90357 100194 90423 100197
rect 91200 100194 92000 100224
rect 90357 100192 92000 100194
rect 90357 100136 90362 100192
rect 90418 100136 92000 100192
rect 90357 100134 92000 100136
rect 90357 100131 90423 100134
rect 1944 100128 2264 100129
rect 1944 100064 1952 100128
rect 2016 100064 2032 100128
rect 2096 100064 2112 100128
rect 2176 100064 2192 100128
rect 2256 100064 2264 100128
rect 1944 100063 2264 100064
rect 85944 100128 86264 100129
rect 85944 100064 85952 100128
rect 86016 100064 86032 100128
rect 86096 100064 86112 100128
rect 86176 100064 86192 100128
rect 86256 100064 86264 100128
rect 85944 100063 86264 100064
rect 89944 100128 90264 100129
rect 89944 100064 89952 100128
rect 90016 100064 90032 100128
rect 90096 100064 90112 100128
rect 90176 100064 90192 100128
rect 90256 100064 90264 100128
rect 91200 100104 92000 100134
rect 89944 100063 90264 100064
rect 86861 99786 86927 99789
rect 86861 99784 87154 99786
rect 86861 99728 86866 99784
rect 86922 99728 87154 99784
rect 86861 99726 87154 99728
rect 86861 99723 86927 99726
rect 3944 99584 4264 99585
rect 3944 99520 3952 99584
rect 4016 99520 4032 99584
rect 4096 99520 4112 99584
rect 4176 99520 4192 99584
rect 4256 99520 4264 99584
rect 3944 99519 4264 99520
rect 84193 99514 84259 99517
rect 84510 99514 84516 99516
rect 84193 99512 84516 99514
rect 84193 99456 84198 99512
rect 84254 99456 84516 99512
rect 84193 99454 84516 99456
rect 84193 99451 84259 99454
rect 84510 99452 84516 99454
rect 84580 99452 84586 99516
rect 85113 99514 85179 99517
rect 85430 99514 85436 99516
rect 85113 99512 85436 99514
rect 85113 99456 85118 99512
rect 85174 99456 85436 99512
rect 85113 99454 85436 99456
rect 85113 99451 85179 99454
rect 85430 99452 85436 99454
rect 85500 99452 85506 99516
rect 86677 99514 86743 99517
rect 86902 99514 86908 99516
rect 86677 99512 86908 99514
rect 86677 99456 86682 99512
rect 86738 99456 86908 99512
rect 86677 99454 86908 99456
rect 86677 99451 86743 99454
rect 86902 99452 86908 99454
rect 86972 99452 86978 99516
rect 87094 99393 87154 99726
rect 87944 99584 88264 99585
rect 87944 99520 87952 99584
rect 88016 99520 88032 99584
rect 88096 99520 88112 99584
rect 88176 99520 88192 99584
rect 88256 99520 88264 99584
rect 87944 99519 88264 99520
rect 87094 99388 87203 99393
rect 84510 99316 84516 99380
rect 84580 99378 84586 99380
rect 85113 99378 85179 99381
rect 84580 99376 85179 99378
rect 84580 99320 85118 99376
rect 85174 99320 85179 99376
rect 84580 99318 85179 99320
rect 84580 99316 84586 99318
rect 85113 99315 85179 99318
rect 86493 99378 86559 99381
rect 86718 99378 86724 99380
rect 86493 99376 86724 99378
rect 86493 99320 86498 99376
rect 86554 99320 86724 99376
rect 86493 99318 86724 99320
rect 86493 99315 86559 99318
rect 86718 99316 86724 99318
rect 86788 99316 86794 99380
rect 87094 99332 87142 99388
rect 87198 99332 87203 99388
rect 87094 99330 87203 99332
rect 87137 99327 87203 99330
rect 85389 99108 85455 99109
rect 85389 99106 85436 99108
rect 85344 99104 85436 99106
rect 85344 99048 85394 99104
rect 85344 99046 85436 99048
rect 85389 99044 85436 99046
rect 85500 99044 85506 99108
rect 85389 99043 85455 99044
rect 1944 99040 2264 99041
rect 1944 98976 1952 99040
rect 2016 98976 2032 99040
rect 2096 98976 2112 99040
rect 2176 98976 2192 99040
rect 2256 98976 2264 99040
rect 1944 98975 2264 98976
rect 85944 99040 86264 99041
rect 85944 98976 85952 99040
rect 86016 98976 86032 99040
rect 86096 98976 86112 99040
rect 86176 98976 86192 99040
rect 86256 98976 86264 99040
rect 85944 98975 86264 98976
rect 89944 99040 90264 99041
rect 89944 98976 89952 99040
rect 90016 98976 90032 99040
rect 90096 98976 90112 99040
rect 90176 98976 90192 99040
rect 90256 98976 90264 99040
rect 89944 98975 90264 98976
rect 91200 98970 92000 99000
rect 90406 98910 92000 98970
rect 87597 98834 87663 98837
rect 90406 98834 90466 98910
rect 91200 98880 92000 98910
rect 87597 98832 90466 98834
rect 87597 98776 87602 98832
rect 87658 98776 90466 98832
rect 87597 98774 90466 98776
rect 87597 98771 87663 98774
rect 3944 98496 4264 98497
rect 3944 98432 3952 98496
rect 4016 98432 4032 98496
rect 4096 98432 4112 98496
rect 4176 98432 4192 98496
rect 4256 98432 4264 98496
rect 3944 98431 4264 98432
rect 87944 98496 88264 98497
rect 87944 98432 87952 98496
rect 88016 98432 88032 98496
rect 88096 98432 88112 98496
rect 88176 98432 88192 98496
rect 88256 98432 88264 98496
rect 87944 98431 88264 98432
rect 89110 98092 89116 98156
rect 89180 98154 89186 98156
rect 90582 98154 90588 98156
rect 89180 98094 90588 98154
rect 89180 98092 89186 98094
rect 90582 98092 90588 98094
rect 90652 98092 90658 98156
rect 1944 97952 2264 97953
rect 1944 97888 1952 97952
rect 2016 97888 2032 97952
rect 2096 97888 2112 97952
rect 2176 97888 2192 97952
rect 2256 97888 2264 97952
rect 1944 97887 2264 97888
rect 85944 97952 86264 97953
rect 85944 97888 85952 97952
rect 86016 97888 86032 97952
rect 86096 97888 86112 97952
rect 86176 97888 86192 97952
rect 86256 97888 86264 97952
rect 85944 97887 86264 97888
rect 89944 97952 90264 97953
rect 89944 97888 89952 97952
rect 90016 97888 90032 97952
rect 90096 97888 90112 97952
rect 90176 97888 90192 97952
rect 90256 97888 90264 97952
rect 89944 97887 90264 97888
rect 87229 97882 87295 97885
rect 89294 97882 89300 97884
rect 87229 97880 89300 97882
rect 87229 97824 87234 97880
rect 87290 97824 89300 97880
rect 87229 97822 89300 97824
rect 87229 97819 87295 97822
rect 89294 97820 89300 97822
rect 89364 97820 89370 97884
rect 86953 97746 87019 97749
rect 91200 97746 92000 97776
rect 86953 97744 92000 97746
rect 86953 97688 86958 97744
rect 87014 97688 92000 97744
rect 86953 97686 92000 97688
rect 86953 97683 87019 97686
rect 91200 97656 92000 97686
rect 82813 97610 82879 97613
rect 88701 97610 88767 97613
rect 82813 97608 88767 97610
rect 82813 97552 82818 97608
rect 82874 97552 88706 97608
rect 88762 97552 88767 97608
rect 82813 97550 88767 97552
rect 82813 97547 82879 97550
rect 88701 97547 88767 97550
rect 84745 97474 84811 97477
rect 85021 97474 85087 97477
rect 84745 97472 85087 97474
rect 84745 97416 84750 97472
rect 84806 97416 85026 97472
rect 85082 97416 85087 97472
rect 84745 97414 85087 97416
rect 84745 97411 84811 97414
rect 85021 97411 85087 97414
rect 3944 97408 4264 97409
rect 3944 97344 3952 97408
rect 4016 97344 4032 97408
rect 4096 97344 4112 97408
rect 4176 97344 4192 97408
rect 4256 97344 4264 97408
rect 3944 97343 4264 97344
rect 87944 97408 88264 97409
rect 87944 97344 87952 97408
rect 88016 97344 88032 97408
rect 88096 97344 88112 97408
rect 88176 97344 88192 97408
rect 88256 97344 88264 97408
rect 87944 97343 88264 97344
rect 85246 97338 85252 97340
rect 40358 97278 85252 97338
rect 21909 97202 21975 97205
rect 22645 97204 22711 97205
rect 40358 97204 40418 97278
rect 85246 97276 85252 97278
rect 85316 97276 85322 97340
rect 22645 97202 22692 97204
rect 21909 97200 22692 97202
rect 21909 97144 21914 97200
rect 21970 97144 22650 97200
rect 21909 97142 22692 97144
rect 21909 97139 21975 97142
rect 22645 97140 22692 97142
rect 22756 97140 22762 97204
rect 40350 97140 40356 97204
rect 40420 97140 40426 97204
rect 78949 97202 79015 97205
rect 79910 97202 79916 97204
rect 40910 97142 78874 97202
rect 22645 97139 22711 97140
rect 14641 97068 14707 97069
rect 14590 97066 14596 97068
rect 14550 97006 14596 97066
rect 14660 97064 14707 97068
rect 14702 97008 14707 97064
rect 14590 97004 14596 97006
rect 14660 97004 14707 97008
rect 14641 97003 14707 97004
rect 17125 97068 17191 97069
rect 18045 97068 18111 97069
rect 24301 97068 24367 97069
rect 25405 97068 25471 97069
rect 30097 97068 30163 97069
rect 17125 97064 17172 97068
rect 17236 97066 17242 97068
rect 17125 97008 17130 97064
rect 17125 97004 17172 97008
rect 17236 97006 17282 97066
rect 18045 97064 18092 97068
rect 18156 97066 18162 97068
rect 18045 97008 18050 97064
rect 17236 97004 17242 97006
rect 18045 97004 18092 97008
rect 18156 97006 18202 97066
rect 24301 97064 24348 97068
rect 24412 97066 24418 97068
rect 24301 97008 24306 97064
rect 18156 97004 18162 97006
rect 24301 97004 24348 97008
rect 24412 97006 24458 97066
rect 25405 97064 25452 97068
rect 25516 97066 25522 97068
rect 30046 97066 30052 97068
rect 25405 97008 25410 97064
rect 24412 97004 24418 97006
rect 25405 97004 25452 97008
rect 25516 97006 25562 97066
rect 30006 97006 30052 97066
rect 30116 97064 30163 97068
rect 30158 97008 30163 97064
rect 25516 97004 25522 97006
rect 30046 97004 30052 97006
rect 30116 97004 30163 97008
rect 17125 97003 17191 97004
rect 18045 97003 18111 97004
rect 24301 97003 24367 97004
rect 25405 97003 25471 97004
rect 30097 97003 30163 97004
rect 32029 97068 32095 97069
rect 33133 97068 33199 97069
rect 32029 97064 32076 97068
rect 32140 97066 32146 97068
rect 32029 97008 32034 97064
rect 32029 97004 32076 97008
rect 32140 97006 32186 97066
rect 33133 97064 33180 97068
rect 33244 97066 33250 97068
rect 33133 97008 33138 97064
rect 32140 97004 32146 97006
rect 33133 97004 33180 97008
rect 33244 97006 33290 97066
rect 33244 97004 33250 97006
rect 32029 97003 32095 97004
rect 33133 97003 33199 97004
rect 5717 96930 5783 96933
rect 6177 96930 6243 96933
rect 35934 96930 35940 96932
rect 5717 96928 35940 96930
rect 5717 96872 5722 96928
rect 5778 96872 6182 96928
rect 6238 96872 35940 96928
rect 5717 96870 35940 96872
rect 5717 96867 5783 96870
rect 6177 96867 6243 96870
rect 35934 96868 35940 96870
rect 36004 96930 36010 96932
rect 40910 96930 40970 97142
rect 42926 97004 42932 97068
rect 42996 97066 43002 97068
rect 77385 97066 77451 97069
rect 78673 97066 78739 97069
rect 42996 97006 77310 97066
rect 42996 97004 43002 97006
rect 54150 96930 54156 96932
rect 36004 96870 40970 96930
rect 51030 96870 54156 96930
rect 36004 96868 36010 96870
rect 1944 96864 2264 96865
rect 1944 96800 1952 96864
rect 2016 96800 2032 96864
rect 2096 96800 2112 96864
rect 2176 96800 2192 96864
rect 2256 96800 2264 96864
rect 1944 96799 2264 96800
rect 5901 96794 5967 96797
rect 6361 96794 6427 96797
rect 40534 96794 40540 96796
rect 5901 96792 40540 96794
rect 5901 96736 5906 96792
rect 5962 96736 6366 96792
rect 6422 96736 40540 96792
rect 5901 96734 40540 96736
rect 5901 96731 5967 96734
rect 6361 96731 6427 96734
rect 40534 96732 40540 96734
rect 40604 96732 40610 96796
rect 47158 96732 47164 96796
rect 47228 96794 47234 96796
rect 51030 96794 51090 96870
rect 54150 96868 54156 96870
rect 54220 96868 54226 96932
rect 54845 96930 54911 96933
rect 60457 96930 60523 96933
rect 54845 96928 60523 96930
rect 54845 96872 54850 96928
rect 54906 96872 60462 96928
rect 60518 96872 60523 96928
rect 54845 96870 60523 96872
rect 54845 96867 54911 96870
rect 60457 96867 60523 96870
rect 60641 96930 60707 96933
rect 77109 96930 77175 96933
rect 60641 96928 77175 96930
rect 60641 96872 60646 96928
rect 60702 96872 77114 96928
rect 77170 96872 77175 96928
rect 60641 96870 77175 96872
rect 77250 96930 77310 97006
rect 77385 97064 78739 97066
rect 77385 97008 77390 97064
rect 77446 97008 78678 97064
rect 78734 97008 78739 97064
rect 77385 97006 78739 97008
rect 78814 97066 78874 97142
rect 78949 97200 79916 97202
rect 78949 97144 78954 97200
rect 79010 97144 79916 97200
rect 78949 97142 79916 97144
rect 78949 97139 79015 97142
rect 79910 97140 79916 97142
rect 79980 97140 79986 97204
rect 80145 97202 80211 97205
rect 87270 97202 87276 97204
rect 80145 97200 87276 97202
rect 80145 97144 80150 97200
rect 80206 97144 87276 97200
rect 80145 97142 87276 97144
rect 80145 97139 80211 97142
rect 87270 97140 87276 97142
rect 87340 97140 87346 97204
rect 83273 97066 83339 97069
rect 87454 97066 87460 97068
rect 78814 97064 83339 97066
rect 78814 97008 83278 97064
rect 83334 97008 83339 97064
rect 78814 97006 83339 97008
rect 77385 97003 77451 97006
rect 78673 97003 78739 97006
rect 83273 97003 83339 97006
rect 85070 97006 87460 97066
rect 84878 96930 84884 96932
rect 77250 96870 84884 96930
rect 60641 96867 60707 96870
rect 77109 96867 77175 96870
rect 84878 96868 84884 96870
rect 84948 96868 84954 96932
rect 61561 96796 61627 96797
rect 61745 96796 61811 96797
rect 47228 96734 51090 96794
rect 47228 96732 47234 96734
rect 52126 96732 52132 96796
rect 52196 96794 52202 96796
rect 60590 96794 60596 96796
rect 52196 96734 60596 96794
rect 52196 96732 52202 96734
rect 60590 96732 60596 96734
rect 60660 96732 60666 96796
rect 61510 96794 61516 96796
rect 61470 96734 61516 96794
rect 61580 96792 61627 96796
rect 61622 96736 61627 96792
rect 61510 96732 61516 96734
rect 61580 96732 61627 96736
rect 61694 96732 61700 96796
rect 61764 96794 61811 96796
rect 61929 96794 61995 96797
rect 79501 96794 79567 96797
rect 61764 96792 61856 96794
rect 61806 96736 61856 96792
rect 61764 96734 61856 96736
rect 61929 96792 79426 96794
rect 61929 96736 61934 96792
rect 61990 96736 79426 96792
rect 61929 96734 79426 96736
rect 61764 96732 61811 96734
rect 61561 96731 61627 96732
rect 61745 96731 61811 96732
rect 61929 96731 61995 96734
rect 5809 96658 5875 96661
rect 42742 96658 42748 96660
rect 5809 96656 42748 96658
rect 5809 96600 5814 96656
rect 5870 96600 42748 96656
rect 5809 96598 42748 96600
rect 5809 96595 5875 96598
rect 42742 96596 42748 96598
rect 42812 96596 42818 96660
rect 53741 96658 53807 96661
rect 57605 96658 57671 96661
rect 57881 96660 57947 96661
rect 58065 96660 58131 96661
rect 57830 96658 57836 96660
rect 53741 96656 57671 96658
rect 53741 96600 53746 96656
rect 53802 96600 57610 96656
rect 57666 96600 57671 96656
rect 53741 96598 57671 96600
rect 57790 96598 57836 96658
rect 57900 96656 57947 96660
rect 57942 96600 57947 96656
rect 53741 96595 53807 96598
rect 57605 96595 57671 96598
rect 57830 96596 57836 96598
rect 57900 96596 57947 96600
rect 58014 96596 58020 96660
rect 58084 96658 58131 96660
rect 58084 96656 58176 96658
rect 58126 96600 58176 96656
rect 58084 96598 58176 96600
rect 58084 96596 58131 96598
rect 58382 96596 58388 96660
rect 58452 96658 58458 96660
rect 59537 96658 59603 96661
rect 59721 96660 59787 96661
rect 58452 96656 59603 96658
rect 58452 96600 59542 96656
rect 59598 96600 59603 96656
rect 58452 96598 59603 96600
rect 58452 96596 58458 96598
rect 57881 96595 57947 96596
rect 58065 96595 58131 96596
rect 59537 96595 59603 96598
rect 59670 96596 59676 96660
rect 59740 96658 59787 96660
rect 59905 96658 59971 96661
rect 60222 96658 60228 96660
rect 59740 96656 59832 96658
rect 59782 96600 59832 96656
rect 59740 96598 59832 96600
rect 59905 96656 60228 96658
rect 59905 96600 59910 96656
rect 59966 96600 60228 96656
rect 59905 96598 60228 96600
rect 59740 96596 59787 96598
rect 59721 96595 59787 96596
rect 59905 96595 59971 96598
rect 60222 96596 60228 96598
rect 60292 96596 60298 96660
rect 60457 96658 60523 96661
rect 76925 96658 76991 96661
rect 60457 96656 76991 96658
rect 60457 96600 60462 96656
rect 60518 96600 76930 96656
rect 76986 96600 76991 96656
rect 60457 96598 76991 96600
rect 60457 96595 60523 96598
rect 76925 96595 76991 96598
rect 77109 96658 77175 96661
rect 79225 96658 79291 96661
rect 77109 96656 79291 96658
rect 77109 96600 77114 96656
rect 77170 96600 79230 96656
rect 79286 96600 79291 96656
rect 77109 96598 79291 96600
rect 79366 96658 79426 96734
rect 79501 96792 82370 96794
rect 79501 96736 79506 96792
rect 79562 96736 82370 96792
rect 79501 96734 82370 96736
rect 79501 96731 79567 96734
rect 82169 96658 82235 96661
rect 79366 96656 82235 96658
rect 79366 96600 82174 96656
rect 82230 96600 82235 96656
rect 79366 96598 82235 96600
rect 82310 96658 82370 96734
rect 82486 96732 82492 96796
rect 82556 96794 82562 96796
rect 82629 96794 82695 96797
rect 82556 96792 82695 96794
rect 82556 96736 82634 96792
rect 82690 96736 82695 96792
rect 82556 96734 82695 96736
rect 82556 96732 82562 96734
rect 82629 96731 82695 96734
rect 82905 96794 82971 96797
rect 85070 96794 85130 97006
rect 87454 97004 87460 97006
rect 87524 97004 87530 97068
rect 85944 96864 86264 96865
rect 85944 96800 85952 96864
rect 86016 96800 86032 96864
rect 86096 96800 86112 96864
rect 86176 96800 86192 96864
rect 86256 96800 86264 96864
rect 85944 96799 86264 96800
rect 89944 96864 90264 96865
rect 89944 96800 89952 96864
rect 90016 96800 90032 96864
rect 90096 96800 90112 96864
rect 90176 96800 90192 96864
rect 90256 96800 90264 96864
rect 89944 96799 90264 96800
rect 87638 96794 87644 96796
rect 82905 96792 85130 96794
rect 82905 96736 82910 96792
rect 82966 96736 85130 96792
rect 82905 96734 85130 96736
rect 86358 96734 87644 96794
rect 82905 96731 82971 96734
rect 86358 96658 86418 96734
rect 87638 96732 87644 96734
rect 87708 96732 87714 96796
rect 82310 96598 86418 96658
rect 86953 96658 87019 96661
rect 91200 96658 92000 96688
rect 86953 96656 92000 96658
rect 86953 96600 86958 96656
rect 87014 96600 92000 96656
rect 86953 96598 92000 96600
rect 77109 96595 77175 96598
rect 79225 96595 79291 96598
rect 82169 96595 82235 96598
rect 86953 96595 87019 96598
rect 91200 96568 92000 96598
rect 16481 96524 16547 96525
rect 16430 96522 16436 96524
rect 16390 96462 16436 96522
rect 16500 96520 16547 96524
rect 85798 96522 85804 96524
rect 16542 96464 16547 96520
rect 16430 96460 16436 96462
rect 16500 96460 16547 96464
rect 16481 96459 16547 96460
rect 28950 96462 85804 96522
rect 15745 96388 15811 96389
rect 15694 96386 15700 96388
rect 15654 96326 15700 96386
rect 15764 96384 15811 96388
rect 15806 96328 15811 96384
rect 15694 96324 15700 96326
rect 15764 96324 15811 96328
rect 21214 96324 21220 96388
rect 21284 96386 21290 96388
rect 28950 96386 29010 96462
rect 85798 96460 85804 96462
rect 85868 96460 85874 96524
rect 21284 96326 29010 96386
rect 46841 96386 46907 96389
rect 50337 96386 50403 96389
rect 46841 96384 50403 96386
rect 46841 96328 46846 96384
rect 46902 96328 50342 96384
rect 50398 96328 50403 96384
rect 46841 96326 50403 96328
rect 21284 96324 21290 96326
rect 15745 96323 15811 96324
rect 46841 96323 46907 96326
rect 50337 96323 50403 96326
rect 50470 96324 50476 96388
rect 50540 96386 50546 96388
rect 51022 96386 51028 96388
rect 50540 96326 51028 96386
rect 50540 96324 50546 96326
rect 51022 96324 51028 96326
rect 51092 96324 51098 96388
rect 51165 96386 51231 96389
rect 80145 96386 80211 96389
rect 87321 96386 87387 96389
rect 51165 96384 80211 96386
rect 51165 96328 51170 96384
rect 51226 96328 80150 96384
rect 80206 96328 80211 96384
rect 51165 96326 80211 96328
rect 51165 96323 51231 96326
rect 80145 96323 80211 96326
rect 80286 96384 87387 96386
rect 80286 96328 87326 96384
rect 87382 96328 87387 96384
rect 80286 96326 87387 96328
rect 3944 96320 4264 96321
rect 3944 96256 3952 96320
rect 4016 96256 4032 96320
rect 4096 96256 4112 96320
rect 4176 96256 4192 96320
rect 4256 96256 4264 96320
rect 3944 96255 4264 96256
rect 9581 96252 9647 96253
rect 22093 96252 22159 96253
rect 27981 96252 28047 96253
rect 29177 96252 29243 96253
rect 9581 96248 9628 96252
rect 9692 96250 9698 96252
rect 9581 96192 9586 96248
rect 9581 96188 9628 96192
rect 9692 96190 9738 96250
rect 22093 96248 22140 96252
rect 22204 96250 22210 96252
rect 22093 96192 22098 96248
rect 9692 96188 9698 96190
rect 22093 96188 22140 96192
rect 22204 96190 22250 96250
rect 22204 96188 22210 96190
rect 27978 96188 27984 96252
rect 28048 96250 28054 96252
rect 29146 96250 29152 96252
rect 28048 96190 28138 96250
rect 29086 96190 29152 96250
rect 29216 96248 29243 96252
rect 29238 96192 29243 96248
rect 28048 96188 28054 96190
rect 29146 96188 29152 96190
rect 29216 96188 29243 96192
rect 9581 96187 9647 96188
rect 22093 96187 22159 96188
rect 27981 96187 28047 96188
rect 29177 96187 29243 96188
rect 41965 96252 42031 96253
rect 41965 96248 42000 96252
rect 42064 96250 42070 96252
rect 44173 96250 44239 96253
rect 80286 96250 80346 96326
rect 87321 96323 87387 96326
rect 87944 96320 88264 96321
rect 87944 96256 87952 96320
rect 88016 96256 88032 96320
rect 88096 96256 88112 96320
rect 88176 96256 88192 96320
rect 88256 96256 88264 96320
rect 87944 96255 88264 96256
rect 41965 96192 41970 96248
rect 41965 96188 42000 96192
rect 42064 96190 42122 96250
rect 44173 96248 80346 96250
rect 44173 96192 44178 96248
rect 44234 96192 80346 96248
rect 44173 96190 80346 96192
rect 80513 96250 80579 96253
rect 84009 96250 84075 96253
rect 80513 96248 84075 96250
rect 80513 96192 80518 96248
rect 80574 96192 84014 96248
rect 84070 96192 84075 96248
rect 80513 96190 84075 96192
rect 42064 96188 42070 96190
rect 41965 96187 42062 96188
rect 44173 96187 44239 96190
rect 80513 96187 80579 96190
rect 84009 96187 84075 96190
rect 20989 96116 21055 96117
rect 20970 96114 20976 96116
rect 20898 96054 20976 96114
rect 21040 96112 21055 96116
rect 21050 96056 21055 96112
rect 20970 96052 20976 96054
rect 21040 96052 21055 96056
rect 20989 96051 21055 96052
rect 26785 96116 26851 96117
rect 31477 96116 31543 96117
rect 34973 96116 35039 96117
rect 26785 96112 26816 96116
rect 26880 96114 26886 96116
rect 26785 96056 26790 96112
rect 26785 96052 26816 96056
rect 26880 96054 26942 96114
rect 31477 96112 31488 96116
rect 31552 96114 31558 96116
rect 31477 96056 31482 96112
rect 26880 96052 26886 96054
rect 31477 96052 31488 96056
rect 31552 96054 31634 96114
rect 34973 96112 34992 96116
rect 35056 96114 35062 96116
rect 42002 96114 42062 96187
rect 79501 96114 79567 96117
rect 34973 96056 34978 96112
rect 31552 96052 31558 96054
rect 34973 96052 34992 96056
rect 35056 96054 35130 96114
rect 42002 96112 79567 96114
rect 42002 96056 79506 96112
rect 79562 96056 79567 96112
rect 42002 96054 79567 96056
rect 35056 96052 35062 96054
rect 26785 96051 26851 96052
rect 31477 96051 31543 96052
rect 34973 96051 35039 96052
rect 79501 96051 79567 96054
rect 79685 96114 79751 96117
rect 83549 96114 83615 96117
rect 79685 96112 83615 96114
rect 79685 96056 79690 96112
rect 79746 96056 83554 96112
rect 83610 96056 83615 96112
rect 79685 96054 83615 96056
rect 79685 96051 79751 96054
rect 83549 96051 83615 96054
rect 39573 95980 39639 95981
rect 39573 95978 39620 95980
rect 39492 95976 39620 95978
rect 39684 95978 39690 95980
rect 74625 95978 74691 95981
rect 39684 95976 74691 95978
rect 39492 95920 39578 95976
rect 39684 95920 74630 95976
rect 74686 95920 74691 95976
rect 39492 95918 39620 95920
rect 39573 95916 39620 95918
rect 39684 95918 74691 95920
rect 39684 95916 39690 95918
rect 39573 95915 39639 95916
rect 74625 95915 74691 95918
rect 74809 95978 74875 95981
rect 76833 95978 76899 95981
rect 74809 95976 76899 95978
rect 74809 95920 74814 95976
rect 74870 95920 76838 95976
rect 76894 95920 76899 95976
rect 74809 95918 76899 95920
rect 74809 95915 74875 95918
rect 76833 95915 76899 95918
rect 77017 95978 77083 95981
rect 80237 95978 80303 95981
rect 77017 95976 80303 95978
rect 77017 95920 77022 95976
rect 77078 95920 80242 95976
rect 80298 95920 80303 95976
rect 77017 95918 80303 95920
rect 77017 95915 77083 95918
rect 80237 95915 80303 95918
rect 80421 95978 80487 95981
rect 87781 95978 87847 95981
rect 80421 95976 87847 95978
rect 80421 95920 80426 95976
rect 80482 95920 87786 95976
rect 87842 95920 87847 95976
rect 80421 95918 87847 95920
rect 80421 95915 80487 95918
rect 87781 95915 87847 95918
rect 38469 95844 38535 95845
rect 38469 95842 38516 95844
rect 38388 95840 38516 95842
rect 38580 95842 38586 95844
rect 83365 95842 83431 95845
rect 38580 95840 83431 95842
rect 38388 95784 38474 95840
rect 38580 95784 83370 95840
rect 83426 95784 83431 95840
rect 38388 95782 38516 95784
rect 38469 95780 38516 95782
rect 38580 95782 83431 95784
rect 38580 95780 38586 95782
rect 38469 95779 38535 95780
rect 83365 95779 83431 95782
rect 1944 95776 2264 95777
rect 1944 95712 1952 95776
rect 2016 95712 2032 95776
rect 2096 95712 2112 95776
rect 2176 95712 2192 95776
rect 2256 95712 2264 95776
rect 1944 95711 2264 95712
rect 85944 95776 86264 95777
rect 85944 95712 85952 95776
rect 86016 95712 86032 95776
rect 86096 95712 86112 95776
rect 86176 95712 86192 95776
rect 86256 95712 86264 95776
rect 85944 95711 86264 95712
rect 89944 95776 90264 95777
rect 89944 95712 89952 95776
rect 90016 95712 90032 95776
rect 90096 95712 90112 95776
rect 90176 95712 90192 95776
rect 90256 95712 90264 95776
rect 89944 95711 90264 95712
rect 32990 95644 32996 95708
rect 33060 95706 33066 95708
rect 74809 95706 74875 95709
rect 82445 95706 82511 95709
rect 33060 95704 74875 95706
rect 33060 95648 74814 95704
rect 74870 95648 74875 95704
rect 33060 95646 74875 95648
rect 33060 95644 33066 95646
rect 74809 95643 74875 95646
rect 74950 95704 82511 95706
rect 74950 95648 82450 95704
rect 82506 95648 82511 95704
rect 74950 95646 82511 95648
rect 28758 95508 28764 95572
rect 28828 95570 28834 95572
rect 74950 95570 75010 95646
rect 82445 95643 82511 95646
rect 75177 95572 75243 95573
rect 75126 95570 75132 95572
rect 28828 95510 75010 95570
rect 75086 95510 75132 95570
rect 75196 95568 75243 95572
rect 75238 95512 75243 95568
rect 28828 95508 28834 95510
rect 75126 95508 75132 95510
rect 75196 95508 75243 95512
rect 75177 95507 75243 95508
rect 76097 95570 76163 95573
rect 79174 95570 79180 95572
rect 76097 95568 79180 95570
rect 76097 95512 76102 95568
rect 76158 95512 79180 95568
rect 76097 95510 79180 95512
rect 76097 95507 76163 95510
rect 79174 95508 79180 95510
rect 79244 95508 79250 95572
rect 86769 95570 86835 95573
rect 79366 95568 86835 95570
rect 79366 95512 86774 95568
rect 86830 95512 86835 95568
rect 79366 95510 86835 95512
rect 23974 95372 23980 95436
rect 24044 95434 24050 95436
rect 79366 95434 79426 95510
rect 86769 95507 86835 95510
rect 24044 95374 79426 95434
rect 79501 95434 79567 95437
rect 85573 95434 85639 95437
rect 79501 95432 85639 95434
rect 79501 95376 79506 95432
rect 79562 95376 85578 95432
rect 85634 95376 85639 95432
rect 79501 95374 85639 95376
rect 24044 95372 24050 95374
rect 79501 95371 79567 95374
rect 85573 95371 85639 95374
rect 86953 95434 87019 95437
rect 91200 95434 92000 95464
rect 86953 95432 92000 95434
rect 86953 95376 86958 95432
rect 87014 95376 92000 95432
rect 86953 95374 92000 95376
rect 86953 95371 87019 95374
rect 91200 95344 92000 95374
rect 24577 95300 24643 95301
rect 37825 95300 37891 95301
rect 41137 95300 41203 95301
rect 45369 95300 45435 95301
rect 47945 95300 48011 95301
rect 24526 95298 24532 95300
rect 24486 95238 24532 95298
rect 24596 95296 24643 95300
rect 37774 95298 37780 95300
rect 24638 95240 24643 95296
rect 24526 95236 24532 95238
rect 24596 95236 24643 95240
rect 37734 95238 37780 95298
rect 37844 95296 37891 95300
rect 41086 95298 41092 95300
rect 37886 95240 37891 95296
rect 37774 95236 37780 95238
rect 37844 95236 37891 95240
rect 41046 95238 41092 95298
rect 41156 95296 41203 95300
rect 45318 95298 45324 95300
rect 41198 95240 41203 95296
rect 41086 95236 41092 95238
rect 41156 95236 41203 95240
rect 45278 95238 45324 95298
rect 45388 95296 45435 95300
rect 45430 95240 45435 95296
rect 45318 95236 45324 95238
rect 45388 95236 45435 95240
rect 47894 95236 47900 95300
rect 47964 95298 48011 95300
rect 48221 95298 48287 95301
rect 63953 95298 64019 95301
rect 64137 95300 64203 95301
rect 47964 95296 48056 95298
rect 48006 95240 48056 95296
rect 47964 95238 48056 95240
rect 48221 95296 64019 95298
rect 48221 95240 48226 95296
rect 48282 95240 63958 95296
rect 64014 95240 64019 95296
rect 48221 95238 64019 95240
rect 47964 95236 48011 95238
rect 24577 95235 24643 95236
rect 37825 95235 37891 95236
rect 41137 95235 41203 95236
rect 45369 95235 45435 95236
rect 47945 95235 48011 95236
rect 48221 95235 48287 95238
rect 63953 95235 64019 95238
rect 64086 95236 64092 95300
rect 64156 95298 64203 95300
rect 64321 95298 64387 95301
rect 85614 95298 85620 95300
rect 64156 95296 64248 95298
rect 64198 95240 64248 95296
rect 64156 95238 64248 95240
rect 64321 95296 85620 95298
rect 64321 95240 64326 95296
rect 64382 95240 85620 95296
rect 64321 95238 85620 95240
rect 64156 95236 64203 95238
rect 64137 95235 64203 95236
rect 64321 95235 64387 95238
rect 85614 95236 85620 95238
rect 85684 95236 85690 95300
rect 3944 95232 4264 95233
rect 3944 95168 3952 95232
rect 4016 95168 4032 95232
rect 4096 95168 4112 95232
rect 4176 95168 4192 95232
rect 4256 95168 4264 95232
rect 3944 95167 4264 95168
rect 87944 95232 88264 95233
rect 87944 95168 87952 95232
rect 88016 95168 88032 95232
rect 88096 95168 88112 95232
rect 88176 95168 88192 95232
rect 88256 95168 88264 95232
rect 87944 95167 88264 95168
rect 12801 95164 12867 95165
rect 12750 95162 12756 95164
rect 12710 95102 12756 95162
rect 12820 95160 12867 95164
rect 12862 95104 12867 95160
rect 12750 95100 12756 95102
rect 12820 95100 12867 95104
rect 12801 95099 12867 95100
rect 19333 95164 19399 95165
rect 24761 95164 24827 95165
rect 19333 95160 19380 95164
rect 19444 95162 19450 95164
rect 19333 95104 19338 95160
rect 19333 95100 19380 95104
rect 19444 95102 19490 95162
rect 19444 95100 19450 95102
rect 24710 95100 24716 95164
rect 24780 95162 24827 95164
rect 24780 95160 24872 95162
rect 24822 95104 24872 95160
rect 24780 95102 24872 95104
rect 24780 95100 24827 95102
rect 25814 95100 25820 95164
rect 25884 95162 25890 95164
rect 25957 95162 26023 95165
rect 25884 95160 26023 95162
rect 25884 95104 25962 95160
rect 26018 95104 26023 95160
rect 25884 95102 26023 95104
rect 25884 95100 25890 95102
rect 19333 95099 19399 95100
rect 24761 95099 24827 95100
rect 25957 95099 26023 95102
rect 27470 95100 27476 95164
rect 27540 95162 27546 95164
rect 27540 95102 35910 95162
rect 27540 95100 27546 95102
rect 22870 94964 22876 95028
rect 22940 95026 22946 95028
rect 23381 95026 23447 95029
rect 22940 95024 23447 95026
rect 22940 94968 23386 95024
rect 23442 94968 23447 95024
rect 22940 94966 23447 94968
rect 22940 94964 22946 94966
rect 23381 94963 23447 94966
rect 29862 94964 29868 95028
rect 29932 95026 29938 95028
rect 30281 95026 30347 95029
rect 29932 95024 30347 95026
rect 29932 94968 30286 95024
rect 30342 94968 30347 95024
rect 29932 94966 30347 94968
rect 29932 94964 29938 94966
rect 30281 94963 30347 94966
rect 30966 94964 30972 95028
rect 31036 95026 31042 95028
rect 31661 95026 31727 95029
rect 31036 95024 31727 95026
rect 31036 94968 31666 95024
rect 31722 94968 31727 95024
rect 31036 94966 31727 94968
rect 35850 95026 35910 95102
rect 37958 95100 37964 95164
rect 38028 95162 38034 95164
rect 38561 95162 38627 95165
rect 38028 95160 38627 95162
rect 38028 95104 38566 95160
rect 38622 95104 38627 95160
rect 38028 95102 38627 95104
rect 38028 95100 38034 95102
rect 38561 95099 38627 95102
rect 43846 95100 43852 95164
rect 43916 95162 43922 95164
rect 44081 95162 44147 95165
rect 43916 95160 44147 95162
rect 43916 95104 44086 95160
rect 44142 95104 44147 95160
rect 43916 95102 44147 95104
rect 43916 95100 43922 95102
rect 44081 95099 44147 95102
rect 44398 95100 44404 95164
rect 44468 95162 44474 95164
rect 45185 95162 45251 95165
rect 45553 95164 45619 95165
rect 46657 95164 46723 95165
rect 48129 95164 48195 95165
rect 44468 95160 45251 95162
rect 44468 95104 45190 95160
rect 45246 95104 45251 95160
rect 44468 95102 45251 95104
rect 44468 95100 44474 95102
rect 45185 95099 45251 95102
rect 45502 95100 45508 95164
rect 45572 95162 45619 95164
rect 46606 95162 46612 95164
rect 45572 95160 45664 95162
rect 45614 95104 45664 95160
rect 45572 95102 45664 95104
rect 46566 95102 46612 95162
rect 46676 95160 46723 95164
rect 46718 95104 46723 95160
rect 45572 95100 45619 95102
rect 46606 95100 46612 95102
rect 46676 95100 46723 95104
rect 48078 95100 48084 95164
rect 48148 95162 48195 95164
rect 50797 95162 50863 95165
rect 83733 95162 83799 95165
rect 48148 95160 48240 95162
rect 48190 95104 48240 95160
rect 48148 95102 48240 95104
rect 50797 95160 83799 95162
rect 50797 95104 50802 95160
rect 50858 95104 83738 95160
rect 83794 95104 83799 95160
rect 50797 95102 83799 95104
rect 48148 95100 48195 95102
rect 45553 95099 45619 95100
rect 46657 95099 46723 95100
rect 48129 95099 48195 95100
rect 50797 95099 50863 95102
rect 83733 95099 83799 95102
rect 79501 95026 79567 95029
rect 35850 95024 79567 95026
rect 35850 94968 79506 95024
rect 79562 94968 79567 95024
rect 35850 94966 79567 94968
rect 31036 94964 31042 94966
rect 31661 94963 31727 94966
rect 79501 94963 79567 94966
rect 79726 94964 79732 95028
rect 79796 95026 79802 95028
rect 80053 95026 80119 95029
rect 80513 95028 80579 95029
rect 79796 95024 80119 95026
rect 79796 94968 80058 95024
rect 80114 94968 80119 95024
rect 79796 94966 80119 94968
rect 79796 94964 79802 94966
rect 80053 94963 80119 94966
rect 80462 94964 80468 95028
rect 80532 95026 80579 95028
rect 81433 95026 81499 95029
rect 82905 95026 82971 95029
rect 80532 95024 80624 95026
rect 80574 94968 80624 95024
rect 80532 94966 80624 94968
rect 81433 95024 82971 95026
rect 81433 94968 81438 95024
rect 81494 94968 82910 95024
rect 82966 94968 82971 95024
rect 81433 94966 82971 94968
rect 80532 94964 80579 94966
rect 80513 94963 80579 94964
rect 81433 94963 81499 94966
rect 82905 94963 82971 94966
rect 19926 94828 19932 94892
rect 19996 94890 20002 94892
rect 20621 94890 20687 94893
rect 19996 94888 20687 94890
rect 19996 94832 20626 94888
rect 20682 94832 20687 94888
rect 19996 94830 20687 94832
rect 19996 94828 20002 94830
rect 20621 94827 20687 94830
rect 31702 94828 31708 94892
rect 31772 94890 31778 94892
rect 83774 94890 83780 94892
rect 31772 94830 83780 94890
rect 31772 94828 31778 94830
rect 83774 94828 83780 94830
rect 83844 94828 83850 94892
rect 34462 94692 34468 94756
rect 34532 94754 34538 94756
rect 84101 94754 84167 94757
rect 34532 94752 84167 94754
rect 34532 94696 84106 94752
rect 84162 94696 84167 94752
rect 34532 94694 84167 94696
rect 34532 94692 34538 94694
rect 84101 94691 84167 94694
rect 1944 94688 2264 94689
rect 1944 94624 1952 94688
rect 2016 94624 2032 94688
rect 2096 94624 2112 94688
rect 2176 94624 2192 94688
rect 2256 94624 2264 94688
rect 1944 94623 2264 94624
rect 85944 94688 86264 94689
rect 85944 94624 85952 94688
rect 86016 94624 86032 94688
rect 86096 94624 86112 94688
rect 86176 94624 86192 94688
rect 86256 94624 86264 94688
rect 85944 94623 86264 94624
rect 89944 94688 90264 94689
rect 89944 94624 89952 94688
rect 90016 94624 90032 94688
rect 90096 94624 90112 94688
rect 90176 94624 90192 94688
rect 90256 94624 90264 94688
rect 89944 94623 90264 94624
rect 37273 94620 37339 94621
rect 37222 94556 37228 94620
rect 37292 94618 37339 94620
rect 82169 94618 82235 94621
rect 37292 94616 37384 94618
rect 37334 94560 37384 94616
rect 37292 94558 37384 94560
rect 40910 94616 82235 94618
rect 40910 94560 82174 94616
rect 82230 94560 82235 94616
rect 40910 94558 82235 94560
rect 37292 94556 37339 94558
rect 37273 94555 37339 94556
rect 36854 94420 36860 94484
rect 36924 94482 36930 94484
rect 40910 94482 40970 94558
rect 82169 94555 82235 94558
rect 82353 94618 82419 94621
rect 82353 94616 84210 94618
rect 82353 94560 82358 94616
rect 82414 94560 84210 94616
rect 82353 94558 84210 94560
rect 82353 94555 82419 94558
rect 36924 94422 40970 94482
rect 36924 94420 36930 94422
rect 42558 94420 42564 94484
rect 42628 94482 42634 94484
rect 42701 94482 42767 94485
rect 42628 94480 42767 94482
rect 42628 94424 42706 94480
rect 42762 94424 42767 94480
rect 42628 94422 42767 94424
rect 42628 94420 42634 94422
rect 42701 94419 42767 94422
rect 44950 94420 44956 94484
rect 45020 94482 45026 94484
rect 45093 94482 45159 94485
rect 45020 94480 45159 94482
rect 45020 94424 45098 94480
rect 45154 94424 45159 94480
rect 45020 94422 45159 94424
rect 45020 94420 45026 94422
rect 45093 94419 45159 94422
rect 46238 94420 46244 94484
rect 46308 94482 46314 94484
rect 49877 94482 49943 94485
rect 46308 94480 49943 94482
rect 46308 94424 49882 94480
rect 49938 94424 49943 94480
rect 46308 94422 49943 94424
rect 46308 94420 46314 94422
rect 49877 94419 49943 94422
rect 50153 94482 50219 94485
rect 84009 94482 84075 94485
rect 84150 94484 84210 94558
rect 50153 94480 84075 94482
rect 50153 94424 50158 94480
rect 50214 94424 84014 94480
rect 84070 94424 84075 94480
rect 50153 94422 84075 94424
rect 50153 94419 50219 94422
rect 84009 94419 84075 94422
rect 84142 94420 84148 94484
rect 84212 94482 84218 94484
rect 84929 94482 84995 94485
rect 84212 94480 84995 94482
rect 84212 94424 84934 94480
rect 84990 94424 84995 94480
rect 84212 94422 84995 94424
rect 84212 94420 84218 94422
rect 84929 94419 84995 94422
rect 39982 94284 39988 94348
rect 40052 94346 40058 94348
rect 83590 94346 83596 94348
rect 40052 94286 83596 94346
rect 40052 94284 40058 94286
rect 83590 94284 83596 94286
rect 83660 94284 83666 94348
rect 86953 94346 87019 94349
rect 86953 94344 89730 94346
rect 86953 94288 86958 94344
rect 87014 94288 89730 94344
rect 86953 94286 89730 94288
rect 86953 94283 87019 94286
rect 39246 94148 39252 94212
rect 39316 94210 39322 94212
rect 50153 94210 50219 94213
rect 83406 94210 83412 94212
rect 39316 94208 50219 94210
rect 39316 94152 50158 94208
rect 50214 94152 50219 94208
rect 39316 94150 50219 94152
rect 39316 94148 39322 94150
rect 50153 94147 50219 94150
rect 50340 94150 83412 94210
rect 3944 94144 4264 94145
rect 3944 94080 3952 94144
rect 4016 94080 4032 94144
rect 4096 94080 4112 94144
rect 4176 94080 4192 94144
rect 4256 94080 4264 94144
rect 3944 94079 4264 94080
rect 41270 94012 41276 94076
rect 41340 94074 41346 94076
rect 50340 94074 50400 94150
rect 83406 94148 83412 94150
rect 83476 94148 83482 94212
rect 89670 94210 89730 94286
rect 91200 94210 92000 94240
rect 89670 94150 92000 94210
rect 87944 94144 88264 94145
rect 87944 94080 87952 94144
rect 88016 94080 88032 94144
rect 88096 94080 88112 94144
rect 88176 94080 88192 94144
rect 88256 94080 88264 94144
rect 91200 94120 92000 94150
rect 87944 94079 88264 94080
rect 41340 94014 50400 94074
rect 50981 94074 51047 94077
rect 79225 94074 79291 94077
rect 86534 94074 86540 94076
rect 50981 94072 79291 94074
rect 50981 94016 50986 94072
rect 51042 94016 79230 94072
rect 79286 94016 79291 94072
rect 50981 94014 79291 94016
rect 41340 94012 41346 94014
rect 50981 94011 51047 94014
rect 79225 94011 79291 94014
rect 79366 94014 86540 94074
rect 19190 93876 19196 93940
rect 19260 93938 19266 93940
rect 79366 93938 79426 94014
rect 86534 94012 86540 94014
rect 86604 94012 86610 94076
rect 19260 93878 79426 93938
rect 79501 93938 79567 93941
rect 86350 93938 86356 93940
rect 79501 93936 86356 93938
rect 79501 93880 79506 93936
rect 79562 93880 86356 93936
rect 79501 93878 86356 93880
rect 19260 93876 19266 93878
rect 79501 93875 79567 93878
rect 86350 93876 86356 93878
rect 86420 93876 86426 93940
rect 35750 93740 35756 93804
rect 35820 93802 35826 93804
rect 82486 93802 82492 93804
rect 35820 93742 82492 93802
rect 35820 93740 35826 93742
rect 82486 93740 82492 93742
rect 82556 93740 82562 93804
rect 82629 93802 82695 93805
rect 83406 93802 83412 93804
rect 82629 93800 83412 93802
rect 82629 93744 82634 93800
rect 82690 93744 83412 93800
rect 82629 93742 83412 93744
rect 82629 93739 82695 93742
rect 83406 93740 83412 93742
rect 83476 93802 83482 93804
rect 83476 93742 85130 93802
rect 83476 93740 83482 93742
rect 85070 93669 85130 93742
rect 31702 93604 31708 93668
rect 31772 93666 31778 93668
rect 40861 93666 40927 93669
rect 42609 93668 42675 93669
rect 44081 93668 44147 93669
rect 46657 93668 46723 93669
rect 47945 93668 48011 93669
rect 31772 93664 40927 93666
rect 31772 93608 40866 93664
rect 40922 93608 40927 93664
rect 31772 93606 40927 93608
rect 31772 93604 31778 93606
rect 40861 93603 40927 93606
rect 42558 93604 42564 93668
rect 42628 93666 42675 93668
rect 42628 93664 42720 93666
rect 42670 93608 42720 93664
rect 42628 93606 42720 93608
rect 42628 93604 42675 93606
rect 44030 93604 44036 93668
rect 44100 93666 44147 93668
rect 44100 93664 44192 93666
rect 44142 93608 44192 93664
rect 44100 93606 44192 93608
rect 44100 93604 44147 93606
rect 46606 93604 46612 93668
rect 46676 93666 46723 93668
rect 46676 93664 46768 93666
rect 46718 93608 46768 93664
rect 46676 93606 46768 93608
rect 46676 93604 46723 93606
rect 47894 93604 47900 93668
rect 47964 93666 48011 93668
rect 47964 93664 48056 93666
rect 48006 93608 48056 93664
rect 47964 93606 48056 93608
rect 47964 93604 48011 93606
rect 48262 93604 48268 93668
rect 48332 93666 48338 93668
rect 48773 93666 48839 93669
rect 49049 93668 49115 93669
rect 48998 93666 49004 93668
rect 48332 93664 48839 93666
rect 48332 93608 48778 93664
rect 48834 93608 48839 93664
rect 48332 93606 48839 93608
rect 48958 93606 49004 93666
rect 49068 93664 49115 93668
rect 49110 93608 49115 93664
rect 48332 93604 48338 93606
rect 42609 93603 42675 93604
rect 44081 93603 44147 93604
rect 46657 93603 46723 93604
rect 47945 93603 48011 93604
rect 48773 93603 48839 93606
rect 48998 93604 49004 93606
rect 49068 93604 49115 93608
rect 49182 93604 49188 93668
rect 49252 93666 49258 93668
rect 49601 93666 49667 93669
rect 49969 93668 50035 93669
rect 49918 93666 49924 93668
rect 49252 93664 49667 93666
rect 49252 93608 49606 93664
rect 49662 93608 49667 93664
rect 49252 93606 49667 93608
rect 49878 93606 49924 93666
rect 49988 93664 50035 93668
rect 50030 93608 50035 93664
rect 49252 93604 49258 93606
rect 49049 93603 49115 93604
rect 49601 93603 49667 93606
rect 49918 93604 49924 93606
rect 49988 93604 50035 93608
rect 50286 93604 50292 93668
rect 50356 93666 50362 93668
rect 50613 93666 50679 93669
rect 51257 93668 51323 93669
rect 51441 93668 51507 93669
rect 52177 93668 52243 93669
rect 52545 93668 52611 93669
rect 53281 93668 53347 93669
rect 51206 93666 51212 93668
rect 50356 93664 50679 93666
rect 50356 93608 50618 93664
rect 50674 93608 50679 93664
rect 50356 93606 50679 93608
rect 51166 93606 51212 93666
rect 51276 93664 51323 93668
rect 51318 93608 51323 93664
rect 50356 93604 50362 93606
rect 49969 93603 50035 93604
rect 50613 93603 50679 93606
rect 51206 93604 51212 93606
rect 51276 93604 51323 93608
rect 51390 93604 51396 93668
rect 51460 93666 51507 93668
rect 52126 93666 52132 93668
rect 51460 93664 51552 93666
rect 51502 93608 51552 93664
rect 51460 93606 51552 93608
rect 52086 93606 52132 93666
rect 52196 93664 52243 93668
rect 52238 93608 52243 93664
rect 51460 93604 51507 93606
rect 52126 93604 52132 93606
rect 52196 93604 52243 93608
rect 52494 93604 52500 93668
rect 52564 93666 52611 93668
rect 53230 93666 53236 93668
rect 52564 93664 52656 93666
rect 52606 93608 52656 93664
rect 52564 93606 52656 93608
rect 53190 93606 53236 93666
rect 53300 93664 53347 93668
rect 53741 93668 53807 93669
rect 54017 93668 54083 93669
rect 53741 93666 53788 93668
rect 53342 93608 53347 93664
rect 52564 93604 52611 93606
rect 53230 93604 53236 93606
rect 53300 93604 53347 93608
rect 53696 93664 53788 93666
rect 53696 93608 53746 93664
rect 53696 93606 53788 93608
rect 51257 93603 51323 93604
rect 51441 93603 51507 93604
rect 52177 93603 52243 93604
rect 52545 93603 52611 93604
rect 53281 93603 53347 93604
rect 53741 93604 53788 93606
rect 53852 93604 53858 93668
rect 53966 93604 53972 93668
rect 54036 93666 54083 93668
rect 54201 93666 54267 93669
rect 54569 93668 54635 93669
rect 54937 93668 55003 93669
rect 54334 93666 54340 93668
rect 54036 93664 54128 93666
rect 54078 93608 54128 93664
rect 54036 93606 54128 93608
rect 54201 93664 54340 93666
rect 54201 93608 54206 93664
rect 54262 93608 54340 93664
rect 54201 93606 54340 93608
rect 54036 93604 54083 93606
rect 53741 93603 53807 93604
rect 54017 93603 54083 93604
rect 54201 93603 54267 93606
rect 54334 93604 54340 93606
rect 54404 93604 54410 93668
rect 54518 93666 54524 93668
rect 54478 93606 54524 93666
rect 54588 93664 54635 93668
rect 54630 93608 54635 93664
rect 54518 93604 54524 93606
rect 54588 93604 54635 93608
rect 54886 93604 54892 93668
rect 54956 93666 55003 93668
rect 54956 93664 55048 93666
rect 54998 93608 55048 93664
rect 54956 93606 55048 93608
rect 54956 93604 55003 93606
rect 55254 93604 55260 93668
rect 55324 93666 55330 93668
rect 77017 93666 77083 93669
rect 55324 93664 77083 93666
rect 55324 93608 77022 93664
rect 77078 93608 77083 93664
rect 55324 93606 77083 93608
rect 55324 93604 55330 93606
rect 54569 93603 54635 93604
rect 54937 93603 55003 93604
rect 77017 93603 77083 93606
rect 77293 93666 77359 93669
rect 79041 93666 79107 93669
rect 85070 93668 85179 93669
rect 84326 93666 84332 93668
rect 77293 93664 79107 93666
rect 77293 93608 77298 93664
rect 77354 93608 79046 93664
rect 79102 93608 79107 93664
rect 77293 93606 79107 93608
rect 77293 93603 77359 93606
rect 79041 93603 79107 93606
rect 79228 93606 84332 93666
rect 1944 93600 2264 93601
rect 1944 93536 1952 93600
rect 2016 93536 2032 93600
rect 2096 93536 2112 93600
rect 2176 93536 2192 93600
rect 2256 93536 2264 93600
rect 1944 93535 2264 93536
rect 4429 93530 4495 93533
rect 79228 93530 79288 93606
rect 84326 93604 84332 93606
rect 84396 93604 84402 93668
rect 85062 93604 85068 93668
rect 85132 93666 85179 93668
rect 85132 93664 85224 93666
rect 85174 93608 85224 93664
rect 85132 93606 85224 93608
rect 85132 93604 85179 93606
rect 85113 93603 85179 93604
rect 85944 93600 86264 93601
rect 85944 93536 85952 93600
rect 86016 93536 86032 93600
rect 86096 93536 86112 93600
rect 86176 93536 86192 93600
rect 86256 93536 86264 93600
rect 85944 93535 86264 93536
rect 89944 93600 90264 93601
rect 89944 93536 89952 93600
rect 90016 93536 90032 93600
rect 90096 93536 90112 93600
rect 90176 93536 90192 93600
rect 90256 93536 90264 93600
rect 89944 93535 90264 93536
rect 85021 93530 85087 93533
rect 4429 93528 79288 93530
rect 4429 93472 4434 93528
rect 4490 93472 79288 93528
rect 4429 93470 79288 93472
rect 79366 93528 85087 93530
rect 79366 93472 85026 93528
rect 85082 93472 85087 93528
rect 79366 93470 85087 93472
rect 4429 93467 4495 93470
rect 30230 93332 30236 93396
rect 30300 93394 30306 93396
rect 40861 93394 40927 93397
rect 79366 93394 79426 93470
rect 85021 93467 85087 93470
rect 30300 93334 40786 93394
rect 30300 93332 30306 93334
rect 27470 93196 27476 93260
rect 27540 93258 27546 93260
rect 40585 93258 40651 93261
rect 27540 93256 40651 93258
rect 27540 93200 40590 93256
rect 40646 93200 40651 93256
rect 27540 93198 40651 93200
rect 40726 93258 40786 93334
rect 40861 93392 79426 93394
rect 40861 93336 40866 93392
rect 40922 93336 79426 93392
rect 40861 93334 79426 93336
rect 79501 93394 79567 93397
rect 83774 93394 83780 93396
rect 79501 93392 83780 93394
rect 79501 93336 79506 93392
rect 79562 93336 83780 93392
rect 79501 93334 83780 93336
rect 40861 93331 40927 93334
rect 79501 93331 79567 93334
rect 83774 93332 83780 93334
rect 83844 93332 83850 93396
rect 84561 93258 84627 93261
rect 40726 93256 84627 93258
rect 40726 93200 84566 93256
rect 84622 93200 84627 93256
rect 40726 93198 84627 93200
rect 27540 93196 27546 93198
rect 40585 93195 40651 93198
rect 84561 93195 84627 93198
rect 28942 93060 28948 93124
rect 29012 93122 29018 93124
rect 77477 93122 77543 93125
rect 29012 93120 77543 93122
rect 29012 93064 77482 93120
rect 77538 93064 77543 93120
rect 29012 93062 77543 93064
rect 29012 93060 29018 93062
rect 77477 93059 77543 93062
rect 77661 93122 77727 93125
rect 83590 93122 83596 93124
rect 77661 93120 83596 93122
rect 77661 93064 77666 93120
rect 77722 93064 83596 93120
rect 77661 93062 83596 93064
rect 77661 93059 77727 93062
rect 83590 93060 83596 93062
rect 83660 93060 83666 93124
rect 3944 93056 4264 93057
rect 3944 92992 3952 93056
rect 4016 92992 4032 93056
rect 4096 92992 4112 93056
rect 4176 92992 4192 93056
rect 4256 92992 4264 93056
rect 3944 92991 4264 92992
rect 87944 93056 88264 93057
rect 87944 92992 87952 93056
rect 88016 92992 88032 93056
rect 88096 92992 88112 93056
rect 88176 92992 88192 93056
rect 88256 92992 88264 93056
rect 87944 92991 88264 92992
rect 26182 92924 26188 92988
rect 26252 92986 26258 92988
rect 82721 92986 82787 92989
rect 91200 92986 92000 93016
rect 26252 92984 82787 92986
rect 26252 92928 82726 92984
rect 82782 92928 82787 92984
rect 26252 92926 82787 92928
rect 26252 92924 26258 92926
rect 82721 92923 82787 92926
rect 89670 92926 92000 92986
rect 32857 92852 32923 92853
rect 34145 92852 34211 92853
rect 35249 92852 35315 92853
rect 36721 92852 36787 92853
rect 38377 92852 38443 92853
rect 32806 92788 32812 92852
rect 32876 92850 32923 92852
rect 32876 92848 32968 92850
rect 32918 92792 32968 92848
rect 32876 92790 32968 92792
rect 32876 92788 32923 92790
rect 34094 92788 34100 92852
rect 34164 92850 34211 92852
rect 34164 92848 34256 92850
rect 34206 92792 34256 92848
rect 34164 92790 34256 92792
rect 34164 92788 34211 92790
rect 35198 92788 35204 92852
rect 35268 92850 35315 92852
rect 35268 92848 35360 92850
rect 35310 92792 35360 92848
rect 35268 92790 35360 92792
rect 35268 92788 35315 92790
rect 36670 92788 36676 92852
rect 36740 92850 36787 92852
rect 36740 92848 36832 92850
rect 36782 92792 36832 92848
rect 36740 92790 36832 92792
rect 36740 92788 36787 92790
rect 38326 92788 38332 92852
rect 38396 92850 38443 92852
rect 39941 92852 40007 92853
rect 39941 92850 39988 92852
rect 38396 92848 38488 92850
rect 38438 92792 38488 92848
rect 38396 92790 38488 92792
rect 39896 92848 39988 92850
rect 39896 92792 39946 92848
rect 39896 92790 39988 92792
rect 38396 92788 38443 92790
rect 32857 92787 32923 92788
rect 34145 92787 34211 92788
rect 35249 92787 35315 92788
rect 36721 92787 36787 92788
rect 38377 92787 38443 92788
rect 39941 92788 39988 92790
rect 40052 92788 40058 92852
rect 40585 92850 40651 92853
rect 77661 92850 77727 92853
rect 40585 92848 77727 92850
rect 40585 92792 40590 92848
rect 40646 92792 77666 92848
rect 77722 92792 77727 92848
rect 40585 92790 77727 92792
rect 39941 92787 40007 92788
rect 40585 92787 40651 92790
rect 77661 92787 77727 92790
rect 80094 92788 80100 92852
rect 80164 92850 80170 92852
rect 82077 92850 82143 92853
rect 80164 92848 82143 92850
rect 80164 92792 82082 92848
rect 82138 92792 82143 92848
rect 80164 92790 82143 92792
rect 80164 92788 80170 92790
rect 82077 92787 82143 92790
rect 87270 92788 87276 92852
rect 87340 92850 87346 92852
rect 89670 92850 89730 92926
rect 91200 92896 92000 92926
rect 87340 92790 89730 92850
rect 87340 92788 87346 92790
rect 1944 92512 2264 92513
rect 1944 92448 1952 92512
rect 2016 92448 2032 92512
rect 2096 92448 2112 92512
rect 2176 92448 2192 92512
rect 2256 92448 2264 92512
rect 1944 92447 2264 92448
rect 85944 92512 86264 92513
rect 85944 92448 85952 92512
rect 86016 92448 86032 92512
rect 86096 92448 86112 92512
rect 86176 92448 86192 92512
rect 86256 92448 86264 92512
rect 85944 92447 86264 92448
rect 89944 92512 90264 92513
rect 89944 92448 89952 92512
rect 90016 92448 90032 92512
rect 90096 92448 90112 92512
rect 90176 92448 90192 92512
rect 90256 92448 90264 92512
rect 89944 92447 90264 92448
rect 4705 92442 4771 92445
rect 4838 92442 4844 92444
rect 4705 92440 4844 92442
rect 4705 92384 4710 92440
rect 4766 92384 4844 92440
rect 4705 92382 4844 92384
rect 4705 92379 4771 92382
rect 4838 92380 4844 92382
rect 4908 92380 4914 92444
rect 83230 92034 83290 92044
rect 85573 92034 85639 92037
rect 83230 92032 85639 92034
rect 83230 91976 85578 92032
rect 85634 91976 85639 92032
rect 83230 91974 85639 91976
rect 85573 91971 85639 91974
rect 3944 91968 4264 91969
rect 3944 91904 3952 91968
rect 4016 91904 4032 91968
rect 4096 91904 4112 91968
rect 4176 91904 4192 91968
rect 4256 91904 4264 91968
rect 3944 91903 4264 91904
rect 87944 91968 88264 91969
rect 87944 91904 87952 91968
rect 88016 91904 88032 91968
rect 88096 91904 88112 91968
rect 88176 91904 88192 91968
rect 88256 91904 88264 91968
rect 87944 91903 88264 91904
rect 86902 91700 86908 91764
rect 86972 91762 86978 91764
rect 91200 91762 92000 91792
rect 86972 91702 92000 91762
rect 86972 91700 86978 91702
rect 91200 91672 92000 91702
rect 1944 91424 2264 91425
rect 1944 91360 1952 91424
rect 2016 91360 2032 91424
rect 2096 91360 2112 91424
rect 2176 91360 2192 91424
rect 2256 91360 2264 91424
rect 1944 91359 2264 91360
rect 85944 91424 86264 91425
rect 85944 91360 85952 91424
rect 86016 91360 86032 91424
rect 86096 91360 86112 91424
rect 86176 91360 86192 91424
rect 86256 91360 86264 91424
rect 85944 91359 86264 91360
rect 89944 91424 90264 91425
rect 89944 91360 89952 91424
rect 90016 91360 90032 91424
rect 90096 91360 90112 91424
rect 90176 91360 90192 91424
rect 90256 91360 90264 91424
rect 89944 91359 90264 91360
rect 4705 91082 4771 91085
rect 5073 91082 5139 91085
rect 4705 91080 5139 91082
rect 4705 91024 4710 91080
rect 4766 91024 5078 91080
rect 5134 91024 5139 91080
rect 4705 91022 5139 91024
rect 4705 91019 4771 91022
rect 5073 91019 5139 91022
rect 3944 90880 4264 90881
rect 3944 90816 3952 90880
rect 4016 90816 4032 90880
rect 4096 90816 4112 90880
rect 4176 90816 4192 90880
rect 4256 90816 4264 90880
rect 3944 90815 4264 90816
rect 87944 90880 88264 90881
rect 87944 90816 87952 90880
rect 88016 90816 88032 90880
rect 88096 90816 88112 90880
rect 88176 90816 88192 90880
rect 88256 90816 88264 90880
rect 87944 90815 88264 90816
rect 86902 90476 86908 90540
rect 86972 90538 86978 90540
rect 91200 90538 92000 90568
rect 86972 90478 92000 90538
rect 86972 90476 86978 90478
rect 91200 90448 92000 90478
rect 1944 90336 2264 90337
rect 1944 90272 1952 90336
rect 2016 90272 2032 90336
rect 2096 90272 2112 90336
rect 2176 90272 2192 90336
rect 2256 90272 2264 90336
rect 1944 90271 2264 90272
rect 85944 90336 86264 90337
rect 85944 90272 85952 90336
rect 86016 90272 86032 90336
rect 86096 90272 86112 90336
rect 86176 90272 86192 90336
rect 86256 90272 86264 90336
rect 85944 90271 86264 90272
rect 89944 90336 90264 90337
rect 89944 90272 89952 90336
rect 90016 90272 90032 90336
rect 90096 90272 90112 90336
rect 90176 90272 90192 90336
rect 90256 90272 90264 90336
rect 89944 90271 90264 90272
rect 87505 89858 87571 89861
rect 87278 89856 87571 89858
rect 87278 89800 87510 89856
rect 87566 89800 87571 89856
rect 87278 89798 87571 89800
rect 3944 89792 4264 89793
rect 3944 89728 3952 89792
rect 4016 89728 4032 89792
rect 4096 89728 4112 89792
rect 4176 89728 4192 89792
rect 4256 89728 4264 89792
rect 3944 89727 4264 89728
rect 86677 89586 86743 89589
rect 86861 89586 86927 89589
rect 86677 89584 86927 89586
rect 86677 89528 86682 89584
rect 86738 89528 86866 89584
rect 86922 89528 86927 89584
rect 86677 89526 86927 89528
rect 86677 89523 86743 89526
rect 86861 89523 86927 89526
rect 87045 89586 87111 89589
rect 87278 89586 87338 89798
rect 87505 89795 87571 89798
rect 87944 89792 88264 89793
rect 87944 89728 87952 89792
rect 88016 89728 88032 89792
rect 88096 89728 88112 89792
rect 88176 89728 88192 89792
rect 88256 89728 88264 89792
rect 87944 89727 88264 89728
rect 87045 89584 87338 89586
rect 87045 89528 87050 89584
rect 87106 89528 87338 89584
rect 87045 89526 87338 89528
rect 87045 89523 87111 89526
rect 5165 89452 5231 89453
rect 5165 89448 5212 89452
rect 5276 89450 5282 89452
rect 5165 89392 5170 89448
rect 5165 89388 5212 89392
rect 5276 89390 5322 89450
rect 5276 89388 5282 89390
rect 5165 89387 5231 89388
rect 4705 89314 4771 89317
rect 91200 89314 92000 89344
rect 4705 89312 4906 89314
rect 4705 89256 4710 89312
rect 4766 89256 4906 89312
rect 4705 89254 4906 89256
rect 4705 89251 4771 89254
rect 1944 89248 2264 89249
rect 1944 89184 1952 89248
rect 2016 89184 2032 89248
rect 2096 89184 2112 89248
rect 2176 89184 2192 89248
rect 2256 89184 2264 89248
rect 1944 89183 2264 89184
rect 4846 89178 4906 89254
rect 90406 89254 92000 89314
rect 85944 89248 86264 89249
rect 85944 89184 85952 89248
rect 86016 89184 86032 89248
rect 86096 89184 86112 89248
rect 86176 89184 86192 89248
rect 86256 89184 86264 89248
rect 85944 89183 86264 89184
rect 89944 89248 90264 89249
rect 89944 89184 89952 89248
rect 90016 89184 90032 89248
rect 90096 89184 90112 89248
rect 90176 89184 90192 89248
rect 90256 89184 90264 89248
rect 89944 89183 90264 89184
rect 5073 89178 5139 89181
rect 5574 89178 5580 89180
rect 4846 89176 5580 89178
rect 4846 89120 5078 89176
rect 5134 89120 5580 89176
rect 4846 89118 5580 89120
rect 5073 89115 5139 89118
rect 5574 89116 5580 89118
rect 5644 89116 5650 89180
rect 4797 89042 4863 89045
rect 4797 89040 5642 89042
rect 4797 88984 4802 89040
rect 4858 88984 5642 89040
rect 4797 88982 5642 88984
rect 4797 88979 4863 88982
rect 5582 88978 5642 88982
rect 86902 88980 86908 89044
rect 86972 89042 86978 89044
rect 90406 89042 90466 89254
rect 91200 89224 92000 89254
rect 86972 88982 90466 89042
rect 86972 88980 86978 88982
rect 5582 88918 6164 88978
rect 4797 88908 4863 88909
rect 4797 88904 4844 88908
rect 4908 88906 4914 88908
rect 4797 88848 4802 88904
rect 4797 88844 4844 88848
rect 4908 88846 4954 88906
rect 4908 88844 4914 88846
rect 4797 88843 4863 88844
rect 5257 88772 5323 88773
rect 5206 88708 5212 88772
rect 5276 88770 5323 88772
rect 5276 88768 5368 88770
rect 5318 88712 5368 88768
rect 5276 88710 5368 88712
rect 5276 88708 5323 88710
rect 5257 88707 5323 88708
rect 3944 88704 4264 88705
rect 3944 88640 3952 88704
rect 4016 88640 4032 88704
rect 4096 88640 4112 88704
rect 4176 88640 4192 88704
rect 4256 88640 4264 88704
rect 3944 88639 4264 88640
rect 87944 88704 88264 88705
rect 87944 88640 87952 88704
rect 88016 88640 88032 88704
rect 88096 88640 88112 88704
rect 88176 88640 88192 88704
rect 88256 88640 88264 88704
rect 87944 88639 88264 88640
rect 1944 88160 2264 88161
rect 1944 88096 1952 88160
rect 2016 88096 2032 88160
rect 2096 88096 2112 88160
rect 2176 88096 2192 88160
rect 2256 88096 2264 88160
rect 1944 88095 2264 88096
rect 85944 88160 86264 88161
rect 85944 88096 85952 88160
rect 86016 88096 86032 88160
rect 86096 88096 86112 88160
rect 86176 88096 86192 88160
rect 86256 88096 86264 88160
rect 85944 88095 86264 88096
rect 89944 88160 90264 88161
rect 89944 88096 89952 88160
rect 90016 88096 90032 88160
rect 90096 88096 90112 88160
rect 90176 88096 90192 88160
rect 90256 88096 90264 88160
rect 89944 88095 90264 88096
rect 91200 88090 92000 88120
rect 90406 88030 92000 88090
rect 87965 87954 88031 87957
rect 90406 87954 90466 88030
rect 91200 88000 92000 88030
rect 87965 87952 90466 87954
rect 87965 87896 87970 87952
rect 88026 87896 90466 87952
rect 87965 87894 90466 87896
rect 87965 87891 88031 87894
rect 4981 87818 5047 87821
rect 6134 87818 6194 87820
rect 4981 87816 6194 87818
rect 4981 87760 4986 87816
rect 5042 87760 6194 87816
rect 4981 87758 6194 87760
rect 4981 87755 5047 87758
rect 3944 87616 4264 87617
rect 3944 87552 3952 87616
rect 4016 87552 4032 87616
rect 4096 87552 4112 87616
rect 4176 87552 4192 87616
rect 4256 87552 4264 87616
rect 3944 87551 4264 87552
rect 87944 87616 88264 87617
rect 87944 87552 87952 87616
rect 88016 87552 88032 87616
rect 88096 87552 88112 87616
rect 88176 87552 88192 87616
rect 88256 87552 88264 87616
rect 87944 87551 88264 87552
rect 1944 87072 2264 87073
rect 1944 87008 1952 87072
rect 2016 87008 2032 87072
rect 2096 87008 2112 87072
rect 2176 87008 2192 87072
rect 2256 87008 2264 87072
rect 1944 87007 2264 87008
rect 85944 87072 86264 87073
rect 85944 87008 85952 87072
rect 86016 87008 86032 87072
rect 86096 87008 86112 87072
rect 86176 87008 86192 87072
rect 86256 87008 86264 87072
rect 85944 87007 86264 87008
rect 89944 87072 90264 87073
rect 89944 87008 89952 87072
rect 90016 87008 90032 87072
rect 90096 87008 90112 87072
rect 90176 87008 90192 87072
rect 90256 87008 90264 87072
rect 89944 87007 90264 87008
rect 86677 86866 86743 86869
rect 91200 86866 92000 86896
rect 86677 86864 92000 86866
rect 86677 86808 86682 86864
rect 86738 86808 92000 86864
rect 86677 86806 92000 86808
rect 86677 86803 86743 86806
rect 91200 86776 92000 86806
rect 4705 86730 4771 86733
rect 5390 86730 5396 86732
rect 4705 86728 5396 86730
rect 4705 86672 4710 86728
rect 4766 86672 5396 86728
rect 4705 86670 5396 86672
rect 4705 86667 4771 86670
rect 5390 86668 5396 86670
rect 5460 86668 5466 86732
rect 3944 86528 4264 86529
rect 3944 86464 3952 86528
rect 4016 86464 4032 86528
rect 4096 86464 4112 86528
rect 4176 86464 4192 86528
rect 4256 86464 4264 86528
rect 3944 86463 4264 86464
rect 87944 86528 88264 86529
rect 87944 86464 87952 86528
rect 88016 86464 88032 86528
rect 88096 86464 88112 86528
rect 88176 86464 88192 86528
rect 88256 86464 88264 86528
rect 87944 86463 88264 86464
rect 5165 86322 5231 86325
rect 5165 86320 6194 86322
rect 5165 86264 5170 86320
rect 5226 86264 6194 86320
rect 5165 86262 6194 86264
rect 5165 86259 5231 86262
rect 6134 86120 6194 86262
rect 1944 85984 2264 85985
rect 1944 85920 1952 85984
rect 2016 85920 2032 85984
rect 2096 85920 2112 85984
rect 2176 85920 2192 85984
rect 2256 85920 2264 85984
rect 1944 85919 2264 85920
rect 85944 85984 86264 85985
rect 85944 85920 85952 85984
rect 86016 85920 86032 85984
rect 86096 85920 86112 85984
rect 86176 85920 86192 85984
rect 86256 85920 86264 85984
rect 85944 85919 86264 85920
rect 89944 85984 90264 85985
rect 89944 85920 89952 85984
rect 90016 85920 90032 85984
rect 90096 85920 90112 85984
rect 90176 85920 90192 85984
rect 90256 85920 90264 85984
rect 89944 85919 90264 85920
rect 87965 85642 88031 85645
rect 91200 85642 92000 85672
rect 87965 85640 92000 85642
rect 87965 85584 87970 85640
rect 88026 85584 92000 85640
rect 87965 85582 92000 85584
rect 87965 85579 88031 85582
rect 91200 85552 92000 85582
rect 3944 85440 4264 85441
rect 3944 85376 3952 85440
rect 4016 85376 4032 85440
rect 4096 85376 4112 85440
rect 4176 85376 4192 85440
rect 4256 85376 4264 85440
rect 3944 85375 4264 85376
rect 87944 85440 88264 85441
rect 87944 85376 87952 85440
rect 88016 85376 88032 85440
rect 88096 85376 88112 85440
rect 88176 85376 88192 85440
rect 88256 85376 88264 85440
rect 87944 85375 88264 85376
rect 85021 85370 85087 85373
rect 85021 85368 85130 85370
rect 85021 85312 85026 85368
rect 85082 85312 85130 85368
rect 85021 85307 85130 85312
rect 4705 85234 4771 85237
rect 4705 85232 6194 85234
rect 4705 85176 4710 85232
rect 4766 85176 6194 85232
rect 4705 85174 6194 85176
rect 4705 85171 4771 85174
rect 6134 84992 6194 85174
rect 85070 84965 85130 85307
rect 87689 85234 87755 85237
rect 87278 85232 87755 85234
rect 87278 85176 87694 85232
rect 87750 85176 87755 85232
rect 87278 85174 87755 85176
rect 85389 85098 85455 85101
rect 85021 84960 85130 84965
rect 85021 84904 85026 84960
rect 85082 84904 85130 84960
rect 85021 84902 85130 84904
rect 85254 85096 85455 85098
rect 85254 85040 85394 85096
rect 85450 85040 85455 85096
rect 85254 85038 85455 85040
rect 85021 84899 85087 84902
rect 1944 84896 2264 84897
rect 1944 84832 1952 84896
rect 2016 84832 2032 84896
rect 2096 84832 2112 84896
rect 2176 84832 2192 84896
rect 2256 84832 2264 84896
rect 1944 84831 2264 84832
rect 85021 84690 85087 84693
rect 85254 84690 85314 85038
rect 85389 85035 85455 85038
rect 87045 85098 87111 85101
rect 87045 85096 87154 85098
rect 87045 85040 87050 85096
rect 87106 85040 87154 85096
rect 87045 85035 87154 85040
rect 85944 84896 86264 84897
rect 85944 84832 85952 84896
rect 86016 84832 86032 84896
rect 86096 84832 86112 84896
rect 86176 84832 86192 84896
rect 86256 84832 86264 84896
rect 85944 84831 86264 84832
rect 85021 84688 85314 84690
rect 85021 84632 85026 84688
rect 85082 84632 85314 84688
rect 85021 84630 85314 84632
rect 85021 84627 85087 84630
rect 87094 84554 87154 85035
rect 87278 84693 87338 85174
rect 87689 85171 87755 85174
rect 87413 85096 87479 85101
rect 87413 85040 87418 85096
rect 87474 85040 87479 85096
rect 87413 85035 87479 85040
rect 87416 84826 87476 85035
rect 89944 84896 90264 84897
rect 89944 84832 89952 84896
rect 90016 84832 90032 84896
rect 90096 84832 90112 84896
rect 90176 84832 90192 84896
rect 90256 84832 90264 84896
rect 89944 84831 90264 84832
rect 87781 84826 87847 84829
rect 87416 84824 87847 84826
rect 87416 84768 87786 84824
rect 87842 84768 87847 84824
rect 87416 84766 87847 84768
rect 87781 84763 87847 84766
rect 87229 84688 87338 84693
rect 87229 84632 87234 84688
rect 87290 84632 87338 84688
rect 87229 84630 87338 84632
rect 87229 84627 87295 84630
rect 87321 84554 87387 84557
rect 87094 84552 87387 84554
rect 87094 84496 87326 84552
rect 87382 84496 87387 84552
rect 87094 84494 87387 84496
rect 87321 84491 87387 84494
rect 87965 84554 88031 84557
rect 87965 84552 89730 84554
rect 87965 84496 87970 84552
rect 88026 84496 89730 84552
rect 87965 84494 89730 84496
rect 87965 84491 88031 84494
rect 89670 84418 89730 84494
rect 91200 84418 92000 84448
rect 89670 84358 92000 84418
rect 3944 84352 4264 84353
rect 3944 84288 3952 84352
rect 4016 84288 4032 84352
rect 4096 84288 4112 84352
rect 4176 84288 4192 84352
rect 4256 84288 4264 84352
rect 3944 84287 4264 84288
rect 87944 84352 88264 84353
rect 87944 84288 87952 84352
rect 88016 84288 88032 84352
rect 88096 84288 88112 84352
rect 88176 84288 88192 84352
rect 88256 84288 88264 84352
rect 91200 84328 92000 84358
rect 87944 84287 88264 84288
rect 1944 83808 2264 83809
rect 1944 83744 1952 83808
rect 2016 83744 2032 83808
rect 2096 83744 2112 83808
rect 2176 83744 2192 83808
rect 2256 83744 2264 83808
rect 1944 83743 2264 83744
rect 85944 83808 86264 83809
rect 85944 83744 85952 83808
rect 86016 83744 86032 83808
rect 86096 83744 86112 83808
rect 86176 83744 86192 83808
rect 86256 83744 86264 83808
rect 85944 83743 86264 83744
rect 89944 83808 90264 83809
rect 89944 83744 89952 83808
rect 90016 83744 90032 83808
rect 90096 83744 90112 83808
rect 90176 83744 90192 83808
rect 90256 83744 90264 83808
rect 89944 83743 90264 83744
rect 87965 83466 88031 83469
rect 87965 83464 89730 83466
rect 87965 83408 87970 83464
rect 88026 83408 89730 83464
rect 87965 83406 89730 83408
rect 87965 83403 88031 83406
rect 4797 83330 4863 83333
rect 4797 83328 6194 83330
rect 4797 83272 4802 83328
rect 4858 83272 6194 83328
rect 4797 83270 6194 83272
rect 4797 83267 4863 83270
rect 3944 83264 4264 83265
rect 3944 83200 3952 83264
rect 4016 83200 4032 83264
rect 4096 83200 4112 83264
rect 4176 83200 4192 83264
rect 4256 83200 4264 83264
rect 3944 83199 4264 83200
rect 87944 83264 88264 83265
rect 87944 83200 87952 83264
rect 88016 83200 88032 83264
rect 88096 83200 88112 83264
rect 88176 83200 88192 83264
rect 88256 83200 88264 83264
rect 87944 83199 88264 83200
rect 89670 83194 89730 83406
rect 91200 83194 92000 83224
rect 89670 83134 92000 83194
rect 91200 83104 92000 83134
rect 1944 82720 2264 82721
rect 1944 82656 1952 82720
rect 2016 82656 2032 82720
rect 2096 82656 2112 82720
rect 2176 82656 2192 82720
rect 2256 82656 2264 82720
rect 1944 82655 2264 82656
rect 85944 82720 86264 82721
rect 85944 82656 85952 82720
rect 86016 82656 86032 82720
rect 86096 82656 86112 82720
rect 86176 82656 86192 82720
rect 86256 82656 86264 82720
rect 85944 82655 86264 82656
rect 89944 82720 90264 82721
rect 89944 82656 89952 82720
rect 90016 82656 90032 82720
rect 90096 82656 90112 82720
rect 90176 82656 90192 82720
rect 90256 82656 90264 82720
rect 89944 82655 90264 82656
rect 4797 82242 4863 82245
rect 5165 82242 5231 82245
rect 4797 82240 6194 82242
rect 4797 82184 4802 82240
rect 4858 82184 5170 82240
rect 5226 82184 6194 82240
rect 4797 82182 6194 82184
rect 4797 82179 4863 82182
rect 5165 82179 5231 82182
rect 3944 82176 4264 82177
rect 3944 82112 3952 82176
rect 4016 82112 4032 82176
rect 4096 82112 4112 82176
rect 4176 82112 4192 82176
rect 4256 82112 4264 82176
rect 6134 82164 6194 82182
rect 87944 82176 88264 82177
rect 3944 82111 4264 82112
rect 87944 82112 87952 82176
rect 88016 82112 88032 82176
rect 88096 82112 88112 82176
rect 88176 82112 88192 82176
rect 88256 82112 88264 82176
rect 87944 82111 88264 82112
rect 87965 81970 88031 81973
rect 91200 81970 92000 82000
rect 87965 81968 92000 81970
rect 87965 81912 87970 81968
rect 88026 81912 92000 81968
rect 87965 81910 92000 81912
rect 87965 81907 88031 81910
rect 91200 81880 92000 81910
rect 1944 81632 2264 81633
rect 1944 81568 1952 81632
rect 2016 81568 2032 81632
rect 2096 81568 2112 81632
rect 2176 81568 2192 81632
rect 2256 81568 2264 81632
rect 1944 81567 2264 81568
rect 85944 81632 86264 81633
rect 85944 81568 85952 81632
rect 86016 81568 86032 81632
rect 86096 81568 86112 81632
rect 86176 81568 86192 81632
rect 86256 81568 86264 81632
rect 85944 81567 86264 81568
rect 89944 81632 90264 81633
rect 89944 81568 89952 81632
rect 90016 81568 90032 81632
rect 90096 81568 90112 81632
rect 90176 81568 90192 81632
rect 90256 81568 90264 81632
rect 89944 81567 90264 81568
rect 3944 81088 4264 81089
rect 3944 81024 3952 81088
rect 4016 81024 4032 81088
rect 4096 81024 4112 81088
rect 4176 81024 4192 81088
rect 4256 81024 4264 81088
rect 3944 81023 4264 81024
rect 87944 81088 88264 81089
rect 87944 81024 87952 81088
rect 88016 81024 88032 81088
rect 88096 81024 88112 81088
rect 88176 81024 88192 81088
rect 88256 81024 88264 81088
rect 87944 81023 88264 81024
rect 87965 80746 88031 80749
rect 91200 80746 92000 80776
rect 87965 80744 92000 80746
rect 87965 80688 87970 80744
rect 88026 80688 92000 80744
rect 87965 80686 92000 80688
rect 87965 80683 88031 80686
rect 91200 80656 92000 80686
rect 1944 80544 2264 80545
rect 1944 80480 1952 80544
rect 2016 80480 2032 80544
rect 2096 80480 2112 80544
rect 2176 80480 2192 80544
rect 2256 80480 2264 80544
rect 1944 80479 2264 80480
rect 85944 80544 86264 80545
rect 85944 80480 85952 80544
rect 86016 80480 86032 80544
rect 86096 80480 86112 80544
rect 86176 80480 86192 80544
rect 86256 80480 86264 80544
rect 85944 80479 86264 80480
rect 89944 80544 90264 80545
rect 89944 80480 89952 80544
rect 90016 80480 90032 80544
rect 90096 80480 90112 80544
rect 90176 80480 90192 80544
rect 90256 80480 90264 80544
rect 89944 80479 90264 80480
rect 4797 80474 4863 80477
rect 5257 80474 5323 80477
rect 4797 80472 6194 80474
rect 4797 80416 4802 80472
rect 4858 80416 5262 80472
rect 5318 80416 6194 80472
rect 4797 80414 6194 80416
rect 4797 80411 4863 80414
rect 5257 80411 5323 80414
rect 86861 80202 86927 80205
rect 86861 80200 87338 80202
rect 86861 80144 86866 80200
rect 86922 80144 87338 80200
rect 86861 80142 87338 80144
rect 86861 80139 86927 80142
rect 87278 80073 87338 80142
rect 86953 80066 87019 80069
rect 87278 80068 87387 80073
rect 86953 80064 87154 80066
rect 86953 80008 86958 80064
rect 87014 80008 87154 80064
rect 87278 80012 87326 80068
rect 87382 80012 87387 80068
rect 87278 80010 87387 80012
rect 86953 80006 87154 80008
rect 87321 80007 87387 80010
rect 86953 80003 87019 80006
rect 3944 80000 4264 80001
rect 3944 79936 3952 80000
rect 4016 79936 4032 80000
rect 4096 79936 4112 80000
rect 4176 79936 4192 80000
rect 4256 79936 4264 80000
rect 3944 79935 4264 79936
rect 87094 79930 87154 80006
rect 87944 80000 88264 80001
rect 87944 79936 87952 80000
rect 88016 79936 88032 80000
rect 88096 79936 88112 80000
rect 88176 79936 88192 80000
rect 88256 79936 88264 80000
rect 87944 79935 88264 79936
rect 87413 79930 87479 79933
rect 87094 79928 87479 79930
rect 87094 79872 87418 79928
rect 87474 79872 87479 79928
rect 87094 79870 87479 79872
rect 87413 79867 87479 79870
rect 88241 79658 88307 79661
rect 88241 79656 90466 79658
rect 88241 79600 88246 79656
rect 88302 79600 90466 79656
rect 88241 79598 90466 79600
rect 88241 79595 88307 79598
rect 90406 79522 90466 79598
rect 91200 79522 92000 79552
rect 90406 79462 92000 79522
rect 1944 79456 2264 79457
rect 1944 79392 1952 79456
rect 2016 79392 2032 79456
rect 2096 79392 2112 79456
rect 2176 79392 2192 79456
rect 2256 79392 2264 79456
rect 1944 79391 2264 79392
rect 85944 79456 86264 79457
rect 85944 79392 85952 79456
rect 86016 79392 86032 79456
rect 86096 79392 86112 79456
rect 86176 79392 86192 79456
rect 86256 79392 86264 79456
rect 85944 79391 86264 79392
rect 89944 79456 90264 79457
rect 89944 79392 89952 79456
rect 90016 79392 90032 79456
rect 90096 79392 90112 79456
rect 90176 79392 90192 79456
rect 90256 79392 90264 79456
rect 91200 79432 92000 79462
rect 89944 79391 90264 79392
rect 3944 78912 4264 78913
rect 3944 78848 3952 78912
rect 4016 78848 4032 78912
rect 4096 78848 4112 78912
rect 4176 78848 4192 78912
rect 4256 78848 4264 78912
rect 3944 78847 4264 78848
rect 87944 78912 88264 78913
rect 87944 78848 87952 78912
rect 88016 78848 88032 78912
rect 88096 78848 88112 78912
rect 88176 78848 88192 78912
rect 88256 78848 88264 78912
rect 87944 78847 88264 78848
rect 87045 78570 87111 78573
rect 87045 78568 90466 78570
rect 87045 78512 87050 78568
rect 87106 78512 90466 78568
rect 87045 78510 90466 78512
rect 87045 78507 87111 78510
rect 1944 78368 2264 78369
rect 1944 78304 1952 78368
rect 2016 78304 2032 78368
rect 2096 78304 2112 78368
rect 2176 78304 2192 78368
rect 2256 78304 2264 78368
rect 1944 78303 2264 78304
rect 85944 78368 86264 78369
rect 85944 78304 85952 78368
rect 86016 78304 86032 78368
rect 86096 78304 86112 78368
rect 86176 78304 86192 78368
rect 86256 78304 86264 78368
rect 85944 78303 86264 78304
rect 89944 78368 90264 78369
rect 89944 78304 89952 78368
rect 90016 78304 90032 78368
rect 90096 78304 90112 78368
rect 90176 78304 90192 78368
rect 90256 78304 90264 78368
rect 89944 78303 90264 78304
rect 90406 78298 90466 78510
rect 91200 78298 92000 78328
rect 90406 78238 92000 78298
rect 91200 78208 92000 78238
rect 3944 77824 4264 77825
rect 3944 77760 3952 77824
rect 4016 77760 4032 77824
rect 4096 77760 4112 77824
rect 4176 77760 4192 77824
rect 4256 77760 4264 77824
rect 3944 77759 4264 77760
rect 87944 77824 88264 77825
rect 87944 77760 87952 77824
rect 88016 77760 88032 77824
rect 88096 77760 88112 77824
rect 88176 77760 88192 77824
rect 88256 77760 88264 77824
rect 87944 77759 88264 77760
rect 1944 77280 2264 77281
rect 1944 77216 1952 77280
rect 2016 77216 2032 77280
rect 2096 77216 2112 77280
rect 2176 77216 2192 77280
rect 2256 77216 2264 77280
rect 1944 77215 2264 77216
rect 85944 77280 86264 77281
rect 85944 77216 85952 77280
rect 86016 77216 86032 77280
rect 86096 77216 86112 77280
rect 86176 77216 86192 77280
rect 86256 77216 86264 77280
rect 85944 77215 86264 77216
rect 89944 77280 90264 77281
rect 89944 77216 89952 77280
rect 90016 77216 90032 77280
rect 90096 77216 90112 77280
rect 90176 77216 90192 77280
rect 90256 77216 90264 77280
rect 89944 77215 90264 77216
rect 91200 77210 92000 77240
rect 90406 77150 92000 77210
rect 87137 77074 87203 77077
rect 90406 77074 90466 77150
rect 91200 77120 92000 77150
rect 87137 77072 90466 77074
rect 87137 77016 87142 77072
rect 87198 77016 90466 77072
rect 87137 77014 90466 77016
rect 87137 77011 87203 77014
rect 3944 76736 4264 76737
rect 3944 76672 3952 76736
rect 4016 76672 4032 76736
rect 4096 76672 4112 76736
rect 4176 76672 4192 76736
rect 4256 76672 4264 76736
rect 3944 76671 4264 76672
rect 87944 76736 88264 76737
rect 87944 76672 87952 76736
rect 88016 76672 88032 76736
rect 88096 76672 88112 76736
rect 88176 76672 88192 76736
rect 88256 76672 88264 76736
rect 87944 76671 88264 76672
rect 1944 76192 2264 76193
rect 1944 76128 1952 76192
rect 2016 76128 2032 76192
rect 2096 76128 2112 76192
rect 2176 76128 2192 76192
rect 2256 76128 2264 76192
rect 1944 76127 2264 76128
rect 85944 76192 86264 76193
rect 85944 76128 85952 76192
rect 86016 76128 86032 76192
rect 86096 76128 86112 76192
rect 86176 76128 86192 76192
rect 86256 76128 86264 76192
rect 85944 76127 86264 76128
rect 89944 76192 90264 76193
rect 89944 76128 89952 76192
rect 90016 76128 90032 76192
rect 90096 76128 90112 76192
rect 90176 76128 90192 76192
rect 90256 76128 90264 76192
rect 89944 76127 90264 76128
rect 87045 75986 87111 75989
rect 91200 75986 92000 76016
rect 87045 75984 92000 75986
rect 87045 75928 87050 75984
rect 87106 75928 92000 75984
rect 87045 75926 92000 75928
rect 87045 75923 87111 75926
rect 91200 75896 92000 75926
rect 3944 75648 4264 75649
rect 3944 75584 3952 75648
rect 4016 75584 4032 75648
rect 4096 75584 4112 75648
rect 4176 75584 4192 75648
rect 4256 75584 4264 75648
rect 3944 75583 4264 75584
rect 87944 75648 88264 75649
rect 87944 75584 87952 75648
rect 88016 75584 88032 75648
rect 88096 75584 88112 75648
rect 88176 75584 88192 75648
rect 88256 75584 88264 75648
rect 87944 75583 88264 75584
rect 1944 75104 2264 75105
rect 1944 75040 1952 75104
rect 2016 75040 2032 75104
rect 2096 75040 2112 75104
rect 2176 75040 2192 75104
rect 2256 75040 2264 75104
rect 1944 75039 2264 75040
rect 85944 75104 86264 75105
rect 85944 75040 85952 75104
rect 86016 75040 86032 75104
rect 86096 75040 86112 75104
rect 86176 75040 86192 75104
rect 86256 75040 86264 75104
rect 85944 75039 86264 75040
rect 89944 75104 90264 75105
rect 89944 75040 89952 75104
rect 90016 75040 90032 75104
rect 90096 75040 90112 75104
rect 90176 75040 90192 75104
rect 90256 75040 90264 75104
rect 89944 75039 90264 75040
rect 86953 74762 87019 74765
rect 91200 74762 92000 74792
rect 86953 74760 92000 74762
rect 86953 74704 86958 74760
rect 87014 74704 92000 74760
rect 86953 74702 92000 74704
rect 86953 74699 87019 74702
rect 91200 74672 92000 74702
rect 3944 74560 4264 74561
rect 3944 74496 3952 74560
rect 4016 74496 4032 74560
rect 4096 74496 4112 74560
rect 4176 74496 4192 74560
rect 4256 74496 4264 74560
rect 3944 74495 4264 74496
rect 87944 74560 88264 74561
rect 87944 74496 87952 74560
rect 88016 74496 88032 74560
rect 88096 74496 88112 74560
rect 88176 74496 88192 74560
rect 88256 74496 88264 74560
rect 87944 74495 88264 74496
rect 1944 74016 2264 74017
rect 1944 73952 1952 74016
rect 2016 73952 2032 74016
rect 2096 73952 2112 74016
rect 2176 73952 2192 74016
rect 2256 73952 2264 74016
rect 1944 73951 2264 73952
rect 85944 74016 86264 74017
rect 85944 73952 85952 74016
rect 86016 73952 86032 74016
rect 86096 73952 86112 74016
rect 86176 73952 86192 74016
rect 86256 73952 86264 74016
rect 85944 73951 86264 73952
rect 89944 74016 90264 74017
rect 89944 73952 89952 74016
rect 90016 73952 90032 74016
rect 90096 73952 90112 74016
rect 90176 73952 90192 74016
rect 90256 73952 90264 74016
rect 89944 73951 90264 73952
rect 86953 73674 87019 73677
rect 86953 73672 89730 73674
rect 86953 73616 86958 73672
rect 87014 73616 89730 73672
rect 86953 73614 89730 73616
rect 86953 73611 87019 73614
rect 89670 73538 89730 73614
rect 91200 73538 92000 73568
rect 89670 73478 92000 73538
rect 3944 73472 4264 73473
rect 3944 73408 3952 73472
rect 4016 73408 4032 73472
rect 4096 73408 4112 73472
rect 4176 73408 4192 73472
rect 4256 73408 4264 73472
rect 3944 73407 4264 73408
rect 87944 73472 88264 73473
rect 87944 73408 87952 73472
rect 88016 73408 88032 73472
rect 88096 73408 88112 73472
rect 88176 73408 88192 73472
rect 88256 73408 88264 73472
rect 91200 73448 92000 73478
rect 87944 73407 88264 73408
rect 1944 72928 2264 72929
rect 1944 72864 1952 72928
rect 2016 72864 2032 72928
rect 2096 72864 2112 72928
rect 2176 72864 2192 72928
rect 2256 72864 2264 72928
rect 1944 72863 2264 72864
rect 85944 72928 86264 72929
rect 85944 72864 85952 72928
rect 86016 72864 86032 72928
rect 86096 72864 86112 72928
rect 86176 72864 86192 72928
rect 86256 72864 86264 72928
rect 85944 72863 86264 72864
rect 89944 72928 90264 72929
rect 89944 72864 89952 72928
rect 90016 72864 90032 72928
rect 90096 72864 90112 72928
rect 90176 72864 90192 72928
rect 90256 72864 90264 72928
rect 89944 72863 90264 72864
rect 87229 72586 87295 72589
rect 87229 72584 89730 72586
rect 87229 72528 87234 72584
rect 87290 72528 89730 72584
rect 87229 72526 89730 72528
rect 87229 72523 87295 72526
rect 3944 72384 4264 72385
rect 3944 72320 3952 72384
rect 4016 72320 4032 72384
rect 4096 72320 4112 72384
rect 4176 72320 4192 72384
rect 4256 72320 4264 72384
rect 3944 72319 4264 72320
rect 87944 72384 88264 72385
rect 87944 72320 87952 72384
rect 88016 72320 88032 72384
rect 88096 72320 88112 72384
rect 88176 72320 88192 72384
rect 88256 72320 88264 72384
rect 87944 72319 88264 72320
rect 89670 72314 89730 72526
rect 91200 72314 92000 72344
rect 89670 72254 92000 72314
rect 91200 72224 92000 72254
rect 1944 71840 2264 71841
rect 1944 71776 1952 71840
rect 2016 71776 2032 71840
rect 2096 71776 2112 71840
rect 2176 71776 2192 71840
rect 2256 71776 2264 71840
rect 1944 71775 2264 71776
rect 85944 71840 86264 71841
rect 85944 71776 85952 71840
rect 86016 71776 86032 71840
rect 86096 71776 86112 71840
rect 86176 71776 86192 71840
rect 86256 71776 86264 71840
rect 85944 71775 86264 71776
rect 89944 71840 90264 71841
rect 89944 71776 89952 71840
rect 90016 71776 90032 71840
rect 90096 71776 90112 71840
rect 90176 71776 90192 71840
rect 90256 71776 90264 71840
rect 89944 71775 90264 71776
rect 3944 71296 4264 71297
rect 3944 71232 3952 71296
rect 4016 71232 4032 71296
rect 4096 71232 4112 71296
rect 4176 71232 4192 71296
rect 4256 71232 4264 71296
rect 3944 71231 4264 71232
rect 87944 71296 88264 71297
rect 87944 71232 87952 71296
rect 88016 71232 88032 71296
rect 88096 71232 88112 71296
rect 88176 71232 88192 71296
rect 88256 71232 88264 71296
rect 87944 71231 88264 71232
rect 87137 71090 87203 71093
rect 91200 71090 92000 71120
rect 87137 71088 92000 71090
rect 87137 71032 87142 71088
rect 87198 71032 92000 71088
rect 87137 71030 92000 71032
rect 87137 71027 87203 71030
rect 91200 71000 92000 71030
rect 1944 70752 2264 70753
rect 1944 70688 1952 70752
rect 2016 70688 2032 70752
rect 2096 70688 2112 70752
rect 2176 70688 2192 70752
rect 2256 70688 2264 70752
rect 1944 70687 2264 70688
rect 85944 70752 86264 70753
rect 85944 70688 85952 70752
rect 86016 70688 86032 70752
rect 86096 70688 86112 70752
rect 86176 70688 86192 70752
rect 86256 70688 86264 70752
rect 85944 70687 86264 70688
rect 89944 70752 90264 70753
rect 89944 70688 89952 70752
rect 90016 70688 90032 70752
rect 90096 70688 90112 70752
rect 90176 70688 90192 70752
rect 90256 70688 90264 70752
rect 89944 70687 90264 70688
rect 3944 70208 4264 70209
rect 3944 70144 3952 70208
rect 4016 70144 4032 70208
rect 4096 70144 4112 70208
rect 4176 70144 4192 70208
rect 4256 70144 4264 70208
rect 3944 70143 4264 70144
rect 87944 70208 88264 70209
rect 87944 70144 87952 70208
rect 88016 70144 88032 70208
rect 88096 70144 88112 70208
rect 88176 70144 88192 70208
rect 88256 70144 88264 70208
rect 87944 70143 88264 70144
rect 87781 69866 87847 69869
rect 91200 69866 92000 69896
rect 87781 69864 92000 69866
rect 87781 69808 87786 69864
rect 87842 69808 92000 69864
rect 87781 69806 92000 69808
rect 87781 69803 87847 69806
rect 91200 69776 92000 69806
rect 1944 69664 2264 69665
rect 1944 69600 1952 69664
rect 2016 69600 2032 69664
rect 2096 69600 2112 69664
rect 2176 69600 2192 69664
rect 2256 69600 2264 69664
rect 1944 69599 2264 69600
rect 85944 69664 86264 69665
rect 85944 69600 85952 69664
rect 86016 69600 86032 69664
rect 86096 69600 86112 69664
rect 86176 69600 86192 69664
rect 86256 69600 86264 69664
rect 85944 69599 86264 69600
rect 89944 69664 90264 69665
rect 89944 69600 89952 69664
rect 90016 69600 90032 69664
rect 90096 69600 90112 69664
rect 90176 69600 90192 69664
rect 90256 69600 90264 69664
rect 89944 69599 90264 69600
rect 3944 69120 4264 69121
rect 3944 69056 3952 69120
rect 4016 69056 4032 69120
rect 4096 69056 4112 69120
rect 4176 69056 4192 69120
rect 4256 69056 4264 69120
rect 3944 69055 4264 69056
rect 87944 69120 88264 69121
rect 87944 69056 87952 69120
rect 88016 69056 88032 69120
rect 88096 69056 88112 69120
rect 88176 69056 88192 69120
rect 88256 69056 88264 69120
rect 87944 69055 88264 69056
rect 87137 68778 87203 68781
rect 87137 68776 90466 68778
rect 87137 68720 87142 68776
rect 87198 68720 90466 68776
rect 87137 68718 90466 68720
rect 87137 68715 87203 68718
rect 90406 68642 90466 68718
rect 91200 68642 92000 68672
rect 90406 68582 92000 68642
rect 1944 68576 2264 68577
rect 1944 68512 1952 68576
rect 2016 68512 2032 68576
rect 2096 68512 2112 68576
rect 2176 68512 2192 68576
rect 2256 68512 2264 68576
rect 1944 68511 2264 68512
rect 85944 68576 86264 68577
rect 85944 68512 85952 68576
rect 86016 68512 86032 68576
rect 86096 68512 86112 68576
rect 86176 68512 86192 68576
rect 86256 68512 86264 68576
rect 85944 68511 86264 68512
rect 89944 68576 90264 68577
rect 89944 68512 89952 68576
rect 90016 68512 90032 68576
rect 90096 68512 90112 68576
rect 90176 68512 90192 68576
rect 90256 68512 90264 68576
rect 91200 68552 92000 68582
rect 89944 68511 90264 68512
rect 3944 68032 4264 68033
rect 3944 67968 3952 68032
rect 4016 67968 4032 68032
rect 4096 67968 4112 68032
rect 4176 67968 4192 68032
rect 4256 67968 4264 68032
rect 3944 67967 4264 67968
rect 87944 68032 88264 68033
rect 87944 67968 87952 68032
rect 88016 67968 88032 68032
rect 88096 67968 88112 68032
rect 88176 67968 88192 68032
rect 88256 67968 88264 68032
rect 87944 67967 88264 67968
rect 1944 67488 2264 67489
rect 1944 67424 1952 67488
rect 2016 67424 2032 67488
rect 2096 67424 2112 67488
rect 2176 67424 2192 67488
rect 2256 67424 2264 67488
rect 1944 67423 2264 67424
rect 85944 67488 86264 67489
rect 85944 67424 85952 67488
rect 86016 67424 86032 67488
rect 86096 67424 86112 67488
rect 86176 67424 86192 67488
rect 86256 67424 86264 67488
rect 85944 67423 86264 67424
rect 89944 67488 90264 67489
rect 89944 67424 89952 67488
rect 90016 67424 90032 67488
rect 90096 67424 90112 67488
rect 90176 67424 90192 67488
rect 90256 67424 90264 67488
rect 89944 67423 90264 67424
rect 91200 67418 92000 67448
rect 90406 67358 92000 67418
rect 87321 67282 87387 67285
rect 90406 67282 90466 67358
rect 91200 67328 92000 67358
rect 87321 67280 90466 67282
rect 87321 67224 87326 67280
rect 87382 67224 90466 67280
rect 87321 67222 90466 67224
rect 87321 67219 87387 67222
rect 3944 66944 4264 66945
rect 3944 66880 3952 66944
rect 4016 66880 4032 66944
rect 4096 66880 4112 66944
rect 4176 66880 4192 66944
rect 4256 66880 4264 66944
rect 3944 66879 4264 66880
rect 87944 66944 88264 66945
rect 87944 66880 87952 66944
rect 88016 66880 88032 66944
rect 88096 66880 88112 66944
rect 88176 66880 88192 66944
rect 88256 66880 88264 66944
rect 87944 66879 88264 66880
rect 1944 66400 2264 66401
rect 1944 66336 1952 66400
rect 2016 66336 2032 66400
rect 2096 66336 2112 66400
rect 2176 66336 2192 66400
rect 2256 66336 2264 66400
rect 1944 66335 2264 66336
rect 85944 66400 86264 66401
rect 85944 66336 85952 66400
rect 86016 66336 86032 66400
rect 86096 66336 86112 66400
rect 86176 66336 86192 66400
rect 86256 66336 86264 66400
rect 85944 66335 86264 66336
rect 89944 66400 90264 66401
rect 89944 66336 89952 66400
rect 90016 66336 90032 66400
rect 90096 66336 90112 66400
rect 90176 66336 90192 66400
rect 90256 66336 90264 66400
rect 89944 66335 90264 66336
rect 87781 66194 87847 66197
rect 91200 66194 92000 66224
rect 87781 66192 92000 66194
rect 87781 66136 87786 66192
rect 87842 66136 92000 66192
rect 87781 66134 92000 66136
rect 87781 66131 87847 66134
rect 91200 66104 92000 66134
rect 3944 65856 4264 65857
rect 3944 65792 3952 65856
rect 4016 65792 4032 65856
rect 4096 65792 4112 65856
rect 4176 65792 4192 65856
rect 4256 65792 4264 65856
rect 3944 65791 4264 65792
rect 87944 65856 88264 65857
rect 87944 65792 87952 65856
rect 88016 65792 88032 65856
rect 88096 65792 88112 65856
rect 88176 65792 88192 65856
rect 88256 65792 88264 65856
rect 87944 65791 88264 65792
rect 1944 65312 2264 65313
rect 1944 65248 1952 65312
rect 2016 65248 2032 65312
rect 2096 65248 2112 65312
rect 2176 65248 2192 65312
rect 2256 65248 2264 65312
rect 1944 65247 2264 65248
rect 85944 65312 86264 65313
rect 85944 65248 85952 65312
rect 86016 65248 86032 65312
rect 86096 65248 86112 65312
rect 86176 65248 86192 65312
rect 86256 65248 86264 65312
rect 85944 65247 86264 65248
rect 89944 65312 90264 65313
rect 89944 65248 89952 65312
rect 90016 65248 90032 65312
rect 90096 65248 90112 65312
rect 90176 65248 90192 65312
rect 90256 65248 90264 65312
rect 89944 65247 90264 65248
rect 87321 64970 87387 64973
rect 91200 64970 92000 65000
rect 87321 64968 92000 64970
rect 87321 64912 87326 64968
rect 87382 64912 92000 64968
rect 87321 64910 92000 64912
rect 87321 64907 87387 64910
rect 91200 64880 92000 64910
rect 3944 64768 4264 64769
rect 3944 64704 3952 64768
rect 4016 64704 4032 64768
rect 4096 64704 4112 64768
rect 4176 64704 4192 64768
rect 4256 64704 4264 64768
rect 3944 64703 4264 64704
rect 87944 64768 88264 64769
rect 87944 64704 87952 64768
rect 88016 64704 88032 64768
rect 88096 64704 88112 64768
rect 88176 64704 88192 64768
rect 88256 64704 88264 64768
rect 87944 64703 88264 64704
rect 1944 64224 2264 64225
rect 1944 64160 1952 64224
rect 2016 64160 2032 64224
rect 2096 64160 2112 64224
rect 2176 64160 2192 64224
rect 2256 64160 2264 64224
rect 1944 64159 2264 64160
rect 85944 64224 86264 64225
rect 85944 64160 85952 64224
rect 86016 64160 86032 64224
rect 86096 64160 86112 64224
rect 86176 64160 86192 64224
rect 86256 64160 86264 64224
rect 85944 64159 86264 64160
rect 89944 64224 90264 64225
rect 89944 64160 89952 64224
rect 90016 64160 90032 64224
rect 90096 64160 90112 64224
rect 90176 64160 90192 64224
rect 90256 64160 90264 64224
rect 89944 64159 90264 64160
rect 87505 63882 87571 63885
rect 87505 63880 88442 63882
rect 87505 63824 87510 63880
rect 87566 63824 88442 63880
rect 87505 63822 88442 63824
rect 87505 63819 87571 63822
rect 88382 63746 88442 63822
rect 91200 63746 92000 63776
rect 88382 63686 92000 63746
rect 3944 63680 4264 63681
rect 3944 63616 3952 63680
rect 4016 63616 4032 63680
rect 4096 63616 4112 63680
rect 4176 63616 4192 63680
rect 4256 63616 4264 63680
rect 3944 63615 4264 63616
rect 87944 63680 88264 63681
rect 87944 63616 87952 63680
rect 88016 63616 88032 63680
rect 88096 63616 88112 63680
rect 88176 63616 88192 63680
rect 88256 63616 88264 63680
rect 91200 63656 92000 63686
rect 87944 63615 88264 63616
rect 1944 63136 2264 63137
rect 1944 63072 1952 63136
rect 2016 63072 2032 63136
rect 2096 63072 2112 63136
rect 2176 63072 2192 63136
rect 2256 63072 2264 63136
rect 1944 63071 2264 63072
rect 85944 63136 86264 63137
rect 85944 63072 85952 63136
rect 86016 63072 86032 63136
rect 86096 63072 86112 63136
rect 86176 63072 86192 63136
rect 86256 63072 86264 63136
rect 85944 63071 86264 63072
rect 89944 63136 90264 63137
rect 89944 63072 89952 63136
rect 90016 63072 90032 63136
rect 90096 63072 90112 63136
rect 90176 63072 90192 63136
rect 90256 63072 90264 63136
rect 89944 63071 90264 63072
rect 87781 62794 87847 62797
rect 87781 62792 88442 62794
rect 87781 62736 87786 62792
rect 87842 62736 88442 62792
rect 87781 62734 88442 62736
rect 87781 62731 87847 62734
rect 3944 62592 4264 62593
rect 3944 62528 3952 62592
rect 4016 62528 4032 62592
rect 4096 62528 4112 62592
rect 4176 62528 4192 62592
rect 4256 62528 4264 62592
rect 3944 62527 4264 62528
rect 87944 62592 88264 62593
rect 87944 62528 87952 62592
rect 88016 62528 88032 62592
rect 88096 62528 88112 62592
rect 88176 62528 88192 62592
rect 88256 62528 88264 62592
rect 87944 62527 88264 62528
rect 88382 62522 88442 62734
rect 91200 62522 92000 62552
rect 88382 62462 92000 62522
rect 91200 62432 92000 62462
rect 1944 62048 2264 62049
rect 1944 61984 1952 62048
rect 2016 61984 2032 62048
rect 2096 61984 2112 62048
rect 2176 61984 2192 62048
rect 2256 61984 2264 62048
rect 1944 61983 2264 61984
rect 85944 62048 86264 62049
rect 85944 61984 85952 62048
rect 86016 61984 86032 62048
rect 86096 61984 86112 62048
rect 86176 61984 86192 62048
rect 86256 61984 86264 62048
rect 85944 61983 86264 61984
rect 89944 62048 90264 62049
rect 89944 61984 89952 62048
rect 90016 61984 90032 62048
rect 90096 61984 90112 62048
rect 90176 61984 90192 62048
rect 90256 61984 90264 62048
rect 89944 61983 90264 61984
rect 3944 61504 4264 61505
rect 3944 61440 3952 61504
rect 4016 61440 4032 61504
rect 4096 61440 4112 61504
rect 4176 61440 4192 61504
rect 4256 61440 4264 61504
rect 3944 61439 4264 61440
rect 87944 61504 88264 61505
rect 87944 61440 87952 61504
rect 88016 61440 88032 61504
rect 88096 61440 88112 61504
rect 88176 61440 88192 61504
rect 88256 61440 88264 61504
rect 87944 61439 88264 61440
rect 87781 61298 87847 61301
rect 91200 61298 92000 61328
rect 87781 61296 92000 61298
rect 87781 61240 87786 61296
rect 87842 61240 92000 61296
rect 87781 61238 92000 61240
rect 87781 61235 87847 61238
rect 91200 61208 92000 61238
rect 1944 60960 2264 60961
rect 1944 60896 1952 60960
rect 2016 60896 2032 60960
rect 2096 60896 2112 60960
rect 2176 60896 2192 60960
rect 2256 60896 2264 60960
rect 1944 60895 2264 60896
rect 85944 60960 86264 60961
rect 85944 60896 85952 60960
rect 86016 60896 86032 60960
rect 86096 60896 86112 60960
rect 86176 60896 86192 60960
rect 86256 60896 86264 60960
rect 85944 60895 86264 60896
rect 89944 60960 90264 60961
rect 89944 60896 89952 60960
rect 90016 60896 90032 60960
rect 90096 60896 90112 60960
rect 90176 60896 90192 60960
rect 90256 60896 90264 60960
rect 89944 60895 90264 60896
rect 3944 60416 4264 60417
rect 3944 60352 3952 60416
rect 4016 60352 4032 60416
rect 4096 60352 4112 60416
rect 4176 60352 4192 60416
rect 4256 60352 4264 60416
rect 3944 60351 4264 60352
rect 87944 60416 88264 60417
rect 87944 60352 87952 60416
rect 88016 60352 88032 60416
rect 88096 60352 88112 60416
rect 88176 60352 88192 60416
rect 88256 60352 88264 60416
rect 87944 60351 88264 60352
rect 87689 60074 87755 60077
rect 91200 60074 92000 60104
rect 87689 60072 92000 60074
rect 87689 60016 87694 60072
rect 87750 60016 92000 60072
rect 87689 60014 92000 60016
rect 87689 60011 87755 60014
rect 91200 59984 92000 60014
rect 1944 59872 2264 59873
rect 1944 59808 1952 59872
rect 2016 59808 2032 59872
rect 2096 59808 2112 59872
rect 2176 59808 2192 59872
rect 2256 59808 2264 59872
rect 1944 59807 2264 59808
rect 85944 59872 86264 59873
rect 85944 59808 85952 59872
rect 86016 59808 86032 59872
rect 86096 59808 86112 59872
rect 86176 59808 86192 59872
rect 86256 59808 86264 59872
rect 85944 59807 86264 59808
rect 89944 59872 90264 59873
rect 89944 59808 89952 59872
rect 90016 59808 90032 59872
rect 90096 59808 90112 59872
rect 90176 59808 90192 59872
rect 90256 59808 90264 59872
rect 89944 59807 90264 59808
rect 3944 59328 4264 59329
rect 3944 59264 3952 59328
rect 4016 59264 4032 59328
rect 4096 59264 4112 59328
rect 4176 59264 4192 59328
rect 4256 59264 4264 59328
rect 3944 59263 4264 59264
rect 87944 59328 88264 59329
rect 87944 59264 87952 59328
rect 88016 59264 88032 59328
rect 88096 59264 88112 59328
rect 88176 59264 88192 59328
rect 88256 59264 88264 59328
rect 87944 59263 88264 59264
rect 87413 58986 87479 58989
rect 87413 58984 90466 58986
rect 87413 58928 87418 58984
rect 87474 58928 90466 58984
rect 87413 58926 90466 58928
rect 87413 58923 87479 58926
rect 90406 58850 90466 58926
rect 91200 58850 92000 58880
rect 90406 58790 92000 58850
rect 1944 58784 2264 58785
rect 1944 58720 1952 58784
rect 2016 58720 2032 58784
rect 2096 58720 2112 58784
rect 2176 58720 2192 58784
rect 2256 58720 2264 58784
rect 1944 58719 2264 58720
rect 85944 58784 86264 58785
rect 85944 58720 85952 58784
rect 86016 58720 86032 58784
rect 86096 58720 86112 58784
rect 86176 58720 86192 58784
rect 86256 58720 86264 58784
rect 85944 58719 86264 58720
rect 89944 58784 90264 58785
rect 89944 58720 89952 58784
rect 90016 58720 90032 58784
rect 90096 58720 90112 58784
rect 90176 58720 90192 58784
rect 90256 58720 90264 58784
rect 91200 58760 92000 58790
rect 89944 58719 90264 58720
rect 3944 58240 4264 58241
rect 3944 58176 3952 58240
rect 4016 58176 4032 58240
rect 4096 58176 4112 58240
rect 4176 58176 4192 58240
rect 4256 58176 4264 58240
rect 3944 58175 4264 58176
rect 87944 58240 88264 58241
rect 87944 58176 87952 58240
rect 88016 58176 88032 58240
rect 88096 58176 88112 58240
rect 88176 58176 88192 58240
rect 88256 58176 88264 58240
rect 87944 58175 88264 58176
rect 86953 57898 87019 57901
rect 86953 57896 90466 57898
rect 86953 57840 86958 57896
rect 87014 57840 90466 57896
rect 86953 57838 90466 57840
rect 86953 57835 87019 57838
rect 90406 57762 90466 57838
rect 91200 57762 92000 57792
rect 90406 57702 92000 57762
rect 1944 57696 2264 57697
rect 1944 57632 1952 57696
rect 2016 57632 2032 57696
rect 2096 57632 2112 57696
rect 2176 57632 2192 57696
rect 2256 57632 2264 57696
rect 1944 57631 2264 57632
rect 85944 57696 86264 57697
rect 85944 57632 85952 57696
rect 86016 57632 86032 57696
rect 86096 57632 86112 57696
rect 86176 57632 86192 57696
rect 86256 57632 86264 57696
rect 85944 57631 86264 57632
rect 89944 57696 90264 57697
rect 89944 57632 89952 57696
rect 90016 57632 90032 57696
rect 90096 57632 90112 57696
rect 90176 57632 90192 57696
rect 90256 57632 90264 57696
rect 91200 57672 92000 57702
rect 89944 57631 90264 57632
rect 3944 57152 4264 57153
rect 3944 57088 3952 57152
rect 4016 57088 4032 57152
rect 4096 57088 4112 57152
rect 4176 57088 4192 57152
rect 4256 57088 4264 57152
rect 3944 57087 4264 57088
rect 87944 57152 88264 57153
rect 87944 57088 87952 57152
rect 88016 57088 88032 57152
rect 88096 57088 88112 57152
rect 88176 57088 88192 57152
rect 88256 57088 88264 57152
rect 87944 57087 88264 57088
rect 1944 56608 2264 56609
rect 1944 56544 1952 56608
rect 2016 56544 2032 56608
rect 2096 56544 2112 56608
rect 2176 56544 2192 56608
rect 2256 56544 2264 56608
rect 1944 56543 2264 56544
rect 85944 56608 86264 56609
rect 85944 56544 85952 56608
rect 86016 56544 86032 56608
rect 86096 56544 86112 56608
rect 86176 56544 86192 56608
rect 86256 56544 86264 56608
rect 85944 56543 86264 56544
rect 89944 56608 90264 56609
rect 89944 56544 89952 56608
rect 90016 56544 90032 56608
rect 90096 56544 90112 56608
rect 90176 56544 90192 56608
rect 90256 56544 90264 56608
rect 89944 56543 90264 56544
rect 91200 56538 92000 56568
rect 90406 56478 92000 56538
rect 87045 56402 87111 56405
rect 90406 56402 90466 56478
rect 91200 56448 92000 56478
rect 87045 56400 90466 56402
rect 87045 56344 87050 56400
rect 87106 56344 90466 56400
rect 87045 56342 90466 56344
rect 87045 56339 87111 56342
rect 3944 56064 4264 56065
rect 3944 56000 3952 56064
rect 4016 56000 4032 56064
rect 4096 56000 4112 56064
rect 4176 56000 4192 56064
rect 4256 56000 4264 56064
rect 3944 55999 4264 56000
rect 87944 56064 88264 56065
rect 87944 56000 87952 56064
rect 88016 56000 88032 56064
rect 88096 56000 88112 56064
rect 88176 56000 88192 56064
rect 88256 56000 88264 56064
rect 87944 55999 88264 56000
rect 1944 55520 2264 55521
rect 1944 55456 1952 55520
rect 2016 55456 2032 55520
rect 2096 55456 2112 55520
rect 2176 55456 2192 55520
rect 2256 55456 2264 55520
rect 1944 55455 2264 55456
rect 85944 55520 86264 55521
rect 85944 55456 85952 55520
rect 86016 55456 86032 55520
rect 86096 55456 86112 55520
rect 86176 55456 86192 55520
rect 86256 55456 86264 55520
rect 85944 55455 86264 55456
rect 89944 55520 90264 55521
rect 89944 55456 89952 55520
rect 90016 55456 90032 55520
rect 90096 55456 90112 55520
rect 90176 55456 90192 55520
rect 90256 55456 90264 55520
rect 89944 55455 90264 55456
rect 82445 55314 82511 55317
rect 84142 55314 84148 55316
rect 82445 55312 84148 55314
rect 82445 55256 82450 55312
rect 82506 55256 84148 55312
rect 82445 55254 84148 55256
rect 82445 55251 82511 55254
rect 84142 55252 84148 55254
rect 84212 55252 84218 55316
rect 86953 55314 87019 55317
rect 91200 55314 92000 55344
rect 86953 55312 92000 55314
rect 86953 55256 86958 55312
rect 87014 55256 92000 55312
rect 86953 55254 92000 55256
rect 86953 55251 87019 55254
rect 91200 55224 92000 55254
rect 3944 54976 4264 54977
rect 3944 54912 3952 54976
rect 4016 54912 4032 54976
rect 4096 54912 4112 54976
rect 4176 54912 4192 54976
rect 4256 54912 4264 54976
rect 3944 54911 4264 54912
rect 87944 54976 88264 54977
rect 87944 54912 87952 54976
rect 88016 54912 88032 54976
rect 88096 54912 88112 54976
rect 88176 54912 88192 54976
rect 88256 54912 88264 54976
rect 87944 54911 88264 54912
rect 1944 54432 2264 54433
rect 1944 54368 1952 54432
rect 2016 54368 2032 54432
rect 2096 54368 2112 54432
rect 2176 54368 2192 54432
rect 2256 54368 2264 54432
rect 1944 54367 2264 54368
rect 85944 54432 86264 54433
rect 85944 54368 85952 54432
rect 86016 54368 86032 54432
rect 86096 54368 86112 54432
rect 86176 54368 86192 54432
rect 86256 54368 86264 54432
rect 85944 54367 86264 54368
rect 89944 54432 90264 54433
rect 89944 54368 89952 54432
rect 90016 54368 90032 54432
rect 90096 54368 90112 54432
rect 90176 54368 90192 54432
rect 90256 54368 90264 54432
rect 89944 54367 90264 54368
rect 86953 54090 87019 54093
rect 91200 54090 92000 54120
rect 86953 54088 92000 54090
rect 86953 54032 86958 54088
rect 87014 54032 92000 54088
rect 86953 54030 92000 54032
rect 86953 54027 87019 54030
rect 91200 54000 92000 54030
rect 3944 53888 4264 53889
rect 3944 53824 3952 53888
rect 4016 53824 4032 53888
rect 4096 53824 4112 53888
rect 4176 53824 4192 53888
rect 4256 53824 4264 53888
rect 3944 53823 4264 53824
rect 87944 53888 88264 53889
rect 87944 53824 87952 53888
rect 88016 53824 88032 53888
rect 88096 53824 88112 53888
rect 88176 53824 88192 53888
rect 88256 53824 88264 53888
rect 87944 53823 88264 53824
rect 1944 53344 2264 53345
rect 1944 53280 1952 53344
rect 2016 53280 2032 53344
rect 2096 53280 2112 53344
rect 2176 53280 2192 53344
rect 2256 53280 2264 53344
rect 1944 53279 2264 53280
rect 85944 53344 86264 53345
rect 85944 53280 85952 53344
rect 86016 53280 86032 53344
rect 86096 53280 86112 53344
rect 86176 53280 86192 53344
rect 86256 53280 86264 53344
rect 85944 53279 86264 53280
rect 89944 53344 90264 53345
rect 89944 53280 89952 53344
rect 90016 53280 90032 53344
rect 90096 53280 90112 53344
rect 90176 53280 90192 53344
rect 90256 53280 90264 53344
rect 89944 53279 90264 53280
rect 86953 53002 87019 53005
rect 86953 53000 88442 53002
rect 86953 52944 86958 53000
rect 87014 52944 88442 53000
rect 86953 52942 88442 52944
rect 86953 52939 87019 52942
rect 88382 52866 88442 52942
rect 91200 52866 92000 52896
rect 88382 52806 92000 52866
rect 3944 52800 4264 52801
rect 3944 52736 3952 52800
rect 4016 52736 4032 52800
rect 4096 52736 4112 52800
rect 4176 52736 4192 52800
rect 4256 52736 4264 52800
rect 3944 52735 4264 52736
rect 87944 52800 88264 52801
rect 87944 52736 87952 52800
rect 88016 52736 88032 52800
rect 88096 52736 88112 52800
rect 88176 52736 88192 52800
rect 88256 52736 88264 52800
rect 91200 52776 92000 52806
rect 87944 52735 88264 52736
rect 1944 52256 2264 52257
rect 1944 52192 1952 52256
rect 2016 52192 2032 52256
rect 2096 52192 2112 52256
rect 2176 52192 2192 52256
rect 2256 52192 2264 52256
rect 1944 52191 2264 52192
rect 85944 52256 86264 52257
rect 85944 52192 85952 52256
rect 86016 52192 86032 52256
rect 86096 52192 86112 52256
rect 86176 52192 86192 52256
rect 86256 52192 86264 52256
rect 85944 52191 86264 52192
rect 89944 52256 90264 52257
rect 89944 52192 89952 52256
rect 90016 52192 90032 52256
rect 90096 52192 90112 52256
rect 90176 52192 90192 52256
rect 90256 52192 90264 52256
rect 89944 52191 90264 52192
rect 3944 51712 4264 51713
rect 3944 51648 3952 51712
rect 4016 51648 4032 51712
rect 4096 51648 4112 51712
rect 4176 51648 4192 51712
rect 4256 51648 4264 51712
rect 3944 51647 4264 51648
rect 87944 51712 88264 51713
rect 87944 51648 87952 51712
rect 88016 51648 88032 51712
rect 88096 51648 88112 51712
rect 88176 51648 88192 51712
rect 88256 51648 88264 51712
rect 87944 51647 88264 51648
rect 91200 51642 92000 51672
rect 88382 51582 92000 51642
rect 83774 51308 83780 51372
rect 83844 51370 83850 51372
rect 88382 51370 88442 51582
rect 91200 51552 92000 51582
rect 83844 51310 88442 51370
rect 83844 51308 83850 51310
rect 1944 51168 2264 51169
rect 1944 51104 1952 51168
rect 2016 51104 2032 51168
rect 2096 51104 2112 51168
rect 2176 51104 2192 51168
rect 2256 51104 2264 51168
rect 1944 51103 2264 51104
rect 85944 51168 86264 51169
rect 85944 51104 85952 51168
rect 86016 51104 86032 51168
rect 86096 51104 86112 51168
rect 86176 51104 86192 51168
rect 86256 51104 86264 51168
rect 85944 51103 86264 51104
rect 89944 51168 90264 51169
rect 89944 51104 89952 51168
rect 90016 51104 90032 51168
rect 90096 51104 90112 51168
rect 90176 51104 90192 51168
rect 90256 51104 90264 51168
rect 89944 51103 90264 51104
rect 3944 50624 4264 50625
rect 3944 50560 3952 50624
rect 4016 50560 4032 50624
rect 4096 50560 4112 50624
rect 4176 50560 4192 50624
rect 4256 50560 4264 50624
rect 3944 50559 4264 50560
rect 87944 50624 88264 50625
rect 87944 50560 87952 50624
rect 88016 50560 88032 50624
rect 88096 50560 88112 50624
rect 88176 50560 88192 50624
rect 88256 50560 88264 50624
rect 87944 50559 88264 50560
rect 91200 50418 92000 50448
rect 84150 50358 92000 50418
rect 1944 50080 2264 50081
rect 1944 50016 1952 50080
rect 2016 50016 2032 50080
rect 2096 50016 2112 50080
rect 2176 50016 2192 50080
rect 2256 50016 2264 50080
rect 1944 50015 2264 50016
rect 83590 49676 83596 49740
rect 83660 49738 83666 49740
rect 84150 49738 84210 50358
rect 91200 50328 92000 50358
rect 85944 50080 86264 50081
rect 85944 50016 85952 50080
rect 86016 50016 86032 50080
rect 86096 50016 86112 50080
rect 86176 50016 86192 50080
rect 86256 50016 86264 50080
rect 85944 50015 86264 50016
rect 89944 50080 90264 50081
rect 89944 50016 89952 50080
rect 90016 50016 90032 50080
rect 90096 50016 90112 50080
rect 90176 50016 90192 50080
rect 90256 50016 90264 50080
rect 89944 50015 90264 50016
rect 83660 49678 84210 49738
rect 83660 49676 83666 49678
rect 3944 49536 4264 49537
rect 3944 49472 3952 49536
rect 4016 49472 4032 49536
rect 4096 49472 4112 49536
rect 4176 49472 4192 49536
rect 4256 49472 4264 49536
rect 3944 49471 4264 49472
rect 87944 49536 88264 49537
rect 87944 49472 87952 49536
rect 88016 49472 88032 49536
rect 88096 49472 88112 49536
rect 88176 49472 88192 49536
rect 88256 49472 88264 49536
rect 87944 49471 88264 49472
rect 87689 49194 87755 49197
rect 91200 49194 92000 49224
rect 87689 49192 92000 49194
rect 87689 49136 87694 49192
rect 87750 49136 92000 49192
rect 87689 49134 92000 49136
rect 87689 49131 87755 49134
rect 91200 49104 92000 49134
rect 1944 48992 2264 48993
rect 1944 48928 1952 48992
rect 2016 48928 2032 48992
rect 2096 48928 2112 48992
rect 2176 48928 2192 48992
rect 2256 48928 2264 48992
rect 1944 48927 2264 48928
rect 85944 48992 86264 48993
rect 85944 48928 85952 48992
rect 86016 48928 86032 48992
rect 86096 48928 86112 48992
rect 86176 48928 86192 48992
rect 86256 48928 86264 48992
rect 85944 48927 86264 48928
rect 89944 48992 90264 48993
rect 89944 48928 89952 48992
rect 90016 48928 90032 48992
rect 90096 48928 90112 48992
rect 90176 48928 90192 48992
rect 90256 48928 90264 48992
rect 89944 48927 90264 48928
rect 3944 48448 4264 48449
rect 3944 48384 3952 48448
rect 4016 48384 4032 48448
rect 4096 48384 4112 48448
rect 4176 48384 4192 48448
rect 4256 48384 4264 48448
rect 3944 48383 4264 48384
rect 87944 48448 88264 48449
rect 87944 48384 87952 48448
rect 88016 48384 88032 48448
rect 88096 48384 88112 48448
rect 88176 48384 88192 48448
rect 88256 48384 88264 48448
rect 87944 48383 88264 48384
rect 87597 48106 87663 48109
rect 87597 48104 90466 48106
rect 87597 48048 87602 48104
rect 87658 48048 90466 48104
rect 87597 48046 90466 48048
rect 87597 48043 87663 48046
rect 90406 47970 90466 48046
rect 91200 47970 92000 48000
rect 90406 47910 92000 47970
rect 1944 47904 2264 47905
rect 1944 47840 1952 47904
rect 2016 47840 2032 47904
rect 2096 47840 2112 47904
rect 2176 47840 2192 47904
rect 2256 47840 2264 47904
rect 1944 47839 2264 47840
rect 85944 47904 86264 47905
rect 85944 47840 85952 47904
rect 86016 47840 86032 47904
rect 86096 47840 86112 47904
rect 86176 47840 86192 47904
rect 86256 47840 86264 47904
rect 85944 47839 86264 47840
rect 89944 47904 90264 47905
rect 89944 47840 89952 47904
rect 90016 47840 90032 47904
rect 90096 47840 90112 47904
rect 90176 47840 90192 47904
rect 90256 47840 90264 47904
rect 91200 47880 92000 47910
rect 89944 47839 90264 47840
rect 3944 47360 4264 47361
rect 3944 47296 3952 47360
rect 4016 47296 4032 47360
rect 4096 47296 4112 47360
rect 4176 47296 4192 47360
rect 4256 47296 4264 47360
rect 3944 47295 4264 47296
rect 87944 47360 88264 47361
rect 87944 47296 87952 47360
rect 88016 47296 88032 47360
rect 88096 47296 88112 47360
rect 88176 47296 88192 47360
rect 88256 47296 88264 47360
rect 87944 47295 88264 47296
rect 1944 46816 2264 46817
rect 1944 46752 1952 46816
rect 2016 46752 2032 46816
rect 2096 46752 2112 46816
rect 2176 46752 2192 46816
rect 2256 46752 2264 46816
rect 1944 46751 2264 46752
rect 85944 46816 86264 46817
rect 85944 46752 85952 46816
rect 86016 46752 86032 46816
rect 86096 46752 86112 46816
rect 86176 46752 86192 46816
rect 86256 46752 86264 46816
rect 85944 46751 86264 46752
rect 89944 46816 90264 46817
rect 89944 46752 89952 46816
rect 90016 46752 90032 46816
rect 90096 46752 90112 46816
rect 90176 46752 90192 46816
rect 90256 46752 90264 46816
rect 89944 46751 90264 46752
rect 91200 46746 92000 46776
rect 90406 46686 92000 46746
rect 87689 46610 87755 46613
rect 90406 46610 90466 46686
rect 91200 46656 92000 46686
rect 87689 46608 90466 46610
rect 87689 46552 87694 46608
rect 87750 46552 90466 46608
rect 87689 46550 90466 46552
rect 87689 46547 87755 46550
rect 3944 46272 4264 46273
rect 3944 46208 3952 46272
rect 4016 46208 4032 46272
rect 4096 46208 4112 46272
rect 4176 46208 4192 46272
rect 4256 46208 4264 46272
rect 3944 46207 4264 46208
rect 87944 46272 88264 46273
rect 87944 46208 87952 46272
rect 88016 46208 88032 46272
rect 88096 46208 88112 46272
rect 88176 46208 88192 46272
rect 88256 46208 88264 46272
rect 87944 46207 88264 46208
rect 1944 45728 2264 45729
rect 1944 45664 1952 45728
rect 2016 45664 2032 45728
rect 2096 45664 2112 45728
rect 2176 45664 2192 45728
rect 2256 45664 2264 45728
rect 1944 45663 2264 45664
rect 85944 45728 86264 45729
rect 85944 45664 85952 45728
rect 86016 45664 86032 45728
rect 86096 45664 86112 45728
rect 86176 45664 86192 45728
rect 86256 45664 86264 45728
rect 85944 45663 86264 45664
rect 89944 45728 90264 45729
rect 89944 45664 89952 45728
rect 90016 45664 90032 45728
rect 90096 45664 90112 45728
rect 90176 45664 90192 45728
rect 90256 45664 90264 45728
rect 89944 45663 90264 45664
rect 82445 45522 82511 45525
rect 83406 45522 83412 45524
rect 82445 45520 83412 45522
rect 82445 45464 82450 45520
rect 82506 45464 83412 45520
rect 82445 45462 83412 45464
rect 82445 45459 82511 45462
rect 83406 45460 83412 45462
rect 83476 45460 83482 45524
rect 87597 45522 87663 45525
rect 91200 45522 92000 45552
rect 87597 45520 92000 45522
rect 87597 45464 87602 45520
rect 87658 45464 92000 45520
rect 87597 45462 92000 45464
rect 87597 45459 87663 45462
rect 91200 45432 92000 45462
rect 3944 45184 4264 45185
rect 3944 45120 3952 45184
rect 4016 45120 4032 45184
rect 4096 45120 4112 45184
rect 4176 45120 4192 45184
rect 4256 45120 4264 45184
rect 3944 45119 4264 45120
rect 87944 45184 88264 45185
rect 87944 45120 87952 45184
rect 88016 45120 88032 45184
rect 88096 45120 88112 45184
rect 88176 45120 88192 45184
rect 88256 45120 88264 45184
rect 87944 45119 88264 45120
rect 1944 44640 2264 44641
rect 1944 44576 1952 44640
rect 2016 44576 2032 44640
rect 2096 44576 2112 44640
rect 2176 44576 2192 44640
rect 2256 44576 2264 44640
rect 1944 44575 2264 44576
rect 85944 44640 86264 44641
rect 85944 44576 85952 44640
rect 86016 44576 86032 44640
rect 86096 44576 86112 44640
rect 86176 44576 86192 44640
rect 86256 44576 86264 44640
rect 85944 44575 86264 44576
rect 89944 44640 90264 44641
rect 89944 44576 89952 44640
rect 90016 44576 90032 44640
rect 90096 44576 90112 44640
rect 90176 44576 90192 44640
rect 90256 44576 90264 44640
rect 89944 44575 90264 44576
rect 87689 44298 87755 44301
rect 91200 44298 92000 44328
rect 87689 44296 92000 44298
rect 87689 44240 87694 44296
rect 87750 44240 92000 44296
rect 87689 44238 92000 44240
rect 87689 44235 87755 44238
rect 91200 44208 92000 44238
rect 3944 44096 4264 44097
rect 3944 44032 3952 44096
rect 4016 44032 4032 44096
rect 4096 44032 4112 44096
rect 4176 44032 4192 44096
rect 4256 44032 4264 44096
rect 3944 44031 4264 44032
rect 87944 44096 88264 44097
rect 87944 44032 87952 44096
rect 88016 44032 88032 44096
rect 88096 44032 88112 44096
rect 88176 44032 88192 44096
rect 88256 44032 88264 44096
rect 87944 44031 88264 44032
rect 1944 43552 2264 43553
rect 1944 43488 1952 43552
rect 2016 43488 2032 43552
rect 2096 43488 2112 43552
rect 2176 43488 2192 43552
rect 2256 43488 2264 43552
rect 1944 43487 2264 43488
rect 85944 43552 86264 43553
rect 85944 43488 85952 43552
rect 86016 43488 86032 43552
rect 86096 43488 86112 43552
rect 86176 43488 86192 43552
rect 86256 43488 86264 43552
rect 85944 43487 86264 43488
rect 89944 43552 90264 43553
rect 89944 43488 89952 43552
rect 90016 43488 90032 43552
rect 90096 43488 90112 43552
rect 90176 43488 90192 43552
rect 90256 43488 90264 43552
rect 89944 43487 90264 43488
rect 87689 43210 87755 43213
rect 87689 43208 88442 43210
rect 87689 43152 87694 43208
rect 87750 43152 88442 43208
rect 87689 43150 88442 43152
rect 87689 43147 87755 43150
rect 88382 43074 88442 43150
rect 91200 43074 92000 43104
rect 88382 43014 92000 43074
rect 3944 43008 4264 43009
rect 3944 42944 3952 43008
rect 4016 42944 4032 43008
rect 4096 42944 4112 43008
rect 4176 42944 4192 43008
rect 4256 42944 4264 43008
rect 3944 42943 4264 42944
rect 87944 43008 88264 43009
rect 87944 42944 87952 43008
rect 88016 42944 88032 43008
rect 88096 42944 88112 43008
rect 88176 42944 88192 43008
rect 88256 42944 88264 43008
rect 91200 42984 92000 43014
rect 87944 42943 88264 42944
rect 1944 42464 2264 42465
rect 1944 42400 1952 42464
rect 2016 42400 2032 42464
rect 2096 42400 2112 42464
rect 2176 42400 2192 42464
rect 2256 42400 2264 42464
rect 1944 42399 2264 42400
rect 85944 42464 86264 42465
rect 85944 42400 85952 42464
rect 86016 42400 86032 42464
rect 86096 42400 86112 42464
rect 86176 42400 86192 42464
rect 86256 42400 86264 42464
rect 85944 42399 86264 42400
rect 89944 42464 90264 42465
rect 89944 42400 89952 42464
rect 90016 42400 90032 42464
rect 90096 42400 90112 42464
rect 90176 42400 90192 42464
rect 90256 42400 90264 42464
rect 89944 42399 90264 42400
rect 3944 41920 4264 41921
rect 3944 41856 3952 41920
rect 4016 41856 4032 41920
rect 4096 41856 4112 41920
rect 4176 41856 4192 41920
rect 4256 41856 4264 41920
rect 3944 41855 4264 41856
rect 87944 41920 88264 41921
rect 87944 41856 87952 41920
rect 88016 41856 88032 41920
rect 88096 41856 88112 41920
rect 88176 41856 88192 41920
rect 88256 41856 88264 41920
rect 87944 41855 88264 41856
rect 91200 41850 92000 41880
rect 88382 41790 92000 41850
rect 87781 41714 87847 41717
rect 88382 41714 88442 41790
rect 91200 41760 92000 41790
rect 87781 41712 88442 41714
rect 87781 41656 87786 41712
rect 87842 41656 88442 41712
rect 87781 41654 88442 41656
rect 87781 41651 87847 41654
rect 1944 41376 2264 41377
rect 1944 41312 1952 41376
rect 2016 41312 2032 41376
rect 2096 41312 2112 41376
rect 2176 41312 2192 41376
rect 2256 41312 2264 41376
rect 1944 41311 2264 41312
rect 85944 41376 86264 41377
rect 85944 41312 85952 41376
rect 86016 41312 86032 41376
rect 86096 41312 86112 41376
rect 86176 41312 86192 41376
rect 86256 41312 86264 41376
rect 85944 41311 86264 41312
rect 89944 41376 90264 41377
rect 89944 41312 89952 41376
rect 90016 41312 90032 41376
rect 90096 41312 90112 41376
rect 90176 41312 90192 41376
rect 90256 41312 90264 41376
rect 89944 41311 90264 41312
rect 3944 40832 4264 40833
rect 3944 40768 3952 40832
rect 4016 40768 4032 40832
rect 4096 40768 4112 40832
rect 4176 40768 4192 40832
rect 4256 40768 4264 40832
rect 3944 40767 4264 40768
rect 87944 40832 88264 40833
rect 87944 40768 87952 40832
rect 88016 40768 88032 40832
rect 88096 40768 88112 40832
rect 88176 40768 88192 40832
rect 88256 40768 88264 40832
rect 87944 40767 88264 40768
rect 87873 40626 87939 40629
rect 91200 40626 92000 40656
rect 87873 40624 92000 40626
rect 87873 40568 87878 40624
rect 87934 40568 92000 40624
rect 87873 40566 92000 40568
rect 87873 40563 87939 40566
rect 91200 40536 92000 40566
rect 1944 40288 2264 40289
rect 1944 40224 1952 40288
rect 2016 40224 2032 40288
rect 2096 40224 2112 40288
rect 2176 40224 2192 40288
rect 2256 40224 2264 40288
rect 1944 40223 2264 40224
rect 85944 40288 86264 40289
rect 85944 40224 85952 40288
rect 86016 40224 86032 40288
rect 86096 40224 86112 40288
rect 86176 40224 86192 40288
rect 86256 40224 86264 40288
rect 85944 40223 86264 40224
rect 89944 40288 90264 40289
rect 89944 40224 89952 40288
rect 90016 40224 90032 40288
rect 90096 40224 90112 40288
rect 90176 40224 90192 40288
rect 90256 40224 90264 40288
rect 89944 40223 90264 40224
rect 3944 39744 4264 39745
rect 3944 39680 3952 39744
rect 4016 39680 4032 39744
rect 4096 39680 4112 39744
rect 4176 39680 4192 39744
rect 4256 39680 4264 39744
rect 3944 39679 4264 39680
rect 87944 39744 88264 39745
rect 87944 39680 87952 39744
rect 88016 39680 88032 39744
rect 88096 39680 88112 39744
rect 88176 39680 88192 39744
rect 88256 39680 88264 39744
rect 87944 39679 88264 39680
rect 87505 39402 87571 39405
rect 91200 39402 92000 39432
rect 87505 39400 92000 39402
rect 87505 39344 87510 39400
rect 87566 39344 92000 39400
rect 87505 39342 92000 39344
rect 87505 39339 87571 39342
rect 91200 39312 92000 39342
rect 1944 39200 2264 39201
rect 1944 39136 1952 39200
rect 2016 39136 2032 39200
rect 2096 39136 2112 39200
rect 2176 39136 2192 39200
rect 2256 39136 2264 39200
rect 1944 39135 2264 39136
rect 85944 39200 86264 39201
rect 85944 39136 85952 39200
rect 86016 39136 86032 39200
rect 86096 39136 86112 39200
rect 86176 39136 86192 39200
rect 86256 39136 86264 39200
rect 85944 39135 86264 39136
rect 89944 39200 90264 39201
rect 89944 39136 89952 39200
rect 90016 39136 90032 39200
rect 90096 39136 90112 39200
rect 90176 39136 90192 39200
rect 90256 39136 90264 39200
rect 89944 39135 90264 39136
rect 3944 38656 4264 38657
rect 3944 38592 3952 38656
rect 4016 38592 4032 38656
rect 4096 38592 4112 38656
rect 4176 38592 4192 38656
rect 4256 38592 4264 38656
rect 3944 38591 4264 38592
rect 87944 38656 88264 38657
rect 87944 38592 87952 38656
rect 88016 38592 88032 38656
rect 88096 38592 88112 38656
rect 88176 38592 88192 38656
rect 88256 38592 88264 38656
rect 87944 38591 88264 38592
rect 86677 38314 86743 38317
rect 91200 38314 92000 38344
rect 86677 38312 92000 38314
rect 86677 38256 86682 38312
rect 86738 38256 92000 38312
rect 86677 38254 92000 38256
rect 86677 38251 86743 38254
rect 91200 38224 92000 38254
rect 1944 38112 2264 38113
rect 1944 38048 1952 38112
rect 2016 38048 2032 38112
rect 2096 38048 2112 38112
rect 2176 38048 2192 38112
rect 2256 38048 2264 38112
rect 1944 38047 2264 38048
rect 85944 38112 86264 38113
rect 85944 38048 85952 38112
rect 86016 38048 86032 38112
rect 86096 38048 86112 38112
rect 86176 38048 86192 38112
rect 86256 38048 86264 38112
rect 85944 38047 86264 38048
rect 89944 38112 90264 38113
rect 89944 38048 89952 38112
rect 90016 38048 90032 38112
rect 90096 38048 90112 38112
rect 90176 38048 90192 38112
rect 90256 38048 90264 38112
rect 89944 38047 90264 38048
rect 3944 37568 4264 37569
rect 3944 37504 3952 37568
rect 4016 37504 4032 37568
rect 4096 37504 4112 37568
rect 4176 37504 4192 37568
rect 4256 37504 4264 37568
rect 3944 37503 4264 37504
rect 87944 37568 88264 37569
rect 87944 37504 87952 37568
rect 88016 37504 88032 37568
rect 88096 37504 88112 37568
rect 88176 37504 88192 37568
rect 88256 37504 88264 37568
rect 87944 37503 88264 37504
rect 91200 37090 92000 37120
rect 90406 37030 92000 37090
rect 1944 37024 2264 37025
rect 1944 36960 1952 37024
rect 2016 36960 2032 37024
rect 2096 36960 2112 37024
rect 2176 36960 2192 37024
rect 2256 36960 2264 37024
rect 1944 36959 2264 36960
rect 85944 37024 86264 37025
rect 85944 36960 85952 37024
rect 86016 36960 86032 37024
rect 86096 36960 86112 37024
rect 86176 36960 86192 37024
rect 86256 36960 86264 37024
rect 85944 36959 86264 36960
rect 89944 37024 90264 37025
rect 89944 36960 89952 37024
rect 90016 36960 90032 37024
rect 90096 36960 90112 37024
rect 90176 36960 90192 37024
rect 90256 36960 90264 37024
rect 89944 36959 90264 36960
rect 86953 36818 87019 36821
rect 90406 36818 90466 37030
rect 91200 37000 92000 37030
rect 86953 36816 90466 36818
rect 86953 36760 86958 36816
rect 87014 36760 90466 36816
rect 86953 36758 90466 36760
rect 86953 36755 87019 36758
rect 3944 36480 4264 36481
rect 3944 36416 3952 36480
rect 4016 36416 4032 36480
rect 4096 36416 4112 36480
rect 4176 36416 4192 36480
rect 4256 36416 4264 36480
rect 3944 36415 4264 36416
rect 87944 36480 88264 36481
rect 87944 36416 87952 36480
rect 88016 36416 88032 36480
rect 88096 36416 88112 36480
rect 88176 36416 88192 36480
rect 88256 36416 88264 36480
rect 87944 36415 88264 36416
rect 1944 35936 2264 35937
rect 1944 35872 1952 35936
rect 2016 35872 2032 35936
rect 2096 35872 2112 35936
rect 2176 35872 2192 35936
rect 2256 35872 2264 35936
rect 1944 35871 2264 35872
rect 85944 35936 86264 35937
rect 85944 35872 85952 35936
rect 86016 35872 86032 35936
rect 86096 35872 86112 35936
rect 86176 35872 86192 35936
rect 86256 35872 86264 35936
rect 85944 35871 86264 35872
rect 89944 35936 90264 35937
rect 89944 35872 89952 35936
rect 90016 35872 90032 35936
rect 90096 35872 90112 35936
rect 90176 35872 90192 35936
rect 90256 35872 90264 35936
rect 89944 35871 90264 35872
rect 91200 35866 92000 35896
rect 90406 35806 92000 35866
rect 87321 35730 87387 35733
rect 90406 35730 90466 35806
rect 91200 35776 92000 35806
rect 87321 35728 90466 35730
rect 87321 35672 87326 35728
rect 87382 35672 90466 35728
rect 87321 35670 90466 35672
rect 87321 35667 87387 35670
rect 3944 35392 4264 35393
rect 3944 35328 3952 35392
rect 4016 35328 4032 35392
rect 4096 35328 4112 35392
rect 4176 35328 4192 35392
rect 4256 35328 4264 35392
rect 3944 35327 4264 35328
rect 87944 35392 88264 35393
rect 87944 35328 87952 35392
rect 88016 35328 88032 35392
rect 88096 35328 88112 35392
rect 88176 35328 88192 35392
rect 88256 35328 88264 35392
rect 87944 35327 88264 35328
rect 1944 34848 2264 34849
rect 1944 34784 1952 34848
rect 2016 34784 2032 34848
rect 2096 34784 2112 34848
rect 2176 34784 2192 34848
rect 2256 34784 2264 34848
rect 1944 34783 2264 34784
rect 85944 34848 86264 34849
rect 85944 34784 85952 34848
rect 86016 34784 86032 34848
rect 86096 34784 86112 34848
rect 86176 34784 86192 34848
rect 86256 34784 86264 34848
rect 85944 34783 86264 34784
rect 89944 34848 90264 34849
rect 89944 34784 89952 34848
rect 90016 34784 90032 34848
rect 90096 34784 90112 34848
rect 90176 34784 90192 34848
rect 90256 34784 90264 34848
rect 89944 34783 90264 34784
rect 86953 34642 87019 34645
rect 91200 34642 92000 34672
rect 86953 34640 92000 34642
rect 86953 34584 86958 34640
rect 87014 34584 92000 34640
rect 86953 34582 92000 34584
rect 86953 34579 87019 34582
rect 91200 34552 92000 34582
rect 3944 34304 4264 34305
rect 3944 34240 3952 34304
rect 4016 34240 4032 34304
rect 4096 34240 4112 34304
rect 4176 34240 4192 34304
rect 4256 34240 4264 34304
rect 3944 34239 4264 34240
rect 87944 34304 88264 34305
rect 87944 34240 87952 34304
rect 88016 34240 88032 34304
rect 88096 34240 88112 34304
rect 88176 34240 88192 34304
rect 88256 34240 88264 34304
rect 87944 34239 88264 34240
rect 83406 33764 83412 33828
rect 83476 33826 83482 33828
rect 83958 33826 83964 33828
rect 83476 33766 83964 33826
rect 83476 33764 83482 33766
rect 83958 33764 83964 33766
rect 84028 33764 84034 33828
rect 1944 33760 2264 33761
rect 1944 33696 1952 33760
rect 2016 33696 2032 33760
rect 2096 33696 2112 33760
rect 2176 33696 2192 33760
rect 2256 33696 2264 33760
rect 1944 33695 2264 33696
rect 85944 33760 86264 33761
rect 85944 33696 85952 33760
rect 86016 33696 86032 33760
rect 86096 33696 86112 33760
rect 86176 33696 86192 33760
rect 86256 33696 86264 33760
rect 85944 33695 86264 33696
rect 89944 33760 90264 33761
rect 89944 33696 89952 33760
rect 90016 33696 90032 33760
rect 90096 33696 90112 33760
rect 90176 33696 90192 33760
rect 90256 33696 90264 33760
rect 89944 33695 90264 33696
rect 86769 33418 86835 33421
rect 91200 33418 92000 33448
rect 86769 33416 92000 33418
rect 86769 33360 86774 33416
rect 86830 33360 92000 33416
rect 86769 33358 92000 33360
rect 86769 33355 86835 33358
rect 91200 33328 92000 33358
rect 3944 33216 4264 33217
rect 3944 33152 3952 33216
rect 4016 33152 4032 33216
rect 4096 33152 4112 33216
rect 4176 33152 4192 33216
rect 4256 33152 4264 33216
rect 3944 33151 4264 33152
rect 87944 33216 88264 33217
rect 87944 33152 87952 33216
rect 88016 33152 88032 33216
rect 88096 33152 88112 33216
rect 88176 33152 88192 33216
rect 88256 33152 88264 33216
rect 87944 33151 88264 33152
rect 1944 32672 2264 32673
rect 1944 32608 1952 32672
rect 2016 32608 2032 32672
rect 2096 32608 2112 32672
rect 2176 32608 2192 32672
rect 2256 32608 2264 32672
rect 1944 32607 2264 32608
rect 85944 32672 86264 32673
rect 85944 32608 85952 32672
rect 86016 32608 86032 32672
rect 86096 32608 86112 32672
rect 86176 32608 86192 32672
rect 86256 32608 86264 32672
rect 85944 32607 86264 32608
rect 89944 32672 90264 32673
rect 89944 32608 89952 32672
rect 90016 32608 90032 32672
rect 90096 32608 90112 32672
rect 90176 32608 90192 32672
rect 90256 32608 90264 32672
rect 89944 32607 90264 32608
rect 91200 32194 92000 32224
rect 88382 32134 92000 32194
rect 3944 32128 4264 32129
rect 3944 32064 3952 32128
rect 4016 32064 4032 32128
rect 4096 32064 4112 32128
rect 4176 32064 4192 32128
rect 4256 32064 4264 32128
rect 3944 32063 4264 32064
rect 87944 32128 88264 32129
rect 87944 32064 87952 32128
rect 88016 32064 88032 32128
rect 88096 32064 88112 32128
rect 88176 32064 88192 32128
rect 88256 32064 88264 32128
rect 87944 32063 88264 32064
rect 84745 32058 84811 32061
rect 83230 32056 84811 32058
rect 83230 32000 84750 32056
rect 84806 32000 84811 32056
rect 83230 31998 84811 32000
rect 83230 31773 83290 31998
rect 84745 31995 84811 31998
rect 86953 31922 87019 31925
rect 88382 31922 88442 32134
rect 91200 32104 92000 32134
rect 86953 31920 88442 31922
rect 86953 31864 86958 31920
rect 87014 31864 88442 31920
rect 86953 31862 88442 31864
rect 86953 31859 87019 31862
rect 1944 31584 2264 31585
rect 1944 31520 1952 31584
rect 2016 31520 2032 31584
rect 2096 31520 2112 31584
rect 2176 31520 2192 31584
rect 2256 31520 2264 31584
rect 1944 31519 2264 31520
rect 85944 31584 86264 31585
rect 85944 31520 85952 31584
rect 86016 31520 86032 31584
rect 86096 31520 86112 31584
rect 86176 31520 86192 31584
rect 86256 31520 86264 31584
rect 85944 31519 86264 31520
rect 89944 31584 90264 31585
rect 89944 31520 89952 31584
rect 90016 31520 90032 31584
rect 90096 31520 90112 31584
rect 90176 31520 90192 31584
rect 90256 31520 90264 31584
rect 89944 31519 90264 31520
rect 3944 31040 4264 31041
rect 3944 30976 3952 31040
rect 4016 30976 4032 31040
rect 4096 30976 4112 31040
rect 4176 30976 4192 31040
rect 4256 30976 4264 31040
rect 3944 30975 4264 30976
rect 87944 31040 88264 31041
rect 87944 30976 87952 31040
rect 88016 30976 88032 31040
rect 88096 30976 88112 31040
rect 88176 30976 88192 31040
rect 88256 30976 88264 31040
rect 87944 30975 88264 30976
rect 91200 30970 92000 31000
rect 89670 30910 92000 30970
rect 86585 30834 86651 30837
rect 89670 30834 89730 30910
rect 91200 30880 92000 30910
rect 86585 30832 89730 30834
rect 86585 30776 86590 30832
rect 86646 30776 89730 30832
rect 86585 30774 89730 30776
rect 86585 30771 86651 30774
rect 1944 30496 2264 30497
rect 1944 30432 1952 30496
rect 2016 30432 2032 30496
rect 2096 30432 2112 30496
rect 2176 30432 2192 30496
rect 2256 30432 2264 30496
rect 1944 30431 2264 30432
rect 85944 30496 86264 30497
rect 85944 30432 85952 30496
rect 86016 30432 86032 30496
rect 86096 30432 86112 30496
rect 86176 30432 86192 30496
rect 86256 30432 86264 30496
rect 85944 30431 86264 30432
rect 89944 30496 90264 30497
rect 89944 30432 89952 30496
rect 90016 30432 90032 30496
rect 90096 30432 90112 30496
rect 90176 30432 90192 30496
rect 90256 30432 90264 30496
rect 89944 30431 90264 30432
rect 84745 30290 84811 30293
rect 83230 30288 84811 30290
rect 83230 30232 84750 30288
rect 84806 30232 84811 30288
rect 83230 30230 84811 30232
rect 83230 30073 83290 30230
rect 84745 30227 84811 30230
rect 3944 29952 4264 29953
rect 3944 29888 3952 29952
rect 4016 29888 4032 29952
rect 4096 29888 4112 29952
rect 4176 29888 4192 29952
rect 4256 29888 4264 29952
rect 3944 29887 4264 29888
rect 87944 29952 88264 29953
rect 87944 29888 87952 29952
rect 88016 29888 88032 29952
rect 88096 29888 88112 29952
rect 88176 29888 88192 29952
rect 88256 29888 88264 29952
rect 87944 29887 88264 29888
rect 86953 29746 87019 29749
rect 91200 29746 92000 29776
rect 86953 29744 92000 29746
rect 86953 29688 86958 29744
rect 87014 29688 92000 29744
rect 86953 29686 92000 29688
rect 86953 29683 87019 29686
rect 91200 29656 92000 29686
rect 1944 29408 2264 29409
rect 1944 29344 1952 29408
rect 2016 29344 2032 29408
rect 2096 29344 2112 29408
rect 2176 29344 2192 29408
rect 2256 29344 2264 29408
rect 1944 29343 2264 29344
rect 85944 29408 86264 29409
rect 85944 29344 85952 29408
rect 86016 29344 86032 29408
rect 86096 29344 86112 29408
rect 86176 29344 86192 29408
rect 86256 29344 86264 29408
rect 85944 29343 86264 29344
rect 89944 29408 90264 29409
rect 89944 29344 89952 29408
rect 90016 29344 90032 29408
rect 90096 29344 90112 29408
rect 90176 29344 90192 29408
rect 90256 29344 90264 29408
rect 89944 29343 90264 29344
rect 83230 28930 83290 28945
rect 84561 28930 84627 28933
rect 83230 28928 84627 28930
rect 83230 28872 84566 28928
rect 84622 28872 84627 28928
rect 83230 28870 84627 28872
rect 84561 28867 84627 28870
rect 3944 28864 4264 28865
rect 3944 28800 3952 28864
rect 4016 28800 4032 28864
rect 4096 28800 4112 28864
rect 4176 28800 4192 28864
rect 4256 28800 4264 28864
rect 3944 28799 4264 28800
rect 87944 28864 88264 28865
rect 87944 28800 87952 28864
rect 88016 28800 88032 28864
rect 88096 28800 88112 28864
rect 88176 28800 88192 28864
rect 88256 28800 88264 28864
rect 87944 28799 88264 28800
rect 86953 28522 87019 28525
rect 91200 28522 92000 28552
rect 86953 28520 92000 28522
rect 86953 28464 86958 28520
rect 87014 28464 92000 28520
rect 86953 28462 92000 28464
rect 86953 28459 87019 28462
rect 91200 28432 92000 28462
rect 1944 28320 2264 28321
rect 1944 28256 1952 28320
rect 2016 28256 2032 28320
rect 2096 28256 2112 28320
rect 2176 28256 2192 28320
rect 2256 28256 2264 28320
rect 1944 28255 2264 28256
rect 85944 28320 86264 28321
rect 85944 28256 85952 28320
rect 86016 28256 86032 28320
rect 86096 28256 86112 28320
rect 86176 28256 86192 28320
rect 86256 28256 86264 28320
rect 85944 28255 86264 28256
rect 89944 28320 90264 28321
rect 89944 28256 89952 28320
rect 90016 28256 90032 28320
rect 90096 28256 90112 28320
rect 90176 28256 90192 28320
rect 90256 28256 90264 28320
rect 89944 28255 90264 28256
rect 3944 27776 4264 27777
rect 3944 27712 3952 27776
rect 4016 27712 4032 27776
rect 4096 27712 4112 27776
rect 4176 27712 4192 27776
rect 4256 27712 4264 27776
rect 3944 27711 4264 27712
rect 87944 27776 88264 27777
rect 87944 27712 87952 27776
rect 88016 27712 88032 27776
rect 88096 27712 88112 27776
rect 88176 27712 88192 27776
rect 88256 27712 88264 27776
rect 87944 27711 88264 27712
rect 84561 27570 84627 27573
rect 83230 27568 84627 27570
rect 83230 27512 84566 27568
rect 84622 27512 84627 27568
rect 83230 27510 84627 27512
rect 83230 27245 83290 27510
rect 84561 27507 84627 27510
rect 91200 27298 92000 27328
rect 90406 27238 92000 27298
rect 1944 27232 2264 27233
rect 1944 27168 1952 27232
rect 2016 27168 2032 27232
rect 2096 27168 2112 27232
rect 2176 27168 2192 27232
rect 2256 27168 2264 27232
rect 1944 27167 2264 27168
rect 85944 27232 86264 27233
rect 85944 27168 85952 27232
rect 86016 27168 86032 27232
rect 86096 27168 86112 27232
rect 86176 27168 86192 27232
rect 86256 27168 86264 27232
rect 85944 27167 86264 27168
rect 89944 27232 90264 27233
rect 89944 27168 89952 27232
rect 90016 27168 90032 27232
rect 90096 27168 90112 27232
rect 90176 27168 90192 27232
rect 90256 27168 90264 27232
rect 89944 27167 90264 27168
rect 86953 27026 87019 27029
rect 90406 27026 90466 27238
rect 91200 27208 92000 27238
rect 86953 27024 90466 27026
rect 86953 26968 86958 27024
rect 87014 26968 90466 27024
rect 86953 26966 90466 26968
rect 86953 26963 87019 26966
rect 3944 26688 4264 26689
rect 3944 26624 3952 26688
rect 4016 26624 4032 26688
rect 4096 26624 4112 26688
rect 4176 26624 4192 26688
rect 4256 26624 4264 26688
rect 3944 26623 4264 26624
rect 87944 26688 88264 26689
rect 87944 26624 87952 26688
rect 88016 26624 88032 26688
rect 88096 26624 88112 26688
rect 88176 26624 88192 26688
rect 88256 26624 88264 26688
rect 87944 26623 88264 26624
rect 84561 26210 84627 26213
rect 83782 26208 84627 26210
rect 83782 26152 84566 26208
rect 84622 26152 84627 26208
rect 83782 26150 84627 26152
rect 83782 26147 83842 26150
rect 84561 26147 84627 26150
rect 1944 26144 2264 26145
rect 1944 26080 1952 26144
rect 2016 26080 2032 26144
rect 2096 26080 2112 26144
rect 2176 26080 2192 26144
rect 2256 26080 2264 26144
rect 83260 26087 83842 26147
rect 85944 26144 86264 26145
rect 1944 26079 2264 26080
rect 85944 26080 85952 26144
rect 86016 26080 86032 26144
rect 86096 26080 86112 26144
rect 86176 26080 86192 26144
rect 86256 26080 86264 26144
rect 85944 26079 86264 26080
rect 89944 26144 90264 26145
rect 89944 26080 89952 26144
rect 90016 26080 90032 26144
rect 90096 26080 90112 26144
rect 90176 26080 90192 26144
rect 90256 26080 90264 26144
rect 89944 26079 90264 26080
rect 91200 26074 92000 26104
rect 90406 26014 92000 26074
rect 87229 25938 87295 25941
rect 90406 25938 90466 26014
rect 91200 25984 92000 26014
rect 87229 25936 90466 25938
rect 87229 25880 87234 25936
rect 87290 25880 90466 25936
rect 87229 25878 90466 25880
rect 87229 25875 87295 25878
rect 3944 25600 4264 25601
rect 3944 25536 3952 25600
rect 4016 25536 4032 25600
rect 4096 25536 4112 25600
rect 4176 25536 4192 25600
rect 4256 25536 4264 25600
rect 3944 25535 4264 25536
rect 87944 25600 88264 25601
rect 87944 25536 87952 25600
rect 88016 25536 88032 25600
rect 88096 25536 88112 25600
rect 88176 25536 88192 25600
rect 88256 25536 88264 25600
rect 87944 25535 88264 25536
rect 1944 25056 2264 25057
rect 1944 24992 1952 25056
rect 2016 24992 2032 25056
rect 2096 24992 2112 25056
rect 2176 24992 2192 25056
rect 2256 24992 2264 25056
rect 1944 24991 2264 24992
rect 85944 25056 86264 25057
rect 85944 24992 85952 25056
rect 86016 24992 86032 25056
rect 86096 24992 86112 25056
rect 86176 24992 86192 25056
rect 86256 24992 86264 25056
rect 85944 24991 86264 24992
rect 89944 25056 90264 25057
rect 89944 24992 89952 25056
rect 90016 24992 90032 25056
rect 90096 24992 90112 25056
rect 90176 24992 90192 25056
rect 90256 24992 90264 25056
rect 89944 24991 90264 24992
rect 86953 24850 87019 24853
rect 91200 24850 92000 24880
rect 86953 24848 92000 24850
rect 86953 24792 86958 24848
rect 87014 24792 92000 24848
rect 86953 24790 92000 24792
rect 86953 24787 87019 24790
rect 91200 24760 92000 24790
rect 3944 24512 4264 24513
rect 3944 24448 3952 24512
rect 4016 24448 4032 24512
rect 4096 24448 4112 24512
rect 4176 24448 4192 24512
rect 4256 24448 4264 24512
rect 3944 24447 4264 24448
rect 87944 24512 88264 24513
rect 87944 24448 87952 24512
rect 88016 24448 88032 24512
rect 88096 24448 88112 24512
rect 88176 24448 88192 24512
rect 88256 24448 88264 24512
rect 87944 24447 88264 24448
rect 84285 24442 84351 24445
rect 83230 24440 84351 24442
rect 83230 24384 84290 24440
rect 84346 24384 84351 24440
rect 83230 24382 84351 24384
rect 84285 24379 84351 24382
rect 1944 23968 2264 23969
rect 1944 23904 1952 23968
rect 2016 23904 2032 23968
rect 2096 23904 2112 23968
rect 2176 23904 2192 23968
rect 2256 23904 2264 23968
rect 1944 23903 2264 23904
rect 85944 23968 86264 23969
rect 85944 23904 85952 23968
rect 86016 23904 86032 23968
rect 86096 23904 86112 23968
rect 86176 23904 86192 23968
rect 86256 23904 86264 23968
rect 85944 23903 86264 23904
rect 89944 23968 90264 23969
rect 89944 23904 89952 23968
rect 90016 23904 90032 23968
rect 90096 23904 90112 23968
rect 90176 23904 90192 23968
rect 90256 23904 90264 23968
rect 89944 23903 90264 23904
rect 87045 23626 87111 23629
rect 91200 23626 92000 23656
rect 87045 23624 92000 23626
rect 87045 23568 87050 23624
rect 87106 23568 92000 23624
rect 87045 23566 92000 23568
rect 87045 23563 87111 23566
rect 91200 23536 92000 23566
rect 3944 23424 4264 23425
rect 3944 23360 3952 23424
rect 4016 23360 4032 23424
rect 4096 23360 4112 23424
rect 4176 23360 4192 23424
rect 4256 23360 4264 23424
rect 3944 23359 4264 23360
rect 87944 23424 88264 23425
rect 87944 23360 87952 23424
rect 88016 23360 88032 23424
rect 88096 23360 88112 23424
rect 88176 23360 88192 23424
rect 88256 23360 88264 23424
rect 87944 23359 88264 23360
rect 84285 23354 84351 23357
rect 83230 23352 84351 23354
rect 83230 23296 84290 23352
rect 84346 23296 84351 23352
rect 83230 23294 84351 23296
rect 83230 23289 83290 23294
rect 84285 23291 84351 23294
rect 1944 22880 2264 22881
rect 1944 22816 1952 22880
rect 2016 22816 2032 22880
rect 2096 22816 2112 22880
rect 2176 22816 2192 22880
rect 2256 22816 2264 22880
rect 1944 22815 2264 22816
rect 85944 22880 86264 22881
rect 85944 22816 85952 22880
rect 86016 22816 86032 22880
rect 86096 22816 86112 22880
rect 86176 22816 86192 22880
rect 86256 22816 86264 22880
rect 85944 22815 86264 22816
rect 89944 22880 90264 22881
rect 89944 22816 89952 22880
rect 90016 22816 90032 22880
rect 90096 22816 90112 22880
rect 90176 22816 90192 22880
rect 90256 22816 90264 22880
rect 89944 22815 90264 22816
rect 4705 22402 4771 22405
rect 6318 22402 6378 22616
rect 87137 22538 87203 22541
rect 87137 22536 89730 22538
rect 87137 22480 87142 22536
rect 87198 22480 89730 22536
rect 87137 22478 89730 22480
rect 87137 22475 87203 22478
rect 4705 22400 6378 22402
rect 4705 22344 4710 22400
rect 4766 22344 6378 22400
rect 4705 22342 6378 22344
rect 89670 22402 89730 22478
rect 91200 22402 92000 22432
rect 89670 22342 92000 22402
rect 4705 22339 4771 22342
rect 3944 22336 4264 22337
rect 3944 22272 3952 22336
rect 4016 22272 4032 22336
rect 4096 22272 4112 22336
rect 4176 22272 4192 22336
rect 4256 22272 4264 22336
rect 3944 22271 4264 22272
rect 87944 22336 88264 22337
rect 87944 22272 87952 22336
rect 88016 22272 88032 22336
rect 88096 22272 88112 22336
rect 88176 22272 88192 22336
rect 88256 22272 88264 22336
rect 91200 22312 92000 22342
rect 87944 22271 88264 22272
rect 1944 21792 2264 21793
rect 1944 21728 1952 21792
rect 2016 21728 2032 21792
rect 2096 21728 2112 21792
rect 2176 21728 2192 21792
rect 2256 21728 2264 21792
rect 1944 21727 2264 21728
rect 85944 21792 86264 21793
rect 85944 21728 85952 21792
rect 86016 21728 86032 21792
rect 86096 21728 86112 21792
rect 86176 21728 86192 21792
rect 86256 21728 86264 21792
rect 85944 21727 86264 21728
rect 89944 21792 90264 21793
rect 89944 21728 89952 21792
rect 90016 21728 90032 21792
rect 90096 21728 90112 21792
rect 90176 21728 90192 21792
rect 90256 21728 90264 21792
rect 89944 21727 90264 21728
rect 3944 21248 4264 21249
rect 3944 21184 3952 21248
rect 4016 21184 4032 21248
rect 4096 21184 4112 21248
rect 4176 21184 4192 21248
rect 4256 21184 4264 21248
rect 3944 21183 4264 21184
rect 87944 21248 88264 21249
rect 87944 21184 87952 21248
rect 88016 21184 88032 21248
rect 88096 21184 88112 21248
rect 88176 21184 88192 21248
rect 88256 21184 88264 21248
rect 87944 21183 88264 21184
rect 91200 21178 92000 21208
rect 88382 21118 92000 21178
rect 87873 21042 87939 21045
rect 88382 21042 88442 21118
rect 91200 21088 92000 21118
rect 87873 21040 88442 21042
rect 87873 20984 87878 21040
rect 87934 20984 88442 21040
rect 87873 20982 88442 20984
rect 87873 20979 87939 20982
rect 4797 20906 4863 20909
rect 6134 20906 6194 20916
rect 4797 20904 6194 20906
rect 4797 20848 4802 20904
rect 4858 20848 6194 20904
rect 4797 20846 6194 20848
rect 4797 20843 4863 20846
rect 1944 20704 2264 20705
rect 1944 20640 1952 20704
rect 2016 20640 2032 20704
rect 2096 20640 2112 20704
rect 2176 20640 2192 20704
rect 2256 20640 2264 20704
rect 1944 20639 2264 20640
rect 85944 20704 86264 20705
rect 85944 20640 85952 20704
rect 86016 20640 86032 20704
rect 86096 20640 86112 20704
rect 86176 20640 86192 20704
rect 86256 20640 86264 20704
rect 85944 20639 86264 20640
rect 89944 20704 90264 20705
rect 89944 20640 89952 20704
rect 90016 20640 90032 20704
rect 90096 20640 90112 20704
rect 90176 20640 90192 20704
rect 90256 20640 90264 20704
rect 89944 20639 90264 20640
rect 3944 20160 4264 20161
rect 3944 20096 3952 20160
rect 4016 20096 4032 20160
rect 4096 20096 4112 20160
rect 4176 20096 4192 20160
rect 4256 20096 4264 20160
rect 3944 20095 4264 20096
rect 87944 20160 88264 20161
rect 87944 20096 87952 20160
rect 88016 20096 88032 20160
rect 88096 20096 88112 20160
rect 88176 20096 88192 20160
rect 88256 20096 88264 20160
rect 87944 20095 88264 20096
rect 86309 19954 86375 19957
rect 91200 19954 92000 19984
rect 86309 19952 92000 19954
rect 86309 19896 86314 19952
rect 86370 19896 92000 19952
rect 86309 19894 92000 19896
rect 86309 19891 86375 19894
rect 91200 19864 92000 19894
rect 1944 19616 2264 19617
rect 1944 19552 1952 19616
rect 2016 19552 2032 19616
rect 2096 19552 2112 19616
rect 2176 19552 2192 19616
rect 2256 19552 2264 19616
rect 1944 19551 2264 19552
rect 85944 19616 86264 19617
rect 85944 19552 85952 19616
rect 86016 19552 86032 19616
rect 86096 19552 86112 19616
rect 86176 19552 86192 19616
rect 86256 19552 86264 19616
rect 85944 19551 86264 19552
rect 89944 19616 90264 19617
rect 89944 19552 89952 19616
rect 90016 19552 90032 19616
rect 90096 19552 90112 19616
rect 90176 19552 90192 19616
rect 90256 19552 90264 19616
rect 89944 19551 90264 19552
rect 3944 19072 4264 19073
rect 3944 19008 3952 19072
rect 4016 19008 4032 19072
rect 4096 19008 4112 19072
rect 4176 19008 4192 19072
rect 4256 19008 4264 19072
rect 3944 19007 4264 19008
rect 87944 19072 88264 19073
rect 87944 19008 87952 19072
rect 88016 19008 88032 19072
rect 88096 19008 88112 19072
rect 88176 19008 88192 19072
rect 88256 19008 88264 19072
rect 87944 19007 88264 19008
rect 87137 18866 87203 18869
rect 91200 18866 92000 18896
rect 87137 18864 92000 18866
rect 87137 18808 87142 18864
rect 87198 18808 92000 18864
rect 87137 18806 92000 18808
rect 87137 18803 87203 18806
rect 91200 18776 92000 18806
rect 1944 18528 2264 18529
rect 1944 18464 1952 18528
rect 2016 18464 2032 18528
rect 2096 18464 2112 18528
rect 2176 18464 2192 18528
rect 2256 18464 2264 18528
rect 1944 18463 2264 18464
rect 85944 18528 86264 18529
rect 85944 18464 85952 18528
rect 86016 18464 86032 18528
rect 86096 18464 86112 18528
rect 86176 18464 86192 18528
rect 86256 18464 86264 18528
rect 85944 18463 86264 18464
rect 89944 18528 90264 18529
rect 89944 18464 89952 18528
rect 90016 18464 90032 18528
rect 90096 18464 90112 18528
rect 90176 18464 90192 18528
rect 90256 18464 90264 18528
rect 89944 18463 90264 18464
rect 3944 17984 4264 17985
rect 3944 17920 3952 17984
rect 4016 17920 4032 17984
rect 4096 17920 4112 17984
rect 4176 17920 4192 17984
rect 4256 17920 4264 17984
rect 3944 17919 4264 17920
rect 87944 17984 88264 17985
rect 87944 17920 87952 17984
rect 88016 17920 88032 17984
rect 88096 17920 88112 17984
rect 88176 17920 88192 17984
rect 88256 17920 88264 17984
rect 87944 17919 88264 17920
rect 87229 17642 87295 17645
rect 91200 17642 92000 17672
rect 87229 17640 92000 17642
rect 87229 17584 87234 17640
rect 87290 17584 92000 17640
rect 87229 17582 92000 17584
rect 87229 17579 87295 17582
rect 91200 17552 92000 17582
rect 1944 17440 2264 17441
rect 1944 17376 1952 17440
rect 2016 17376 2032 17440
rect 2096 17376 2112 17440
rect 2176 17376 2192 17440
rect 2256 17376 2264 17440
rect 1944 17375 2264 17376
rect 85944 17440 86264 17441
rect 85944 17376 85952 17440
rect 86016 17376 86032 17440
rect 86096 17376 86112 17440
rect 86176 17376 86192 17440
rect 86256 17376 86264 17440
rect 85944 17375 86264 17376
rect 89944 17440 90264 17441
rect 89944 17376 89952 17440
rect 90016 17376 90032 17440
rect 90096 17376 90112 17440
rect 90176 17376 90192 17440
rect 90256 17376 90264 17440
rect 89944 17375 90264 17376
rect 3944 16896 4264 16897
rect 3944 16832 3952 16896
rect 4016 16832 4032 16896
rect 4096 16832 4112 16896
rect 4176 16832 4192 16896
rect 4256 16832 4264 16896
rect 3944 16831 4264 16832
rect 87944 16896 88264 16897
rect 87944 16832 87952 16896
rect 88016 16832 88032 16896
rect 88096 16832 88112 16896
rect 88176 16832 88192 16896
rect 88256 16832 88264 16896
rect 87944 16831 88264 16832
rect 82445 16690 82511 16693
rect 84142 16690 84148 16692
rect 82445 16688 84148 16690
rect 82445 16632 82450 16688
rect 82506 16632 84148 16688
rect 82445 16630 84148 16632
rect 82445 16627 82511 16630
rect 84142 16628 84148 16630
rect 84212 16628 84218 16692
rect 91200 16418 92000 16448
rect 90406 16358 92000 16418
rect 1944 16352 2264 16353
rect 1944 16288 1952 16352
rect 2016 16288 2032 16352
rect 2096 16288 2112 16352
rect 2176 16288 2192 16352
rect 2256 16288 2264 16352
rect 1944 16287 2264 16288
rect 85944 16352 86264 16353
rect 85944 16288 85952 16352
rect 86016 16288 86032 16352
rect 86096 16288 86112 16352
rect 86176 16288 86192 16352
rect 86256 16288 86264 16352
rect 85944 16287 86264 16288
rect 89944 16352 90264 16353
rect 89944 16288 89952 16352
rect 90016 16288 90032 16352
rect 90096 16288 90112 16352
rect 90176 16288 90192 16352
rect 90256 16288 90264 16352
rect 89944 16287 90264 16288
rect 87137 16146 87203 16149
rect 90406 16146 90466 16358
rect 91200 16328 92000 16358
rect 87137 16144 90466 16146
rect 87137 16088 87142 16144
rect 87198 16088 90466 16144
rect 87137 16086 90466 16088
rect 87137 16083 87203 16086
rect 3944 15808 4264 15809
rect 3944 15744 3952 15808
rect 4016 15744 4032 15808
rect 4096 15744 4112 15808
rect 4176 15744 4192 15808
rect 4256 15744 4264 15808
rect 3944 15743 4264 15744
rect 87944 15808 88264 15809
rect 87944 15744 87952 15808
rect 88016 15744 88032 15808
rect 88096 15744 88112 15808
rect 88176 15744 88192 15808
rect 88256 15744 88264 15808
rect 87944 15743 88264 15744
rect 1944 15264 2264 15265
rect 1944 15200 1952 15264
rect 2016 15200 2032 15264
rect 2096 15200 2112 15264
rect 2176 15200 2192 15264
rect 2256 15200 2264 15264
rect 1944 15199 2264 15200
rect 85944 15264 86264 15265
rect 85944 15200 85952 15264
rect 86016 15200 86032 15264
rect 86096 15200 86112 15264
rect 86176 15200 86192 15264
rect 86256 15200 86264 15264
rect 85944 15199 86264 15200
rect 89944 15264 90264 15265
rect 89944 15200 89952 15264
rect 90016 15200 90032 15264
rect 90096 15200 90112 15264
rect 90176 15200 90192 15264
rect 90256 15200 90264 15264
rect 89944 15199 90264 15200
rect 91200 15194 92000 15224
rect 90406 15134 92000 15194
rect 87137 15058 87203 15061
rect 90406 15058 90466 15134
rect 91200 15104 92000 15134
rect 87137 15056 90466 15058
rect 87137 15000 87142 15056
rect 87198 15000 90466 15056
rect 87137 14998 90466 15000
rect 87137 14995 87203 14998
rect 3944 14720 4264 14721
rect 3944 14656 3952 14720
rect 4016 14656 4032 14720
rect 4096 14656 4112 14720
rect 4176 14656 4192 14720
rect 4256 14656 4264 14720
rect 3944 14655 4264 14656
rect 87944 14720 88264 14721
rect 87944 14656 87952 14720
rect 88016 14656 88032 14720
rect 88096 14656 88112 14720
rect 88176 14656 88192 14720
rect 88256 14656 88264 14720
rect 87944 14655 88264 14656
rect 1944 14176 2264 14177
rect 1944 14112 1952 14176
rect 2016 14112 2032 14176
rect 2096 14112 2112 14176
rect 2176 14112 2192 14176
rect 2256 14112 2264 14176
rect 1944 14111 2264 14112
rect 85944 14176 86264 14177
rect 85944 14112 85952 14176
rect 86016 14112 86032 14176
rect 86096 14112 86112 14176
rect 86176 14112 86192 14176
rect 86256 14112 86264 14176
rect 85944 14111 86264 14112
rect 89944 14176 90264 14177
rect 89944 14112 89952 14176
rect 90016 14112 90032 14176
rect 90096 14112 90112 14176
rect 90176 14112 90192 14176
rect 90256 14112 90264 14176
rect 89944 14111 90264 14112
rect 86401 13970 86467 13973
rect 91200 13970 92000 14000
rect 86401 13968 92000 13970
rect 86401 13912 86406 13968
rect 86462 13912 92000 13968
rect 86401 13910 92000 13912
rect 86401 13907 86467 13910
rect 91200 13880 92000 13910
rect 3944 13632 4264 13633
rect 3944 13568 3952 13632
rect 4016 13568 4032 13632
rect 4096 13568 4112 13632
rect 4176 13568 4192 13632
rect 4256 13568 4264 13632
rect 3944 13567 4264 13568
rect 87944 13632 88264 13633
rect 87944 13568 87952 13632
rect 88016 13568 88032 13632
rect 88096 13568 88112 13632
rect 88176 13568 88192 13632
rect 88256 13568 88264 13632
rect 87944 13567 88264 13568
rect 1944 13088 2264 13089
rect 1944 13024 1952 13088
rect 2016 13024 2032 13088
rect 2096 13024 2112 13088
rect 2176 13024 2192 13088
rect 2256 13024 2264 13088
rect 1944 13023 2264 13024
rect 85944 13088 86264 13089
rect 85944 13024 85952 13088
rect 86016 13024 86032 13088
rect 86096 13024 86112 13088
rect 86176 13024 86192 13088
rect 86256 13024 86264 13088
rect 85944 13023 86264 13024
rect 89944 13088 90264 13089
rect 89944 13024 89952 13088
rect 90016 13024 90032 13088
rect 90096 13024 90112 13088
rect 90176 13024 90192 13088
rect 90256 13024 90264 13088
rect 89944 13023 90264 13024
rect 86953 12746 87019 12749
rect 91200 12746 92000 12776
rect 86953 12744 92000 12746
rect 86953 12688 86958 12744
rect 87014 12688 92000 12744
rect 86953 12686 92000 12688
rect 86953 12683 87019 12686
rect 91200 12656 92000 12686
rect 3944 12544 4264 12545
rect 3944 12480 3952 12544
rect 4016 12480 4032 12544
rect 4096 12480 4112 12544
rect 4176 12480 4192 12544
rect 4256 12480 4264 12544
rect 3944 12479 4264 12480
rect 87944 12544 88264 12545
rect 87944 12480 87952 12544
rect 88016 12480 88032 12544
rect 88096 12480 88112 12544
rect 88176 12480 88192 12544
rect 88256 12480 88264 12544
rect 87944 12479 88264 12480
rect 1944 12000 2264 12001
rect 1944 11936 1952 12000
rect 2016 11936 2032 12000
rect 2096 11936 2112 12000
rect 2176 11936 2192 12000
rect 2256 11936 2264 12000
rect 1944 11935 2264 11936
rect 85944 12000 86264 12001
rect 85944 11936 85952 12000
rect 86016 11936 86032 12000
rect 86096 11936 86112 12000
rect 86176 11936 86192 12000
rect 86256 11936 86264 12000
rect 85944 11935 86264 11936
rect 89944 12000 90264 12001
rect 89944 11936 89952 12000
rect 90016 11936 90032 12000
rect 90096 11936 90112 12000
rect 90176 11936 90192 12000
rect 90256 11936 90264 12000
rect 89944 11935 90264 11936
rect 91200 11522 92000 11552
rect 89670 11462 92000 11522
rect 3944 11456 4264 11457
rect 3944 11392 3952 11456
rect 4016 11392 4032 11456
rect 4096 11392 4112 11456
rect 4176 11392 4192 11456
rect 4256 11392 4264 11456
rect 3944 11391 4264 11392
rect 87944 11456 88264 11457
rect 87944 11392 87952 11456
rect 88016 11392 88032 11456
rect 88096 11392 88112 11456
rect 88176 11392 88192 11456
rect 88256 11392 88264 11456
rect 87944 11391 88264 11392
rect 86953 11250 87019 11253
rect 89670 11250 89730 11462
rect 91200 11432 92000 11462
rect 86953 11248 89730 11250
rect 86953 11192 86958 11248
rect 87014 11192 89730 11248
rect 86953 11190 89730 11192
rect 86953 11187 87019 11190
rect 1944 10912 2264 10913
rect 1944 10848 1952 10912
rect 2016 10848 2032 10912
rect 2096 10848 2112 10912
rect 2176 10848 2192 10912
rect 2256 10848 2264 10912
rect 1944 10847 2264 10848
rect 85944 10912 86264 10913
rect 85944 10848 85952 10912
rect 86016 10848 86032 10912
rect 86096 10848 86112 10912
rect 86176 10848 86192 10912
rect 86256 10848 86264 10912
rect 85944 10847 86264 10848
rect 89944 10912 90264 10913
rect 89944 10848 89952 10912
rect 90016 10848 90032 10912
rect 90096 10848 90112 10912
rect 90176 10848 90192 10912
rect 90256 10848 90264 10912
rect 89944 10847 90264 10848
rect 3944 10368 4264 10369
rect 3944 10304 3952 10368
rect 4016 10304 4032 10368
rect 4096 10304 4112 10368
rect 4176 10304 4192 10368
rect 4256 10304 4264 10368
rect 3944 10303 4264 10304
rect 87944 10368 88264 10369
rect 87944 10304 87952 10368
rect 88016 10304 88032 10368
rect 88096 10304 88112 10368
rect 88176 10304 88192 10368
rect 88256 10304 88264 10368
rect 87944 10303 88264 10304
rect 91200 10298 92000 10328
rect 89670 10238 92000 10298
rect 4429 10164 4495 10165
rect 4429 10162 4476 10164
rect 4384 10160 4476 10162
rect 4384 10104 4434 10160
rect 4384 10102 4476 10104
rect 4429 10100 4476 10102
rect 4540 10100 4546 10164
rect 86493 10162 86559 10165
rect 89670 10162 89730 10238
rect 91200 10208 92000 10238
rect 86493 10160 89730 10162
rect 86493 10104 86498 10160
rect 86554 10104 89730 10160
rect 86493 10102 89730 10104
rect 4429 10099 4495 10100
rect 86493 10099 86559 10102
rect 1944 9824 2264 9825
rect 1944 9760 1952 9824
rect 2016 9760 2032 9824
rect 2096 9760 2112 9824
rect 2176 9760 2192 9824
rect 2256 9760 2264 9824
rect 1944 9759 2264 9760
rect 85944 9824 86264 9825
rect 85944 9760 85952 9824
rect 86016 9760 86032 9824
rect 86096 9760 86112 9824
rect 86176 9760 86192 9824
rect 86256 9760 86264 9824
rect 85944 9759 86264 9760
rect 89944 9824 90264 9825
rect 89944 9760 89952 9824
rect 90016 9760 90032 9824
rect 90096 9760 90112 9824
rect 90176 9760 90192 9824
rect 90256 9760 90264 9824
rect 89944 9759 90264 9760
rect 3944 9280 4264 9281
rect 3944 9216 3952 9280
rect 4016 9216 4032 9280
rect 4096 9216 4112 9280
rect 4176 9216 4192 9280
rect 4256 9216 4264 9280
rect 3944 9215 4264 9216
rect 87944 9280 88264 9281
rect 87944 9216 87952 9280
rect 88016 9216 88032 9280
rect 88096 9216 88112 9280
rect 88176 9216 88192 9280
rect 88256 9216 88264 9280
rect 87944 9215 88264 9216
rect 86953 9074 87019 9077
rect 91200 9074 92000 9104
rect 86953 9072 92000 9074
rect 86953 9016 86958 9072
rect 87014 9016 92000 9072
rect 86953 9014 92000 9016
rect 86953 9011 87019 9014
rect 91200 8984 92000 9014
rect 1944 8736 2264 8737
rect 1944 8672 1952 8736
rect 2016 8672 2032 8736
rect 2096 8672 2112 8736
rect 2176 8672 2192 8736
rect 2256 8672 2264 8736
rect 1944 8671 2264 8672
rect 85944 8736 86264 8737
rect 85944 8672 85952 8736
rect 86016 8672 86032 8736
rect 86096 8672 86112 8736
rect 86176 8672 86192 8736
rect 86256 8672 86264 8736
rect 85944 8671 86264 8672
rect 89944 8736 90264 8737
rect 89944 8672 89952 8736
rect 90016 8672 90032 8736
rect 90096 8672 90112 8736
rect 90176 8672 90192 8736
rect 90256 8672 90264 8736
rect 89944 8671 90264 8672
rect 3944 8192 4264 8193
rect 3944 8128 3952 8192
rect 4016 8128 4032 8192
rect 4096 8128 4112 8192
rect 4176 8128 4192 8192
rect 4256 8128 4264 8192
rect 3944 8127 4264 8128
rect 87944 8192 88264 8193
rect 87944 8128 87952 8192
rect 88016 8128 88032 8192
rect 88096 8128 88112 8192
rect 88176 8128 88192 8192
rect 88256 8128 88264 8192
rect 87944 8127 88264 8128
rect 87873 7850 87939 7853
rect 91200 7850 92000 7880
rect 87873 7848 92000 7850
rect 87873 7792 87878 7848
rect 87934 7792 92000 7848
rect 87873 7790 92000 7792
rect 87873 7787 87939 7790
rect 91200 7760 92000 7790
rect 1944 7648 2264 7649
rect 1944 7584 1952 7648
rect 2016 7584 2032 7648
rect 2096 7584 2112 7648
rect 2176 7584 2192 7648
rect 2256 7584 2264 7648
rect 1944 7583 2264 7584
rect 85944 7648 86264 7649
rect 85944 7584 85952 7648
rect 86016 7584 86032 7648
rect 86096 7584 86112 7648
rect 86176 7584 86192 7648
rect 86256 7584 86264 7648
rect 85944 7583 86264 7584
rect 89944 7648 90264 7649
rect 89944 7584 89952 7648
rect 90016 7584 90032 7648
rect 90096 7584 90112 7648
rect 90176 7584 90192 7648
rect 90256 7584 90264 7648
rect 89944 7583 90264 7584
rect 3944 7104 4264 7105
rect 3944 7040 3952 7104
rect 4016 7040 4032 7104
rect 4096 7040 4112 7104
rect 4176 7040 4192 7104
rect 4256 7040 4264 7104
rect 3944 7039 4264 7040
rect 87944 7104 88264 7105
rect 87944 7040 87952 7104
rect 88016 7040 88032 7104
rect 88096 7040 88112 7104
rect 88176 7040 88192 7104
rect 88256 7040 88264 7104
rect 87944 7039 88264 7040
rect 91200 6626 92000 6656
rect 90406 6566 92000 6626
rect 1944 6560 2264 6561
rect 1944 6496 1952 6560
rect 2016 6496 2032 6560
rect 2096 6496 2112 6560
rect 2176 6496 2192 6560
rect 2256 6496 2264 6560
rect 1944 6495 2264 6496
rect 85944 6560 86264 6561
rect 85944 6496 85952 6560
rect 86016 6496 86032 6560
rect 86096 6496 86112 6560
rect 86176 6496 86192 6560
rect 86256 6496 86264 6560
rect 85944 6495 86264 6496
rect 89944 6560 90264 6561
rect 89944 6496 89952 6560
rect 90016 6496 90032 6560
rect 90096 6496 90112 6560
rect 90176 6496 90192 6560
rect 90256 6496 90264 6560
rect 89944 6495 90264 6496
rect 87321 6354 87387 6357
rect 90406 6354 90466 6566
rect 91200 6536 92000 6566
rect 87321 6352 90466 6354
rect 87321 6296 87326 6352
rect 87382 6296 90466 6352
rect 87321 6294 90466 6296
rect 87321 6291 87387 6294
rect 3944 6016 4264 6017
rect 3944 5952 3952 6016
rect 4016 5952 4032 6016
rect 4096 5952 4112 6016
rect 4176 5952 4192 6016
rect 4256 5952 4264 6016
rect 3944 5951 4264 5952
rect 87944 6016 88264 6017
rect 87944 5952 87952 6016
rect 88016 5952 88032 6016
rect 88096 5952 88112 6016
rect 88176 5952 88192 6016
rect 88256 5952 88264 6016
rect 87944 5951 88264 5952
rect 1944 5472 2264 5473
rect 1944 5408 1952 5472
rect 2016 5408 2032 5472
rect 2096 5408 2112 5472
rect 2176 5408 2192 5472
rect 2256 5408 2264 5472
rect 1944 5407 2264 5408
rect 85944 5472 86264 5473
rect 85944 5408 85952 5472
rect 86016 5408 86032 5472
rect 86096 5408 86112 5472
rect 86176 5408 86192 5472
rect 86256 5408 86264 5472
rect 85944 5407 86264 5408
rect 89944 5472 90264 5473
rect 89944 5408 89952 5472
rect 90016 5408 90032 5472
rect 90096 5408 90112 5472
rect 90176 5408 90192 5472
rect 90256 5408 90264 5472
rect 89944 5407 90264 5408
rect 91200 5402 92000 5432
rect 90406 5342 92000 5402
rect 87045 5266 87111 5269
rect 90406 5266 90466 5342
rect 91200 5312 92000 5342
rect 87045 5264 90466 5266
rect 87045 5208 87050 5264
rect 87106 5208 90466 5264
rect 87045 5206 90466 5208
rect 87045 5203 87111 5206
rect 3944 4928 4264 4929
rect 3944 4864 3952 4928
rect 4016 4864 4032 4928
rect 4096 4864 4112 4928
rect 4176 4864 4192 4928
rect 4256 4864 4264 4928
rect 3944 4863 4264 4864
rect 87944 4928 88264 4929
rect 87944 4864 87952 4928
rect 88016 4864 88032 4928
rect 88096 4864 88112 4928
rect 88176 4864 88192 4928
rect 88256 4864 88264 4928
rect 87944 4863 88264 4864
rect 1944 4384 2264 4385
rect 1944 4320 1952 4384
rect 2016 4320 2032 4384
rect 2096 4320 2112 4384
rect 2176 4320 2192 4384
rect 2256 4320 2264 4384
rect 1944 4319 2264 4320
rect 85944 4384 86264 4385
rect 85944 4320 85952 4384
rect 86016 4320 86032 4384
rect 86096 4320 86112 4384
rect 86176 4320 86192 4384
rect 86256 4320 86264 4384
rect 85944 4319 86264 4320
rect 89944 4384 90264 4385
rect 89944 4320 89952 4384
rect 90016 4320 90032 4384
rect 90096 4320 90112 4384
rect 90176 4320 90192 4384
rect 90256 4320 90264 4384
rect 89944 4319 90264 4320
rect 87597 4178 87663 4181
rect 91200 4178 92000 4208
rect 87597 4176 92000 4178
rect 87597 4120 87602 4176
rect 87658 4120 92000 4176
rect 87597 4118 92000 4120
rect 87597 4115 87663 4118
rect 91200 4088 92000 4118
rect 4797 3908 4863 3909
rect 4797 3906 4844 3908
rect 4752 3904 4844 3906
rect 4752 3848 4802 3904
rect 4752 3846 4844 3848
rect 4797 3844 4844 3846
rect 4908 3844 4914 3908
rect 4797 3843 4863 3844
rect 3944 3840 4264 3841
rect 3944 3776 3952 3840
rect 4016 3776 4032 3840
rect 4096 3776 4112 3840
rect 4176 3776 4192 3840
rect 4256 3776 4264 3840
rect 3944 3775 4264 3776
rect 87944 3840 88264 3841
rect 87944 3776 87952 3840
rect 88016 3776 88032 3840
rect 88096 3776 88112 3840
rect 88176 3776 88192 3840
rect 88256 3776 88264 3840
rect 87944 3775 88264 3776
rect 3509 3362 3575 3365
rect 5901 3362 5967 3365
rect 3509 3360 5967 3362
rect 3509 3304 3514 3360
rect 3570 3304 5906 3360
rect 5962 3304 5967 3360
rect 3509 3302 5967 3304
rect 3509 3299 3575 3302
rect 5901 3299 5967 3302
rect 1944 3296 2264 3297
rect 1944 3232 1952 3296
rect 2016 3232 2032 3296
rect 2096 3232 2112 3296
rect 2176 3232 2192 3296
rect 2256 3232 2264 3296
rect 1944 3231 2264 3232
rect 85944 3296 86264 3297
rect 85944 3232 85952 3296
rect 86016 3232 86032 3296
rect 86096 3232 86112 3296
rect 86176 3232 86192 3296
rect 86256 3232 86264 3296
rect 85944 3231 86264 3232
rect 89944 3296 90264 3297
rect 89944 3232 89952 3296
rect 90016 3232 90032 3296
rect 90096 3232 90112 3296
rect 90176 3232 90192 3296
rect 90256 3232 90264 3296
rect 89944 3231 90264 3232
rect 4337 3226 4403 3229
rect 4613 3226 4679 3229
rect 47761 3228 47827 3229
rect 39062 3226 39068 3228
rect 4337 3224 39068 3226
rect 4337 3168 4342 3224
rect 4398 3168 4618 3224
rect 4674 3168 39068 3224
rect 4337 3166 39068 3168
rect 4337 3163 4403 3166
rect 4613 3163 4679 3166
rect 39062 3164 39068 3166
rect 39132 3164 39138 3228
rect 45318 3164 45324 3228
rect 45388 3226 45394 3228
rect 45388 3166 45570 3226
rect 45388 3164 45394 3166
rect 3785 3090 3851 3093
rect 4889 3090 4955 3093
rect 3785 3088 4955 3090
rect 3785 3032 3790 3088
rect 3846 3032 4894 3088
rect 4950 3032 4955 3088
rect 3785 3030 4955 3032
rect 3785 3027 3851 3030
rect 4889 3027 4955 3030
rect 5717 3090 5783 3093
rect 40166 3090 40172 3092
rect 5717 3088 40172 3090
rect 5717 3032 5722 3088
rect 5778 3032 40172 3088
rect 5717 3030 40172 3032
rect 5717 3027 5783 3030
rect 40166 3028 40172 3030
rect 40236 3028 40242 3092
rect 45510 3090 45570 3166
rect 47710 3164 47716 3228
rect 47780 3226 47827 3228
rect 48681 3226 48747 3229
rect 83181 3226 83247 3229
rect 47780 3224 47872 3226
rect 47822 3168 47872 3224
rect 47780 3166 47872 3168
rect 48681 3224 83247 3226
rect 48681 3168 48686 3224
rect 48742 3168 83186 3224
rect 83242 3168 83247 3224
rect 48681 3166 83247 3168
rect 47780 3164 47827 3166
rect 47761 3163 47827 3164
rect 48681 3163 48747 3166
rect 83181 3163 83247 3166
rect 83457 3090 83523 3093
rect 45510 3088 83523 3090
rect 45510 3032 83462 3088
rect 83518 3032 83523 3088
rect 45510 3030 83523 3032
rect 83457 3027 83523 3030
rect 3601 2954 3667 2957
rect 5625 2954 5691 2957
rect 6545 2954 6611 2957
rect 37958 2954 37964 2956
rect 3601 2952 4538 2954
rect 3601 2896 3606 2952
rect 3662 2896 4538 2952
rect 3601 2894 4538 2896
rect 3601 2891 3667 2894
rect 4478 2818 4538 2894
rect 5625 2952 37964 2954
rect 5625 2896 5630 2952
rect 5686 2896 6550 2952
rect 6606 2896 37964 2952
rect 5625 2894 37964 2896
rect 5625 2891 5691 2894
rect 6545 2891 6611 2894
rect 37958 2892 37964 2894
rect 38028 2892 38034 2956
rect 44030 2892 44036 2956
rect 44100 2954 44106 2956
rect 48681 2954 48747 2957
rect 49969 2956 50035 2957
rect 53465 2956 53531 2957
rect 49918 2954 49924 2956
rect 44100 2952 48747 2954
rect 44100 2896 48686 2952
rect 48742 2896 48747 2952
rect 44100 2894 48747 2896
rect 49878 2894 49924 2954
rect 49988 2952 50035 2956
rect 50030 2896 50035 2952
rect 44100 2892 44106 2894
rect 48681 2891 48747 2894
rect 49918 2892 49924 2894
rect 49988 2892 50035 2896
rect 53414 2892 53420 2956
rect 53484 2954 53531 2956
rect 82997 2954 83063 2957
rect 53484 2952 53576 2954
rect 53526 2896 53576 2952
rect 53484 2894 53576 2896
rect 55170 2952 83063 2954
rect 55170 2896 83002 2952
rect 83058 2896 83063 2952
rect 55170 2894 83063 2896
rect 53484 2892 53531 2894
rect 49969 2891 50035 2892
rect 53465 2891 53531 2892
rect 5349 2818 5415 2821
rect 25998 2818 26004 2820
rect 4478 2816 26004 2818
rect 4478 2760 5354 2816
rect 5410 2760 26004 2816
rect 4478 2758 26004 2760
rect 5349 2755 5415 2758
rect 25998 2756 26004 2758
rect 26068 2756 26074 2820
rect 46238 2756 46244 2820
rect 46308 2818 46314 2820
rect 55170 2818 55230 2894
rect 82997 2891 83063 2894
rect 87045 2954 87111 2957
rect 91200 2954 92000 2984
rect 87045 2952 92000 2954
rect 87045 2896 87050 2952
rect 87106 2896 92000 2952
rect 87045 2894 92000 2896
rect 87045 2891 87111 2894
rect 91200 2864 92000 2894
rect 46308 2758 55230 2818
rect 82905 2818 82971 2821
rect 83181 2818 83247 2821
rect 82905 2816 83247 2818
rect 82905 2760 82910 2816
rect 82966 2760 83186 2816
rect 83242 2760 83247 2816
rect 82905 2758 83247 2760
rect 46308 2756 46314 2758
rect 82905 2755 82971 2758
rect 83181 2755 83247 2758
rect 3944 2752 4264 2753
rect 3944 2688 3952 2752
rect 4016 2688 4032 2752
rect 4096 2688 4112 2752
rect 4176 2688 4192 2752
rect 4256 2688 4264 2752
rect 3944 2687 4264 2688
rect 87944 2752 88264 2753
rect 87944 2688 87952 2752
rect 88016 2688 88032 2752
rect 88096 2688 88112 2752
rect 88176 2688 88192 2752
rect 88256 2688 88264 2752
rect 87944 2687 88264 2688
rect 8109 2684 8175 2685
rect 15285 2684 15351 2685
rect 20713 2684 20779 2685
rect 8109 2682 8156 2684
rect 8064 2680 8156 2682
rect 8064 2624 8114 2680
rect 8064 2622 8156 2624
rect 8109 2620 8156 2622
rect 8220 2620 8226 2684
rect 15285 2680 15332 2684
rect 15396 2682 15402 2684
rect 15285 2624 15290 2680
rect 15285 2620 15332 2624
rect 15396 2622 15442 2682
rect 15396 2620 15402 2622
rect 20662 2620 20668 2684
rect 20732 2682 20779 2684
rect 25037 2684 25103 2685
rect 25037 2682 25084 2684
rect 20732 2680 20824 2682
rect 20774 2624 20824 2680
rect 20732 2622 20824 2624
rect 24992 2680 25084 2682
rect 24992 2624 25042 2680
rect 24992 2622 25084 2624
rect 20732 2620 20779 2622
rect 8109 2619 8175 2620
rect 15285 2619 15351 2620
rect 20713 2619 20779 2620
rect 25037 2620 25084 2622
rect 25148 2620 25154 2684
rect 25037 2619 25103 2620
rect 22645 2548 22711 2549
rect 22645 2546 22692 2548
rect 22600 2544 22692 2546
rect 22600 2488 22650 2544
rect 22600 2486 22692 2488
rect 22645 2484 22692 2486
rect 22756 2484 22762 2548
rect 22645 2483 22711 2484
rect 9765 2276 9831 2277
rect 13905 2276 13971 2277
rect 16297 2276 16363 2277
rect 22093 2276 22159 2277
rect 9765 2272 9801 2276
rect 9865 2274 9871 2276
rect 9765 2216 9770 2272
rect 9765 2212 9801 2216
rect 9865 2214 9922 2274
rect 13905 2272 13968 2276
rect 13905 2216 13910 2272
rect 13966 2216 13968 2272
rect 9865 2212 9871 2214
rect 13905 2212 13968 2216
rect 14032 2274 14038 2276
rect 14032 2214 14062 2274
rect 16297 2272 16304 2276
rect 16368 2274 16374 2276
rect 16297 2216 16302 2272
rect 14032 2212 14038 2214
rect 16297 2212 16304 2216
rect 16368 2214 16454 2274
rect 22093 2272 22144 2276
rect 22208 2274 22214 2276
rect 24117 2274 24183 2277
rect 32673 2276 32739 2277
rect 36169 2276 36235 2277
rect 37457 2276 37523 2277
rect 51349 2276 51415 2277
rect 52545 2276 52611 2277
rect 24474 2274 24480 2276
rect 22093 2216 22098 2272
rect 16368 2212 16374 2214
rect 22093 2212 22144 2216
rect 22208 2214 22250 2274
rect 24117 2272 24480 2274
rect 24117 2216 24122 2272
rect 24178 2216 24480 2272
rect 24117 2214 24480 2216
rect 22208 2212 22214 2214
rect 9765 2211 9831 2212
rect 13905 2211 13971 2212
rect 16297 2211 16363 2212
rect 22093 2211 22159 2212
rect 24117 2211 24183 2214
rect 24474 2212 24480 2214
rect 24544 2212 24550 2276
rect 32650 2212 32656 2276
rect 32720 2274 32739 2276
rect 32720 2272 32812 2274
rect 32734 2216 32812 2272
rect 32720 2214 32812 2216
rect 32720 2212 32739 2214
rect 36154 2212 36160 2276
rect 36224 2274 36235 2276
rect 36224 2272 36316 2274
rect 36230 2216 36316 2272
rect 36224 2214 36316 2216
rect 36224 2212 36235 2214
rect 37446 2212 37452 2276
rect 37516 2274 37523 2276
rect 37516 2272 37608 2274
rect 37518 2216 37608 2272
rect 37516 2214 37608 2216
rect 37516 2212 37523 2214
rect 51338 2212 51344 2276
rect 51408 2274 51415 2276
rect 52506 2274 52512 2276
rect 51408 2272 51500 2274
rect 51410 2216 51500 2272
rect 51408 2214 51500 2216
rect 52454 2214 52512 2274
rect 52576 2272 52611 2276
rect 52606 2216 52611 2272
rect 51408 2212 51415 2214
rect 52506 2212 52512 2214
rect 52576 2212 52611 2216
rect 32673 2211 32739 2212
rect 36169 2211 36235 2212
rect 37457 2211 37523 2212
rect 51349 2211 51415 2212
rect 52545 2211 52611 2212
rect 1944 2208 2264 2209
rect 1944 2144 1952 2208
rect 2016 2144 2032 2208
rect 2096 2144 2112 2208
rect 2176 2144 2192 2208
rect 2256 2144 2264 2208
rect 1944 2143 2264 2144
rect 85944 2208 86264 2209
rect 85944 2144 85952 2208
rect 86016 2144 86032 2208
rect 86096 2144 86112 2208
rect 86176 2144 86192 2208
rect 86256 2144 86264 2208
rect 85944 2143 86264 2144
rect 89944 2208 90264 2209
rect 89944 2144 89952 2208
rect 90016 2144 90032 2208
rect 90096 2144 90112 2208
rect 90176 2144 90192 2208
rect 90256 2144 90264 2208
rect 89944 2143 90264 2144
rect 32765 2140 32831 2141
rect 33961 2140 34027 2141
rect 32765 2138 32780 2140
rect 32688 2136 32780 2138
rect 32688 2080 32770 2136
rect 32688 2078 32780 2080
rect 32765 2076 32780 2078
rect 32844 2076 32850 2140
rect 33942 2076 33948 2140
rect 34012 2138 34027 2140
rect 36261 2140 36327 2141
rect 36261 2138 36284 2140
rect 34012 2136 34104 2138
rect 34022 2080 34104 2136
rect 34012 2078 34104 2080
rect 36192 2136 36284 2138
rect 36192 2080 36266 2136
rect 36192 2078 36284 2080
rect 34012 2076 34027 2078
rect 32765 2075 32831 2076
rect 33961 2075 34027 2076
rect 36261 2076 36284 2078
rect 36348 2076 36354 2140
rect 36261 2075 36327 2076
rect 29085 2004 29151 2005
rect 30465 2004 30531 2005
rect 31661 2004 31727 2005
rect 29085 2002 29152 2004
rect 29060 2000 29152 2002
rect 29060 1944 29090 2000
rect 29146 1944 29152 2000
rect 29060 1942 29152 1944
rect 29085 1940 29152 1942
rect 29216 1940 29222 2004
rect 30438 1940 30444 2004
rect 30508 2002 30531 2004
rect 31606 2002 31612 2004
rect 30508 2000 30600 2002
rect 30526 1944 30600 2000
rect 30508 1942 30600 1944
rect 31570 1942 31612 2002
rect 31676 2000 31727 2004
rect 31722 1944 31727 2000
rect 30508 1940 30531 1942
rect 31606 1940 31612 1942
rect 31676 1940 31727 1944
rect 29085 1939 29151 1940
rect 30465 1939 30531 1940
rect 31661 1939 31727 1940
rect 17493 1868 17559 1869
rect 17466 1866 17472 1868
rect 17402 1806 17472 1866
rect 17536 1864 17559 1868
rect 21081 1868 21147 1869
rect 22277 1868 22343 1869
rect 25773 1868 25839 1869
rect 26969 1868 27035 1869
rect 28165 1868 28231 1869
rect 21081 1866 21100 1868
rect 17554 1808 17559 1864
rect 17466 1804 17472 1806
rect 17536 1804 17559 1808
rect 21008 1864 21100 1866
rect 21008 1808 21086 1864
rect 21008 1806 21100 1808
rect 17493 1803 17559 1804
rect 21081 1804 21100 1806
rect 21164 1804 21170 1868
rect 22262 1804 22268 1868
rect 22332 1866 22343 1868
rect 22332 1864 22424 1866
rect 22338 1808 22424 1864
rect 22332 1806 22424 1808
rect 22332 1804 22343 1806
rect 25766 1804 25772 1868
rect 25836 1866 25842 1868
rect 25836 1806 25928 1866
rect 25836 1804 25842 1806
rect 26934 1804 26940 1868
rect 27004 1866 27035 1868
rect 27004 1864 27096 1866
rect 27030 1808 27096 1864
rect 27004 1806 27096 1808
rect 27004 1804 27035 1806
rect 28102 1804 28108 1868
rect 28172 1866 28231 1868
rect 28172 1864 28264 1866
rect 28226 1808 28264 1864
rect 28172 1806 28264 1808
rect 28172 1804 28231 1806
rect 21081 1803 21147 1804
rect 22277 1803 22343 1804
rect 25773 1803 25839 1804
rect 26969 1803 27035 1804
rect 28165 1803 28231 1804
rect 86861 1730 86927 1733
rect 91200 1730 92000 1760
rect 86861 1728 92000 1730
rect 86861 1672 86866 1728
rect 86922 1672 92000 1728
rect 86861 1670 92000 1672
rect 86861 1667 86927 1670
rect 91200 1640 92000 1670
rect 48998 1532 49004 1596
rect 49068 1594 49074 1596
rect 83549 1594 83615 1597
rect 49068 1592 83615 1594
rect 49068 1536 83554 1592
rect 83610 1536 83615 1592
rect 49068 1534 83615 1536
rect 49068 1532 49074 1534
rect 83549 1531 83615 1534
rect 9765 1458 9831 1461
rect 83406 1458 83412 1460
rect 9765 1456 83412 1458
rect 9765 1400 9770 1456
rect 9826 1400 83412 1456
rect 9765 1398 83412 1400
rect 9765 1395 9831 1398
rect 83406 1396 83412 1398
rect 83476 1396 83482 1460
rect 12433 1322 12499 1325
rect 12750 1322 12756 1324
rect 12433 1320 12756 1322
rect 12433 1264 12438 1320
rect 12494 1264 12756 1320
rect 12433 1262 12756 1264
rect 12433 1259 12499 1262
rect 12750 1260 12756 1262
rect 12820 1260 12826 1324
rect 18822 1260 18828 1324
rect 18892 1322 18898 1324
rect 19241 1322 19307 1325
rect 18892 1320 19307 1322
rect 18892 1264 19246 1320
rect 19302 1264 19307 1320
rect 18892 1262 19307 1264
rect 18892 1260 18898 1262
rect 19241 1259 19307 1262
rect 29310 1260 29316 1324
rect 29380 1322 29386 1324
rect 30281 1322 30347 1325
rect 29380 1320 30347 1322
rect 29380 1264 30286 1320
rect 30342 1264 30347 1320
rect 29380 1262 30347 1264
rect 29380 1260 29386 1262
rect 30281 1259 30347 1262
rect 35198 1260 35204 1324
rect 35268 1322 35274 1324
rect 35525 1322 35591 1325
rect 35268 1320 35591 1322
rect 35268 1264 35530 1320
rect 35586 1264 35591 1320
rect 35268 1262 35591 1264
rect 35268 1260 35274 1262
rect 35525 1259 35591 1262
rect 39246 1260 39252 1324
rect 39316 1322 39322 1324
rect 39849 1322 39915 1325
rect 39316 1320 39915 1322
rect 39316 1264 39854 1320
rect 39910 1264 39915 1320
rect 39316 1262 39915 1264
rect 39316 1260 39322 1262
rect 39849 1259 39915 1262
rect 44766 1260 44772 1324
rect 44836 1322 44842 1324
rect 44909 1322 44975 1325
rect 44836 1320 44975 1322
rect 44836 1264 44914 1320
rect 44970 1264 44975 1320
rect 44836 1262 44975 1264
rect 44836 1260 44842 1262
rect 44909 1259 44975 1262
rect 48078 1260 48084 1324
rect 48148 1322 48154 1324
rect 48221 1322 48287 1325
rect 48148 1320 48287 1322
rect 48148 1264 48226 1320
rect 48282 1264 48287 1320
rect 48148 1262 48287 1264
rect 48148 1260 48154 1262
rect 48221 1259 48287 1262
rect 17953 1186 18019 1189
rect 18638 1186 18644 1188
rect 17953 1184 18644 1186
rect 17953 1128 17958 1184
rect 18014 1128 18644 1184
rect 17953 1126 18644 1128
rect 17953 1123 18019 1126
rect 18638 1124 18644 1126
rect 18708 1124 18714 1188
rect 19333 1186 19399 1189
rect 19742 1186 19748 1188
rect 19333 1184 19748 1186
rect 19333 1128 19338 1184
rect 19394 1128 19748 1184
rect 19333 1126 19748 1128
rect 19333 1123 19399 1126
rect 19742 1124 19748 1126
rect 19812 1124 19818 1188
rect 28993 1186 29059 1189
rect 29678 1186 29684 1188
rect 28993 1184 29684 1186
rect 28993 1128 28998 1184
rect 29054 1128 29684 1184
rect 28993 1126 29684 1128
rect 28993 1123 29059 1126
rect 29678 1124 29684 1126
rect 29748 1124 29754 1188
rect 34513 1186 34579 1189
rect 34830 1186 34836 1188
rect 34513 1184 34836 1186
rect 34513 1128 34518 1184
rect 34574 1128 34836 1184
rect 34513 1126 34836 1128
rect 34513 1123 34579 1126
rect 34830 1124 34836 1126
rect 34900 1124 34906 1188
rect 39798 1124 39804 1188
rect 39868 1186 39874 1188
rect 39941 1186 40007 1189
rect 39868 1184 40007 1186
rect 39868 1128 39946 1184
rect 40002 1128 40007 1184
rect 39868 1126 40007 1128
rect 39868 1124 39874 1126
rect 39941 1123 40007 1126
rect 52126 1124 52132 1188
rect 52196 1186 52202 1188
rect 52361 1186 52427 1189
rect 52196 1184 52427 1186
rect 52196 1128 52366 1184
rect 52422 1128 52427 1184
rect 52196 1126 52427 1128
rect 52196 1124 52202 1126
rect 52361 1123 52427 1126
rect 24761 1052 24827 1053
rect 24710 988 24716 1052
rect 24780 1050 24827 1052
rect 30373 1050 30439 1053
rect 41321 1052 41387 1053
rect 30966 1050 30972 1052
rect 24780 1048 24872 1050
rect 24822 992 24872 1048
rect 24780 990 24872 992
rect 30373 1048 30972 1050
rect 30373 992 30378 1048
rect 30434 992 30972 1048
rect 30373 990 30972 992
rect 24780 988 24827 990
rect 24761 987 24827 988
rect 30373 987 30439 990
rect 30966 988 30972 990
rect 31036 988 31042 1052
rect 41270 988 41276 1052
rect 41340 1050 41387 1052
rect 41340 1048 41432 1050
rect 41382 992 41432 1048
rect 41340 990 41432 992
rect 41340 988 41387 990
rect 42558 988 42564 1052
rect 42628 1050 42634 1052
rect 42701 1050 42767 1053
rect 42628 1048 42767 1050
rect 42628 992 42706 1048
rect 42762 992 42767 1048
rect 42628 990 42767 992
rect 42628 988 42634 990
rect 41321 987 41387 988
rect 42701 987 42767 990
rect 45686 988 45692 1052
rect 45756 1050 45762 1052
rect 46749 1050 46815 1053
rect 45756 1048 46815 1050
rect 45756 992 46754 1048
rect 46810 992 46815 1048
rect 45756 990 46815 992
rect 45756 988 45762 990
rect 46749 987 46815 990
rect 49182 988 49188 1052
rect 49252 1050 49258 1052
rect 49601 1050 49667 1053
rect 49252 1048 49667 1050
rect 49252 992 49606 1048
rect 49662 992 49667 1048
rect 49252 990 49667 992
rect 49252 988 49258 990
rect 49601 987 49667 990
rect 53782 988 53788 1052
rect 53852 1050 53858 1052
rect 54661 1050 54727 1053
rect 53852 1048 54727 1050
rect 53852 992 54666 1048
rect 54722 992 54727 1048
rect 53852 990 54727 992
rect 53852 988 53858 990
rect 54661 987 54727 990
rect 27613 916 27679 917
rect 27613 914 27660 916
rect 27568 912 27660 914
rect 27568 856 27618 912
rect 27568 854 27660 856
rect 27613 852 27660 854
rect 27724 852 27730 916
rect 42793 914 42859 917
rect 43110 914 43116 916
rect 42793 912 43116 914
rect 42793 856 42798 912
rect 42854 856 43116 912
rect 42793 854 43116 856
rect 27613 851 27679 852
rect 42793 851 42859 854
rect 43110 852 43116 854
rect 43180 852 43186 916
rect 43294 852 43300 916
rect 43364 914 43370 916
rect 44081 914 44147 917
rect 46841 916 46907 917
rect 43364 912 44147 914
rect 43364 856 44086 912
rect 44142 856 44147 912
rect 43364 854 44147 856
rect 43364 852 43370 854
rect 44081 851 44147 854
rect 46790 852 46796 916
rect 46860 914 46907 916
rect 46860 912 46952 914
rect 46902 856 46952 912
rect 46860 854 46952 856
rect 46860 852 46907 854
rect 46841 851 46907 852
rect 23422 716 23428 780
rect 23492 778 23498 780
rect 24761 778 24827 781
rect 23492 776 24827 778
rect 23492 720 24766 776
rect 24822 720 24827 776
rect 23492 718 24827 720
rect 23492 716 23498 718
rect 24761 715 24827 718
rect 33133 778 33199 781
rect 33726 778 33732 780
rect 33133 776 33732 778
rect 33133 720 33138 776
rect 33194 720 33732 776
rect 33133 718 33732 720
rect 33133 715 33199 718
rect 33726 716 33732 718
rect 33796 716 33802 780
rect 50286 716 50292 780
rect 50356 778 50362 780
rect 50981 778 51047 781
rect 50356 776 51047 778
rect 50356 720 50986 776
rect 51042 720 51047 776
rect 50356 718 51047 720
rect 50356 716 50362 718
rect 50981 715 51047 718
rect 54702 716 54708 780
rect 54772 778 54778 780
rect 55029 778 55095 781
rect 54772 776 55095 778
rect 54772 720 55034 776
rect 55090 720 55095 776
rect 54772 718 55095 720
rect 54772 716 54778 718
rect 55029 715 55095 718
rect 86953 642 87019 645
rect 91200 642 92000 672
rect 86953 640 92000 642
rect 86953 584 86958 640
rect 87014 584 92000 640
rect 86953 582 92000 584
rect 86953 579 87019 582
rect 91200 552 92000 582
rect 52678 444 52684 508
rect 52748 506 52754 508
rect 53741 506 53807 509
rect 55121 508 55187 509
rect 55070 506 55076 508
rect 52748 504 53807 506
rect 52748 448 53746 504
rect 53802 448 53807 504
rect 52748 446 53807 448
rect 55030 446 55076 506
rect 55140 504 55187 508
rect 55182 448 55187 504
rect 52748 444 52754 446
rect 53741 443 53807 446
rect 55070 444 55076 446
rect 55140 444 55187 448
rect 55121 443 55187 444
rect 19926 172 19932 236
rect 19996 234 20002 236
rect 20621 234 20687 237
rect 19996 232 20687 234
rect 19996 176 20626 232
rect 20682 176 20687 232
rect 19996 174 20687 176
rect 19996 172 20002 174
rect 20621 171 20687 174
<< via3 >>
rect 89300 191388 89364 191452
rect 88932 190164 88996 190228
rect 1952 189340 2016 189344
rect 1952 189284 1956 189340
rect 1956 189284 2012 189340
rect 2012 189284 2016 189340
rect 1952 189280 2016 189284
rect 2032 189340 2096 189344
rect 2032 189284 2036 189340
rect 2036 189284 2092 189340
rect 2092 189284 2096 189340
rect 2032 189280 2096 189284
rect 2112 189340 2176 189344
rect 2112 189284 2116 189340
rect 2116 189284 2172 189340
rect 2172 189284 2176 189340
rect 2112 189280 2176 189284
rect 2192 189340 2256 189344
rect 2192 189284 2196 189340
rect 2196 189284 2252 189340
rect 2252 189284 2256 189340
rect 2192 189280 2256 189284
rect 85952 189340 86016 189344
rect 85952 189284 85956 189340
rect 85956 189284 86012 189340
rect 86012 189284 86016 189340
rect 85952 189280 86016 189284
rect 86032 189340 86096 189344
rect 86032 189284 86036 189340
rect 86036 189284 86092 189340
rect 86092 189284 86096 189340
rect 86032 189280 86096 189284
rect 86112 189340 86176 189344
rect 86112 189284 86116 189340
rect 86116 189284 86172 189340
rect 86172 189284 86176 189340
rect 86112 189280 86176 189284
rect 86192 189340 86256 189344
rect 86192 189284 86196 189340
rect 86196 189284 86252 189340
rect 86252 189284 86256 189340
rect 86192 189280 86256 189284
rect 89952 189340 90016 189344
rect 89952 189284 89956 189340
rect 89956 189284 90012 189340
rect 90012 189284 90016 189340
rect 89952 189280 90016 189284
rect 90032 189340 90096 189344
rect 90032 189284 90036 189340
rect 90036 189284 90092 189340
rect 90092 189284 90096 189340
rect 90032 189280 90096 189284
rect 90112 189340 90176 189344
rect 90112 189284 90116 189340
rect 90116 189284 90172 189340
rect 90172 189284 90176 189340
rect 90112 189280 90176 189284
rect 90192 189340 90256 189344
rect 90192 189284 90196 189340
rect 90196 189284 90252 189340
rect 90252 189284 90256 189340
rect 90192 189280 90256 189284
rect 75132 189076 75196 189140
rect 89116 188940 89180 189004
rect 3952 188796 4016 188800
rect 3952 188740 3956 188796
rect 3956 188740 4012 188796
rect 4012 188740 4016 188796
rect 3952 188736 4016 188740
rect 4032 188796 4096 188800
rect 4032 188740 4036 188796
rect 4036 188740 4092 188796
rect 4092 188740 4096 188796
rect 4032 188736 4096 188740
rect 4112 188796 4176 188800
rect 4112 188740 4116 188796
rect 4116 188740 4172 188796
rect 4172 188740 4176 188796
rect 4112 188736 4176 188740
rect 4192 188796 4256 188800
rect 4192 188740 4196 188796
rect 4196 188740 4252 188796
rect 4252 188740 4256 188796
rect 4192 188736 4256 188740
rect 87952 188796 88016 188800
rect 87952 188740 87956 188796
rect 87956 188740 88012 188796
rect 88012 188740 88016 188796
rect 87952 188736 88016 188740
rect 88032 188796 88096 188800
rect 88032 188740 88036 188796
rect 88036 188740 88092 188796
rect 88092 188740 88096 188796
rect 88032 188736 88096 188740
rect 88112 188796 88176 188800
rect 88112 188740 88116 188796
rect 88116 188740 88172 188796
rect 88172 188740 88176 188796
rect 88112 188736 88176 188740
rect 88192 188796 88256 188800
rect 88192 188740 88196 188796
rect 88196 188740 88252 188796
rect 88252 188740 88256 188796
rect 88192 188736 88256 188740
rect 1952 188252 2016 188256
rect 1952 188196 1956 188252
rect 1956 188196 2012 188252
rect 2012 188196 2016 188252
rect 1952 188192 2016 188196
rect 2032 188252 2096 188256
rect 2032 188196 2036 188252
rect 2036 188196 2092 188252
rect 2092 188196 2096 188252
rect 2032 188192 2096 188196
rect 2112 188252 2176 188256
rect 2112 188196 2116 188252
rect 2116 188196 2172 188252
rect 2172 188196 2176 188252
rect 2112 188192 2176 188196
rect 2192 188252 2256 188256
rect 2192 188196 2196 188252
rect 2196 188196 2252 188252
rect 2252 188196 2256 188252
rect 2192 188192 2256 188196
rect 85952 188252 86016 188256
rect 85952 188196 85956 188252
rect 85956 188196 86012 188252
rect 86012 188196 86016 188252
rect 85952 188192 86016 188196
rect 86032 188252 86096 188256
rect 86032 188196 86036 188252
rect 86036 188196 86092 188252
rect 86092 188196 86096 188252
rect 86032 188192 86096 188196
rect 86112 188252 86176 188256
rect 86112 188196 86116 188252
rect 86116 188196 86172 188252
rect 86172 188196 86176 188252
rect 86112 188192 86176 188196
rect 86192 188252 86256 188256
rect 86192 188196 86196 188252
rect 86196 188196 86252 188252
rect 86252 188196 86256 188252
rect 86192 188192 86256 188196
rect 89952 188252 90016 188256
rect 89952 188196 89956 188252
rect 89956 188196 90012 188252
rect 90012 188196 90016 188252
rect 89952 188192 90016 188196
rect 90032 188252 90096 188256
rect 90032 188196 90036 188252
rect 90036 188196 90092 188252
rect 90092 188196 90096 188252
rect 90032 188192 90096 188196
rect 90112 188252 90176 188256
rect 90112 188196 90116 188252
rect 90116 188196 90172 188252
rect 90172 188196 90176 188252
rect 90112 188192 90176 188196
rect 90192 188252 90256 188256
rect 90192 188196 90196 188252
rect 90196 188196 90252 188252
rect 90252 188196 90256 188252
rect 90192 188192 90256 188196
rect 89484 187716 89548 187780
rect 3952 187708 4016 187712
rect 3952 187652 3956 187708
rect 3956 187652 4012 187708
rect 4012 187652 4016 187708
rect 3952 187648 4016 187652
rect 4032 187708 4096 187712
rect 4032 187652 4036 187708
rect 4036 187652 4092 187708
rect 4092 187652 4096 187708
rect 4032 187648 4096 187652
rect 4112 187708 4176 187712
rect 4112 187652 4116 187708
rect 4116 187652 4172 187708
rect 4172 187652 4176 187708
rect 4112 187648 4176 187652
rect 4192 187708 4256 187712
rect 4192 187652 4196 187708
rect 4196 187652 4252 187708
rect 4252 187652 4256 187708
rect 4192 187648 4256 187652
rect 87952 187708 88016 187712
rect 87952 187652 87956 187708
rect 87956 187652 88012 187708
rect 88012 187652 88016 187708
rect 87952 187648 88016 187652
rect 88032 187708 88096 187712
rect 88032 187652 88036 187708
rect 88036 187652 88092 187708
rect 88092 187652 88096 187708
rect 88032 187648 88096 187652
rect 88112 187708 88176 187712
rect 88112 187652 88116 187708
rect 88116 187652 88172 187708
rect 88172 187652 88176 187708
rect 88112 187648 88176 187652
rect 88192 187708 88256 187712
rect 88192 187652 88196 187708
rect 88196 187652 88252 187708
rect 88252 187652 88256 187708
rect 88192 187648 88256 187652
rect 1952 187164 2016 187168
rect 1952 187108 1956 187164
rect 1956 187108 2012 187164
rect 2012 187108 2016 187164
rect 1952 187104 2016 187108
rect 2032 187164 2096 187168
rect 2032 187108 2036 187164
rect 2036 187108 2092 187164
rect 2092 187108 2096 187164
rect 2032 187104 2096 187108
rect 2112 187164 2176 187168
rect 2112 187108 2116 187164
rect 2116 187108 2172 187164
rect 2172 187108 2176 187164
rect 2112 187104 2176 187108
rect 2192 187164 2256 187168
rect 2192 187108 2196 187164
rect 2196 187108 2252 187164
rect 2252 187108 2256 187164
rect 2192 187104 2256 187108
rect 85952 187164 86016 187168
rect 85952 187108 85956 187164
rect 85956 187108 86012 187164
rect 86012 187108 86016 187164
rect 85952 187104 86016 187108
rect 86032 187164 86096 187168
rect 86032 187108 86036 187164
rect 86036 187108 86092 187164
rect 86092 187108 86096 187164
rect 86032 187104 86096 187108
rect 86112 187164 86176 187168
rect 86112 187108 86116 187164
rect 86116 187108 86172 187164
rect 86172 187108 86176 187164
rect 86112 187104 86176 187108
rect 86192 187164 86256 187168
rect 86192 187108 86196 187164
rect 86196 187108 86252 187164
rect 86252 187108 86256 187164
rect 86192 187104 86256 187108
rect 89952 187164 90016 187168
rect 89952 187108 89956 187164
rect 89956 187108 90012 187164
rect 90012 187108 90016 187164
rect 89952 187104 90016 187108
rect 90032 187164 90096 187168
rect 90032 187108 90036 187164
rect 90036 187108 90092 187164
rect 90092 187108 90096 187164
rect 90032 187104 90096 187108
rect 90112 187164 90176 187168
rect 90112 187108 90116 187164
rect 90116 187108 90172 187164
rect 90172 187108 90176 187164
rect 90112 187104 90176 187108
rect 90192 187164 90256 187168
rect 90192 187108 90196 187164
rect 90196 187108 90252 187164
rect 90252 187108 90256 187164
rect 90192 187104 90256 187108
rect 79364 187096 79428 187100
rect 79364 187040 79378 187096
rect 79378 187040 79428 187096
rect 79364 187036 79428 187040
rect 3952 186620 4016 186624
rect 3952 186564 3956 186620
rect 3956 186564 4012 186620
rect 4012 186564 4016 186620
rect 3952 186560 4016 186564
rect 4032 186620 4096 186624
rect 4032 186564 4036 186620
rect 4036 186564 4092 186620
rect 4092 186564 4096 186620
rect 4032 186560 4096 186564
rect 4112 186620 4176 186624
rect 4112 186564 4116 186620
rect 4116 186564 4172 186620
rect 4172 186564 4176 186620
rect 4112 186560 4176 186564
rect 4192 186620 4256 186624
rect 4192 186564 4196 186620
rect 4196 186564 4252 186620
rect 4252 186564 4256 186620
rect 4192 186560 4256 186564
rect 87952 186620 88016 186624
rect 87952 186564 87956 186620
rect 87956 186564 88012 186620
rect 88012 186564 88016 186620
rect 87952 186560 88016 186564
rect 88032 186620 88096 186624
rect 88032 186564 88036 186620
rect 88036 186564 88092 186620
rect 88092 186564 88096 186620
rect 88032 186560 88096 186564
rect 88112 186620 88176 186624
rect 88112 186564 88116 186620
rect 88116 186564 88172 186620
rect 88172 186564 88176 186620
rect 88112 186560 88176 186564
rect 88192 186620 88256 186624
rect 88192 186564 88196 186620
rect 88196 186564 88252 186620
rect 88252 186564 88256 186620
rect 88192 186560 88256 186564
rect 88748 186492 88812 186556
rect 1952 186076 2016 186080
rect 1952 186020 1956 186076
rect 1956 186020 2012 186076
rect 2012 186020 2016 186076
rect 1952 186016 2016 186020
rect 2032 186076 2096 186080
rect 2032 186020 2036 186076
rect 2036 186020 2092 186076
rect 2092 186020 2096 186076
rect 2032 186016 2096 186020
rect 2112 186076 2176 186080
rect 2112 186020 2116 186076
rect 2116 186020 2172 186076
rect 2172 186020 2176 186076
rect 2112 186016 2176 186020
rect 2192 186076 2256 186080
rect 2192 186020 2196 186076
rect 2196 186020 2252 186076
rect 2252 186020 2256 186076
rect 2192 186016 2256 186020
rect 85952 186076 86016 186080
rect 85952 186020 85956 186076
rect 85956 186020 86012 186076
rect 86012 186020 86016 186076
rect 85952 186016 86016 186020
rect 86032 186076 86096 186080
rect 86032 186020 86036 186076
rect 86036 186020 86092 186076
rect 86092 186020 86096 186076
rect 86032 186016 86096 186020
rect 86112 186076 86176 186080
rect 86112 186020 86116 186076
rect 86116 186020 86172 186076
rect 86172 186020 86176 186076
rect 86112 186016 86176 186020
rect 86192 186076 86256 186080
rect 86192 186020 86196 186076
rect 86196 186020 86252 186076
rect 86252 186020 86256 186076
rect 86192 186016 86256 186020
rect 89952 186076 90016 186080
rect 89952 186020 89956 186076
rect 89956 186020 90012 186076
rect 90012 186020 90016 186076
rect 89952 186016 90016 186020
rect 90032 186076 90096 186080
rect 90032 186020 90036 186076
rect 90036 186020 90092 186076
rect 90092 186020 90096 186076
rect 90032 186016 90096 186020
rect 90112 186076 90176 186080
rect 90112 186020 90116 186076
rect 90116 186020 90172 186076
rect 90172 186020 90176 186076
rect 90112 186016 90176 186020
rect 90192 186076 90256 186080
rect 90192 186020 90196 186076
rect 90196 186020 90252 186076
rect 90252 186020 90256 186076
rect 90192 186016 90256 186020
rect 3952 185532 4016 185536
rect 3952 185476 3956 185532
rect 3956 185476 4012 185532
rect 4012 185476 4016 185532
rect 3952 185472 4016 185476
rect 4032 185532 4096 185536
rect 4032 185476 4036 185532
rect 4036 185476 4092 185532
rect 4092 185476 4096 185532
rect 4032 185472 4096 185476
rect 4112 185532 4176 185536
rect 4112 185476 4116 185532
rect 4116 185476 4172 185532
rect 4172 185476 4176 185532
rect 4112 185472 4176 185476
rect 4192 185532 4256 185536
rect 4192 185476 4196 185532
rect 4196 185476 4252 185532
rect 4252 185476 4256 185532
rect 4192 185472 4256 185476
rect 87952 185532 88016 185536
rect 87952 185476 87956 185532
rect 87956 185476 88012 185532
rect 88012 185476 88016 185532
rect 87952 185472 88016 185476
rect 88032 185532 88096 185536
rect 88032 185476 88036 185532
rect 88036 185476 88092 185532
rect 88092 185476 88096 185532
rect 88032 185472 88096 185476
rect 88112 185532 88176 185536
rect 88112 185476 88116 185532
rect 88116 185476 88172 185532
rect 88172 185476 88176 185532
rect 88112 185472 88176 185476
rect 88192 185532 88256 185536
rect 88192 185476 88196 185532
rect 88196 185476 88252 185532
rect 88252 185476 88256 185532
rect 88192 185472 88256 185476
rect 88380 185268 88444 185332
rect 1952 184988 2016 184992
rect 1952 184932 1956 184988
rect 1956 184932 2012 184988
rect 2012 184932 2016 184988
rect 1952 184928 2016 184932
rect 2032 184988 2096 184992
rect 2032 184932 2036 184988
rect 2036 184932 2092 184988
rect 2092 184932 2096 184988
rect 2032 184928 2096 184932
rect 2112 184988 2176 184992
rect 2112 184932 2116 184988
rect 2116 184932 2172 184988
rect 2172 184932 2176 184988
rect 2112 184928 2176 184932
rect 2192 184988 2256 184992
rect 2192 184932 2196 184988
rect 2196 184932 2252 184988
rect 2252 184932 2256 184988
rect 2192 184928 2256 184932
rect 85952 184988 86016 184992
rect 85952 184932 85956 184988
rect 85956 184932 86012 184988
rect 86012 184932 86016 184988
rect 85952 184928 86016 184932
rect 86032 184988 86096 184992
rect 86032 184932 86036 184988
rect 86036 184932 86092 184988
rect 86092 184932 86096 184988
rect 86032 184928 86096 184932
rect 86112 184988 86176 184992
rect 86112 184932 86116 184988
rect 86116 184932 86172 184988
rect 86172 184932 86176 184988
rect 86112 184928 86176 184932
rect 86192 184988 86256 184992
rect 86192 184932 86196 184988
rect 86196 184932 86252 184988
rect 86252 184932 86256 184988
rect 86192 184928 86256 184932
rect 89952 184988 90016 184992
rect 89952 184932 89956 184988
rect 89956 184932 90012 184988
rect 90012 184932 90016 184988
rect 89952 184928 90016 184932
rect 90032 184988 90096 184992
rect 90032 184932 90036 184988
rect 90036 184932 90092 184988
rect 90092 184932 90096 184988
rect 90032 184928 90096 184932
rect 90112 184988 90176 184992
rect 90112 184932 90116 184988
rect 90116 184932 90172 184988
rect 90172 184932 90176 184988
rect 90112 184928 90176 184932
rect 90192 184988 90256 184992
rect 90192 184932 90196 184988
rect 90196 184932 90252 184988
rect 90252 184932 90256 184988
rect 90192 184928 90256 184932
rect 3952 184444 4016 184448
rect 3952 184388 3956 184444
rect 3956 184388 4012 184444
rect 4012 184388 4016 184444
rect 3952 184384 4016 184388
rect 4032 184444 4096 184448
rect 4032 184388 4036 184444
rect 4036 184388 4092 184444
rect 4092 184388 4096 184444
rect 4032 184384 4096 184388
rect 4112 184444 4176 184448
rect 4112 184388 4116 184444
rect 4116 184388 4172 184444
rect 4172 184388 4176 184444
rect 4112 184384 4176 184388
rect 4192 184444 4256 184448
rect 4192 184388 4196 184444
rect 4196 184388 4252 184444
rect 4252 184388 4256 184444
rect 4192 184384 4256 184388
rect 87952 184444 88016 184448
rect 87952 184388 87956 184444
rect 87956 184388 88012 184444
rect 88012 184388 88016 184444
rect 87952 184384 88016 184388
rect 88032 184444 88096 184448
rect 88032 184388 88036 184444
rect 88036 184388 88092 184444
rect 88092 184388 88096 184444
rect 88032 184384 88096 184388
rect 88112 184444 88176 184448
rect 88112 184388 88116 184444
rect 88116 184388 88172 184444
rect 88172 184388 88176 184444
rect 88112 184384 88176 184388
rect 88192 184444 88256 184448
rect 88192 184388 88196 184444
rect 88196 184388 88252 184444
rect 88252 184388 88256 184444
rect 88192 184384 88256 184388
rect 87460 184044 87524 184108
rect 1952 183900 2016 183904
rect 1952 183844 1956 183900
rect 1956 183844 2012 183900
rect 2012 183844 2016 183900
rect 1952 183840 2016 183844
rect 2032 183900 2096 183904
rect 2032 183844 2036 183900
rect 2036 183844 2092 183900
rect 2092 183844 2096 183900
rect 2032 183840 2096 183844
rect 2112 183900 2176 183904
rect 2112 183844 2116 183900
rect 2116 183844 2172 183900
rect 2172 183844 2176 183900
rect 2112 183840 2176 183844
rect 2192 183900 2256 183904
rect 2192 183844 2196 183900
rect 2196 183844 2252 183900
rect 2252 183844 2256 183900
rect 2192 183840 2256 183844
rect 85952 183900 86016 183904
rect 85952 183844 85956 183900
rect 85956 183844 86012 183900
rect 86012 183844 86016 183900
rect 85952 183840 86016 183844
rect 86032 183900 86096 183904
rect 86032 183844 86036 183900
rect 86036 183844 86092 183900
rect 86092 183844 86096 183900
rect 86032 183840 86096 183844
rect 86112 183900 86176 183904
rect 86112 183844 86116 183900
rect 86116 183844 86172 183900
rect 86172 183844 86176 183900
rect 86112 183840 86176 183844
rect 86192 183900 86256 183904
rect 86192 183844 86196 183900
rect 86196 183844 86252 183900
rect 86252 183844 86256 183900
rect 86192 183840 86256 183844
rect 89952 183900 90016 183904
rect 89952 183844 89956 183900
rect 89956 183844 90012 183900
rect 90012 183844 90016 183900
rect 89952 183840 90016 183844
rect 90032 183900 90096 183904
rect 90032 183844 90036 183900
rect 90036 183844 90092 183900
rect 90092 183844 90096 183900
rect 90032 183840 90096 183844
rect 90112 183900 90176 183904
rect 90112 183844 90116 183900
rect 90116 183844 90172 183900
rect 90172 183844 90176 183900
rect 90112 183840 90176 183844
rect 90192 183900 90256 183904
rect 90192 183844 90196 183900
rect 90196 183844 90252 183900
rect 90252 183844 90256 183900
rect 90192 183840 90256 183844
rect 3952 183356 4016 183360
rect 3952 183300 3956 183356
rect 3956 183300 4012 183356
rect 4012 183300 4016 183356
rect 3952 183296 4016 183300
rect 4032 183356 4096 183360
rect 4032 183300 4036 183356
rect 4036 183300 4092 183356
rect 4092 183300 4096 183356
rect 4032 183296 4096 183300
rect 4112 183356 4176 183360
rect 4112 183300 4116 183356
rect 4116 183300 4172 183356
rect 4172 183300 4176 183356
rect 4112 183296 4176 183300
rect 4192 183356 4256 183360
rect 4192 183300 4196 183356
rect 4196 183300 4252 183356
rect 4252 183300 4256 183356
rect 4192 183296 4256 183300
rect 87952 183356 88016 183360
rect 87952 183300 87956 183356
rect 87956 183300 88012 183356
rect 88012 183300 88016 183356
rect 87952 183296 88016 183300
rect 88032 183356 88096 183360
rect 88032 183300 88036 183356
rect 88036 183300 88092 183356
rect 88092 183300 88096 183356
rect 88032 183296 88096 183300
rect 88112 183356 88176 183360
rect 88112 183300 88116 183356
rect 88116 183300 88172 183356
rect 88172 183300 88176 183356
rect 88112 183296 88176 183300
rect 88192 183356 88256 183360
rect 88192 183300 88196 183356
rect 88196 183300 88252 183356
rect 88252 183300 88256 183356
rect 88192 183296 88256 183300
rect 1952 182812 2016 182816
rect 1952 182756 1956 182812
rect 1956 182756 2012 182812
rect 2012 182756 2016 182812
rect 1952 182752 2016 182756
rect 2032 182812 2096 182816
rect 2032 182756 2036 182812
rect 2036 182756 2092 182812
rect 2092 182756 2096 182812
rect 2032 182752 2096 182756
rect 2112 182812 2176 182816
rect 2112 182756 2116 182812
rect 2116 182756 2172 182812
rect 2172 182756 2176 182812
rect 2112 182752 2176 182756
rect 2192 182812 2256 182816
rect 2192 182756 2196 182812
rect 2196 182756 2252 182812
rect 2252 182756 2256 182812
rect 2192 182752 2256 182756
rect 85952 182812 86016 182816
rect 85952 182756 85956 182812
rect 85956 182756 86012 182812
rect 86012 182756 86016 182812
rect 85952 182752 86016 182756
rect 86032 182812 86096 182816
rect 86032 182756 86036 182812
rect 86036 182756 86092 182812
rect 86092 182756 86096 182812
rect 86032 182752 86096 182756
rect 86112 182812 86176 182816
rect 86112 182756 86116 182812
rect 86116 182756 86172 182812
rect 86172 182756 86176 182812
rect 86112 182752 86176 182756
rect 86192 182812 86256 182816
rect 86192 182756 86196 182812
rect 86196 182756 86252 182812
rect 86252 182756 86256 182812
rect 86192 182752 86256 182756
rect 89952 182812 90016 182816
rect 89952 182756 89956 182812
rect 89956 182756 90012 182812
rect 90012 182756 90016 182812
rect 89952 182752 90016 182756
rect 90032 182812 90096 182816
rect 90032 182756 90036 182812
rect 90036 182756 90092 182812
rect 90092 182756 90096 182812
rect 90032 182752 90096 182756
rect 90112 182812 90176 182816
rect 90112 182756 90116 182812
rect 90116 182756 90172 182812
rect 90172 182756 90176 182812
rect 90112 182752 90176 182756
rect 90192 182812 90256 182816
rect 90192 182756 90196 182812
rect 90196 182756 90252 182812
rect 90252 182756 90256 182812
rect 90192 182752 90256 182756
rect 87092 182548 87156 182612
rect 3952 182268 4016 182272
rect 3952 182212 3956 182268
rect 3956 182212 4012 182268
rect 4012 182212 4016 182268
rect 3952 182208 4016 182212
rect 4032 182268 4096 182272
rect 4032 182212 4036 182268
rect 4036 182212 4092 182268
rect 4092 182212 4096 182268
rect 4032 182208 4096 182212
rect 4112 182268 4176 182272
rect 4112 182212 4116 182268
rect 4116 182212 4172 182268
rect 4172 182212 4176 182268
rect 4112 182208 4176 182212
rect 4192 182268 4256 182272
rect 4192 182212 4196 182268
rect 4196 182212 4252 182268
rect 4252 182212 4256 182268
rect 4192 182208 4256 182212
rect 87952 182268 88016 182272
rect 87952 182212 87956 182268
rect 87956 182212 88012 182268
rect 88012 182212 88016 182268
rect 87952 182208 88016 182212
rect 88032 182268 88096 182272
rect 88032 182212 88036 182268
rect 88036 182212 88092 182268
rect 88092 182212 88096 182268
rect 88032 182208 88096 182212
rect 88112 182268 88176 182272
rect 88112 182212 88116 182268
rect 88116 182212 88172 182268
rect 88172 182212 88176 182268
rect 88112 182208 88176 182212
rect 88192 182268 88256 182272
rect 88192 182212 88196 182268
rect 88196 182212 88252 182268
rect 88252 182212 88256 182268
rect 88192 182208 88256 182212
rect 1952 181724 2016 181728
rect 1952 181668 1956 181724
rect 1956 181668 2012 181724
rect 2012 181668 2016 181724
rect 1952 181664 2016 181668
rect 2032 181724 2096 181728
rect 2032 181668 2036 181724
rect 2036 181668 2092 181724
rect 2092 181668 2096 181724
rect 2032 181664 2096 181668
rect 2112 181724 2176 181728
rect 2112 181668 2116 181724
rect 2116 181668 2172 181724
rect 2172 181668 2176 181724
rect 2112 181664 2176 181668
rect 2192 181724 2256 181728
rect 2192 181668 2196 181724
rect 2196 181668 2252 181724
rect 2252 181668 2256 181724
rect 2192 181664 2256 181668
rect 85952 181724 86016 181728
rect 85952 181668 85956 181724
rect 85956 181668 86012 181724
rect 86012 181668 86016 181724
rect 85952 181664 86016 181668
rect 86032 181724 86096 181728
rect 86032 181668 86036 181724
rect 86036 181668 86092 181724
rect 86092 181668 86096 181724
rect 86032 181664 86096 181668
rect 86112 181724 86176 181728
rect 86112 181668 86116 181724
rect 86116 181668 86172 181724
rect 86172 181668 86176 181724
rect 86112 181664 86176 181668
rect 86192 181724 86256 181728
rect 86192 181668 86196 181724
rect 86196 181668 86252 181724
rect 86252 181668 86256 181724
rect 86192 181664 86256 181668
rect 89952 181724 90016 181728
rect 89952 181668 89956 181724
rect 89956 181668 90012 181724
rect 90012 181668 90016 181724
rect 89952 181664 90016 181668
rect 90032 181724 90096 181728
rect 90032 181668 90036 181724
rect 90036 181668 90092 181724
rect 90092 181668 90096 181724
rect 90032 181664 90096 181668
rect 90112 181724 90176 181728
rect 90112 181668 90116 181724
rect 90116 181668 90172 181724
rect 90172 181668 90176 181724
rect 90112 181664 90176 181668
rect 90192 181724 90256 181728
rect 90192 181668 90196 181724
rect 90196 181668 90252 181724
rect 90252 181668 90256 181724
rect 90192 181664 90256 181668
rect 3952 181180 4016 181184
rect 3952 181124 3956 181180
rect 3956 181124 4012 181180
rect 4012 181124 4016 181180
rect 3952 181120 4016 181124
rect 4032 181180 4096 181184
rect 4032 181124 4036 181180
rect 4036 181124 4092 181180
rect 4092 181124 4096 181180
rect 4032 181120 4096 181124
rect 4112 181180 4176 181184
rect 4112 181124 4116 181180
rect 4116 181124 4172 181180
rect 4172 181124 4176 181180
rect 4112 181120 4176 181124
rect 4192 181180 4256 181184
rect 4192 181124 4196 181180
rect 4196 181124 4252 181180
rect 4252 181124 4256 181180
rect 4192 181120 4256 181124
rect 87952 181180 88016 181184
rect 87952 181124 87956 181180
rect 87956 181124 88012 181180
rect 88012 181124 88016 181180
rect 87952 181120 88016 181124
rect 88032 181180 88096 181184
rect 88032 181124 88036 181180
rect 88036 181124 88092 181180
rect 88092 181124 88096 181180
rect 88032 181120 88096 181124
rect 88112 181180 88176 181184
rect 88112 181124 88116 181180
rect 88116 181124 88172 181180
rect 88172 181124 88176 181180
rect 88112 181120 88176 181124
rect 88192 181180 88256 181184
rect 88192 181124 88196 181180
rect 88196 181124 88252 181180
rect 88252 181124 88256 181180
rect 88192 181120 88256 181124
rect 1952 180636 2016 180640
rect 1952 180580 1956 180636
rect 1956 180580 2012 180636
rect 2012 180580 2016 180636
rect 1952 180576 2016 180580
rect 2032 180636 2096 180640
rect 2032 180580 2036 180636
rect 2036 180580 2092 180636
rect 2092 180580 2096 180636
rect 2032 180576 2096 180580
rect 2112 180636 2176 180640
rect 2112 180580 2116 180636
rect 2116 180580 2172 180636
rect 2172 180580 2176 180636
rect 2112 180576 2176 180580
rect 2192 180636 2256 180640
rect 2192 180580 2196 180636
rect 2196 180580 2252 180636
rect 2252 180580 2256 180636
rect 2192 180576 2256 180580
rect 85952 180636 86016 180640
rect 85952 180580 85956 180636
rect 85956 180580 86012 180636
rect 86012 180580 86016 180636
rect 85952 180576 86016 180580
rect 86032 180636 86096 180640
rect 86032 180580 86036 180636
rect 86036 180580 86092 180636
rect 86092 180580 86096 180636
rect 86032 180576 86096 180580
rect 86112 180636 86176 180640
rect 86112 180580 86116 180636
rect 86116 180580 86172 180636
rect 86172 180580 86176 180636
rect 86112 180576 86176 180580
rect 86192 180636 86256 180640
rect 86192 180580 86196 180636
rect 86196 180580 86252 180636
rect 86252 180580 86256 180636
rect 86192 180576 86256 180580
rect 89952 180636 90016 180640
rect 89952 180580 89956 180636
rect 89956 180580 90012 180636
rect 90012 180580 90016 180636
rect 89952 180576 90016 180580
rect 90032 180636 90096 180640
rect 90032 180580 90036 180636
rect 90036 180580 90092 180636
rect 90092 180580 90096 180636
rect 90032 180576 90096 180580
rect 90112 180636 90176 180640
rect 90112 180580 90116 180636
rect 90116 180580 90172 180636
rect 90172 180580 90176 180636
rect 90112 180576 90176 180580
rect 90192 180636 90256 180640
rect 90192 180580 90196 180636
rect 90196 180580 90252 180636
rect 90252 180580 90256 180636
rect 90192 180576 90256 180580
rect 87644 180372 87708 180436
rect 3952 180092 4016 180096
rect 3952 180036 3956 180092
rect 3956 180036 4012 180092
rect 4012 180036 4016 180092
rect 3952 180032 4016 180036
rect 4032 180092 4096 180096
rect 4032 180036 4036 180092
rect 4036 180036 4092 180092
rect 4092 180036 4096 180092
rect 4032 180032 4096 180036
rect 4112 180092 4176 180096
rect 4112 180036 4116 180092
rect 4116 180036 4172 180092
rect 4172 180036 4176 180092
rect 4112 180032 4176 180036
rect 4192 180092 4256 180096
rect 4192 180036 4196 180092
rect 4196 180036 4252 180092
rect 4252 180036 4256 180092
rect 4192 180032 4256 180036
rect 87952 180092 88016 180096
rect 87952 180036 87956 180092
rect 87956 180036 88012 180092
rect 88012 180036 88016 180092
rect 87952 180032 88016 180036
rect 88032 180092 88096 180096
rect 88032 180036 88036 180092
rect 88036 180036 88092 180092
rect 88092 180036 88096 180092
rect 88032 180032 88096 180036
rect 88112 180092 88176 180096
rect 88112 180036 88116 180092
rect 88116 180036 88172 180092
rect 88172 180036 88176 180092
rect 88112 180032 88176 180036
rect 88192 180092 88256 180096
rect 88192 180036 88196 180092
rect 88196 180036 88252 180092
rect 88252 180036 88256 180092
rect 88192 180032 88256 180036
rect 1952 179548 2016 179552
rect 1952 179492 1956 179548
rect 1956 179492 2012 179548
rect 2012 179492 2016 179548
rect 1952 179488 2016 179492
rect 2032 179548 2096 179552
rect 2032 179492 2036 179548
rect 2036 179492 2092 179548
rect 2092 179492 2096 179548
rect 2032 179488 2096 179492
rect 2112 179548 2176 179552
rect 2112 179492 2116 179548
rect 2116 179492 2172 179548
rect 2172 179492 2176 179548
rect 2112 179488 2176 179492
rect 2192 179548 2256 179552
rect 2192 179492 2196 179548
rect 2196 179492 2252 179548
rect 2252 179492 2256 179548
rect 2192 179488 2256 179492
rect 85952 179548 86016 179552
rect 85952 179492 85956 179548
rect 85956 179492 86012 179548
rect 86012 179492 86016 179548
rect 85952 179488 86016 179492
rect 86032 179548 86096 179552
rect 86032 179492 86036 179548
rect 86036 179492 86092 179548
rect 86092 179492 86096 179548
rect 86032 179488 86096 179492
rect 86112 179548 86176 179552
rect 86112 179492 86116 179548
rect 86116 179492 86172 179548
rect 86172 179492 86176 179548
rect 86112 179488 86176 179492
rect 86192 179548 86256 179552
rect 86192 179492 86196 179548
rect 86196 179492 86252 179548
rect 86252 179492 86256 179548
rect 86192 179488 86256 179492
rect 89952 179548 90016 179552
rect 89952 179492 89956 179548
rect 89956 179492 90012 179548
rect 90012 179492 90016 179548
rect 89952 179488 90016 179492
rect 90032 179548 90096 179552
rect 90032 179492 90036 179548
rect 90036 179492 90092 179548
rect 90092 179492 90096 179548
rect 90032 179488 90096 179492
rect 90112 179548 90176 179552
rect 90112 179492 90116 179548
rect 90116 179492 90172 179548
rect 90172 179492 90176 179548
rect 90112 179488 90176 179492
rect 90192 179548 90256 179552
rect 90192 179492 90196 179548
rect 90196 179492 90252 179548
rect 90252 179492 90256 179548
rect 90192 179488 90256 179492
rect 87276 179148 87340 179212
rect 3952 179004 4016 179008
rect 3952 178948 3956 179004
rect 3956 178948 4012 179004
rect 4012 178948 4016 179004
rect 3952 178944 4016 178948
rect 4032 179004 4096 179008
rect 4032 178948 4036 179004
rect 4036 178948 4092 179004
rect 4092 178948 4096 179004
rect 4032 178944 4096 178948
rect 4112 179004 4176 179008
rect 4112 178948 4116 179004
rect 4116 178948 4172 179004
rect 4172 178948 4176 179004
rect 4112 178944 4176 178948
rect 4192 179004 4256 179008
rect 4192 178948 4196 179004
rect 4196 178948 4252 179004
rect 4252 178948 4256 179004
rect 4192 178944 4256 178948
rect 87952 179004 88016 179008
rect 87952 178948 87956 179004
rect 87956 178948 88012 179004
rect 88012 178948 88016 179004
rect 87952 178944 88016 178948
rect 88032 179004 88096 179008
rect 88032 178948 88036 179004
rect 88036 178948 88092 179004
rect 88092 178948 88096 179004
rect 88032 178944 88096 178948
rect 88112 179004 88176 179008
rect 88112 178948 88116 179004
rect 88116 178948 88172 179004
rect 88172 178948 88176 179004
rect 88112 178944 88176 178948
rect 88192 179004 88256 179008
rect 88192 178948 88196 179004
rect 88196 178948 88252 179004
rect 88252 178948 88256 179004
rect 88192 178944 88256 178948
rect 1952 178460 2016 178464
rect 1952 178404 1956 178460
rect 1956 178404 2012 178460
rect 2012 178404 2016 178460
rect 1952 178400 2016 178404
rect 2032 178460 2096 178464
rect 2032 178404 2036 178460
rect 2036 178404 2092 178460
rect 2092 178404 2096 178460
rect 2032 178400 2096 178404
rect 2112 178460 2176 178464
rect 2112 178404 2116 178460
rect 2116 178404 2172 178460
rect 2172 178404 2176 178460
rect 2112 178400 2176 178404
rect 2192 178460 2256 178464
rect 2192 178404 2196 178460
rect 2196 178404 2252 178460
rect 2252 178404 2256 178460
rect 2192 178400 2256 178404
rect 85952 178460 86016 178464
rect 85952 178404 85956 178460
rect 85956 178404 86012 178460
rect 86012 178404 86016 178460
rect 85952 178400 86016 178404
rect 86032 178460 86096 178464
rect 86032 178404 86036 178460
rect 86036 178404 86092 178460
rect 86092 178404 86096 178460
rect 86032 178400 86096 178404
rect 86112 178460 86176 178464
rect 86112 178404 86116 178460
rect 86116 178404 86172 178460
rect 86172 178404 86176 178460
rect 86112 178400 86176 178404
rect 86192 178460 86256 178464
rect 86192 178404 86196 178460
rect 86196 178404 86252 178460
rect 86252 178404 86256 178460
rect 86192 178400 86256 178404
rect 89952 178460 90016 178464
rect 89952 178404 89956 178460
rect 89956 178404 90012 178460
rect 90012 178404 90016 178460
rect 89952 178400 90016 178404
rect 90032 178460 90096 178464
rect 90032 178404 90036 178460
rect 90036 178404 90092 178460
rect 90092 178404 90096 178460
rect 90032 178400 90096 178404
rect 90112 178460 90176 178464
rect 90112 178404 90116 178460
rect 90116 178404 90172 178460
rect 90172 178404 90176 178460
rect 90112 178400 90176 178404
rect 90192 178460 90256 178464
rect 90192 178404 90196 178460
rect 90196 178404 90252 178460
rect 90252 178404 90256 178460
rect 90192 178400 90256 178404
rect 3952 177916 4016 177920
rect 3952 177860 3956 177916
rect 3956 177860 4012 177916
rect 4012 177860 4016 177916
rect 3952 177856 4016 177860
rect 4032 177916 4096 177920
rect 4032 177860 4036 177916
rect 4036 177860 4092 177916
rect 4092 177860 4096 177916
rect 4032 177856 4096 177860
rect 4112 177916 4176 177920
rect 4112 177860 4116 177916
rect 4116 177860 4172 177916
rect 4172 177860 4176 177916
rect 4112 177856 4176 177860
rect 4192 177916 4256 177920
rect 4192 177860 4196 177916
rect 4196 177860 4252 177916
rect 4252 177860 4256 177916
rect 4192 177856 4256 177860
rect 87952 177916 88016 177920
rect 87952 177860 87956 177916
rect 87956 177860 88012 177916
rect 88012 177860 88016 177916
rect 87952 177856 88016 177860
rect 88032 177916 88096 177920
rect 88032 177860 88036 177916
rect 88036 177860 88092 177916
rect 88092 177860 88096 177916
rect 88032 177856 88096 177860
rect 88112 177916 88176 177920
rect 88112 177860 88116 177916
rect 88116 177860 88172 177916
rect 88172 177860 88176 177916
rect 88112 177856 88176 177860
rect 88192 177916 88256 177920
rect 88192 177860 88196 177916
rect 88196 177860 88252 177916
rect 88252 177860 88256 177916
rect 88192 177856 88256 177860
rect 1952 177372 2016 177376
rect 1952 177316 1956 177372
rect 1956 177316 2012 177372
rect 2012 177316 2016 177372
rect 1952 177312 2016 177316
rect 2032 177372 2096 177376
rect 2032 177316 2036 177372
rect 2036 177316 2092 177372
rect 2092 177316 2096 177372
rect 2032 177312 2096 177316
rect 2112 177372 2176 177376
rect 2112 177316 2116 177372
rect 2116 177316 2172 177372
rect 2172 177316 2176 177372
rect 2112 177312 2176 177316
rect 2192 177372 2256 177376
rect 2192 177316 2196 177372
rect 2196 177316 2252 177372
rect 2252 177316 2256 177372
rect 2192 177312 2256 177316
rect 85952 177372 86016 177376
rect 85952 177316 85956 177372
rect 85956 177316 86012 177372
rect 86012 177316 86016 177372
rect 85952 177312 86016 177316
rect 86032 177372 86096 177376
rect 86032 177316 86036 177372
rect 86036 177316 86092 177372
rect 86092 177316 86096 177372
rect 86032 177312 86096 177316
rect 86112 177372 86176 177376
rect 86112 177316 86116 177372
rect 86116 177316 86172 177372
rect 86172 177316 86176 177372
rect 86112 177312 86176 177316
rect 86192 177372 86256 177376
rect 86192 177316 86196 177372
rect 86196 177316 86252 177372
rect 86252 177316 86256 177372
rect 86192 177312 86256 177316
rect 89952 177372 90016 177376
rect 89952 177316 89956 177372
rect 89956 177316 90012 177372
rect 90012 177316 90016 177372
rect 89952 177312 90016 177316
rect 90032 177372 90096 177376
rect 90032 177316 90036 177372
rect 90036 177316 90092 177372
rect 90092 177316 90096 177372
rect 90032 177312 90096 177316
rect 90112 177372 90176 177376
rect 90112 177316 90116 177372
rect 90116 177316 90172 177372
rect 90172 177316 90176 177372
rect 90112 177312 90176 177316
rect 90192 177372 90256 177376
rect 90192 177316 90196 177372
rect 90196 177316 90252 177372
rect 90252 177316 90256 177372
rect 90192 177312 90256 177316
rect 83412 176972 83476 177036
rect 3952 176828 4016 176832
rect 3952 176772 3956 176828
rect 3956 176772 4012 176828
rect 4012 176772 4016 176828
rect 3952 176768 4016 176772
rect 4032 176828 4096 176832
rect 4032 176772 4036 176828
rect 4036 176772 4092 176828
rect 4092 176772 4096 176828
rect 4032 176768 4096 176772
rect 4112 176828 4176 176832
rect 4112 176772 4116 176828
rect 4116 176772 4172 176828
rect 4172 176772 4176 176828
rect 4112 176768 4176 176772
rect 4192 176828 4256 176832
rect 4192 176772 4196 176828
rect 4196 176772 4252 176828
rect 4252 176772 4256 176828
rect 4192 176768 4256 176772
rect 87952 176828 88016 176832
rect 87952 176772 87956 176828
rect 87956 176772 88012 176828
rect 88012 176772 88016 176828
rect 87952 176768 88016 176772
rect 88032 176828 88096 176832
rect 88032 176772 88036 176828
rect 88036 176772 88092 176828
rect 88092 176772 88096 176828
rect 88032 176768 88096 176772
rect 88112 176828 88176 176832
rect 88112 176772 88116 176828
rect 88116 176772 88172 176828
rect 88172 176772 88176 176828
rect 88112 176768 88176 176772
rect 88192 176828 88256 176832
rect 88192 176772 88196 176828
rect 88196 176772 88252 176828
rect 88252 176772 88256 176828
rect 88192 176768 88256 176772
rect 1952 176284 2016 176288
rect 1952 176228 1956 176284
rect 1956 176228 2012 176284
rect 2012 176228 2016 176284
rect 1952 176224 2016 176228
rect 2032 176284 2096 176288
rect 2032 176228 2036 176284
rect 2036 176228 2092 176284
rect 2092 176228 2096 176284
rect 2032 176224 2096 176228
rect 2112 176284 2176 176288
rect 2112 176228 2116 176284
rect 2116 176228 2172 176284
rect 2172 176228 2176 176284
rect 2112 176224 2176 176228
rect 2192 176284 2256 176288
rect 2192 176228 2196 176284
rect 2196 176228 2252 176284
rect 2252 176228 2256 176284
rect 2192 176224 2256 176228
rect 85952 176284 86016 176288
rect 85952 176228 85956 176284
rect 85956 176228 86012 176284
rect 86012 176228 86016 176284
rect 85952 176224 86016 176228
rect 86032 176284 86096 176288
rect 86032 176228 86036 176284
rect 86036 176228 86092 176284
rect 86092 176228 86096 176284
rect 86032 176224 86096 176228
rect 86112 176284 86176 176288
rect 86112 176228 86116 176284
rect 86116 176228 86172 176284
rect 86172 176228 86176 176284
rect 86112 176224 86176 176228
rect 86192 176284 86256 176288
rect 86192 176228 86196 176284
rect 86196 176228 86252 176284
rect 86252 176228 86256 176284
rect 86192 176224 86256 176228
rect 89952 176284 90016 176288
rect 89952 176228 89956 176284
rect 89956 176228 90012 176284
rect 90012 176228 90016 176284
rect 89952 176224 90016 176228
rect 90032 176284 90096 176288
rect 90032 176228 90036 176284
rect 90036 176228 90092 176284
rect 90092 176228 90096 176284
rect 90032 176224 90096 176228
rect 90112 176284 90176 176288
rect 90112 176228 90116 176284
rect 90116 176228 90172 176284
rect 90172 176228 90176 176284
rect 90112 176224 90176 176228
rect 90192 176284 90256 176288
rect 90192 176228 90196 176284
rect 90196 176228 90252 176284
rect 90252 176228 90256 176284
rect 90192 176224 90256 176228
rect 3952 175740 4016 175744
rect 3952 175684 3956 175740
rect 3956 175684 4012 175740
rect 4012 175684 4016 175740
rect 3952 175680 4016 175684
rect 4032 175740 4096 175744
rect 4032 175684 4036 175740
rect 4036 175684 4092 175740
rect 4092 175684 4096 175740
rect 4032 175680 4096 175684
rect 4112 175740 4176 175744
rect 4112 175684 4116 175740
rect 4116 175684 4172 175740
rect 4172 175684 4176 175740
rect 4112 175680 4176 175684
rect 4192 175740 4256 175744
rect 4192 175684 4196 175740
rect 4196 175684 4252 175740
rect 4252 175684 4256 175740
rect 4192 175680 4256 175684
rect 87952 175740 88016 175744
rect 87952 175684 87956 175740
rect 87956 175684 88012 175740
rect 88012 175684 88016 175740
rect 87952 175680 88016 175684
rect 88032 175740 88096 175744
rect 88032 175684 88036 175740
rect 88036 175684 88092 175740
rect 88092 175684 88096 175740
rect 88032 175680 88096 175684
rect 88112 175740 88176 175744
rect 88112 175684 88116 175740
rect 88116 175684 88172 175740
rect 88172 175684 88176 175740
rect 88112 175680 88176 175684
rect 88192 175740 88256 175744
rect 88192 175684 88196 175740
rect 88196 175684 88252 175740
rect 88252 175684 88256 175740
rect 88192 175680 88256 175684
rect 83596 175340 83660 175404
rect 1952 175196 2016 175200
rect 1952 175140 1956 175196
rect 1956 175140 2012 175196
rect 2012 175140 2016 175196
rect 1952 175136 2016 175140
rect 2032 175196 2096 175200
rect 2032 175140 2036 175196
rect 2036 175140 2092 175196
rect 2092 175140 2096 175196
rect 2032 175136 2096 175140
rect 2112 175196 2176 175200
rect 2112 175140 2116 175196
rect 2116 175140 2172 175196
rect 2172 175140 2176 175196
rect 2112 175136 2176 175140
rect 2192 175196 2256 175200
rect 2192 175140 2196 175196
rect 2196 175140 2252 175196
rect 2252 175140 2256 175196
rect 2192 175136 2256 175140
rect 85952 175196 86016 175200
rect 85952 175140 85956 175196
rect 85956 175140 86012 175196
rect 86012 175140 86016 175196
rect 85952 175136 86016 175140
rect 86032 175196 86096 175200
rect 86032 175140 86036 175196
rect 86036 175140 86092 175196
rect 86092 175140 86096 175196
rect 86032 175136 86096 175140
rect 86112 175196 86176 175200
rect 86112 175140 86116 175196
rect 86116 175140 86172 175196
rect 86172 175140 86176 175196
rect 86112 175136 86176 175140
rect 86192 175196 86256 175200
rect 86192 175140 86196 175196
rect 86196 175140 86252 175196
rect 86252 175140 86256 175196
rect 86192 175136 86256 175140
rect 89952 175196 90016 175200
rect 89952 175140 89956 175196
rect 89956 175140 90012 175196
rect 90012 175140 90016 175196
rect 89952 175136 90016 175140
rect 90032 175196 90096 175200
rect 90032 175140 90036 175196
rect 90036 175140 90092 175196
rect 90092 175140 90096 175196
rect 90032 175136 90096 175140
rect 90112 175196 90176 175200
rect 90112 175140 90116 175196
rect 90116 175140 90172 175196
rect 90172 175140 90176 175196
rect 90112 175136 90176 175140
rect 90192 175196 90256 175200
rect 90192 175140 90196 175196
rect 90196 175140 90252 175196
rect 90252 175140 90256 175196
rect 90192 175136 90256 175140
rect 3952 174652 4016 174656
rect 3952 174596 3956 174652
rect 3956 174596 4012 174652
rect 4012 174596 4016 174652
rect 3952 174592 4016 174596
rect 4032 174652 4096 174656
rect 4032 174596 4036 174652
rect 4036 174596 4092 174652
rect 4092 174596 4096 174652
rect 4032 174592 4096 174596
rect 4112 174652 4176 174656
rect 4112 174596 4116 174652
rect 4116 174596 4172 174652
rect 4172 174596 4176 174652
rect 4112 174592 4176 174596
rect 4192 174652 4256 174656
rect 4192 174596 4196 174652
rect 4196 174596 4252 174652
rect 4252 174596 4256 174652
rect 4192 174592 4256 174596
rect 87952 174652 88016 174656
rect 87952 174596 87956 174652
rect 87956 174596 88012 174652
rect 88012 174596 88016 174652
rect 87952 174592 88016 174596
rect 88032 174652 88096 174656
rect 88032 174596 88036 174652
rect 88036 174596 88092 174652
rect 88092 174596 88096 174652
rect 88032 174592 88096 174596
rect 88112 174652 88176 174656
rect 88112 174596 88116 174652
rect 88116 174596 88172 174652
rect 88172 174596 88176 174652
rect 88112 174592 88176 174596
rect 88192 174652 88256 174656
rect 88192 174596 88196 174652
rect 88196 174596 88252 174652
rect 88252 174596 88256 174652
rect 88192 174592 88256 174596
rect 1952 174108 2016 174112
rect 1952 174052 1956 174108
rect 1956 174052 2012 174108
rect 2012 174052 2016 174108
rect 1952 174048 2016 174052
rect 2032 174108 2096 174112
rect 2032 174052 2036 174108
rect 2036 174052 2092 174108
rect 2092 174052 2096 174108
rect 2032 174048 2096 174052
rect 2112 174108 2176 174112
rect 2112 174052 2116 174108
rect 2116 174052 2172 174108
rect 2172 174052 2176 174108
rect 2112 174048 2176 174052
rect 2192 174108 2256 174112
rect 2192 174052 2196 174108
rect 2196 174052 2252 174108
rect 2252 174052 2256 174108
rect 2192 174048 2256 174052
rect 85952 174108 86016 174112
rect 85952 174052 85956 174108
rect 85956 174052 86012 174108
rect 86012 174052 86016 174108
rect 85952 174048 86016 174052
rect 86032 174108 86096 174112
rect 86032 174052 86036 174108
rect 86036 174052 86092 174108
rect 86092 174052 86096 174108
rect 86032 174048 86096 174052
rect 86112 174108 86176 174112
rect 86112 174052 86116 174108
rect 86116 174052 86172 174108
rect 86172 174052 86176 174108
rect 86112 174048 86176 174052
rect 86192 174108 86256 174112
rect 86192 174052 86196 174108
rect 86196 174052 86252 174108
rect 86252 174052 86256 174108
rect 86192 174048 86256 174052
rect 89952 174108 90016 174112
rect 89952 174052 89956 174108
rect 89956 174052 90012 174108
rect 90012 174052 90016 174108
rect 89952 174048 90016 174052
rect 90032 174108 90096 174112
rect 90032 174052 90036 174108
rect 90036 174052 90092 174108
rect 90092 174052 90096 174108
rect 90032 174048 90096 174052
rect 90112 174108 90176 174112
rect 90112 174052 90116 174108
rect 90116 174052 90172 174108
rect 90172 174052 90176 174108
rect 90112 174048 90176 174052
rect 90192 174108 90256 174112
rect 90192 174052 90196 174108
rect 90196 174052 90252 174108
rect 90252 174052 90256 174108
rect 90192 174048 90256 174052
rect 3952 173564 4016 173568
rect 3952 173508 3956 173564
rect 3956 173508 4012 173564
rect 4012 173508 4016 173564
rect 3952 173504 4016 173508
rect 4032 173564 4096 173568
rect 4032 173508 4036 173564
rect 4036 173508 4092 173564
rect 4092 173508 4096 173564
rect 4032 173504 4096 173508
rect 4112 173564 4176 173568
rect 4112 173508 4116 173564
rect 4116 173508 4172 173564
rect 4172 173508 4176 173564
rect 4112 173504 4176 173508
rect 4192 173564 4256 173568
rect 4192 173508 4196 173564
rect 4196 173508 4252 173564
rect 4252 173508 4256 173564
rect 4192 173504 4256 173508
rect 87952 173564 88016 173568
rect 87952 173508 87956 173564
rect 87956 173508 88012 173564
rect 88012 173508 88016 173564
rect 87952 173504 88016 173508
rect 88032 173564 88096 173568
rect 88032 173508 88036 173564
rect 88036 173508 88092 173564
rect 88092 173508 88096 173564
rect 88032 173504 88096 173508
rect 88112 173564 88176 173568
rect 88112 173508 88116 173564
rect 88116 173508 88172 173564
rect 88172 173508 88176 173564
rect 88112 173504 88176 173508
rect 88192 173564 88256 173568
rect 88192 173508 88196 173564
rect 88196 173508 88252 173564
rect 88252 173508 88256 173564
rect 88192 173504 88256 173508
rect 1952 173020 2016 173024
rect 1952 172964 1956 173020
rect 1956 172964 2012 173020
rect 2012 172964 2016 173020
rect 1952 172960 2016 172964
rect 2032 173020 2096 173024
rect 2032 172964 2036 173020
rect 2036 172964 2092 173020
rect 2092 172964 2096 173020
rect 2032 172960 2096 172964
rect 2112 173020 2176 173024
rect 2112 172964 2116 173020
rect 2116 172964 2172 173020
rect 2172 172964 2176 173020
rect 2112 172960 2176 172964
rect 2192 173020 2256 173024
rect 2192 172964 2196 173020
rect 2196 172964 2252 173020
rect 2252 172964 2256 173020
rect 2192 172960 2256 172964
rect 85952 173020 86016 173024
rect 85952 172964 85956 173020
rect 85956 172964 86012 173020
rect 86012 172964 86016 173020
rect 85952 172960 86016 172964
rect 86032 173020 86096 173024
rect 86032 172964 86036 173020
rect 86036 172964 86092 173020
rect 86092 172964 86096 173020
rect 86032 172960 86096 172964
rect 86112 173020 86176 173024
rect 86112 172964 86116 173020
rect 86116 172964 86172 173020
rect 86172 172964 86176 173020
rect 86112 172960 86176 172964
rect 86192 173020 86256 173024
rect 86192 172964 86196 173020
rect 86196 172964 86252 173020
rect 86252 172964 86256 173020
rect 86192 172960 86256 172964
rect 89952 173020 90016 173024
rect 89952 172964 89956 173020
rect 89956 172964 90012 173020
rect 90012 172964 90016 173020
rect 89952 172960 90016 172964
rect 90032 173020 90096 173024
rect 90032 172964 90036 173020
rect 90036 172964 90092 173020
rect 90092 172964 90096 173020
rect 90032 172960 90096 172964
rect 90112 173020 90176 173024
rect 90112 172964 90116 173020
rect 90116 172964 90172 173020
rect 90172 172964 90176 173020
rect 90112 172960 90176 172964
rect 90192 173020 90256 173024
rect 90192 172964 90196 173020
rect 90196 172964 90252 173020
rect 90252 172964 90256 173020
rect 90192 172960 90256 172964
rect 3952 172476 4016 172480
rect 3952 172420 3956 172476
rect 3956 172420 4012 172476
rect 4012 172420 4016 172476
rect 3952 172416 4016 172420
rect 4032 172476 4096 172480
rect 4032 172420 4036 172476
rect 4036 172420 4092 172476
rect 4092 172420 4096 172476
rect 4032 172416 4096 172420
rect 4112 172476 4176 172480
rect 4112 172420 4116 172476
rect 4116 172420 4172 172476
rect 4172 172420 4176 172476
rect 4112 172416 4176 172420
rect 4192 172476 4256 172480
rect 4192 172420 4196 172476
rect 4196 172420 4252 172476
rect 4252 172420 4256 172476
rect 4192 172416 4256 172420
rect 87952 172476 88016 172480
rect 87952 172420 87956 172476
rect 87956 172420 88012 172476
rect 88012 172420 88016 172476
rect 87952 172416 88016 172420
rect 88032 172476 88096 172480
rect 88032 172420 88036 172476
rect 88036 172420 88092 172476
rect 88092 172420 88096 172476
rect 88032 172416 88096 172420
rect 88112 172476 88176 172480
rect 88112 172420 88116 172476
rect 88116 172420 88172 172476
rect 88172 172420 88176 172476
rect 88112 172416 88176 172420
rect 88192 172476 88256 172480
rect 88192 172420 88196 172476
rect 88196 172420 88252 172476
rect 88252 172420 88256 172476
rect 88192 172416 88256 172420
rect 1952 171932 2016 171936
rect 1952 171876 1956 171932
rect 1956 171876 2012 171932
rect 2012 171876 2016 171932
rect 1952 171872 2016 171876
rect 2032 171932 2096 171936
rect 2032 171876 2036 171932
rect 2036 171876 2092 171932
rect 2092 171876 2096 171932
rect 2032 171872 2096 171876
rect 2112 171932 2176 171936
rect 2112 171876 2116 171932
rect 2116 171876 2172 171932
rect 2172 171876 2176 171932
rect 2112 171872 2176 171876
rect 2192 171932 2256 171936
rect 2192 171876 2196 171932
rect 2196 171876 2252 171932
rect 2252 171876 2256 171932
rect 2192 171872 2256 171876
rect 85952 171932 86016 171936
rect 85952 171876 85956 171932
rect 85956 171876 86012 171932
rect 86012 171876 86016 171932
rect 85952 171872 86016 171876
rect 86032 171932 86096 171936
rect 86032 171876 86036 171932
rect 86036 171876 86092 171932
rect 86092 171876 86096 171932
rect 86032 171872 86096 171876
rect 86112 171932 86176 171936
rect 86112 171876 86116 171932
rect 86116 171876 86172 171932
rect 86172 171876 86176 171932
rect 86112 171872 86176 171876
rect 86192 171932 86256 171936
rect 86192 171876 86196 171932
rect 86196 171876 86252 171932
rect 86252 171876 86256 171932
rect 86192 171872 86256 171876
rect 89952 171932 90016 171936
rect 89952 171876 89956 171932
rect 89956 171876 90012 171932
rect 90012 171876 90016 171932
rect 89952 171872 90016 171876
rect 90032 171932 90096 171936
rect 90032 171876 90036 171932
rect 90036 171876 90092 171932
rect 90092 171876 90096 171932
rect 90032 171872 90096 171876
rect 90112 171932 90176 171936
rect 90112 171876 90116 171932
rect 90116 171876 90172 171932
rect 90172 171876 90176 171932
rect 90112 171872 90176 171876
rect 90192 171932 90256 171936
rect 90192 171876 90196 171932
rect 90196 171876 90252 171932
rect 90252 171876 90256 171932
rect 90192 171872 90256 171876
rect 3952 171388 4016 171392
rect 3952 171332 3956 171388
rect 3956 171332 4012 171388
rect 4012 171332 4016 171388
rect 3952 171328 4016 171332
rect 4032 171388 4096 171392
rect 4032 171332 4036 171388
rect 4036 171332 4092 171388
rect 4092 171332 4096 171388
rect 4032 171328 4096 171332
rect 4112 171388 4176 171392
rect 4112 171332 4116 171388
rect 4116 171332 4172 171388
rect 4172 171332 4176 171388
rect 4112 171328 4176 171332
rect 4192 171388 4256 171392
rect 4192 171332 4196 171388
rect 4196 171332 4252 171388
rect 4252 171332 4256 171388
rect 4192 171328 4256 171332
rect 87952 171388 88016 171392
rect 87952 171332 87956 171388
rect 87956 171332 88012 171388
rect 88012 171332 88016 171388
rect 87952 171328 88016 171332
rect 88032 171388 88096 171392
rect 88032 171332 88036 171388
rect 88036 171332 88092 171388
rect 88092 171332 88096 171388
rect 88032 171328 88096 171332
rect 88112 171388 88176 171392
rect 88112 171332 88116 171388
rect 88116 171332 88172 171388
rect 88172 171332 88176 171388
rect 88112 171328 88176 171332
rect 88192 171388 88256 171392
rect 88192 171332 88196 171388
rect 88196 171332 88252 171388
rect 88252 171332 88256 171388
rect 88192 171328 88256 171332
rect 1952 170844 2016 170848
rect 1952 170788 1956 170844
rect 1956 170788 2012 170844
rect 2012 170788 2016 170844
rect 1952 170784 2016 170788
rect 2032 170844 2096 170848
rect 2032 170788 2036 170844
rect 2036 170788 2092 170844
rect 2092 170788 2096 170844
rect 2032 170784 2096 170788
rect 2112 170844 2176 170848
rect 2112 170788 2116 170844
rect 2116 170788 2172 170844
rect 2172 170788 2176 170844
rect 2112 170784 2176 170788
rect 2192 170844 2256 170848
rect 2192 170788 2196 170844
rect 2196 170788 2252 170844
rect 2252 170788 2256 170844
rect 2192 170784 2256 170788
rect 85952 170844 86016 170848
rect 85952 170788 85956 170844
rect 85956 170788 86012 170844
rect 86012 170788 86016 170844
rect 85952 170784 86016 170788
rect 86032 170844 86096 170848
rect 86032 170788 86036 170844
rect 86036 170788 86092 170844
rect 86092 170788 86096 170844
rect 86032 170784 86096 170788
rect 86112 170844 86176 170848
rect 86112 170788 86116 170844
rect 86116 170788 86172 170844
rect 86172 170788 86176 170844
rect 86112 170784 86176 170788
rect 86192 170844 86256 170848
rect 86192 170788 86196 170844
rect 86196 170788 86252 170844
rect 86252 170788 86256 170844
rect 86192 170784 86256 170788
rect 89952 170844 90016 170848
rect 89952 170788 89956 170844
rect 89956 170788 90012 170844
rect 90012 170788 90016 170844
rect 89952 170784 90016 170788
rect 90032 170844 90096 170848
rect 90032 170788 90036 170844
rect 90036 170788 90092 170844
rect 90092 170788 90096 170844
rect 90032 170784 90096 170788
rect 90112 170844 90176 170848
rect 90112 170788 90116 170844
rect 90116 170788 90172 170844
rect 90172 170788 90176 170844
rect 90112 170784 90176 170788
rect 90192 170844 90256 170848
rect 90192 170788 90196 170844
rect 90196 170788 90252 170844
rect 90252 170788 90256 170844
rect 90192 170784 90256 170788
rect 3952 170300 4016 170304
rect 3952 170244 3956 170300
rect 3956 170244 4012 170300
rect 4012 170244 4016 170300
rect 3952 170240 4016 170244
rect 4032 170300 4096 170304
rect 4032 170244 4036 170300
rect 4036 170244 4092 170300
rect 4092 170244 4096 170300
rect 4032 170240 4096 170244
rect 4112 170300 4176 170304
rect 4112 170244 4116 170300
rect 4116 170244 4172 170300
rect 4172 170244 4176 170300
rect 4112 170240 4176 170244
rect 4192 170300 4256 170304
rect 4192 170244 4196 170300
rect 4196 170244 4252 170300
rect 4252 170244 4256 170300
rect 4192 170240 4256 170244
rect 87952 170300 88016 170304
rect 87952 170244 87956 170300
rect 87956 170244 88012 170300
rect 88012 170244 88016 170300
rect 87952 170240 88016 170244
rect 88032 170300 88096 170304
rect 88032 170244 88036 170300
rect 88036 170244 88092 170300
rect 88092 170244 88096 170300
rect 88032 170240 88096 170244
rect 88112 170300 88176 170304
rect 88112 170244 88116 170300
rect 88116 170244 88172 170300
rect 88172 170244 88176 170300
rect 88112 170240 88176 170244
rect 88192 170300 88256 170304
rect 88192 170244 88196 170300
rect 88196 170244 88252 170300
rect 88252 170244 88256 170300
rect 88192 170240 88256 170244
rect 1952 169756 2016 169760
rect 1952 169700 1956 169756
rect 1956 169700 2012 169756
rect 2012 169700 2016 169756
rect 1952 169696 2016 169700
rect 2032 169756 2096 169760
rect 2032 169700 2036 169756
rect 2036 169700 2092 169756
rect 2092 169700 2096 169756
rect 2032 169696 2096 169700
rect 2112 169756 2176 169760
rect 2112 169700 2116 169756
rect 2116 169700 2172 169756
rect 2172 169700 2176 169756
rect 2112 169696 2176 169700
rect 2192 169756 2256 169760
rect 2192 169700 2196 169756
rect 2196 169700 2252 169756
rect 2252 169700 2256 169756
rect 2192 169696 2256 169700
rect 85952 169756 86016 169760
rect 85952 169700 85956 169756
rect 85956 169700 86012 169756
rect 86012 169700 86016 169756
rect 85952 169696 86016 169700
rect 86032 169756 86096 169760
rect 86032 169700 86036 169756
rect 86036 169700 86092 169756
rect 86092 169700 86096 169756
rect 86032 169696 86096 169700
rect 86112 169756 86176 169760
rect 86112 169700 86116 169756
rect 86116 169700 86172 169756
rect 86172 169700 86176 169756
rect 86112 169696 86176 169700
rect 86192 169756 86256 169760
rect 86192 169700 86196 169756
rect 86196 169700 86252 169756
rect 86252 169700 86256 169756
rect 86192 169696 86256 169700
rect 89952 169756 90016 169760
rect 89952 169700 89956 169756
rect 89956 169700 90012 169756
rect 90012 169700 90016 169756
rect 89952 169696 90016 169700
rect 90032 169756 90096 169760
rect 90032 169700 90036 169756
rect 90036 169700 90092 169756
rect 90092 169700 90096 169756
rect 90032 169696 90096 169700
rect 90112 169756 90176 169760
rect 90112 169700 90116 169756
rect 90116 169700 90172 169756
rect 90172 169700 90176 169756
rect 90112 169696 90176 169700
rect 90192 169756 90256 169760
rect 90192 169700 90196 169756
rect 90196 169700 90252 169756
rect 90252 169700 90256 169756
rect 90192 169696 90256 169700
rect 3952 169212 4016 169216
rect 3952 169156 3956 169212
rect 3956 169156 4012 169212
rect 4012 169156 4016 169212
rect 3952 169152 4016 169156
rect 4032 169212 4096 169216
rect 4032 169156 4036 169212
rect 4036 169156 4092 169212
rect 4092 169156 4096 169212
rect 4032 169152 4096 169156
rect 4112 169212 4176 169216
rect 4112 169156 4116 169212
rect 4116 169156 4172 169212
rect 4172 169156 4176 169212
rect 4112 169152 4176 169156
rect 4192 169212 4256 169216
rect 4192 169156 4196 169212
rect 4196 169156 4252 169212
rect 4252 169156 4256 169212
rect 4192 169152 4256 169156
rect 87952 169212 88016 169216
rect 87952 169156 87956 169212
rect 87956 169156 88012 169212
rect 88012 169156 88016 169212
rect 87952 169152 88016 169156
rect 88032 169212 88096 169216
rect 88032 169156 88036 169212
rect 88036 169156 88092 169212
rect 88092 169156 88096 169212
rect 88032 169152 88096 169156
rect 88112 169212 88176 169216
rect 88112 169156 88116 169212
rect 88116 169156 88172 169212
rect 88172 169156 88176 169212
rect 88112 169152 88176 169156
rect 88192 169212 88256 169216
rect 88192 169156 88196 169212
rect 88196 169156 88252 169212
rect 88252 169156 88256 169212
rect 88192 169152 88256 169156
rect 1952 168668 2016 168672
rect 1952 168612 1956 168668
rect 1956 168612 2012 168668
rect 2012 168612 2016 168668
rect 1952 168608 2016 168612
rect 2032 168668 2096 168672
rect 2032 168612 2036 168668
rect 2036 168612 2092 168668
rect 2092 168612 2096 168668
rect 2032 168608 2096 168612
rect 2112 168668 2176 168672
rect 2112 168612 2116 168668
rect 2116 168612 2172 168668
rect 2172 168612 2176 168668
rect 2112 168608 2176 168612
rect 2192 168668 2256 168672
rect 2192 168612 2196 168668
rect 2196 168612 2252 168668
rect 2252 168612 2256 168668
rect 2192 168608 2256 168612
rect 85952 168668 86016 168672
rect 85952 168612 85956 168668
rect 85956 168612 86012 168668
rect 86012 168612 86016 168668
rect 85952 168608 86016 168612
rect 86032 168668 86096 168672
rect 86032 168612 86036 168668
rect 86036 168612 86092 168668
rect 86092 168612 86096 168668
rect 86032 168608 86096 168612
rect 86112 168668 86176 168672
rect 86112 168612 86116 168668
rect 86116 168612 86172 168668
rect 86172 168612 86176 168668
rect 86112 168608 86176 168612
rect 86192 168668 86256 168672
rect 86192 168612 86196 168668
rect 86196 168612 86252 168668
rect 86252 168612 86256 168668
rect 86192 168608 86256 168612
rect 89952 168668 90016 168672
rect 89952 168612 89956 168668
rect 89956 168612 90012 168668
rect 90012 168612 90016 168668
rect 89952 168608 90016 168612
rect 90032 168668 90096 168672
rect 90032 168612 90036 168668
rect 90036 168612 90092 168668
rect 90092 168612 90096 168668
rect 90032 168608 90096 168612
rect 90112 168668 90176 168672
rect 90112 168612 90116 168668
rect 90116 168612 90172 168668
rect 90172 168612 90176 168668
rect 90112 168608 90176 168612
rect 90192 168668 90256 168672
rect 90192 168612 90196 168668
rect 90196 168612 90252 168668
rect 90252 168612 90256 168668
rect 90192 168608 90256 168612
rect 3952 168124 4016 168128
rect 3952 168068 3956 168124
rect 3956 168068 4012 168124
rect 4012 168068 4016 168124
rect 3952 168064 4016 168068
rect 4032 168124 4096 168128
rect 4032 168068 4036 168124
rect 4036 168068 4092 168124
rect 4092 168068 4096 168124
rect 4032 168064 4096 168068
rect 4112 168124 4176 168128
rect 4112 168068 4116 168124
rect 4116 168068 4172 168124
rect 4172 168068 4176 168124
rect 4112 168064 4176 168068
rect 4192 168124 4256 168128
rect 4192 168068 4196 168124
rect 4196 168068 4252 168124
rect 4252 168068 4256 168124
rect 4192 168064 4256 168068
rect 87952 168124 88016 168128
rect 87952 168068 87956 168124
rect 87956 168068 88012 168124
rect 88012 168068 88016 168124
rect 87952 168064 88016 168068
rect 88032 168124 88096 168128
rect 88032 168068 88036 168124
rect 88036 168068 88092 168124
rect 88092 168068 88096 168124
rect 88032 168064 88096 168068
rect 88112 168124 88176 168128
rect 88112 168068 88116 168124
rect 88116 168068 88172 168124
rect 88172 168068 88176 168124
rect 88112 168064 88176 168068
rect 88192 168124 88256 168128
rect 88192 168068 88196 168124
rect 88196 168068 88252 168124
rect 88252 168068 88256 168124
rect 88192 168064 88256 168068
rect 1952 167580 2016 167584
rect 1952 167524 1956 167580
rect 1956 167524 2012 167580
rect 2012 167524 2016 167580
rect 1952 167520 2016 167524
rect 2032 167580 2096 167584
rect 2032 167524 2036 167580
rect 2036 167524 2092 167580
rect 2092 167524 2096 167580
rect 2032 167520 2096 167524
rect 2112 167580 2176 167584
rect 2112 167524 2116 167580
rect 2116 167524 2172 167580
rect 2172 167524 2176 167580
rect 2112 167520 2176 167524
rect 2192 167580 2256 167584
rect 2192 167524 2196 167580
rect 2196 167524 2252 167580
rect 2252 167524 2256 167580
rect 2192 167520 2256 167524
rect 85952 167580 86016 167584
rect 85952 167524 85956 167580
rect 85956 167524 86012 167580
rect 86012 167524 86016 167580
rect 85952 167520 86016 167524
rect 86032 167580 86096 167584
rect 86032 167524 86036 167580
rect 86036 167524 86092 167580
rect 86092 167524 86096 167580
rect 86032 167520 86096 167524
rect 86112 167580 86176 167584
rect 86112 167524 86116 167580
rect 86116 167524 86172 167580
rect 86172 167524 86176 167580
rect 86112 167520 86176 167524
rect 86192 167580 86256 167584
rect 86192 167524 86196 167580
rect 86196 167524 86252 167580
rect 86252 167524 86256 167580
rect 86192 167520 86256 167524
rect 89952 167580 90016 167584
rect 89952 167524 89956 167580
rect 89956 167524 90012 167580
rect 90012 167524 90016 167580
rect 89952 167520 90016 167524
rect 90032 167580 90096 167584
rect 90032 167524 90036 167580
rect 90036 167524 90092 167580
rect 90092 167524 90096 167580
rect 90032 167520 90096 167524
rect 90112 167580 90176 167584
rect 90112 167524 90116 167580
rect 90116 167524 90172 167580
rect 90172 167524 90176 167580
rect 90112 167520 90176 167524
rect 90192 167580 90256 167584
rect 90192 167524 90196 167580
rect 90196 167524 90252 167580
rect 90252 167524 90256 167580
rect 90192 167520 90256 167524
rect 83780 167316 83844 167380
rect 3952 167036 4016 167040
rect 3952 166980 3956 167036
rect 3956 166980 4012 167036
rect 4012 166980 4016 167036
rect 3952 166976 4016 166980
rect 4032 167036 4096 167040
rect 4032 166980 4036 167036
rect 4036 166980 4092 167036
rect 4092 166980 4096 167036
rect 4032 166976 4096 166980
rect 4112 167036 4176 167040
rect 4112 166980 4116 167036
rect 4116 166980 4172 167036
rect 4172 166980 4176 167036
rect 4112 166976 4176 166980
rect 4192 167036 4256 167040
rect 4192 166980 4196 167036
rect 4196 166980 4252 167036
rect 4252 166980 4256 167036
rect 4192 166976 4256 166980
rect 87952 167036 88016 167040
rect 87952 166980 87956 167036
rect 87956 166980 88012 167036
rect 88012 166980 88016 167036
rect 87952 166976 88016 166980
rect 88032 167036 88096 167040
rect 88032 166980 88036 167036
rect 88036 166980 88092 167036
rect 88092 166980 88096 167036
rect 88032 166976 88096 166980
rect 88112 167036 88176 167040
rect 88112 166980 88116 167036
rect 88116 166980 88172 167036
rect 88172 166980 88176 167036
rect 88112 166976 88176 166980
rect 88192 167036 88256 167040
rect 88192 166980 88196 167036
rect 88196 166980 88252 167036
rect 88252 166980 88256 167036
rect 88192 166976 88256 166980
rect 1952 166492 2016 166496
rect 1952 166436 1956 166492
rect 1956 166436 2012 166492
rect 2012 166436 2016 166492
rect 1952 166432 2016 166436
rect 2032 166492 2096 166496
rect 2032 166436 2036 166492
rect 2036 166436 2092 166492
rect 2092 166436 2096 166492
rect 2032 166432 2096 166436
rect 2112 166492 2176 166496
rect 2112 166436 2116 166492
rect 2116 166436 2172 166492
rect 2172 166436 2176 166492
rect 2112 166432 2176 166436
rect 2192 166492 2256 166496
rect 2192 166436 2196 166492
rect 2196 166436 2252 166492
rect 2252 166436 2256 166492
rect 2192 166432 2256 166436
rect 85952 166492 86016 166496
rect 85952 166436 85956 166492
rect 85956 166436 86012 166492
rect 86012 166436 86016 166492
rect 85952 166432 86016 166436
rect 86032 166492 86096 166496
rect 86032 166436 86036 166492
rect 86036 166436 86092 166492
rect 86092 166436 86096 166492
rect 86032 166432 86096 166436
rect 86112 166492 86176 166496
rect 86112 166436 86116 166492
rect 86116 166436 86172 166492
rect 86172 166436 86176 166492
rect 86112 166432 86176 166436
rect 86192 166492 86256 166496
rect 86192 166436 86196 166492
rect 86196 166436 86252 166492
rect 86252 166436 86256 166492
rect 86192 166432 86256 166436
rect 89952 166492 90016 166496
rect 89952 166436 89956 166492
rect 89956 166436 90012 166492
rect 90012 166436 90016 166492
rect 89952 166432 90016 166436
rect 90032 166492 90096 166496
rect 90032 166436 90036 166492
rect 90036 166436 90092 166492
rect 90092 166436 90096 166492
rect 90032 166432 90096 166436
rect 90112 166492 90176 166496
rect 90112 166436 90116 166492
rect 90116 166436 90172 166492
rect 90172 166436 90176 166492
rect 90112 166432 90176 166436
rect 90192 166492 90256 166496
rect 90192 166436 90196 166492
rect 90196 166436 90252 166492
rect 90252 166436 90256 166492
rect 90192 166432 90256 166436
rect 3952 165948 4016 165952
rect 3952 165892 3956 165948
rect 3956 165892 4012 165948
rect 4012 165892 4016 165948
rect 3952 165888 4016 165892
rect 4032 165948 4096 165952
rect 4032 165892 4036 165948
rect 4036 165892 4092 165948
rect 4092 165892 4096 165948
rect 4032 165888 4096 165892
rect 4112 165948 4176 165952
rect 4112 165892 4116 165948
rect 4116 165892 4172 165948
rect 4172 165892 4176 165948
rect 4112 165888 4176 165892
rect 4192 165948 4256 165952
rect 4192 165892 4196 165948
rect 4196 165892 4252 165948
rect 4252 165892 4256 165948
rect 4192 165888 4256 165892
rect 87952 165948 88016 165952
rect 87952 165892 87956 165948
rect 87956 165892 88012 165948
rect 88012 165892 88016 165948
rect 87952 165888 88016 165892
rect 88032 165948 88096 165952
rect 88032 165892 88036 165948
rect 88036 165892 88092 165948
rect 88092 165892 88096 165948
rect 88032 165888 88096 165892
rect 88112 165948 88176 165952
rect 88112 165892 88116 165948
rect 88116 165892 88172 165948
rect 88172 165892 88176 165948
rect 88112 165888 88176 165892
rect 88192 165948 88256 165952
rect 88192 165892 88196 165948
rect 88196 165892 88252 165948
rect 88252 165892 88256 165948
rect 88192 165888 88256 165892
rect 1952 165404 2016 165408
rect 1952 165348 1956 165404
rect 1956 165348 2012 165404
rect 2012 165348 2016 165404
rect 1952 165344 2016 165348
rect 2032 165404 2096 165408
rect 2032 165348 2036 165404
rect 2036 165348 2092 165404
rect 2092 165348 2096 165404
rect 2032 165344 2096 165348
rect 2112 165404 2176 165408
rect 2112 165348 2116 165404
rect 2116 165348 2172 165404
rect 2172 165348 2176 165404
rect 2112 165344 2176 165348
rect 2192 165404 2256 165408
rect 2192 165348 2196 165404
rect 2196 165348 2252 165404
rect 2252 165348 2256 165404
rect 2192 165344 2256 165348
rect 85952 165404 86016 165408
rect 85952 165348 85956 165404
rect 85956 165348 86012 165404
rect 86012 165348 86016 165404
rect 85952 165344 86016 165348
rect 86032 165404 86096 165408
rect 86032 165348 86036 165404
rect 86036 165348 86092 165404
rect 86092 165348 86096 165404
rect 86032 165344 86096 165348
rect 86112 165404 86176 165408
rect 86112 165348 86116 165404
rect 86116 165348 86172 165404
rect 86172 165348 86176 165404
rect 86112 165344 86176 165348
rect 86192 165404 86256 165408
rect 86192 165348 86196 165404
rect 86196 165348 86252 165404
rect 86252 165348 86256 165404
rect 86192 165344 86256 165348
rect 89952 165404 90016 165408
rect 89952 165348 89956 165404
rect 89956 165348 90012 165404
rect 90012 165348 90016 165404
rect 89952 165344 90016 165348
rect 90032 165404 90096 165408
rect 90032 165348 90036 165404
rect 90036 165348 90092 165404
rect 90092 165348 90096 165404
rect 90032 165344 90096 165348
rect 90112 165404 90176 165408
rect 90112 165348 90116 165404
rect 90116 165348 90172 165404
rect 90172 165348 90176 165404
rect 90112 165344 90176 165348
rect 90192 165404 90256 165408
rect 90192 165348 90196 165404
rect 90196 165348 90252 165404
rect 90252 165348 90256 165404
rect 90192 165344 90256 165348
rect 3952 164860 4016 164864
rect 3952 164804 3956 164860
rect 3956 164804 4012 164860
rect 4012 164804 4016 164860
rect 3952 164800 4016 164804
rect 4032 164860 4096 164864
rect 4032 164804 4036 164860
rect 4036 164804 4092 164860
rect 4092 164804 4096 164860
rect 4032 164800 4096 164804
rect 4112 164860 4176 164864
rect 4112 164804 4116 164860
rect 4116 164804 4172 164860
rect 4172 164804 4176 164860
rect 4112 164800 4176 164804
rect 4192 164860 4256 164864
rect 4192 164804 4196 164860
rect 4196 164804 4252 164860
rect 4252 164804 4256 164860
rect 4192 164800 4256 164804
rect 87952 164860 88016 164864
rect 87952 164804 87956 164860
rect 87956 164804 88012 164860
rect 88012 164804 88016 164860
rect 87952 164800 88016 164804
rect 88032 164860 88096 164864
rect 88032 164804 88036 164860
rect 88036 164804 88092 164860
rect 88092 164804 88096 164860
rect 88032 164800 88096 164804
rect 88112 164860 88176 164864
rect 88112 164804 88116 164860
rect 88116 164804 88172 164860
rect 88172 164804 88176 164860
rect 88112 164800 88176 164804
rect 88192 164860 88256 164864
rect 88192 164804 88196 164860
rect 88196 164804 88252 164860
rect 88252 164804 88256 164860
rect 88192 164800 88256 164804
rect 1952 164316 2016 164320
rect 1952 164260 1956 164316
rect 1956 164260 2012 164316
rect 2012 164260 2016 164316
rect 1952 164256 2016 164260
rect 2032 164316 2096 164320
rect 2032 164260 2036 164316
rect 2036 164260 2092 164316
rect 2092 164260 2096 164316
rect 2032 164256 2096 164260
rect 2112 164316 2176 164320
rect 2112 164260 2116 164316
rect 2116 164260 2172 164316
rect 2172 164260 2176 164316
rect 2112 164256 2176 164260
rect 2192 164316 2256 164320
rect 2192 164260 2196 164316
rect 2196 164260 2252 164316
rect 2252 164260 2256 164316
rect 2192 164256 2256 164260
rect 85952 164316 86016 164320
rect 85952 164260 85956 164316
rect 85956 164260 86012 164316
rect 86012 164260 86016 164316
rect 85952 164256 86016 164260
rect 86032 164316 86096 164320
rect 86032 164260 86036 164316
rect 86036 164260 86092 164316
rect 86092 164260 86096 164316
rect 86032 164256 86096 164260
rect 86112 164316 86176 164320
rect 86112 164260 86116 164316
rect 86116 164260 86172 164316
rect 86172 164260 86176 164316
rect 86112 164256 86176 164260
rect 86192 164316 86256 164320
rect 86192 164260 86196 164316
rect 86196 164260 86252 164316
rect 86252 164260 86256 164316
rect 86192 164256 86256 164260
rect 89952 164316 90016 164320
rect 89952 164260 89956 164316
rect 89956 164260 90012 164316
rect 90012 164260 90016 164316
rect 89952 164256 90016 164260
rect 90032 164316 90096 164320
rect 90032 164260 90036 164316
rect 90036 164260 90092 164316
rect 90092 164260 90096 164316
rect 90032 164256 90096 164260
rect 90112 164316 90176 164320
rect 90112 164260 90116 164316
rect 90116 164260 90172 164316
rect 90172 164260 90176 164316
rect 90112 164256 90176 164260
rect 90192 164316 90256 164320
rect 90192 164260 90196 164316
rect 90196 164260 90252 164316
rect 90252 164260 90256 164316
rect 90192 164256 90256 164260
rect 84332 164052 84396 164116
rect 3952 163772 4016 163776
rect 3952 163716 3956 163772
rect 3956 163716 4012 163772
rect 4012 163716 4016 163772
rect 3952 163712 4016 163716
rect 4032 163772 4096 163776
rect 4032 163716 4036 163772
rect 4036 163716 4092 163772
rect 4092 163716 4096 163772
rect 4032 163712 4096 163716
rect 4112 163772 4176 163776
rect 4112 163716 4116 163772
rect 4116 163716 4172 163772
rect 4172 163716 4176 163772
rect 4112 163712 4176 163716
rect 4192 163772 4256 163776
rect 4192 163716 4196 163772
rect 4196 163716 4252 163772
rect 4252 163716 4256 163772
rect 4192 163712 4256 163716
rect 87952 163772 88016 163776
rect 87952 163716 87956 163772
rect 87956 163716 88012 163772
rect 88012 163716 88016 163772
rect 87952 163712 88016 163716
rect 88032 163772 88096 163776
rect 88032 163716 88036 163772
rect 88036 163716 88092 163772
rect 88092 163716 88096 163772
rect 88032 163712 88096 163716
rect 88112 163772 88176 163776
rect 88112 163716 88116 163772
rect 88116 163716 88172 163772
rect 88172 163716 88176 163772
rect 88112 163712 88176 163716
rect 88192 163772 88256 163776
rect 88192 163716 88196 163772
rect 88196 163716 88252 163772
rect 88252 163716 88256 163772
rect 88192 163712 88256 163716
rect 1952 163228 2016 163232
rect 1952 163172 1956 163228
rect 1956 163172 2012 163228
rect 2012 163172 2016 163228
rect 1952 163168 2016 163172
rect 2032 163228 2096 163232
rect 2032 163172 2036 163228
rect 2036 163172 2092 163228
rect 2092 163172 2096 163228
rect 2032 163168 2096 163172
rect 2112 163228 2176 163232
rect 2112 163172 2116 163228
rect 2116 163172 2172 163228
rect 2172 163172 2176 163228
rect 2112 163168 2176 163172
rect 2192 163228 2256 163232
rect 2192 163172 2196 163228
rect 2196 163172 2252 163228
rect 2252 163172 2256 163228
rect 2192 163168 2256 163172
rect 85952 163228 86016 163232
rect 85952 163172 85956 163228
rect 85956 163172 86012 163228
rect 86012 163172 86016 163228
rect 85952 163168 86016 163172
rect 86032 163228 86096 163232
rect 86032 163172 86036 163228
rect 86036 163172 86092 163228
rect 86092 163172 86096 163228
rect 86032 163168 86096 163172
rect 86112 163228 86176 163232
rect 86112 163172 86116 163228
rect 86116 163172 86172 163228
rect 86172 163172 86176 163228
rect 86112 163168 86176 163172
rect 86192 163228 86256 163232
rect 86192 163172 86196 163228
rect 86196 163172 86252 163228
rect 86252 163172 86256 163228
rect 86192 163168 86256 163172
rect 89952 163228 90016 163232
rect 89952 163172 89956 163228
rect 89956 163172 90012 163228
rect 90012 163172 90016 163228
rect 89952 163168 90016 163172
rect 90032 163228 90096 163232
rect 90032 163172 90036 163228
rect 90036 163172 90092 163228
rect 90092 163172 90096 163228
rect 90032 163168 90096 163172
rect 90112 163228 90176 163232
rect 90112 163172 90116 163228
rect 90116 163172 90172 163228
rect 90172 163172 90176 163228
rect 90112 163168 90176 163172
rect 90192 163228 90256 163232
rect 90192 163172 90196 163228
rect 90196 163172 90252 163228
rect 90252 163172 90256 163228
rect 90192 163168 90256 163172
rect 3952 162684 4016 162688
rect 3952 162628 3956 162684
rect 3956 162628 4012 162684
rect 4012 162628 4016 162684
rect 3952 162624 4016 162628
rect 4032 162684 4096 162688
rect 4032 162628 4036 162684
rect 4036 162628 4092 162684
rect 4092 162628 4096 162684
rect 4032 162624 4096 162628
rect 4112 162684 4176 162688
rect 4112 162628 4116 162684
rect 4116 162628 4172 162684
rect 4172 162628 4176 162684
rect 4112 162624 4176 162628
rect 4192 162684 4256 162688
rect 4192 162628 4196 162684
rect 4196 162628 4252 162684
rect 4252 162628 4256 162684
rect 4192 162624 4256 162628
rect 87952 162684 88016 162688
rect 87952 162628 87956 162684
rect 87956 162628 88012 162684
rect 88012 162628 88016 162684
rect 87952 162624 88016 162628
rect 88032 162684 88096 162688
rect 88032 162628 88036 162684
rect 88036 162628 88092 162684
rect 88092 162628 88096 162684
rect 88032 162624 88096 162628
rect 88112 162684 88176 162688
rect 88112 162628 88116 162684
rect 88116 162628 88172 162684
rect 88172 162628 88176 162684
rect 88112 162624 88176 162628
rect 88192 162684 88256 162688
rect 88192 162628 88196 162684
rect 88196 162628 88252 162684
rect 88252 162628 88256 162684
rect 88192 162624 88256 162628
rect 1952 162140 2016 162144
rect 1952 162084 1956 162140
rect 1956 162084 2012 162140
rect 2012 162084 2016 162140
rect 1952 162080 2016 162084
rect 2032 162140 2096 162144
rect 2032 162084 2036 162140
rect 2036 162084 2092 162140
rect 2092 162084 2096 162140
rect 2032 162080 2096 162084
rect 2112 162140 2176 162144
rect 2112 162084 2116 162140
rect 2116 162084 2172 162140
rect 2172 162084 2176 162140
rect 2112 162080 2176 162084
rect 2192 162140 2256 162144
rect 2192 162084 2196 162140
rect 2196 162084 2252 162140
rect 2252 162084 2256 162140
rect 2192 162080 2256 162084
rect 85952 162140 86016 162144
rect 85952 162084 85956 162140
rect 85956 162084 86012 162140
rect 86012 162084 86016 162140
rect 85952 162080 86016 162084
rect 86032 162140 86096 162144
rect 86032 162084 86036 162140
rect 86036 162084 86092 162140
rect 86092 162084 86096 162140
rect 86032 162080 86096 162084
rect 86112 162140 86176 162144
rect 86112 162084 86116 162140
rect 86116 162084 86172 162140
rect 86172 162084 86176 162140
rect 86112 162080 86176 162084
rect 86192 162140 86256 162144
rect 86192 162084 86196 162140
rect 86196 162084 86252 162140
rect 86252 162084 86256 162140
rect 86192 162080 86256 162084
rect 89952 162140 90016 162144
rect 89952 162084 89956 162140
rect 89956 162084 90012 162140
rect 90012 162084 90016 162140
rect 89952 162080 90016 162084
rect 90032 162140 90096 162144
rect 90032 162084 90036 162140
rect 90036 162084 90092 162140
rect 90092 162084 90096 162140
rect 90032 162080 90096 162084
rect 90112 162140 90176 162144
rect 90112 162084 90116 162140
rect 90116 162084 90172 162140
rect 90172 162084 90176 162140
rect 90112 162080 90176 162084
rect 90192 162140 90256 162144
rect 90192 162084 90196 162140
rect 90196 162084 90252 162140
rect 90252 162084 90256 162140
rect 90192 162080 90256 162084
rect 86356 161876 86420 161940
rect 85068 161800 85132 161804
rect 85068 161744 85118 161800
rect 85118 161744 85132 161800
rect 85068 161740 85132 161744
rect 3952 161596 4016 161600
rect 3952 161540 3956 161596
rect 3956 161540 4012 161596
rect 4012 161540 4016 161596
rect 3952 161536 4016 161540
rect 4032 161596 4096 161600
rect 4032 161540 4036 161596
rect 4036 161540 4092 161596
rect 4092 161540 4096 161596
rect 4032 161536 4096 161540
rect 4112 161596 4176 161600
rect 4112 161540 4116 161596
rect 4116 161540 4172 161596
rect 4172 161540 4176 161596
rect 4112 161536 4176 161540
rect 4192 161596 4256 161600
rect 4192 161540 4196 161596
rect 4196 161540 4252 161596
rect 4252 161540 4256 161596
rect 4192 161536 4256 161540
rect 87952 161596 88016 161600
rect 87952 161540 87956 161596
rect 87956 161540 88012 161596
rect 88012 161540 88016 161596
rect 87952 161536 88016 161540
rect 88032 161596 88096 161600
rect 88032 161540 88036 161596
rect 88036 161540 88092 161596
rect 88092 161540 88096 161596
rect 88032 161536 88096 161540
rect 88112 161596 88176 161600
rect 88112 161540 88116 161596
rect 88116 161540 88172 161596
rect 88172 161540 88176 161596
rect 88112 161536 88176 161540
rect 88192 161596 88256 161600
rect 88192 161540 88196 161596
rect 88196 161540 88252 161596
rect 88252 161540 88256 161596
rect 88192 161536 88256 161540
rect 1952 161052 2016 161056
rect 1952 160996 1956 161052
rect 1956 160996 2012 161052
rect 2012 160996 2016 161052
rect 1952 160992 2016 160996
rect 2032 161052 2096 161056
rect 2032 160996 2036 161052
rect 2036 160996 2092 161052
rect 2092 160996 2096 161052
rect 2032 160992 2096 160996
rect 2112 161052 2176 161056
rect 2112 160996 2116 161052
rect 2116 160996 2172 161052
rect 2172 160996 2176 161052
rect 2112 160992 2176 160996
rect 2192 161052 2256 161056
rect 2192 160996 2196 161052
rect 2196 160996 2252 161052
rect 2252 160996 2256 161052
rect 2192 160992 2256 160996
rect 85952 161052 86016 161056
rect 85952 160996 85956 161052
rect 85956 160996 86012 161052
rect 86012 160996 86016 161052
rect 85952 160992 86016 160996
rect 86032 161052 86096 161056
rect 86032 160996 86036 161052
rect 86036 160996 86092 161052
rect 86092 160996 86096 161052
rect 86032 160992 86096 160996
rect 86112 161052 86176 161056
rect 86112 160996 86116 161052
rect 86116 160996 86172 161052
rect 86172 160996 86176 161052
rect 86112 160992 86176 160996
rect 86192 161052 86256 161056
rect 86192 160996 86196 161052
rect 86196 160996 86252 161052
rect 86252 160996 86256 161052
rect 86192 160992 86256 160996
rect 89952 161052 90016 161056
rect 89952 160996 89956 161052
rect 89956 160996 90012 161052
rect 90012 160996 90016 161052
rect 89952 160992 90016 160996
rect 90032 161052 90096 161056
rect 90032 160996 90036 161052
rect 90036 160996 90092 161052
rect 90092 160996 90096 161052
rect 90032 160992 90096 160996
rect 90112 161052 90176 161056
rect 90112 160996 90116 161052
rect 90116 160996 90172 161052
rect 90172 160996 90176 161052
rect 90112 160992 90176 160996
rect 90192 161052 90256 161056
rect 90192 160996 90196 161052
rect 90196 160996 90252 161052
rect 90252 160996 90256 161052
rect 90192 160992 90256 160996
rect 3952 160508 4016 160512
rect 3952 160452 3956 160508
rect 3956 160452 4012 160508
rect 4012 160452 4016 160508
rect 3952 160448 4016 160452
rect 4032 160508 4096 160512
rect 4032 160452 4036 160508
rect 4036 160452 4092 160508
rect 4092 160452 4096 160508
rect 4032 160448 4096 160452
rect 4112 160508 4176 160512
rect 4112 160452 4116 160508
rect 4116 160452 4172 160508
rect 4172 160452 4176 160508
rect 4112 160448 4176 160452
rect 4192 160508 4256 160512
rect 4192 160452 4196 160508
rect 4196 160452 4252 160508
rect 4252 160452 4256 160508
rect 4192 160448 4256 160452
rect 87952 160508 88016 160512
rect 87952 160452 87956 160508
rect 87956 160452 88012 160508
rect 88012 160452 88016 160508
rect 87952 160448 88016 160452
rect 88032 160508 88096 160512
rect 88032 160452 88036 160508
rect 88036 160452 88092 160508
rect 88092 160452 88096 160508
rect 88032 160448 88096 160452
rect 88112 160508 88176 160512
rect 88112 160452 88116 160508
rect 88116 160452 88172 160508
rect 88172 160452 88176 160508
rect 88112 160448 88176 160452
rect 88192 160508 88256 160512
rect 88192 160452 88196 160508
rect 88196 160452 88252 160508
rect 88252 160452 88256 160508
rect 88192 160448 88256 160452
rect 1952 159964 2016 159968
rect 1952 159908 1956 159964
rect 1956 159908 2012 159964
rect 2012 159908 2016 159964
rect 1952 159904 2016 159908
rect 2032 159964 2096 159968
rect 2032 159908 2036 159964
rect 2036 159908 2092 159964
rect 2092 159908 2096 159964
rect 2032 159904 2096 159908
rect 2112 159964 2176 159968
rect 2112 159908 2116 159964
rect 2116 159908 2172 159964
rect 2172 159908 2176 159964
rect 2112 159904 2176 159908
rect 2192 159964 2256 159968
rect 2192 159908 2196 159964
rect 2196 159908 2252 159964
rect 2252 159908 2256 159964
rect 2192 159904 2256 159908
rect 85952 159964 86016 159968
rect 85952 159908 85956 159964
rect 85956 159908 86012 159964
rect 86012 159908 86016 159964
rect 85952 159904 86016 159908
rect 86032 159964 86096 159968
rect 86032 159908 86036 159964
rect 86036 159908 86092 159964
rect 86092 159908 86096 159964
rect 86032 159904 86096 159908
rect 86112 159964 86176 159968
rect 86112 159908 86116 159964
rect 86116 159908 86172 159964
rect 86172 159908 86176 159964
rect 86112 159904 86176 159908
rect 86192 159964 86256 159968
rect 86192 159908 86196 159964
rect 86196 159908 86252 159964
rect 86252 159908 86256 159964
rect 86192 159904 86256 159908
rect 89952 159964 90016 159968
rect 89952 159908 89956 159964
rect 89956 159908 90012 159964
rect 90012 159908 90016 159964
rect 89952 159904 90016 159908
rect 90032 159964 90096 159968
rect 90032 159908 90036 159964
rect 90036 159908 90092 159964
rect 90092 159908 90096 159964
rect 90032 159904 90096 159908
rect 90112 159964 90176 159968
rect 90112 159908 90116 159964
rect 90116 159908 90172 159964
rect 90172 159908 90176 159964
rect 90112 159904 90176 159908
rect 90192 159964 90256 159968
rect 90192 159908 90196 159964
rect 90196 159908 90252 159964
rect 90252 159908 90256 159964
rect 90192 159904 90256 159908
rect 3952 159420 4016 159424
rect 3952 159364 3956 159420
rect 3956 159364 4012 159420
rect 4012 159364 4016 159420
rect 3952 159360 4016 159364
rect 4032 159420 4096 159424
rect 4032 159364 4036 159420
rect 4036 159364 4092 159420
rect 4092 159364 4096 159420
rect 4032 159360 4096 159364
rect 4112 159420 4176 159424
rect 4112 159364 4116 159420
rect 4116 159364 4172 159420
rect 4172 159364 4176 159420
rect 4112 159360 4176 159364
rect 4192 159420 4256 159424
rect 4192 159364 4196 159420
rect 4196 159364 4252 159420
rect 4252 159364 4256 159420
rect 4192 159360 4256 159364
rect 87952 159420 88016 159424
rect 87952 159364 87956 159420
rect 87956 159364 88012 159420
rect 88012 159364 88016 159420
rect 87952 159360 88016 159364
rect 88032 159420 88096 159424
rect 88032 159364 88036 159420
rect 88036 159364 88092 159420
rect 88092 159364 88096 159420
rect 88032 159360 88096 159364
rect 88112 159420 88176 159424
rect 88112 159364 88116 159420
rect 88116 159364 88172 159420
rect 88172 159364 88176 159420
rect 88112 159360 88176 159364
rect 88192 159420 88256 159424
rect 88192 159364 88196 159420
rect 88196 159364 88252 159420
rect 88252 159364 88256 159420
rect 88192 159360 88256 159364
rect 1952 158876 2016 158880
rect 1952 158820 1956 158876
rect 1956 158820 2012 158876
rect 2012 158820 2016 158876
rect 1952 158816 2016 158820
rect 2032 158876 2096 158880
rect 2032 158820 2036 158876
rect 2036 158820 2092 158876
rect 2092 158820 2096 158876
rect 2032 158816 2096 158820
rect 2112 158876 2176 158880
rect 2112 158820 2116 158876
rect 2116 158820 2172 158876
rect 2172 158820 2176 158876
rect 2112 158816 2176 158820
rect 2192 158876 2256 158880
rect 2192 158820 2196 158876
rect 2196 158820 2252 158876
rect 2252 158820 2256 158876
rect 2192 158816 2256 158820
rect 85952 158876 86016 158880
rect 85952 158820 85956 158876
rect 85956 158820 86012 158876
rect 86012 158820 86016 158876
rect 85952 158816 86016 158820
rect 86032 158876 86096 158880
rect 86032 158820 86036 158876
rect 86036 158820 86092 158876
rect 86092 158820 86096 158876
rect 86032 158816 86096 158820
rect 86112 158876 86176 158880
rect 86112 158820 86116 158876
rect 86116 158820 86172 158876
rect 86172 158820 86176 158876
rect 86112 158816 86176 158820
rect 86192 158876 86256 158880
rect 86192 158820 86196 158876
rect 86196 158820 86252 158876
rect 86252 158820 86256 158876
rect 86192 158816 86256 158820
rect 89952 158876 90016 158880
rect 89952 158820 89956 158876
rect 89956 158820 90012 158876
rect 90012 158820 90016 158876
rect 89952 158816 90016 158820
rect 90032 158876 90096 158880
rect 90032 158820 90036 158876
rect 90036 158820 90092 158876
rect 90092 158820 90096 158876
rect 90032 158816 90096 158820
rect 90112 158876 90176 158880
rect 90112 158820 90116 158876
rect 90116 158820 90172 158876
rect 90172 158820 90176 158876
rect 90112 158816 90176 158820
rect 90192 158876 90256 158880
rect 90192 158820 90196 158876
rect 90196 158820 90252 158876
rect 90252 158820 90256 158876
rect 90192 158816 90256 158820
rect 3952 158332 4016 158336
rect 3952 158276 3956 158332
rect 3956 158276 4012 158332
rect 4012 158276 4016 158332
rect 3952 158272 4016 158276
rect 4032 158332 4096 158336
rect 4032 158276 4036 158332
rect 4036 158276 4092 158332
rect 4092 158276 4096 158332
rect 4032 158272 4096 158276
rect 4112 158332 4176 158336
rect 4112 158276 4116 158332
rect 4116 158276 4172 158332
rect 4172 158276 4176 158332
rect 4112 158272 4176 158276
rect 4192 158332 4256 158336
rect 4192 158276 4196 158332
rect 4196 158276 4252 158332
rect 4252 158276 4256 158332
rect 4192 158272 4256 158276
rect 87952 158332 88016 158336
rect 87952 158276 87956 158332
rect 87956 158276 88012 158332
rect 88012 158276 88016 158332
rect 87952 158272 88016 158276
rect 88032 158332 88096 158336
rect 88032 158276 88036 158332
rect 88036 158276 88092 158332
rect 88092 158276 88096 158332
rect 88032 158272 88096 158276
rect 88112 158332 88176 158336
rect 88112 158276 88116 158332
rect 88116 158276 88172 158332
rect 88172 158276 88176 158332
rect 88112 158272 88176 158276
rect 88192 158332 88256 158336
rect 88192 158276 88196 158332
rect 88196 158276 88252 158332
rect 88252 158276 88256 158332
rect 88192 158272 88256 158276
rect 1952 157788 2016 157792
rect 1952 157732 1956 157788
rect 1956 157732 2012 157788
rect 2012 157732 2016 157788
rect 1952 157728 2016 157732
rect 2032 157788 2096 157792
rect 2032 157732 2036 157788
rect 2036 157732 2092 157788
rect 2092 157732 2096 157788
rect 2032 157728 2096 157732
rect 2112 157788 2176 157792
rect 2112 157732 2116 157788
rect 2116 157732 2172 157788
rect 2172 157732 2176 157788
rect 2112 157728 2176 157732
rect 2192 157788 2256 157792
rect 2192 157732 2196 157788
rect 2196 157732 2252 157788
rect 2252 157732 2256 157788
rect 2192 157728 2256 157732
rect 85952 157788 86016 157792
rect 85952 157732 85956 157788
rect 85956 157732 86012 157788
rect 86012 157732 86016 157788
rect 85952 157728 86016 157732
rect 86032 157788 86096 157792
rect 86032 157732 86036 157788
rect 86036 157732 86092 157788
rect 86092 157732 86096 157788
rect 86032 157728 86096 157732
rect 86112 157788 86176 157792
rect 86112 157732 86116 157788
rect 86116 157732 86172 157788
rect 86172 157732 86176 157788
rect 86112 157728 86176 157732
rect 86192 157788 86256 157792
rect 86192 157732 86196 157788
rect 86196 157732 86252 157788
rect 86252 157732 86256 157788
rect 86192 157728 86256 157732
rect 89952 157788 90016 157792
rect 89952 157732 89956 157788
rect 89956 157732 90012 157788
rect 90012 157732 90016 157788
rect 89952 157728 90016 157732
rect 90032 157788 90096 157792
rect 90032 157732 90036 157788
rect 90036 157732 90092 157788
rect 90092 157732 90096 157788
rect 90032 157728 90096 157732
rect 90112 157788 90176 157792
rect 90112 157732 90116 157788
rect 90116 157732 90172 157788
rect 90172 157732 90176 157788
rect 90112 157728 90176 157732
rect 90192 157788 90256 157792
rect 90192 157732 90196 157788
rect 90196 157732 90252 157788
rect 90252 157732 90256 157788
rect 90192 157728 90256 157732
rect 3952 157244 4016 157248
rect 3952 157188 3956 157244
rect 3956 157188 4012 157244
rect 4012 157188 4016 157244
rect 3952 157184 4016 157188
rect 4032 157244 4096 157248
rect 4032 157188 4036 157244
rect 4036 157188 4092 157244
rect 4092 157188 4096 157244
rect 4032 157184 4096 157188
rect 4112 157244 4176 157248
rect 4112 157188 4116 157244
rect 4116 157188 4172 157244
rect 4172 157188 4176 157244
rect 4112 157184 4176 157188
rect 4192 157244 4256 157248
rect 4192 157188 4196 157244
rect 4196 157188 4252 157244
rect 4252 157188 4256 157244
rect 4192 157184 4256 157188
rect 87952 157244 88016 157248
rect 87952 157188 87956 157244
rect 87956 157188 88012 157244
rect 88012 157188 88016 157244
rect 87952 157184 88016 157188
rect 88032 157244 88096 157248
rect 88032 157188 88036 157244
rect 88036 157188 88092 157244
rect 88092 157188 88096 157244
rect 88032 157184 88096 157188
rect 88112 157244 88176 157248
rect 88112 157188 88116 157244
rect 88116 157188 88172 157244
rect 88172 157188 88176 157244
rect 88112 157184 88176 157188
rect 88192 157244 88256 157248
rect 88192 157188 88196 157244
rect 88196 157188 88252 157244
rect 88252 157188 88256 157244
rect 88192 157184 88256 157188
rect 1952 156700 2016 156704
rect 1952 156644 1956 156700
rect 1956 156644 2012 156700
rect 2012 156644 2016 156700
rect 1952 156640 2016 156644
rect 2032 156700 2096 156704
rect 2032 156644 2036 156700
rect 2036 156644 2092 156700
rect 2092 156644 2096 156700
rect 2032 156640 2096 156644
rect 2112 156700 2176 156704
rect 2112 156644 2116 156700
rect 2116 156644 2172 156700
rect 2172 156644 2176 156700
rect 2112 156640 2176 156644
rect 2192 156700 2256 156704
rect 2192 156644 2196 156700
rect 2196 156644 2252 156700
rect 2252 156644 2256 156700
rect 2192 156640 2256 156644
rect 85952 156700 86016 156704
rect 85952 156644 85956 156700
rect 85956 156644 86012 156700
rect 86012 156644 86016 156700
rect 85952 156640 86016 156644
rect 86032 156700 86096 156704
rect 86032 156644 86036 156700
rect 86036 156644 86092 156700
rect 86092 156644 86096 156700
rect 86032 156640 86096 156644
rect 86112 156700 86176 156704
rect 86112 156644 86116 156700
rect 86116 156644 86172 156700
rect 86172 156644 86176 156700
rect 86112 156640 86176 156644
rect 86192 156700 86256 156704
rect 86192 156644 86196 156700
rect 86196 156644 86252 156700
rect 86252 156644 86256 156700
rect 86192 156640 86256 156644
rect 89952 156700 90016 156704
rect 89952 156644 89956 156700
rect 89956 156644 90012 156700
rect 90012 156644 90016 156700
rect 89952 156640 90016 156644
rect 90032 156700 90096 156704
rect 90032 156644 90036 156700
rect 90036 156644 90092 156700
rect 90092 156644 90096 156700
rect 90032 156640 90096 156644
rect 90112 156700 90176 156704
rect 90112 156644 90116 156700
rect 90116 156644 90172 156700
rect 90172 156644 90176 156700
rect 90112 156640 90176 156644
rect 90192 156700 90256 156704
rect 90192 156644 90196 156700
rect 90196 156644 90252 156700
rect 90252 156644 90256 156700
rect 90192 156640 90256 156644
rect 85804 156300 85868 156364
rect 3952 156156 4016 156160
rect 3952 156100 3956 156156
rect 3956 156100 4012 156156
rect 4012 156100 4016 156156
rect 3952 156096 4016 156100
rect 4032 156156 4096 156160
rect 4032 156100 4036 156156
rect 4036 156100 4092 156156
rect 4092 156100 4096 156156
rect 4032 156096 4096 156100
rect 4112 156156 4176 156160
rect 4112 156100 4116 156156
rect 4116 156100 4172 156156
rect 4172 156100 4176 156156
rect 4112 156096 4176 156100
rect 4192 156156 4256 156160
rect 4192 156100 4196 156156
rect 4196 156100 4252 156156
rect 4252 156100 4256 156156
rect 4192 156096 4256 156100
rect 87952 156156 88016 156160
rect 87952 156100 87956 156156
rect 87956 156100 88012 156156
rect 88012 156100 88016 156156
rect 87952 156096 88016 156100
rect 88032 156156 88096 156160
rect 88032 156100 88036 156156
rect 88036 156100 88092 156156
rect 88092 156100 88096 156156
rect 88032 156096 88096 156100
rect 88112 156156 88176 156160
rect 88112 156100 88116 156156
rect 88116 156100 88172 156156
rect 88172 156100 88176 156156
rect 88112 156096 88176 156100
rect 88192 156156 88256 156160
rect 88192 156100 88196 156156
rect 88196 156100 88252 156156
rect 88252 156100 88256 156156
rect 88192 156096 88256 156100
rect 1952 155612 2016 155616
rect 1952 155556 1956 155612
rect 1956 155556 2012 155612
rect 2012 155556 2016 155612
rect 1952 155552 2016 155556
rect 2032 155612 2096 155616
rect 2032 155556 2036 155612
rect 2036 155556 2092 155612
rect 2092 155556 2096 155612
rect 2032 155552 2096 155556
rect 2112 155612 2176 155616
rect 2112 155556 2116 155612
rect 2116 155556 2172 155612
rect 2172 155556 2176 155612
rect 2112 155552 2176 155556
rect 2192 155612 2256 155616
rect 2192 155556 2196 155612
rect 2196 155556 2252 155612
rect 2252 155556 2256 155612
rect 2192 155552 2256 155556
rect 85952 155612 86016 155616
rect 85952 155556 85956 155612
rect 85956 155556 86012 155612
rect 86012 155556 86016 155612
rect 85952 155552 86016 155556
rect 86032 155612 86096 155616
rect 86032 155556 86036 155612
rect 86036 155556 86092 155612
rect 86092 155556 86096 155612
rect 86032 155552 86096 155556
rect 86112 155612 86176 155616
rect 86112 155556 86116 155612
rect 86116 155556 86172 155612
rect 86172 155556 86176 155612
rect 86112 155552 86176 155556
rect 86192 155612 86256 155616
rect 86192 155556 86196 155612
rect 86196 155556 86252 155612
rect 86252 155556 86256 155612
rect 86192 155552 86256 155556
rect 89952 155612 90016 155616
rect 89952 155556 89956 155612
rect 89956 155556 90012 155612
rect 90012 155556 90016 155612
rect 89952 155552 90016 155556
rect 90032 155612 90096 155616
rect 90032 155556 90036 155612
rect 90036 155556 90092 155612
rect 90092 155556 90096 155612
rect 90032 155552 90096 155556
rect 90112 155612 90176 155616
rect 90112 155556 90116 155612
rect 90116 155556 90172 155612
rect 90172 155556 90176 155612
rect 90112 155552 90176 155556
rect 90192 155612 90256 155616
rect 90192 155556 90196 155612
rect 90196 155556 90252 155612
rect 90252 155556 90256 155612
rect 90192 155552 90256 155556
rect 3952 155068 4016 155072
rect 3952 155012 3956 155068
rect 3956 155012 4012 155068
rect 4012 155012 4016 155068
rect 3952 155008 4016 155012
rect 4032 155068 4096 155072
rect 4032 155012 4036 155068
rect 4036 155012 4092 155068
rect 4092 155012 4096 155068
rect 4032 155008 4096 155012
rect 4112 155068 4176 155072
rect 4112 155012 4116 155068
rect 4116 155012 4172 155068
rect 4172 155012 4176 155068
rect 4112 155008 4176 155012
rect 4192 155068 4256 155072
rect 4192 155012 4196 155068
rect 4196 155012 4252 155068
rect 4252 155012 4256 155068
rect 4192 155008 4256 155012
rect 87952 155068 88016 155072
rect 87952 155012 87956 155068
rect 87956 155012 88012 155068
rect 88012 155012 88016 155068
rect 87952 155008 88016 155012
rect 88032 155068 88096 155072
rect 88032 155012 88036 155068
rect 88036 155012 88092 155068
rect 88092 155012 88096 155068
rect 88032 155008 88096 155012
rect 88112 155068 88176 155072
rect 88112 155012 88116 155068
rect 88116 155012 88172 155068
rect 88172 155012 88176 155068
rect 88112 155008 88176 155012
rect 88192 155068 88256 155072
rect 88192 155012 88196 155068
rect 88196 155012 88252 155068
rect 88252 155012 88256 155068
rect 88192 155008 88256 155012
rect 1952 154524 2016 154528
rect 1952 154468 1956 154524
rect 1956 154468 2012 154524
rect 2012 154468 2016 154524
rect 1952 154464 2016 154468
rect 2032 154524 2096 154528
rect 2032 154468 2036 154524
rect 2036 154468 2092 154524
rect 2092 154468 2096 154524
rect 2032 154464 2096 154468
rect 2112 154524 2176 154528
rect 2112 154468 2116 154524
rect 2116 154468 2172 154524
rect 2172 154468 2176 154524
rect 2112 154464 2176 154468
rect 2192 154524 2256 154528
rect 2192 154468 2196 154524
rect 2196 154468 2252 154524
rect 2252 154468 2256 154524
rect 2192 154464 2256 154468
rect 85952 154524 86016 154528
rect 85952 154468 85956 154524
rect 85956 154468 86012 154524
rect 86012 154468 86016 154524
rect 85952 154464 86016 154468
rect 86032 154524 86096 154528
rect 86032 154468 86036 154524
rect 86036 154468 86092 154524
rect 86092 154468 86096 154524
rect 86032 154464 86096 154468
rect 86112 154524 86176 154528
rect 86112 154468 86116 154524
rect 86116 154468 86172 154524
rect 86172 154468 86176 154524
rect 86112 154464 86176 154468
rect 86192 154524 86256 154528
rect 86192 154468 86196 154524
rect 86196 154468 86252 154524
rect 86252 154468 86256 154524
rect 86192 154464 86256 154468
rect 89952 154524 90016 154528
rect 89952 154468 89956 154524
rect 89956 154468 90012 154524
rect 90012 154468 90016 154524
rect 89952 154464 90016 154468
rect 90032 154524 90096 154528
rect 90032 154468 90036 154524
rect 90036 154468 90092 154524
rect 90092 154468 90096 154524
rect 90032 154464 90096 154468
rect 90112 154524 90176 154528
rect 90112 154468 90116 154524
rect 90116 154468 90172 154524
rect 90172 154468 90176 154524
rect 90112 154464 90176 154468
rect 90192 154524 90256 154528
rect 90192 154468 90196 154524
rect 90196 154468 90252 154524
rect 90252 154468 90256 154524
rect 90192 154464 90256 154468
rect 84332 153988 84396 154052
rect 3952 153980 4016 153984
rect 3952 153924 3956 153980
rect 3956 153924 4012 153980
rect 4012 153924 4016 153980
rect 3952 153920 4016 153924
rect 4032 153980 4096 153984
rect 4032 153924 4036 153980
rect 4036 153924 4092 153980
rect 4092 153924 4096 153980
rect 4032 153920 4096 153924
rect 4112 153980 4176 153984
rect 4112 153924 4116 153980
rect 4116 153924 4172 153980
rect 4172 153924 4176 153980
rect 4112 153920 4176 153924
rect 4192 153980 4256 153984
rect 4192 153924 4196 153980
rect 4196 153924 4252 153980
rect 4252 153924 4256 153980
rect 4192 153920 4256 153924
rect 87952 153980 88016 153984
rect 87952 153924 87956 153980
rect 87956 153924 88012 153980
rect 88012 153924 88016 153980
rect 87952 153920 88016 153924
rect 88032 153980 88096 153984
rect 88032 153924 88036 153980
rect 88036 153924 88092 153980
rect 88092 153924 88096 153980
rect 88032 153920 88096 153924
rect 88112 153980 88176 153984
rect 88112 153924 88116 153980
rect 88116 153924 88172 153980
rect 88172 153924 88176 153980
rect 88112 153920 88176 153924
rect 88192 153980 88256 153984
rect 88192 153924 88196 153980
rect 88196 153924 88252 153980
rect 88252 153924 88256 153980
rect 88192 153920 88256 153924
rect 86540 153716 86604 153780
rect 1952 153436 2016 153440
rect 1952 153380 1956 153436
rect 1956 153380 2012 153436
rect 2012 153380 2016 153436
rect 1952 153376 2016 153380
rect 2032 153436 2096 153440
rect 2032 153380 2036 153436
rect 2036 153380 2092 153436
rect 2092 153380 2096 153436
rect 2032 153376 2096 153380
rect 2112 153436 2176 153440
rect 2112 153380 2116 153436
rect 2116 153380 2172 153436
rect 2172 153380 2176 153436
rect 2112 153376 2176 153380
rect 2192 153436 2256 153440
rect 2192 153380 2196 153436
rect 2196 153380 2252 153436
rect 2252 153380 2256 153436
rect 2192 153376 2256 153380
rect 85952 153436 86016 153440
rect 85952 153380 85956 153436
rect 85956 153380 86012 153436
rect 86012 153380 86016 153436
rect 85952 153376 86016 153380
rect 86032 153436 86096 153440
rect 86032 153380 86036 153436
rect 86036 153380 86092 153436
rect 86092 153380 86096 153436
rect 86032 153376 86096 153380
rect 86112 153436 86176 153440
rect 86112 153380 86116 153436
rect 86116 153380 86172 153436
rect 86172 153380 86176 153436
rect 86112 153376 86176 153380
rect 86192 153436 86256 153440
rect 86192 153380 86196 153436
rect 86196 153380 86252 153436
rect 86252 153380 86256 153436
rect 86192 153376 86256 153380
rect 89952 153436 90016 153440
rect 89952 153380 89956 153436
rect 89956 153380 90012 153436
rect 90012 153380 90016 153436
rect 89952 153376 90016 153380
rect 90032 153436 90096 153440
rect 90032 153380 90036 153436
rect 90036 153380 90092 153436
rect 90092 153380 90096 153436
rect 90032 153376 90096 153380
rect 90112 153436 90176 153440
rect 90112 153380 90116 153436
rect 90116 153380 90172 153436
rect 90172 153380 90176 153436
rect 90112 153376 90176 153380
rect 90192 153436 90256 153440
rect 90192 153380 90196 153436
rect 90196 153380 90252 153436
rect 90252 153380 90256 153436
rect 90192 153376 90256 153380
rect 3952 152892 4016 152896
rect 3952 152836 3956 152892
rect 3956 152836 4012 152892
rect 4012 152836 4016 152892
rect 3952 152832 4016 152836
rect 4032 152892 4096 152896
rect 4032 152836 4036 152892
rect 4036 152836 4092 152892
rect 4092 152836 4096 152892
rect 4032 152832 4096 152836
rect 4112 152892 4176 152896
rect 4112 152836 4116 152892
rect 4116 152836 4172 152892
rect 4172 152836 4176 152892
rect 4112 152832 4176 152836
rect 4192 152892 4256 152896
rect 4192 152836 4196 152892
rect 4196 152836 4252 152892
rect 4252 152836 4256 152892
rect 4192 152832 4256 152836
rect 87952 152892 88016 152896
rect 87952 152836 87956 152892
rect 87956 152836 88012 152892
rect 88012 152836 88016 152892
rect 87952 152832 88016 152836
rect 88032 152892 88096 152896
rect 88032 152836 88036 152892
rect 88036 152836 88092 152892
rect 88092 152836 88096 152892
rect 88032 152832 88096 152836
rect 88112 152892 88176 152896
rect 88112 152836 88116 152892
rect 88116 152836 88172 152892
rect 88172 152836 88176 152892
rect 88112 152832 88176 152836
rect 88192 152892 88256 152896
rect 88192 152836 88196 152892
rect 88196 152836 88252 152892
rect 88252 152836 88256 152892
rect 88192 152832 88256 152836
rect 1952 152348 2016 152352
rect 1952 152292 1956 152348
rect 1956 152292 2012 152348
rect 2012 152292 2016 152348
rect 1952 152288 2016 152292
rect 2032 152348 2096 152352
rect 2032 152292 2036 152348
rect 2036 152292 2092 152348
rect 2092 152292 2096 152348
rect 2032 152288 2096 152292
rect 2112 152348 2176 152352
rect 2112 152292 2116 152348
rect 2116 152292 2172 152348
rect 2172 152292 2176 152348
rect 2112 152288 2176 152292
rect 2192 152348 2256 152352
rect 2192 152292 2196 152348
rect 2196 152292 2252 152348
rect 2252 152292 2256 152348
rect 2192 152288 2256 152292
rect 85952 152348 86016 152352
rect 85952 152292 85956 152348
rect 85956 152292 86012 152348
rect 86012 152292 86016 152348
rect 85952 152288 86016 152292
rect 86032 152348 86096 152352
rect 86032 152292 86036 152348
rect 86036 152292 86092 152348
rect 86092 152292 86096 152348
rect 86032 152288 86096 152292
rect 86112 152348 86176 152352
rect 86112 152292 86116 152348
rect 86116 152292 86172 152348
rect 86172 152292 86176 152348
rect 86112 152288 86176 152292
rect 86192 152348 86256 152352
rect 86192 152292 86196 152348
rect 86196 152292 86252 152348
rect 86252 152292 86256 152348
rect 86192 152288 86256 152292
rect 89952 152348 90016 152352
rect 89952 152292 89956 152348
rect 89956 152292 90012 152348
rect 90012 152292 90016 152348
rect 89952 152288 90016 152292
rect 90032 152348 90096 152352
rect 90032 152292 90036 152348
rect 90036 152292 90092 152348
rect 90092 152292 90096 152348
rect 90032 152288 90096 152292
rect 90112 152348 90176 152352
rect 90112 152292 90116 152348
rect 90116 152292 90172 152348
rect 90172 152292 90176 152348
rect 90112 152288 90176 152292
rect 90192 152348 90256 152352
rect 90192 152292 90196 152348
rect 90196 152292 90252 152348
rect 90252 152292 90256 152348
rect 90192 152288 90256 152292
rect 3952 151804 4016 151808
rect 3952 151748 3956 151804
rect 3956 151748 4012 151804
rect 4012 151748 4016 151804
rect 3952 151744 4016 151748
rect 4032 151804 4096 151808
rect 4032 151748 4036 151804
rect 4036 151748 4092 151804
rect 4092 151748 4096 151804
rect 4032 151744 4096 151748
rect 4112 151804 4176 151808
rect 4112 151748 4116 151804
rect 4116 151748 4172 151804
rect 4172 151748 4176 151804
rect 4112 151744 4176 151748
rect 4192 151804 4256 151808
rect 4192 151748 4196 151804
rect 4196 151748 4252 151804
rect 4252 151748 4256 151804
rect 4192 151744 4256 151748
rect 87952 151804 88016 151808
rect 87952 151748 87956 151804
rect 87956 151748 88012 151804
rect 88012 151748 88016 151804
rect 87952 151744 88016 151748
rect 88032 151804 88096 151808
rect 88032 151748 88036 151804
rect 88036 151748 88092 151804
rect 88092 151748 88096 151804
rect 88032 151744 88096 151748
rect 88112 151804 88176 151808
rect 88112 151748 88116 151804
rect 88116 151748 88172 151804
rect 88172 151748 88176 151804
rect 88112 151744 88176 151748
rect 88192 151804 88256 151808
rect 88192 151748 88196 151804
rect 88196 151748 88252 151804
rect 88252 151748 88256 151804
rect 88192 151744 88256 151748
rect 1952 151260 2016 151264
rect 1952 151204 1956 151260
rect 1956 151204 2012 151260
rect 2012 151204 2016 151260
rect 1952 151200 2016 151204
rect 2032 151260 2096 151264
rect 2032 151204 2036 151260
rect 2036 151204 2092 151260
rect 2092 151204 2096 151260
rect 2032 151200 2096 151204
rect 2112 151260 2176 151264
rect 2112 151204 2116 151260
rect 2116 151204 2172 151260
rect 2172 151204 2176 151260
rect 2112 151200 2176 151204
rect 2192 151260 2256 151264
rect 2192 151204 2196 151260
rect 2196 151204 2252 151260
rect 2252 151204 2256 151260
rect 2192 151200 2256 151204
rect 85952 151260 86016 151264
rect 85952 151204 85956 151260
rect 85956 151204 86012 151260
rect 86012 151204 86016 151260
rect 85952 151200 86016 151204
rect 86032 151260 86096 151264
rect 86032 151204 86036 151260
rect 86036 151204 86092 151260
rect 86092 151204 86096 151260
rect 86032 151200 86096 151204
rect 86112 151260 86176 151264
rect 86112 151204 86116 151260
rect 86116 151204 86172 151260
rect 86172 151204 86176 151260
rect 86112 151200 86176 151204
rect 86192 151260 86256 151264
rect 86192 151204 86196 151260
rect 86196 151204 86252 151260
rect 86252 151204 86256 151260
rect 86192 151200 86256 151204
rect 89952 151260 90016 151264
rect 89952 151204 89956 151260
rect 89956 151204 90012 151260
rect 90012 151204 90016 151260
rect 89952 151200 90016 151204
rect 90032 151260 90096 151264
rect 90032 151204 90036 151260
rect 90036 151204 90092 151260
rect 90092 151204 90096 151260
rect 90032 151200 90096 151204
rect 90112 151260 90176 151264
rect 90112 151204 90116 151260
rect 90116 151204 90172 151260
rect 90172 151204 90176 151260
rect 90112 151200 90176 151204
rect 90192 151260 90256 151264
rect 90192 151204 90196 151260
rect 90196 151204 90252 151260
rect 90252 151204 90256 151260
rect 90192 151200 90256 151204
rect 3952 150716 4016 150720
rect 3952 150660 3956 150716
rect 3956 150660 4012 150716
rect 4012 150660 4016 150716
rect 3952 150656 4016 150660
rect 4032 150716 4096 150720
rect 4032 150660 4036 150716
rect 4036 150660 4092 150716
rect 4092 150660 4096 150716
rect 4032 150656 4096 150660
rect 4112 150716 4176 150720
rect 4112 150660 4116 150716
rect 4116 150660 4172 150716
rect 4172 150660 4176 150716
rect 4112 150656 4176 150660
rect 4192 150716 4256 150720
rect 4192 150660 4196 150716
rect 4196 150660 4252 150716
rect 4252 150660 4256 150716
rect 4192 150656 4256 150660
rect 87952 150716 88016 150720
rect 87952 150660 87956 150716
rect 87956 150660 88012 150716
rect 88012 150660 88016 150716
rect 87952 150656 88016 150660
rect 88032 150716 88096 150720
rect 88032 150660 88036 150716
rect 88036 150660 88092 150716
rect 88092 150660 88096 150716
rect 88032 150656 88096 150660
rect 88112 150716 88176 150720
rect 88112 150660 88116 150716
rect 88116 150660 88172 150716
rect 88172 150660 88176 150716
rect 88112 150656 88176 150660
rect 88192 150716 88256 150720
rect 88192 150660 88196 150716
rect 88196 150660 88252 150716
rect 88252 150660 88256 150716
rect 88192 150656 88256 150660
rect 1952 150172 2016 150176
rect 1952 150116 1956 150172
rect 1956 150116 2012 150172
rect 2012 150116 2016 150172
rect 1952 150112 2016 150116
rect 2032 150172 2096 150176
rect 2032 150116 2036 150172
rect 2036 150116 2092 150172
rect 2092 150116 2096 150172
rect 2032 150112 2096 150116
rect 2112 150172 2176 150176
rect 2112 150116 2116 150172
rect 2116 150116 2172 150172
rect 2172 150116 2176 150172
rect 2112 150112 2176 150116
rect 2192 150172 2256 150176
rect 2192 150116 2196 150172
rect 2196 150116 2252 150172
rect 2252 150116 2256 150172
rect 2192 150112 2256 150116
rect 85952 150172 86016 150176
rect 85952 150116 85956 150172
rect 85956 150116 86012 150172
rect 86012 150116 86016 150172
rect 85952 150112 86016 150116
rect 86032 150172 86096 150176
rect 86032 150116 86036 150172
rect 86036 150116 86092 150172
rect 86092 150116 86096 150172
rect 86032 150112 86096 150116
rect 86112 150172 86176 150176
rect 86112 150116 86116 150172
rect 86116 150116 86172 150172
rect 86172 150116 86176 150172
rect 86112 150112 86176 150116
rect 86192 150172 86256 150176
rect 86192 150116 86196 150172
rect 86196 150116 86252 150172
rect 86252 150116 86256 150172
rect 86192 150112 86256 150116
rect 89952 150172 90016 150176
rect 89952 150116 89956 150172
rect 89956 150116 90012 150172
rect 90012 150116 90016 150172
rect 89952 150112 90016 150116
rect 90032 150172 90096 150176
rect 90032 150116 90036 150172
rect 90036 150116 90092 150172
rect 90092 150116 90096 150172
rect 90032 150112 90096 150116
rect 90112 150172 90176 150176
rect 90112 150116 90116 150172
rect 90116 150116 90172 150172
rect 90172 150116 90176 150172
rect 90112 150112 90176 150116
rect 90192 150172 90256 150176
rect 90192 150116 90196 150172
rect 90196 150116 90252 150172
rect 90252 150116 90256 150172
rect 90192 150112 90256 150116
rect 3952 149628 4016 149632
rect 3952 149572 3956 149628
rect 3956 149572 4012 149628
rect 4012 149572 4016 149628
rect 3952 149568 4016 149572
rect 4032 149628 4096 149632
rect 4032 149572 4036 149628
rect 4036 149572 4092 149628
rect 4092 149572 4096 149628
rect 4032 149568 4096 149572
rect 4112 149628 4176 149632
rect 4112 149572 4116 149628
rect 4116 149572 4172 149628
rect 4172 149572 4176 149628
rect 4112 149568 4176 149572
rect 4192 149628 4256 149632
rect 4192 149572 4196 149628
rect 4196 149572 4252 149628
rect 4252 149572 4256 149628
rect 4192 149568 4256 149572
rect 87952 149628 88016 149632
rect 87952 149572 87956 149628
rect 87956 149572 88012 149628
rect 88012 149572 88016 149628
rect 87952 149568 88016 149572
rect 88032 149628 88096 149632
rect 88032 149572 88036 149628
rect 88036 149572 88092 149628
rect 88092 149572 88096 149628
rect 88032 149568 88096 149572
rect 88112 149628 88176 149632
rect 88112 149572 88116 149628
rect 88116 149572 88172 149628
rect 88172 149572 88176 149628
rect 88112 149568 88176 149572
rect 88192 149628 88256 149632
rect 88192 149572 88196 149628
rect 88196 149572 88252 149628
rect 88252 149572 88256 149628
rect 88192 149568 88256 149572
rect 1952 149084 2016 149088
rect 1952 149028 1956 149084
rect 1956 149028 2012 149084
rect 2012 149028 2016 149084
rect 1952 149024 2016 149028
rect 2032 149084 2096 149088
rect 2032 149028 2036 149084
rect 2036 149028 2092 149084
rect 2092 149028 2096 149084
rect 2032 149024 2096 149028
rect 2112 149084 2176 149088
rect 2112 149028 2116 149084
rect 2116 149028 2172 149084
rect 2172 149028 2176 149084
rect 2112 149024 2176 149028
rect 2192 149084 2256 149088
rect 2192 149028 2196 149084
rect 2196 149028 2252 149084
rect 2252 149028 2256 149084
rect 2192 149024 2256 149028
rect 85952 149084 86016 149088
rect 85952 149028 85956 149084
rect 85956 149028 86012 149084
rect 86012 149028 86016 149084
rect 85952 149024 86016 149028
rect 86032 149084 86096 149088
rect 86032 149028 86036 149084
rect 86036 149028 86092 149084
rect 86092 149028 86096 149084
rect 86032 149024 86096 149028
rect 86112 149084 86176 149088
rect 86112 149028 86116 149084
rect 86116 149028 86172 149084
rect 86172 149028 86176 149084
rect 86112 149024 86176 149028
rect 86192 149084 86256 149088
rect 86192 149028 86196 149084
rect 86196 149028 86252 149084
rect 86252 149028 86256 149084
rect 86192 149024 86256 149028
rect 89952 149084 90016 149088
rect 89952 149028 89956 149084
rect 89956 149028 90012 149084
rect 90012 149028 90016 149084
rect 89952 149024 90016 149028
rect 90032 149084 90096 149088
rect 90032 149028 90036 149084
rect 90036 149028 90092 149084
rect 90092 149028 90096 149084
rect 90032 149024 90096 149028
rect 90112 149084 90176 149088
rect 90112 149028 90116 149084
rect 90116 149028 90172 149084
rect 90172 149028 90176 149084
rect 90112 149024 90176 149028
rect 90192 149084 90256 149088
rect 90192 149028 90196 149084
rect 90196 149028 90252 149084
rect 90252 149028 90256 149084
rect 90192 149024 90256 149028
rect 3952 148540 4016 148544
rect 3952 148484 3956 148540
rect 3956 148484 4012 148540
rect 4012 148484 4016 148540
rect 3952 148480 4016 148484
rect 4032 148540 4096 148544
rect 4032 148484 4036 148540
rect 4036 148484 4092 148540
rect 4092 148484 4096 148540
rect 4032 148480 4096 148484
rect 4112 148540 4176 148544
rect 4112 148484 4116 148540
rect 4116 148484 4172 148540
rect 4172 148484 4176 148540
rect 4112 148480 4176 148484
rect 4192 148540 4256 148544
rect 4192 148484 4196 148540
rect 4196 148484 4252 148540
rect 4252 148484 4256 148540
rect 4192 148480 4256 148484
rect 87952 148540 88016 148544
rect 87952 148484 87956 148540
rect 87956 148484 88012 148540
rect 88012 148484 88016 148540
rect 87952 148480 88016 148484
rect 88032 148540 88096 148544
rect 88032 148484 88036 148540
rect 88036 148484 88092 148540
rect 88092 148484 88096 148540
rect 88032 148480 88096 148484
rect 88112 148540 88176 148544
rect 88112 148484 88116 148540
rect 88116 148484 88172 148540
rect 88172 148484 88176 148540
rect 88112 148480 88176 148484
rect 88192 148540 88256 148544
rect 88192 148484 88196 148540
rect 88196 148484 88252 148540
rect 88252 148484 88256 148540
rect 88192 148480 88256 148484
rect 1952 147996 2016 148000
rect 1952 147940 1956 147996
rect 1956 147940 2012 147996
rect 2012 147940 2016 147996
rect 1952 147936 2016 147940
rect 2032 147996 2096 148000
rect 2032 147940 2036 147996
rect 2036 147940 2092 147996
rect 2092 147940 2096 147996
rect 2032 147936 2096 147940
rect 2112 147996 2176 148000
rect 2112 147940 2116 147996
rect 2116 147940 2172 147996
rect 2172 147940 2176 147996
rect 2112 147936 2176 147940
rect 2192 147996 2256 148000
rect 2192 147940 2196 147996
rect 2196 147940 2252 147996
rect 2252 147940 2256 147996
rect 2192 147936 2256 147940
rect 85952 147996 86016 148000
rect 85952 147940 85956 147996
rect 85956 147940 86012 147996
rect 86012 147940 86016 147996
rect 85952 147936 86016 147940
rect 86032 147996 86096 148000
rect 86032 147940 86036 147996
rect 86036 147940 86092 147996
rect 86092 147940 86096 147996
rect 86032 147936 86096 147940
rect 86112 147996 86176 148000
rect 86112 147940 86116 147996
rect 86116 147940 86172 147996
rect 86172 147940 86176 147996
rect 86112 147936 86176 147940
rect 86192 147996 86256 148000
rect 86192 147940 86196 147996
rect 86196 147940 86252 147996
rect 86252 147940 86256 147996
rect 86192 147936 86256 147940
rect 89952 147996 90016 148000
rect 89952 147940 89956 147996
rect 89956 147940 90012 147996
rect 90012 147940 90016 147996
rect 89952 147936 90016 147940
rect 90032 147996 90096 148000
rect 90032 147940 90036 147996
rect 90036 147940 90092 147996
rect 90092 147940 90096 147996
rect 90032 147936 90096 147940
rect 90112 147996 90176 148000
rect 90112 147940 90116 147996
rect 90116 147940 90172 147996
rect 90172 147940 90176 147996
rect 90112 147936 90176 147940
rect 90192 147996 90256 148000
rect 90192 147940 90196 147996
rect 90196 147940 90252 147996
rect 90252 147940 90256 147996
rect 90192 147936 90256 147940
rect 86908 147596 86972 147660
rect 3952 147452 4016 147456
rect 3952 147396 3956 147452
rect 3956 147396 4012 147452
rect 4012 147396 4016 147452
rect 3952 147392 4016 147396
rect 4032 147452 4096 147456
rect 4032 147396 4036 147452
rect 4036 147396 4092 147452
rect 4092 147396 4096 147452
rect 4032 147392 4096 147396
rect 4112 147452 4176 147456
rect 4112 147396 4116 147452
rect 4116 147396 4172 147452
rect 4172 147396 4176 147452
rect 4112 147392 4176 147396
rect 4192 147452 4256 147456
rect 4192 147396 4196 147452
rect 4196 147396 4252 147452
rect 4252 147396 4256 147452
rect 4192 147392 4256 147396
rect 87952 147452 88016 147456
rect 87952 147396 87956 147452
rect 87956 147396 88012 147452
rect 88012 147396 88016 147452
rect 87952 147392 88016 147396
rect 88032 147452 88096 147456
rect 88032 147396 88036 147452
rect 88036 147396 88092 147452
rect 88092 147396 88096 147452
rect 88032 147392 88096 147396
rect 88112 147452 88176 147456
rect 88112 147396 88116 147452
rect 88116 147396 88172 147452
rect 88172 147396 88176 147452
rect 88112 147392 88176 147396
rect 88192 147452 88256 147456
rect 88192 147396 88196 147452
rect 88196 147396 88252 147452
rect 88252 147396 88256 147452
rect 88192 147392 88256 147396
rect 1952 146908 2016 146912
rect 1952 146852 1956 146908
rect 1956 146852 2012 146908
rect 2012 146852 2016 146908
rect 1952 146848 2016 146852
rect 2032 146908 2096 146912
rect 2032 146852 2036 146908
rect 2036 146852 2092 146908
rect 2092 146852 2096 146908
rect 2032 146848 2096 146852
rect 2112 146908 2176 146912
rect 2112 146852 2116 146908
rect 2116 146852 2172 146908
rect 2172 146852 2176 146908
rect 2112 146848 2176 146852
rect 2192 146908 2256 146912
rect 2192 146852 2196 146908
rect 2196 146852 2252 146908
rect 2252 146852 2256 146908
rect 2192 146848 2256 146852
rect 85952 146908 86016 146912
rect 85952 146852 85956 146908
rect 85956 146852 86012 146908
rect 86012 146852 86016 146908
rect 85952 146848 86016 146852
rect 86032 146908 86096 146912
rect 86032 146852 86036 146908
rect 86036 146852 86092 146908
rect 86092 146852 86096 146908
rect 86032 146848 86096 146852
rect 86112 146908 86176 146912
rect 86112 146852 86116 146908
rect 86116 146852 86172 146908
rect 86172 146852 86176 146908
rect 86112 146848 86176 146852
rect 86192 146908 86256 146912
rect 86192 146852 86196 146908
rect 86196 146852 86252 146908
rect 86252 146852 86256 146908
rect 86192 146848 86256 146852
rect 89952 146908 90016 146912
rect 89952 146852 89956 146908
rect 89956 146852 90012 146908
rect 90012 146852 90016 146908
rect 89952 146848 90016 146852
rect 90032 146908 90096 146912
rect 90032 146852 90036 146908
rect 90036 146852 90092 146908
rect 90092 146852 90096 146908
rect 90032 146848 90096 146852
rect 90112 146908 90176 146912
rect 90112 146852 90116 146908
rect 90116 146852 90172 146908
rect 90172 146852 90176 146908
rect 90112 146848 90176 146852
rect 90192 146908 90256 146912
rect 90192 146852 90196 146908
rect 90196 146852 90252 146908
rect 90252 146852 90256 146908
rect 90192 146848 90256 146852
rect 3952 146364 4016 146368
rect 3952 146308 3956 146364
rect 3956 146308 4012 146364
rect 4012 146308 4016 146364
rect 3952 146304 4016 146308
rect 4032 146364 4096 146368
rect 4032 146308 4036 146364
rect 4036 146308 4092 146364
rect 4092 146308 4096 146364
rect 4032 146304 4096 146308
rect 4112 146364 4176 146368
rect 4112 146308 4116 146364
rect 4116 146308 4172 146364
rect 4172 146308 4176 146364
rect 4112 146304 4176 146308
rect 4192 146364 4256 146368
rect 4192 146308 4196 146364
rect 4196 146308 4252 146364
rect 4252 146308 4256 146364
rect 4192 146304 4256 146308
rect 87952 146364 88016 146368
rect 87952 146308 87956 146364
rect 87956 146308 88012 146364
rect 88012 146308 88016 146364
rect 87952 146304 88016 146308
rect 88032 146364 88096 146368
rect 88032 146308 88036 146364
rect 88036 146308 88092 146364
rect 88092 146308 88096 146364
rect 88032 146304 88096 146308
rect 88112 146364 88176 146368
rect 88112 146308 88116 146364
rect 88116 146308 88172 146364
rect 88172 146308 88176 146364
rect 88112 146304 88176 146308
rect 88192 146364 88256 146368
rect 88192 146308 88196 146364
rect 88196 146308 88252 146364
rect 88252 146308 88256 146364
rect 88192 146304 88256 146308
rect 1952 145820 2016 145824
rect 1952 145764 1956 145820
rect 1956 145764 2012 145820
rect 2012 145764 2016 145820
rect 1952 145760 2016 145764
rect 2032 145820 2096 145824
rect 2032 145764 2036 145820
rect 2036 145764 2092 145820
rect 2092 145764 2096 145820
rect 2032 145760 2096 145764
rect 2112 145820 2176 145824
rect 2112 145764 2116 145820
rect 2116 145764 2172 145820
rect 2172 145764 2176 145820
rect 2112 145760 2176 145764
rect 2192 145820 2256 145824
rect 2192 145764 2196 145820
rect 2196 145764 2252 145820
rect 2252 145764 2256 145820
rect 2192 145760 2256 145764
rect 85952 145820 86016 145824
rect 85952 145764 85956 145820
rect 85956 145764 86012 145820
rect 86012 145764 86016 145820
rect 85952 145760 86016 145764
rect 86032 145820 86096 145824
rect 86032 145764 86036 145820
rect 86036 145764 86092 145820
rect 86092 145764 86096 145820
rect 86032 145760 86096 145764
rect 86112 145820 86176 145824
rect 86112 145764 86116 145820
rect 86116 145764 86172 145820
rect 86172 145764 86176 145820
rect 86112 145760 86176 145764
rect 86192 145820 86256 145824
rect 86192 145764 86196 145820
rect 86196 145764 86252 145820
rect 86252 145764 86256 145820
rect 86192 145760 86256 145764
rect 89952 145820 90016 145824
rect 89952 145764 89956 145820
rect 89956 145764 90012 145820
rect 90012 145764 90016 145820
rect 89952 145760 90016 145764
rect 90032 145820 90096 145824
rect 90032 145764 90036 145820
rect 90036 145764 90092 145820
rect 90092 145764 90096 145820
rect 90032 145760 90096 145764
rect 90112 145820 90176 145824
rect 90112 145764 90116 145820
rect 90116 145764 90172 145820
rect 90172 145764 90176 145820
rect 90112 145760 90176 145764
rect 90192 145820 90256 145824
rect 90192 145764 90196 145820
rect 90196 145764 90252 145820
rect 90252 145764 90256 145820
rect 90192 145760 90256 145764
rect 3952 145276 4016 145280
rect 3952 145220 3956 145276
rect 3956 145220 4012 145276
rect 4012 145220 4016 145276
rect 3952 145216 4016 145220
rect 4032 145276 4096 145280
rect 4032 145220 4036 145276
rect 4036 145220 4092 145276
rect 4092 145220 4096 145276
rect 4032 145216 4096 145220
rect 4112 145276 4176 145280
rect 4112 145220 4116 145276
rect 4116 145220 4172 145276
rect 4172 145220 4176 145276
rect 4112 145216 4176 145220
rect 4192 145276 4256 145280
rect 4192 145220 4196 145276
rect 4196 145220 4252 145276
rect 4252 145220 4256 145276
rect 4192 145216 4256 145220
rect 87952 145276 88016 145280
rect 87952 145220 87956 145276
rect 87956 145220 88012 145276
rect 88012 145220 88016 145276
rect 87952 145216 88016 145220
rect 88032 145276 88096 145280
rect 88032 145220 88036 145276
rect 88036 145220 88092 145276
rect 88092 145220 88096 145276
rect 88032 145216 88096 145220
rect 88112 145276 88176 145280
rect 88112 145220 88116 145276
rect 88116 145220 88172 145276
rect 88172 145220 88176 145276
rect 88112 145216 88176 145220
rect 88192 145276 88256 145280
rect 88192 145220 88196 145276
rect 88196 145220 88252 145276
rect 88252 145220 88256 145276
rect 88192 145216 88256 145220
rect 1952 144732 2016 144736
rect 1952 144676 1956 144732
rect 1956 144676 2012 144732
rect 2012 144676 2016 144732
rect 1952 144672 2016 144676
rect 2032 144732 2096 144736
rect 2032 144676 2036 144732
rect 2036 144676 2092 144732
rect 2092 144676 2096 144732
rect 2032 144672 2096 144676
rect 2112 144732 2176 144736
rect 2112 144676 2116 144732
rect 2116 144676 2172 144732
rect 2172 144676 2176 144732
rect 2112 144672 2176 144676
rect 2192 144732 2256 144736
rect 2192 144676 2196 144732
rect 2196 144676 2252 144732
rect 2252 144676 2256 144732
rect 2192 144672 2256 144676
rect 85952 144732 86016 144736
rect 85952 144676 85956 144732
rect 85956 144676 86012 144732
rect 86012 144676 86016 144732
rect 85952 144672 86016 144676
rect 86032 144732 86096 144736
rect 86032 144676 86036 144732
rect 86036 144676 86092 144732
rect 86092 144676 86096 144732
rect 86032 144672 86096 144676
rect 86112 144732 86176 144736
rect 86112 144676 86116 144732
rect 86116 144676 86172 144732
rect 86172 144676 86176 144732
rect 86112 144672 86176 144676
rect 86192 144732 86256 144736
rect 86192 144676 86196 144732
rect 86196 144676 86252 144732
rect 86252 144676 86256 144732
rect 86192 144672 86256 144676
rect 89952 144732 90016 144736
rect 89952 144676 89956 144732
rect 89956 144676 90012 144732
rect 90012 144676 90016 144732
rect 89952 144672 90016 144676
rect 90032 144732 90096 144736
rect 90032 144676 90036 144732
rect 90036 144676 90092 144732
rect 90092 144676 90096 144732
rect 90032 144672 90096 144676
rect 90112 144732 90176 144736
rect 90112 144676 90116 144732
rect 90116 144676 90172 144732
rect 90172 144676 90176 144732
rect 90112 144672 90176 144676
rect 90192 144732 90256 144736
rect 90192 144676 90196 144732
rect 90196 144676 90252 144732
rect 90252 144676 90256 144732
rect 90192 144672 90256 144676
rect 3952 144188 4016 144192
rect 3952 144132 3956 144188
rect 3956 144132 4012 144188
rect 4012 144132 4016 144188
rect 3952 144128 4016 144132
rect 4032 144188 4096 144192
rect 4032 144132 4036 144188
rect 4036 144132 4092 144188
rect 4092 144132 4096 144188
rect 4032 144128 4096 144132
rect 4112 144188 4176 144192
rect 4112 144132 4116 144188
rect 4116 144132 4172 144188
rect 4172 144132 4176 144188
rect 4112 144128 4176 144132
rect 4192 144188 4256 144192
rect 4192 144132 4196 144188
rect 4196 144132 4252 144188
rect 4252 144132 4256 144188
rect 4192 144128 4256 144132
rect 87952 144188 88016 144192
rect 87952 144132 87956 144188
rect 87956 144132 88012 144188
rect 88012 144132 88016 144188
rect 87952 144128 88016 144132
rect 88032 144188 88096 144192
rect 88032 144132 88036 144188
rect 88036 144132 88092 144188
rect 88092 144132 88096 144188
rect 88032 144128 88096 144132
rect 88112 144188 88176 144192
rect 88112 144132 88116 144188
rect 88116 144132 88172 144188
rect 88172 144132 88176 144188
rect 88112 144128 88176 144132
rect 88192 144188 88256 144192
rect 88192 144132 88196 144188
rect 88196 144132 88252 144188
rect 88252 144132 88256 144188
rect 88192 144128 88256 144132
rect 1952 143644 2016 143648
rect 1952 143588 1956 143644
rect 1956 143588 2012 143644
rect 2012 143588 2016 143644
rect 1952 143584 2016 143588
rect 2032 143644 2096 143648
rect 2032 143588 2036 143644
rect 2036 143588 2092 143644
rect 2092 143588 2096 143644
rect 2032 143584 2096 143588
rect 2112 143644 2176 143648
rect 2112 143588 2116 143644
rect 2116 143588 2172 143644
rect 2172 143588 2176 143644
rect 2112 143584 2176 143588
rect 2192 143644 2256 143648
rect 2192 143588 2196 143644
rect 2196 143588 2252 143644
rect 2252 143588 2256 143644
rect 2192 143584 2256 143588
rect 85952 143644 86016 143648
rect 85952 143588 85956 143644
rect 85956 143588 86012 143644
rect 86012 143588 86016 143644
rect 85952 143584 86016 143588
rect 86032 143644 86096 143648
rect 86032 143588 86036 143644
rect 86036 143588 86092 143644
rect 86092 143588 86096 143644
rect 86032 143584 86096 143588
rect 86112 143644 86176 143648
rect 86112 143588 86116 143644
rect 86116 143588 86172 143644
rect 86172 143588 86176 143644
rect 86112 143584 86176 143588
rect 86192 143644 86256 143648
rect 86192 143588 86196 143644
rect 86196 143588 86252 143644
rect 86252 143588 86256 143644
rect 86192 143584 86256 143588
rect 89952 143644 90016 143648
rect 89952 143588 89956 143644
rect 89956 143588 90012 143644
rect 90012 143588 90016 143644
rect 89952 143584 90016 143588
rect 90032 143644 90096 143648
rect 90032 143588 90036 143644
rect 90036 143588 90092 143644
rect 90092 143588 90096 143644
rect 90032 143584 90096 143588
rect 90112 143644 90176 143648
rect 90112 143588 90116 143644
rect 90116 143588 90172 143644
rect 90172 143588 90176 143644
rect 90112 143584 90176 143588
rect 90192 143644 90256 143648
rect 90192 143588 90196 143644
rect 90196 143588 90252 143644
rect 90252 143588 90256 143644
rect 90192 143584 90256 143588
rect 3952 143100 4016 143104
rect 3952 143044 3956 143100
rect 3956 143044 4012 143100
rect 4012 143044 4016 143100
rect 3952 143040 4016 143044
rect 4032 143100 4096 143104
rect 4032 143044 4036 143100
rect 4036 143044 4092 143100
rect 4092 143044 4096 143100
rect 4032 143040 4096 143044
rect 4112 143100 4176 143104
rect 4112 143044 4116 143100
rect 4116 143044 4172 143100
rect 4172 143044 4176 143100
rect 4112 143040 4176 143044
rect 4192 143100 4256 143104
rect 4192 143044 4196 143100
rect 4196 143044 4252 143100
rect 4252 143044 4256 143100
rect 4192 143040 4256 143044
rect 87952 143100 88016 143104
rect 87952 143044 87956 143100
rect 87956 143044 88012 143100
rect 88012 143044 88016 143100
rect 87952 143040 88016 143044
rect 88032 143100 88096 143104
rect 88032 143044 88036 143100
rect 88036 143044 88092 143100
rect 88092 143044 88096 143100
rect 88032 143040 88096 143044
rect 88112 143100 88176 143104
rect 88112 143044 88116 143100
rect 88116 143044 88172 143100
rect 88172 143044 88176 143100
rect 88112 143040 88176 143044
rect 88192 143100 88256 143104
rect 88192 143044 88196 143100
rect 88196 143044 88252 143100
rect 88252 143044 88256 143100
rect 88192 143040 88256 143044
rect 1952 142556 2016 142560
rect 1952 142500 1956 142556
rect 1956 142500 2012 142556
rect 2012 142500 2016 142556
rect 1952 142496 2016 142500
rect 2032 142556 2096 142560
rect 2032 142500 2036 142556
rect 2036 142500 2092 142556
rect 2092 142500 2096 142556
rect 2032 142496 2096 142500
rect 2112 142556 2176 142560
rect 2112 142500 2116 142556
rect 2116 142500 2172 142556
rect 2172 142500 2176 142556
rect 2112 142496 2176 142500
rect 2192 142556 2256 142560
rect 2192 142500 2196 142556
rect 2196 142500 2252 142556
rect 2252 142500 2256 142556
rect 2192 142496 2256 142500
rect 85952 142556 86016 142560
rect 85952 142500 85956 142556
rect 85956 142500 86012 142556
rect 86012 142500 86016 142556
rect 85952 142496 86016 142500
rect 86032 142556 86096 142560
rect 86032 142500 86036 142556
rect 86036 142500 86092 142556
rect 86092 142500 86096 142556
rect 86032 142496 86096 142500
rect 86112 142556 86176 142560
rect 86112 142500 86116 142556
rect 86116 142500 86172 142556
rect 86172 142500 86176 142556
rect 86112 142496 86176 142500
rect 86192 142556 86256 142560
rect 86192 142500 86196 142556
rect 86196 142500 86252 142556
rect 86252 142500 86256 142556
rect 86192 142496 86256 142500
rect 89952 142556 90016 142560
rect 89952 142500 89956 142556
rect 89956 142500 90012 142556
rect 90012 142500 90016 142556
rect 89952 142496 90016 142500
rect 90032 142556 90096 142560
rect 90032 142500 90036 142556
rect 90036 142500 90092 142556
rect 90092 142500 90096 142556
rect 90032 142496 90096 142500
rect 90112 142556 90176 142560
rect 90112 142500 90116 142556
rect 90116 142500 90172 142556
rect 90172 142500 90176 142556
rect 90112 142496 90176 142500
rect 90192 142556 90256 142560
rect 90192 142500 90196 142556
rect 90196 142500 90252 142556
rect 90252 142500 90256 142556
rect 90192 142496 90256 142500
rect 3952 142012 4016 142016
rect 3952 141956 3956 142012
rect 3956 141956 4012 142012
rect 4012 141956 4016 142012
rect 3952 141952 4016 141956
rect 4032 142012 4096 142016
rect 4032 141956 4036 142012
rect 4036 141956 4092 142012
rect 4092 141956 4096 142012
rect 4032 141952 4096 141956
rect 4112 142012 4176 142016
rect 4112 141956 4116 142012
rect 4116 141956 4172 142012
rect 4172 141956 4176 142012
rect 4112 141952 4176 141956
rect 4192 142012 4256 142016
rect 4192 141956 4196 142012
rect 4196 141956 4252 142012
rect 4252 141956 4256 142012
rect 4192 141952 4256 141956
rect 87952 142012 88016 142016
rect 87952 141956 87956 142012
rect 87956 141956 88012 142012
rect 88012 141956 88016 142012
rect 87952 141952 88016 141956
rect 88032 142012 88096 142016
rect 88032 141956 88036 142012
rect 88036 141956 88092 142012
rect 88092 141956 88096 142012
rect 88032 141952 88096 141956
rect 88112 142012 88176 142016
rect 88112 141956 88116 142012
rect 88116 141956 88172 142012
rect 88172 141956 88176 142012
rect 88112 141952 88176 141956
rect 88192 142012 88256 142016
rect 88192 141956 88196 142012
rect 88196 141956 88252 142012
rect 88252 141956 88256 142012
rect 88192 141952 88256 141956
rect 1952 141468 2016 141472
rect 1952 141412 1956 141468
rect 1956 141412 2012 141468
rect 2012 141412 2016 141468
rect 1952 141408 2016 141412
rect 2032 141468 2096 141472
rect 2032 141412 2036 141468
rect 2036 141412 2092 141468
rect 2092 141412 2096 141468
rect 2032 141408 2096 141412
rect 2112 141468 2176 141472
rect 2112 141412 2116 141468
rect 2116 141412 2172 141468
rect 2172 141412 2176 141468
rect 2112 141408 2176 141412
rect 2192 141468 2256 141472
rect 2192 141412 2196 141468
rect 2196 141412 2252 141468
rect 2252 141412 2256 141468
rect 2192 141408 2256 141412
rect 85952 141468 86016 141472
rect 85952 141412 85956 141468
rect 85956 141412 86012 141468
rect 86012 141412 86016 141468
rect 85952 141408 86016 141412
rect 86032 141468 86096 141472
rect 86032 141412 86036 141468
rect 86036 141412 86092 141468
rect 86092 141412 86096 141468
rect 86032 141408 86096 141412
rect 86112 141468 86176 141472
rect 86112 141412 86116 141468
rect 86116 141412 86172 141468
rect 86172 141412 86176 141468
rect 86112 141408 86176 141412
rect 86192 141468 86256 141472
rect 86192 141412 86196 141468
rect 86196 141412 86252 141468
rect 86252 141412 86256 141468
rect 86192 141408 86256 141412
rect 89952 141468 90016 141472
rect 89952 141412 89956 141468
rect 89956 141412 90012 141468
rect 90012 141412 90016 141468
rect 89952 141408 90016 141412
rect 90032 141468 90096 141472
rect 90032 141412 90036 141468
rect 90036 141412 90092 141468
rect 90092 141412 90096 141468
rect 90032 141408 90096 141412
rect 90112 141468 90176 141472
rect 90112 141412 90116 141468
rect 90116 141412 90172 141468
rect 90172 141412 90176 141468
rect 90112 141408 90176 141412
rect 90192 141468 90256 141472
rect 90192 141412 90196 141468
rect 90196 141412 90252 141468
rect 90252 141412 90256 141468
rect 90192 141408 90256 141412
rect 3952 140924 4016 140928
rect 3952 140868 3956 140924
rect 3956 140868 4012 140924
rect 4012 140868 4016 140924
rect 3952 140864 4016 140868
rect 4032 140924 4096 140928
rect 4032 140868 4036 140924
rect 4036 140868 4092 140924
rect 4092 140868 4096 140924
rect 4032 140864 4096 140868
rect 4112 140924 4176 140928
rect 4112 140868 4116 140924
rect 4116 140868 4172 140924
rect 4172 140868 4176 140924
rect 4112 140864 4176 140868
rect 4192 140924 4256 140928
rect 4192 140868 4196 140924
rect 4196 140868 4252 140924
rect 4252 140868 4256 140924
rect 4192 140864 4256 140868
rect 87952 140924 88016 140928
rect 87952 140868 87956 140924
rect 87956 140868 88012 140924
rect 88012 140868 88016 140924
rect 87952 140864 88016 140868
rect 88032 140924 88096 140928
rect 88032 140868 88036 140924
rect 88036 140868 88092 140924
rect 88092 140868 88096 140924
rect 88032 140864 88096 140868
rect 88112 140924 88176 140928
rect 88112 140868 88116 140924
rect 88116 140868 88172 140924
rect 88172 140868 88176 140924
rect 88112 140864 88176 140868
rect 88192 140924 88256 140928
rect 88192 140868 88196 140924
rect 88196 140868 88252 140924
rect 88252 140868 88256 140924
rect 88192 140864 88256 140868
rect 1952 140380 2016 140384
rect 1952 140324 1956 140380
rect 1956 140324 2012 140380
rect 2012 140324 2016 140380
rect 1952 140320 2016 140324
rect 2032 140380 2096 140384
rect 2032 140324 2036 140380
rect 2036 140324 2092 140380
rect 2092 140324 2096 140380
rect 2032 140320 2096 140324
rect 2112 140380 2176 140384
rect 2112 140324 2116 140380
rect 2116 140324 2172 140380
rect 2172 140324 2176 140380
rect 2112 140320 2176 140324
rect 2192 140380 2256 140384
rect 2192 140324 2196 140380
rect 2196 140324 2252 140380
rect 2252 140324 2256 140380
rect 2192 140320 2256 140324
rect 85952 140380 86016 140384
rect 85952 140324 85956 140380
rect 85956 140324 86012 140380
rect 86012 140324 86016 140380
rect 85952 140320 86016 140324
rect 86032 140380 86096 140384
rect 86032 140324 86036 140380
rect 86036 140324 86092 140380
rect 86092 140324 86096 140380
rect 86032 140320 86096 140324
rect 86112 140380 86176 140384
rect 86112 140324 86116 140380
rect 86116 140324 86172 140380
rect 86172 140324 86176 140380
rect 86112 140320 86176 140324
rect 86192 140380 86256 140384
rect 86192 140324 86196 140380
rect 86196 140324 86252 140380
rect 86252 140324 86256 140380
rect 86192 140320 86256 140324
rect 89952 140380 90016 140384
rect 89952 140324 89956 140380
rect 89956 140324 90012 140380
rect 90012 140324 90016 140380
rect 89952 140320 90016 140324
rect 90032 140380 90096 140384
rect 90032 140324 90036 140380
rect 90036 140324 90092 140380
rect 90092 140324 90096 140380
rect 90032 140320 90096 140324
rect 90112 140380 90176 140384
rect 90112 140324 90116 140380
rect 90116 140324 90172 140380
rect 90172 140324 90176 140380
rect 90112 140320 90176 140324
rect 90192 140380 90256 140384
rect 90192 140324 90196 140380
rect 90196 140324 90252 140380
rect 90252 140324 90256 140380
rect 90192 140320 90256 140324
rect 3952 139836 4016 139840
rect 3952 139780 3956 139836
rect 3956 139780 4012 139836
rect 4012 139780 4016 139836
rect 3952 139776 4016 139780
rect 4032 139836 4096 139840
rect 4032 139780 4036 139836
rect 4036 139780 4092 139836
rect 4092 139780 4096 139836
rect 4032 139776 4096 139780
rect 4112 139836 4176 139840
rect 4112 139780 4116 139836
rect 4116 139780 4172 139836
rect 4172 139780 4176 139836
rect 4112 139776 4176 139780
rect 4192 139836 4256 139840
rect 4192 139780 4196 139836
rect 4196 139780 4252 139836
rect 4252 139780 4256 139836
rect 4192 139776 4256 139780
rect 87952 139836 88016 139840
rect 87952 139780 87956 139836
rect 87956 139780 88012 139836
rect 88012 139780 88016 139836
rect 87952 139776 88016 139780
rect 88032 139836 88096 139840
rect 88032 139780 88036 139836
rect 88036 139780 88092 139836
rect 88092 139780 88096 139836
rect 88032 139776 88096 139780
rect 88112 139836 88176 139840
rect 88112 139780 88116 139836
rect 88116 139780 88172 139836
rect 88172 139780 88176 139836
rect 88112 139776 88176 139780
rect 88192 139836 88256 139840
rect 88192 139780 88196 139836
rect 88196 139780 88252 139836
rect 88252 139780 88256 139836
rect 88192 139776 88256 139780
rect 1952 139292 2016 139296
rect 1952 139236 1956 139292
rect 1956 139236 2012 139292
rect 2012 139236 2016 139292
rect 1952 139232 2016 139236
rect 2032 139292 2096 139296
rect 2032 139236 2036 139292
rect 2036 139236 2092 139292
rect 2092 139236 2096 139292
rect 2032 139232 2096 139236
rect 2112 139292 2176 139296
rect 2112 139236 2116 139292
rect 2116 139236 2172 139292
rect 2172 139236 2176 139292
rect 2112 139232 2176 139236
rect 2192 139292 2256 139296
rect 2192 139236 2196 139292
rect 2196 139236 2252 139292
rect 2252 139236 2256 139292
rect 2192 139232 2256 139236
rect 85952 139292 86016 139296
rect 85952 139236 85956 139292
rect 85956 139236 86012 139292
rect 86012 139236 86016 139292
rect 85952 139232 86016 139236
rect 86032 139292 86096 139296
rect 86032 139236 86036 139292
rect 86036 139236 86092 139292
rect 86092 139236 86096 139292
rect 86032 139232 86096 139236
rect 86112 139292 86176 139296
rect 86112 139236 86116 139292
rect 86116 139236 86172 139292
rect 86172 139236 86176 139292
rect 86112 139232 86176 139236
rect 86192 139292 86256 139296
rect 86192 139236 86196 139292
rect 86196 139236 86252 139292
rect 86252 139236 86256 139292
rect 86192 139232 86256 139236
rect 89952 139292 90016 139296
rect 89952 139236 89956 139292
rect 89956 139236 90012 139292
rect 90012 139236 90016 139292
rect 89952 139232 90016 139236
rect 90032 139292 90096 139296
rect 90032 139236 90036 139292
rect 90036 139236 90092 139292
rect 90092 139236 90096 139292
rect 90032 139232 90096 139236
rect 90112 139292 90176 139296
rect 90112 139236 90116 139292
rect 90116 139236 90172 139292
rect 90172 139236 90176 139292
rect 90112 139232 90176 139236
rect 90192 139292 90256 139296
rect 90192 139236 90196 139292
rect 90196 139236 90252 139292
rect 90252 139236 90256 139292
rect 90192 139232 90256 139236
rect 3952 138748 4016 138752
rect 3952 138692 3956 138748
rect 3956 138692 4012 138748
rect 4012 138692 4016 138748
rect 3952 138688 4016 138692
rect 4032 138748 4096 138752
rect 4032 138692 4036 138748
rect 4036 138692 4092 138748
rect 4092 138692 4096 138748
rect 4032 138688 4096 138692
rect 4112 138748 4176 138752
rect 4112 138692 4116 138748
rect 4116 138692 4172 138748
rect 4172 138692 4176 138748
rect 4112 138688 4176 138692
rect 4192 138748 4256 138752
rect 4192 138692 4196 138748
rect 4196 138692 4252 138748
rect 4252 138692 4256 138748
rect 4192 138688 4256 138692
rect 87952 138748 88016 138752
rect 87952 138692 87956 138748
rect 87956 138692 88012 138748
rect 88012 138692 88016 138748
rect 87952 138688 88016 138692
rect 88032 138748 88096 138752
rect 88032 138692 88036 138748
rect 88036 138692 88092 138748
rect 88092 138692 88096 138748
rect 88032 138688 88096 138692
rect 88112 138748 88176 138752
rect 88112 138692 88116 138748
rect 88116 138692 88172 138748
rect 88172 138692 88176 138748
rect 88112 138688 88176 138692
rect 88192 138748 88256 138752
rect 88192 138692 88196 138748
rect 88196 138692 88252 138748
rect 88252 138692 88256 138748
rect 88192 138688 88256 138692
rect 1952 138204 2016 138208
rect 1952 138148 1956 138204
rect 1956 138148 2012 138204
rect 2012 138148 2016 138204
rect 1952 138144 2016 138148
rect 2032 138204 2096 138208
rect 2032 138148 2036 138204
rect 2036 138148 2092 138204
rect 2092 138148 2096 138204
rect 2032 138144 2096 138148
rect 2112 138204 2176 138208
rect 2112 138148 2116 138204
rect 2116 138148 2172 138204
rect 2172 138148 2176 138204
rect 2112 138144 2176 138148
rect 2192 138204 2256 138208
rect 2192 138148 2196 138204
rect 2196 138148 2252 138204
rect 2252 138148 2256 138204
rect 2192 138144 2256 138148
rect 85952 138204 86016 138208
rect 85952 138148 85956 138204
rect 85956 138148 86012 138204
rect 86012 138148 86016 138204
rect 85952 138144 86016 138148
rect 86032 138204 86096 138208
rect 86032 138148 86036 138204
rect 86036 138148 86092 138204
rect 86092 138148 86096 138204
rect 86032 138144 86096 138148
rect 86112 138204 86176 138208
rect 86112 138148 86116 138204
rect 86116 138148 86172 138204
rect 86172 138148 86176 138204
rect 86112 138144 86176 138148
rect 86192 138204 86256 138208
rect 86192 138148 86196 138204
rect 86196 138148 86252 138204
rect 86252 138148 86256 138204
rect 86192 138144 86256 138148
rect 89952 138204 90016 138208
rect 89952 138148 89956 138204
rect 89956 138148 90012 138204
rect 90012 138148 90016 138204
rect 89952 138144 90016 138148
rect 90032 138204 90096 138208
rect 90032 138148 90036 138204
rect 90036 138148 90092 138204
rect 90092 138148 90096 138204
rect 90032 138144 90096 138148
rect 90112 138204 90176 138208
rect 90112 138148 90116 138204
rect 90116 138148 90172 138204
rect 90172 138148 90176 138204
rect 90112 138144 90176 138148
rect 90192 138204 90256 138208
rect 90192 138148 90196 138204
rect 90196 138148 90252 138204
rect 90252 138148 90256 138204
rect 90192 138144 90256 138148
rect 3952 137660 4016 137664
rect 3952 137604 3956 137660
rect 3956 137604 4012 137660
rect 4012 137604 4016 137660
rect 3952 137600 4016 137604
rect 4032 137660 4096 137664
rect 4032 137604 4036 137660
rect 4036 137604 4092 137660
rect 4092 137604 4096 137660
rect 4032 137600 4096 137604
rect 4112 137660 4176 137664
rect 4112 137604 4116 137660
rect 4116 137604 4172 137660
rect 4172 137604 4176 137660
rect 4112 137600 4176 137604
rect 4192 137660 4256 137664
rect 4192 137604 4196 137660
rect 4196 137604 4252 137660
rect 4252 137604 4256 137660
rect 4192 137600 4256 137604
rect 87952 137660 88016 137664
rect 87952 137604 87956 137660
rect 87956 137604 88012 137660
rect 88012 137604 88016 137660
rect 87952 137600 88016 137604
rect 88032 137660 88096 137664
rect 88032 137604 88036 137660
rect 88036 137604 88092 137660
rect 88092 137604 88096 137660
rect 88032 137600 88096 137604
rect 88112 137660 88176 137664
rect 88112 137604 88116 137660
rect 88116 137604 88172 137660
rect 88172 137604 88176 137660
rect 88112 137600 88176 137604
rect 88192 137660 88256 137664
rect 88192 137604 88196 137660
rect 88196 137604 88252 137660
rect 88252 137604 88256 137660
rect 88192 137600 88256 137604
rect 1952 137116 2016 137120
rect 1952 137060 1956 137116
rect 1956 137060 2012 137116
rect 2012 137060 2016 137116
rect 1952 137056 2016 137060
rect 2032 137116 2096 137120
rect 2032 137060 2036 137116
rect 2036 137060 2092 137116
rect 2092 137060 2096 137116
rect 2032 137056 2096 137060
rect 2112 137116 2176 137120
rect 2112 137060 2116 137116
rect 2116 137060 2172 137116
rect 2172 137060 2176 137116
rect 2112 137056 2176 137060
rect 2192 137116 2256 137120
rect 2192 137060 2196 137116
rect 2196 137060 2252 137116
rect 2252 137060 2256 137116
rect 2192 137056 2256 137060
rect 85952 137116 86016 137120
rect 85952 137060 85956 137116
rect 85956 137060 86012 137116
rect 86012 137060 86016 137116
rect 85952 137056 86016 137060
rect 86032 137116 86096 137120
rect 86032 137060 86036 137116
rect 86036 137060 86092 137116
rect 86092 137060 86096 137116
rect 86032 137056 86096 137060
rect 86112 137116 86176 137120
rect 86112 137060 86116 137116
rect 86116 137060 86172 137116
rect 86172 137060 86176 137116
rect 86112 137056 86176 137060
rect 86192 137116 86256 137120
rect 86192 137060 86196 137116
rect 86196 137060 86252 137116
rect 86252 137060 86256 137116
rect 86192 137056 86256 137060
rect 89952 137116 90016 137120
rect 89952 137060 89956 137116
rect 89956 137060 90012 137116
rect 90012 137060 90016 137116
rect 89952 137056 90016 137060
rect 90032 137116 90096 137120
rect 90032 137060 90036 137116
rect 90036 137060 90092 137116
rect 90092 137060 90096 137116
rect 90032 137056 90096 137060
rect 90112 137116 90176 137120
rect 90112 137060 90116 137116
rect 90116 137060 90172 137116
rect 90172 137060 90176 137116
rect 90112 137056 90176 137060
rect 90192 137116 90256 137120
rect 90192 137060 90196 137116
rect 90196 137060 90252 137116
rect 90252 137060 90256 137116
rect 90192 137056 90256 137060
rect 3952 136572 4016 136576
rect 3952 136516 3956 136572
rect 3956 136516 4012 136572
rect 4012 136516 4016 136572
rect 3952 136512 4016 136516
rect 4032 136572 4096 136576
rect 4032 136516 4036 136572
rect 4036 136516 4092 136572
rect 4092 136516 4096 136572
rect 4032 136512 4096 136516
rect 4112 136572 4176 136576
rect 4112 136516 4116 136572
rect 4116 136516 4172 136572
rect 4172 136516 4176 136572
rect 4112 136512 4176 136516
rect 4192 136572 4256 136576
rect 4192 136516 4196 136572
rect 4196 136516 4252 136572
rect 4252 136516 4256 136572
rect 4192 136512 4256 136516
rect 87952 136572 88016 136576
rect 87952 136516 87956 136572
rect 87956 136516 88012 136572
rect 88012 136516 88016 136572
rect 87952 136512 88016 136516
rect 88032 136572 88096 136576
rect 88032 136516 88036 136572
rect 88036 136516 88092 136572
rect 88092 136516 88096 136572
rect 88032 136512 88096 136516
rect 88112 136572 88176 136576
rect 88112 136516 88116 136572
rect 88116 136516 88172 136572
rect 88172 136516 88176 136572
rect 88112 136512 88176 136516
rect 88192 136572 88256 136576
rect 88192 136516 88196 136572
rect 88196 136516 88252 136572
rect 88252 136516 88256 136572
rect 88192 136512 88256 136516
rect 1952 136028 2016 136032
rect 1952 135972 1956 136028
rect 1956 135972 2012 136028
rect 2012 135972 2016 136028
rect 1952 135968 2016 135972
rect 2032 136028 2096 136032
rect 2032 135972 2036 136028
rect 2036 135972 2092 136028
rect 2092 135972 2096 136028
rect 2032 135968 2096 135972
rect 2112 136028 2176 136032
rect 2112 135972 2116 136028
rect 2116 135972 2172 136028
rect 2172 135972 2176 136028
rect 2112 135968 2176 135972
rect 2192 136028 2256 136032
rect 2192 135972 2196 136028
rect 2196 135972 2252 136028
rect 2252 135972 2256 136028
rect 2192 135968 2256 135972
rect 85952 136028 86016 136032
rect 85952 135972 85956 136028
rect 85956 135972 86012 136028
rect 86012 135972 86016 136028
rect 85952 135968 86016 135972
rect 86032 136028 86096 136032
rect 86032 135972 86036 136028
rect 86036 135972 86092 136028
rect 86092 135972 86096 136028
rect 86032 135968 86096 135972
rect 86112 136028 86176 136032
rect 86112 135972 86116 136028
rect 86116 135972 86172 136028
rect 86172 135972 86176 136028
rect 86112 135968 86176 135972
rect 86192 136028 86256 136032
rect 86192 135972 86196 136028
rect 86196 135972 86252 136028
rect 86252 135972 86256 136028
rect 86192 135968 86256 135972
rect 89952 136028 90016 136032
rect 89952 135972 89956 136028
rect 89956 135972 90012 136028
rect 90012 135972 90016 136028
rect 89952 135968 90016 135972
rect 90032 136028 90096 136032
rect 90032 135972 90036 136028
rect 90036 135972 90092 136028
rect 90092 135972 90096 136028
rect 90032 135968 90096 135972
rect 90112 136028 90176 136032
rect 90112 135972 90116 136028
rect 90116 135972 90172 136028
rect 90172 135972 90176 136028
rect 90112 135968 90176 135972
rect 90192 136028 90256 136032
rect 90192 135972 90196 136028
rect 90196 135972 90252 136028
rect 90252 135972 90256 136028
rect 90192 135968 90256 135972
rect 3952 135484 4016 135488
rect 3952 135428 3956 135484
rect 3956 135428 4012 135484
rect 4012 135428 4016 135484
rect 3952 135424 4016 135428
rect 4032 135484 4096 135488
rect 4032 135428 4036 135484
rect 4036 135428 4092 135484
rect 4092 135428 4096 135484
rect 4032 135424 4096 135428
rect 4112 135484 4176 135488
rect 4112 135428 4116 135484
rect 4116 135428 4172 135484
rect 4172 135428 4176 135484
rect 4112 135424 4176 135428
rect 4192 135484 4256 135488
rect 4192 135428 4196 135484
rect 4196 135428 4252 135484
rect 4252 135428 4256 135484
rect 4192 135424 4256 135428
rect 87952 135484 88016 135488
rect 87952 135428 87956 135484
rect 87956 135428 88012 135484
rect 88012 135428 88016 135484
rect 87952 135424 88016 135428
rect 88032 135484 88096 135488
rect 88032 135428 88036 135484
rect 88036 135428 88092 135484
rect 88092 135428 88096 135484
rect 88032 135424 88096 135428
rect 88112 135484 88176 135488
rect 88112 135428 88116 135484
rect 88116 135428 88172 135484
rect 88172 135428 88176 135484
rect 88112 135424 88176 135428
rect 88192 135484 88256 135488
rect 88192 135428 88196 135484
rect 88196 135428 88252 135484
rect 88252 135428 88256 135484
rect 88192 135424 88256 135428
rect 1952 134940 2016 134944
rect 1952 134884 1956 134940
rect 1956 134884 2012 134940
rect 2012 134884 2016 134940
rect 1952 134880 2016 134884
rect 2032 134940 2096 134944
rect 2032 134884 2036 134940
rect 2036 134884 2092 134940
rect 2092 134884 2096 134940
rect 2032 134880 2096 134884
rect 2112 134940 2176 134944
rect 2112 134884 2116 134940
rect 2116 134884 2172 134940
rect 2172 134884 2176 134940
rect 2112 134880 2176 134884
rect 2192 134940 2256 134944
rect 2192 134884 2196 134940
rect 2196 134884 2252 134940
rect 2252 134884 2256 134940
rect 2192 134880 2256 134884
rect 85952 134940 86016 134944
rect 85952 134884 85956 134940
rect 85956 134884 86012 134940
rect 86012 134884 86016 134940
rect 85952 134880 86016 134884
rect 86032 134940 86096 134944
rect 86032 134884 86036 134940
rect 86036 134884 86092 134940
rect 86092 134884 86096 134940
rect 86032 134880 86096 134884
rect 86112 134940 86176 134944
rect 86112 134884 86116 134940
rect 86116 134884 86172 134940
rect 86172 134884 86176 134940
rect 86112 134880 86176 134884
rect 86192 134940 86256 134944
rect 86192 134884 86196 134940
rect 86196 134884 86252 134940
rect 86252 134884 86256 134940
rect 86192 134880 86256 134884
rect 89952 134940 90016 134944
rect 89952 134884 89956 134940
rect 89956 134884 90012 134940
rect 90012 134884 90016 134940
rect 89952 134880 90016 134884
rect 90032 134940 90096 134944
rect 90032 134884 90036 134940
rect 90036 134884 90092 134940
rect 90092 134884 90096 134940
rect 90032 134880 90096 134884
rect 90112 134940 90176 134944
rect 90112 134884 90116 134940
rect 90116 134884 90172 134940
rect 90172 134884 90176 134940
rect 90112 134880 90176 134884
rect 90192 134940 90256 134944
rect 90192 134884 90196 134940
rect 90196 134884 90252 134940
rect 90252 134884 90256 134940
rect 90192 134880 90256 134884
rect 3952 134396 4016 134400
rect 3952 134340 3956 134396
rect 3956 134340 4012 134396
rect 4012 134340 4016 134396
rect 3952 134336 4016 134340
rect 4032 134396 4096 134400
rect 4032 134340 4036 134396
rect 4036 134340 4092 134396
rect 4092 134340 4096 134396
rect 4032 134336 4096 134340
rect 4112 134396 4176 134400
rect 4112 134340 4116 134396
rect 4116 134340 4172 134396
rect 4172 134340 4176 134396
rect 4112 134336 4176 134340
rect 4192 134396 4256 134400
rect 4192 134340 4196 134396
rect 4196 134340 4252 134396
rect 4252 134340 4256 134396
rect 4192 134336 4256 134340
rect 87952 134396 88016 134400
rect 87952 134340 87956 134396
rect 87956 134340 88012 134396
rect 88012 134340 88016 134396
rect 87952 134336 88016 134340
rect 88032 134396 88096 134400
rect 88032 134340 88036 134396
rect 88036 134340 88092 134396
rect 88092 134340 88096 134396
rect 88032 134336 88096 134340
rect 88112 134396 88176 134400
rect 88112 134340 88116 134396
rect 88116 134340 88172 134396
rect 88172 134340 88176 134396
rect 88112 134336 88176 134340
rect 88192 134396 88256 134400
rect 88192 134340 88196 134396
rect 88196 134340 88252 134396
rect 88252 134340 88256 134396
rect 88192 134336 88256 134340
rect 1952 133852 2016 133856
rect 1952 133796 1956 133852
rect 1956 133796 2012 133852
rect 2012 133796 2016 133852
rect 1952 133792 2016 133796
rect 2032 133852 2096 133856
rect 2032 133796 2036 133852
rect 2036 133796 2092 133852
rect 2092 133796 2096 133852
rect 2032 133792 2096 133796
rect 2112 133852 2176 133856
rect 2112 133796 2116 133852
rect 2116 133796 2172 133852
rect 2172 133796 2176 133852
rect 2112 133792 2176 133796
rect 2192 133852 2256 133856
rect 2192 133796 2196 133852
rect 2196 133796 2252 133852
rect 2252 133796 2256 133852
rect 2192 133792 2256 133796
rect 85952 133852 86016 133856
rect 85952 133796 85956 133852
rect 85956 133796 86012 133852
rect 86012 133796 86016 133852
rect 85952 133792 86016 133796
rect 86032 133852 86096 133856
rect 86032 133796 86036 133852
rect 86036 133796 86092 133852
rect 86092 133796 86096 133852
rect 86032 133792 86096 133796
rect 86112 133852 86176 133856
rect 86112 133796 86116 133852
rect 86116 133796 86172 133852
rect 86172 133796 86176 133852
rect 86112 133792 86176 133796
rect 86192 133852 86256 133856
rect 86192 133796 86196 133852
rect 86196 133796 86252 133852
rect 86252 133796 86256 133852
rect 86192 133792 86256 133796
rect 89952 133852 90016 133856
rect 89952 133796 89956 133852
rect 89956 133796 90012 133852
rect 90012 133796 90016 133852
rect 89952 133792 90016 133796
rect 90032 133852 90096 133856
rect 90032 133796 90036 133852
rect 90036 133796 90092 133852
rect 90092 133796 90096 133852
rect 90032 133792 90096 133796
rect 90112 133852 90176 133856
rect 90112 133796 90116 133852
rect 90116 133796 90172 133852
rect 90172 133796 90176 133852
rect 90112 133792 90176 133796
rect 90192 133852 90256 133856
rect 90192 133796 90196 133852
rect 90196 133796 90252 133852
rect 90252 133796 90256 133852
rect 90192 133792 90256 133796
rect 3952 133308 4016 133312
rect 3952 133252 3956 133308
rect 3956 133252 4012 133308
rect 4012 133252 4016 133308
rect 3952 133248 4016 133252
rect 4032 133308 4096 133312
rect 4032 133252 4036 133308
rect 4036 133252 4092 133308
rect 4092 133252 4096 133308
rect 4032 133248 4096 133252
rect 4112 133308 4176 133312
rect 4112 133252 4116 133308
rect 4116 133252 4172 133308
rect 4172 133252 4176 133308
rect 4112 133248 4176 133252
rect 4192 133308 4256 133312
rect 4192 133252 4196 133308
rect 4196 133252 4252 133308
rect 4252 133252 4256 133308
rect 4192 133248 4256 133252
rect 87952 133308 88016 133312
rect 87952 133252 87956 133308
rect 87956 133252 88012 133308
rect 88012 133252 88016 133308
rect 87952 133248 88016 133252
rect 88032 133308 88096 133312
rect 88032 133252 88036 133308
rect 88036 133252 88092 133308
rect 88092 133252 88096 133308
rect 88032 133248 88096 133252
rect 88112 133308 88176 133312
rect 88112 133252 88116 133308
rect 88116 133252 88172 133308
rect 88172 133252 88176 133308
rect 88112 133248 88176 133252
rect 88192 133308 88256 133312
rect 88192 133252 88196 133308
rect 88196 133252 88252 133308
rect 88252 133252 88256 133308
rect 88192 133248 88256 133252
rect 84884 133044 84948 133108
rect 1952 132764 2016 132768
rect 1952 132708 1956 132764
rect 1956 132708 2012 132764
rect 2012 132708 2016 132764
rect 1952 132704 2016 132708
rect 2032 132764 2096 132768
rect 2032 132708 2036 132764
rect 2036 132708 2092 132764
rect 2092 132708 2096 132764
rect 2032 132704 2096 132708
rect 2112 132764 2176 132768
rect 2112 132708 2116 132764
rect 2116 132708 2172 132764
rect 2172 132708 2176 132764
rect 2112 132704 2176 132708
rect 2192 132764 2256 132768
rect 2192 132708 2196 132764
rect 2196 132708 2252 132764
rect 2252 132708 2256 132764
rect 2192 132704 2256 132708
rect 85952 132764 86016 132768
rect 85952 132708 85956 132764
rect 85956 132708 86012 132764
rect 86012 132708 86016 132764
rect 85952 132704 86016 132708
rect 86032 132764 86096 132768
rect 86032 132708 86036 132764
rect 86036 132708 86092 132764
rect 86092 132708 86096 132764
rect 86032 132704 86096 132708
rect 86112 132764 86176 132768
rect 86112 132708 86116 132764
rect 86116 132708 86172 132764
rect 86172 132708 86176 132764
rect 86112 132704 86176 132708
rect 86192 132764 86256 132768
rect 86192 132708 86196 132764
rect 86196 132708 86252 132764
rect 86252 132708 86256 132764
rect 86192 132704 86256 132708
rect 89952 132764 90016 132768
rect 89952 132708 89956 132764
rect 89956 132708 90012 132764
rect 90012 132708 90016 132764
rect 89952 132704 90016 132708
rect 90032 132764 90096 132768
rect 90032 132708 90036 132764
rect 90036 132708 90092 132764
rect 90092 132708 90096 132764
rect 90032 132704 90096 132708
rect 90112 132764 90176 132768
rect 90112 132708 90116 132764
rect 90116 132708 90172 132764
rect 90172 132708 90176 132764
rect 90112 132704 90176 132708
rect 90192 132764 90256 132768
rect 90192 132708 90196 132764
rect 90196 132708 90252 132764
rect 90252 132708 90256 132764
rect 90192 132704 90256 132708
rect 83412 132364 83476 132428
rect 83964 132364 84028 132428
rect 83412 132228 83476 132292
rect 3952 132220 4016 132224
rect 3952 132164 3956 132220
rect 3956 132164 4012 132220
rect 4012 132164 4016 132220
rect 3952 132160 4016 132164
rect 4032 132220 4096 132224
rect 4032 132164 4036 132220
rect 4036 132164 4092 132220
rect 4092 132164 4096 132220
rect 4032 132160 4096 132164
rect 4112 132220 4176 132224
rect 4112 132164 4116 132220
rect 4116 132164 4172 132220
rect 4172 132164 4176 132220
rect 4112 132160 4176 132164
rect 4192 132220 4256 132224
rect 4192 132164 4196 132220
rect 4196 132164 4252 132220
rect 4252 132164 4256 132220
rect 4192 132160 4256 132164
rect 87952 132220 88016 132224
rect 87952 132164 87956 132220
rect 87956 132164 88012 132220
rect 88012 132164 88016 132220
rect 87952 132160 88016 132164
rect 88032 132220 88096 132224
rect 88032 132164 88036 132220
rect 88036 132164 88092 132220
rect 88092 132164 88096 132220
rect 88032 132160 88096 132164
rect 88112 132220 88176 132224
rect 88112 132164 88116 132220
rect 88116 132164 88172 132220
rect 88172 132164 88176 132220
rect 88112 132160 88176 132164
rect 88192 132220 88256 132224
rect 88192 132164 88196 132220
rect 88196 132164 88252 132220
rect 88252 132164 88256 132220
rect 88192 132160 88256 132164
rect 1952 131676 2016 131680
rect 1952 131620 1956 131676
rect 1956 131620 2012 131676
rect 2012 131620 2016 131676
rect 1952 131616 2016 131620
rect 2032 131676 2096 131680
rect 2032 131620 2036 131676
rect 2036 131620 2092 131676
rect 2092 131620 2096 131676
rect 2032 131616 2096 131620
rect 2112 131676 2176 131680
rect 2112 131620 2116 131676
rect 2116 131620 2172 131676
rect 2172 131620 2176 131676
rect 2112 131616 2176 131620
rect 2192 131676 2256 131680
rect 2192 131620 2196 131676
rect 2196 131620 2252 131676
rect 2252 131620 2256 131676
rect 2192 131616 2256 131620
rect 85952 131676 86016 131680
rect 85952 131620 85956 131676
rect 85956 131620 86012 131676
rect 86012 131620 86016 131676
rect 85952 131616 86016 131620
rect 86032 131676 86096 131680
rect 86032 131620 86036 131676
rect 86036 131620 86092 131676
rect 86092 131620 86096 131676
rect 86032 131616 86096 131620
rect 86112 131676 86176 131680
rect 86112 131620 86116 131676
rect 86116 131620 86172 131676
rect 86172 131620 86176 131676
rect 86112 131616 86176 131620
rect 86192 131676 86256 131680
rect 86192 131620 86196 131676
rect 86196 131620 86252 131676
rect 86252 131620 86256 131676
rect 86192 131616 86256 131620
rect 89952 131676 90016 131680
rect 89952 131620 89956 131676
rect 89956 131620 90012 131676
rect 90012 131620 90016 131676
rect 89952 131616 90016 131620
rect 90032 131676 90096 131680
rect 90032 131620 90036 131676
rect 90036 131620 90092 131676
rect 90092 131620 90096 131676
rect 90032 131616 90096 131620
rect 90112 131676 90176 131680
rect 90112 131620 90116 131676
rect 90116 131620 90172 131676
rect 90172 131620 90176 131676
rect 90112 131616 90176 131620
rect 90192 131676 90256 131680
rect 90192 131620 90196 131676
rect 90196 131620 90252 131676
rect 90252 131620 90256 131676
rect 90192 131616 90256 131620
rect 3952 131132 4016 131136
rect 3952 131076 3956 131132
rect 3956 131076 4012 131132
rect 4012 131076 4016 131132
rect 3952 131072 4016 131076
rect 4032 131132 4096 131136
rect 4032 131076 4036 131132
rect 4036 131076 4092 131132
rect 4092 131076 4096 131132
rect 4032 131072 4096 131076
rect 4112 131132 4176 131136
rect 4112 131076 4116 131132
rect 4116 131076 4172 131132
rect 4172 131076 4176 131132
rect 4112 131072 4176 131076
rect 4192 131132 4256 131136
rect 4192 131076 4196 131132
rect 4196 131076 4252 131132
rect 4252 131076 4256 131132
rect 4192 131072 4256 131076
rect 87952 131132 88016 131136
rect 87952 131076 87956 131132
rect 87956 131076 88012 131132
rect 88012 131076 88016 131132
rect 87952 131072 88016 131076
rect 88032 131132 88096 131136
rect 88032 131076 88036 131132
rect 88036 131076 88092 131132
rect 88092 131076 88096 131132
rect 88032 131072 88096 131076
rect 88112 131132 88176 131136
rect 88112 131076 88116 131132
rect 88116 131076 88172 131132
rect 88172 131076 88176 131132
rect 88112 131072 88176 131076
rect 88192 131132 88256 131136
rect 88192 131076 88196 131132
rect 88196 131076 88252 131132
rect 88252 131076 88256 131132
rect 88192 131072 88256 131076
rect 1952 130588 2016 130592
rect 1952 130532 1956 130588
rect 1956 130532 2012 130588
rect 2012 130532 2016 130588
rect 1952 130528 2016 130532
rect 2032 130588 2096 130592
rect 2032 130532 2036 130588
rect 2036 130532 2092 130588
rect 2092 130532 2096 130588
rect 2032 130528 2096 130532
rect 2112 130588 2176 130592
rect 2112 130532 2116 130588
rect 2116 130532 2172 130588
rect 2172 130532 2176 130588
rect 2112 130528 2176 130532
rect 2192 130588 2256 130592
rect 2192 130532 2196 130588
rect 2196 130532 2252 130588
rect 2252 130532 2256 130588
rect 2192 130528 2256 130532
rect 85952 130588 86016 130592
rect 85952 130532 85956 130588
rect 85956 130532 86012 130588
rect 86012 130532 86016 130588
rect 85952 130528 86016 130532
rect 86032 130588 86096 130592
rect 86032 130532 86036 130588
rect 86036 130532 86092 130588
rect 86092 130532 86096 130588
rect 86032 130528 86096 130532
rect 86112 130588 86176 130592
rect 86112 130532 86116 130588
rect 86116 130532 86172 130588
rect 86172 130532 86176 130588
rect 86112 130528 86176 130532
rect 86192 130588 86256 130592
rect 86192 130532 86196 130588
rect 86196 130532 86252 130588
rect 86252 130532 86256 130588
rect 86192 130528 86256 130532
rect 89952 130588 90016 130592
rect 89952 130532 89956 130588
rect 89956 130532 90012 130588
rect 90012 130532 90016 130588
rect 89952 130528 90016 130532
rect 90032 130588 90096 130592
rect 90032 130532 90036 130588
rect 90036 130532 90092 130588
rect 90092 130532 90096 130588
rect 90032 130528 90096 130532
rect 90112 130588 90176 130592
rect 90112 130532 90116 130588
rect 90116 130532 90172 130588
rect 90172 130532 90176 130588
rect 90112 130528 90176 130532
rect 90192 130588 90256 130592
rect 90192 130532 90196 130588
rect 90196 130532 90252 130588
rect 90252 130532 90256 130588
rect 90192 130528 90256 130532
rect 85252 130324 85316 130388
rect 3952 130044 4016 130048
rect 3952 129988 3956 130044
rect 3956 129988 4012 130044
rect 4012 129988 4016 130044
rect 3952 129984 4016 129988
rect 4032 130044 4096 130048
rect 4032 129988 4036 130044
rect 4036 129988 4092 130044
rect 4092 129988 4096 130044
rect 4032 129984 4096 129988
rect 4112 130044 4176 130048
rect 4112 129988 4116 130044
rect 4116 129988 4172 130044
rect 4172 129988 4176 130044
rect 4112 129984 4176 129988
rect 4192 130044 4256 130048
rect 4192 129988 4196 130044
rect 4196 129988 4252 130044
rect 4252 129988 4256 130044
rect 4192 129984 4256 129988
rect 87952 130044 88016 130048
rect 87952 129988 87956 130044
rect 87956 129988 88012 130044
rect 88012 129988 88016 130044
rect 87952 129984 88016 129988
rect 88032 130044 88096 130048
rect 88032 129988 88036 130044
rect 88036 129988 88092 130044
rect 88092 129988 88096 130044
rect 88032 129984 88096 129988
rect 88112 130044 88176 130048
rect 88112 129988 88116 130044
rect 88116 129988 88172 130044
rect 88172 129988 88176 130044
rect 88112 129984 88176 129988
rect 88192 130044 88256 130048
rect 88192 129988 88196 130044
rect 88196 129988 88252 130044
rect 88252 129988 88256 130044
rect 88192 129984 88256 129988
rect 1952 129500 2016 129504
rect 1952 129444 1956 129500
rect 1956 129444 2012 129500
rect 2012 129444 2016 129500
rect 1952 129440 2016 129444
rect 2032 129500 2096 129504
rect 2032 129444 2036 129500
rect 2036 129444 2092 129500
rect 2092 129444 2096 129500
rect 2032 129440 2096 129444
rect 2112 129500 2176 129504
rect 2112 129444 2116 129500
rect 2116 129444 2172 129500
rect 2172 129444 2176 129500
rect 2112 129440 2176 129444
rect 2192 129500 2256 129504
rect 2192 129444 2196 129500
rect 2196 129444 2252 129500
rect 2252 129444 2256 129500
rect 2192 129440 2256 129444
rect 85952 129500 86016 129504
rect 85952 129444 85956 129500
rect 85956 129444 86012 129500
rect 86012 129444 86016 129500
rect 85952 129440 86016 129444
rect 86032 129500 86096 129504
rect 86032 129444 86036 129500
rect 86036 129444 86092 129500
rect 86092 129444 86096 129500
rect 86032 129440 86096 129444
rect 86112 129500 86176 129504
rect 86112 129444 86116 129500
rect 86116 129444 86172 129500
rect 86172 129444 86176 129500
rect 86112 129440 86176 129444
rect 86192 129500 86256 129504
rect 86192 129444 86196 129500
rect 86196 129444 86252 129500
rect 86252 129444 86256 129500
rect 86192 129440 86256 129444
rect 89952 129500 90016 129504
rect 89952 129444 89956 129500
rect 89956 129444 90012 129500
rect 90012 129444 90016 129500
rect 89952 129440 90016 129444
rect 90032 129500 90096 129504
rect 90032 129444 90036 129500
rect 90036 129444 90092 129500
rect 90092 129444 90096 129500
rect 90032 129440 90096 129444
rect 90112 129500 90176 129504
rect 90112 129444 90116 129500
rect 90116 129444 90172 129500
rect 90172 129444 90176 129500
rect 90112 129440 90176 129444
rect 90192 129500 90256 129504
rect 90192 129444 90196 129500
rect 90196 129444 90252 129500
rect 90252 129444 90256 129500
rect 90192 129440 90256 129444
rect 3952 128956 4016 128960
rect 3952 128900 3956 128956
rect 3956 128900 4012 128956
rect 4012 128900 4016 128956
rect 3952 128896 4016 128900
rect 4032 128956 4096 128960
rect 4032 128900 4036 128956
rect 4036 128900 4092 128956
rect 4092 128900 4096 128956
rect 4032 128896 4096 128900
rect 4112 128956 4176 128960
rect 4112 128900 4116 128956
rect 4116 128900 4172 128956
rect 4172 128900 4176 128956
rect 4112 128896 4176 128900
rect 4192 128956 4256 128960
rect 4192 128900 4196 128956
rect 4196 128900 4252 128956
rect 4252 128900 4256 128956
rect 4192 128896 4256 128900
rect 87952 128956 88016 128960
rect 87952 128900 87956 128956
rect 87956 128900 88012 128956
rect 88012 128900 88016 128956
rect 87952 128896 88016 128900
rect 88032 128956 88096 128960
rect 88032 128900 88036 128956
rect 88036 128900 88092 128956
rect 88092 128900 88096 128956
rect 88032 128896 88096 128900
rect 88112 128956 88176 128960
rect 88112 128900 88116 128956
rect 88116 128900 88172 128956
rect 88172 128900 88176 128956
rect 88112 128896 88176 128900
rect 88192 128956 88256 128960
rect 88192 128900 88196 128956
rect 88196 128900 88252 128956
rect 88252 128900 88256 128956
rect 88192 128896 88256 128900
rect 1952 128412 2016 128416
rect 1952 128356 1956 128412
rect 1956 128356 2012 128412
rect 2012 128356 2016 128412
rect 1952 128352 2016 128356
rect 2032 128412 2096 128416
rect 2032 128356 2036 128412
rect 2036 128356 2092 128412
rect 2092 128356 2096 128412
rect 2032 128352 2096 128356
rect 2112 128412 2176 128416
rect 2112 128356 2116 128412
rect 2116 128356 2172 128412
rect 2172 128356 2176 128412
rect 2112 128352 2176 128356
rect 2192 128412 2256 128416
rect 2192 128356 2196 128412
rect 2196 128356 2252 128412
rect 2252 128356 2256 128412
rect 2192 128352 2256 128356
rect 85952 128412 86016 128416
rect 85952 128356 85956 128412
rect 85956 128356 86012 128412
rect 86012 128356 86016 128412
rect 85952 128352 86016 128356
rect 86032 128412 86096 128416
rect 86032 128356 86036 128412
rect 86036 128356 86092 128412
rect 86092 128356 86096 128412
rect 86032 128352 86096 128356
rect 86112 128412 86176 128416
rect 86112 128356 86116 128412
rect 86116 128356 86172 128412
rect 86172 128356 86176 128412
rect 86112 128352 86176 128356
rect 86192 128412 86256 128416
rect 86192 128356 86196 128412
rect 86196 128356 86252 128412
rect 86252 128356 86256 128412
rect 86192 128352 86256 128356
rect 89952 128412 90016 128416
rect 89952 128356 89956 128412
rect 89956 128356 90012 128412
rect 90012 128356 90016 128412
rect 89952 128352 90016 128356
rect 90032 128412 90096 128416
rect 90032 128356 90036 128412
rect 90036 128356 90092 128412
rect 90092 128356 90096 128412
rect 90032 128352 90096 128356
rect 90112 128412 90176 128416
rect 90112 128356 90116 128412
rect 90116 128356 90172 128412
rect 90172 128356 90176 128412
rect 90112 128352 90176 128356
rect 90192 128412 90256 128416
rect 90192 128356 90196 128412
rect 90196 128356 90252 128412
rect 90252 128356 90256 128412
rect 90192 128352 90256 128356
rect 3952 127868 4016 127872
rect 3952 127812 3956 127868
rect 3956 127812 4012 127868
rect 4012 127812 4016 127868
rect 3952 127808 4016 127812
rect 4032 127868 4096 127872
rect 4032 127812 4036 127868
rect 4036 127812 4092 127868
rect 4092 127812 4096 127868
rect 4032 127808 4096 127812
rect 4112 127868 4176 127872
rect 4112 127812 4116 127868
rect 4116 127812 4172 127868
rect 4172 127812 4176 127868
rect 4112 127808 4176 127812
rect 4192 127868 4256 127872
rect 4192 127812 4196 127868
rect 4196 127812 4252 127868
rect 4252 127812 4256 127868
rect 4192 127808 4256 127812
rect 87952 127868 88016 127872
rect 87952 127812 87956 127868
rect 87956 127812 88012 127868
rect 88012 127812 88016 127868
rect 87952 127808 88016 127812
rect 88032 127868 88096 127872
rect 88032 127812 88036 127868
rect 88036 127812 88092 127868
rect 88092 127812 88096 127868
rect 88032 127808 88096 127812
rect 88112 127868 88176 127872
rect 88112 127812 88116 127868
rect 88116 127812 88172 127868
rect 88172 127812 88176 127868
rect 88112 127808 88176 127812
rect 88192 127868 88256 127872
rect 88192 127812 88196 127868
rect 88196 127812 88252 127868
rect 88252 127812 88256 127868
rect 88192 127808 88256 127812
rect 1952 127324 2016 127328
rect 1952 127268 1956 127324
rect 1956 127268 2012 127324
rect 2012 127268 2016 127324
rect 1952 127264 2016 127268
rect 2032 127324 2096 127328
rect 2032 127268 2036 127324
rect 2036 127268 2092 127324
rect 2092 127268 2096 127324
rect 2032 127264 2096 127268
rect 2112 127324 2176 127328
rect 2112 127268 2116 127324
rect 2116 127268 2172 127324
rect 2172 127268 2176 127324
rect 2112 127264 2176 127268
rect 2192 127324 2256 127328
rect 2192 127268 2196 127324
rect 2196 127268 2252 127324
rect 2252 127268 2256 127324
rect 2192 127264 2256 127268
rect 85952 127324 86016 127328
rect 85952 127268 85956 127324
rect 85956 127268 86012 127324
rect 86012 127268 86016 127324
rect 85952 127264 86016 127268
rect 86032 127324 86096 127328
rect 86032 127268 86036 127324
rect 86036 127268 86092 127324
rect 86092 127268 86096 127324
rect 86032 127264 86096 127268
rect 86112 127324 86176 127328
rect 86112 127268 86116 127324
rect 86116 127268 86172 127324
rect 86172 127268 86176 127324
rect 86112 127264 86176 127268
rect 86192 127324 86256 127328
rect 86192 127268 86196 127324
rect 86196 127268 86252 127324
rect 86252 127268 86256 127324
rect 86192 127264 86256 127268
rect 89952 127324 90016 127328
rect 89952 127268 89956 127324
rect 89956 127268 90012 127324
rect 90012 127268 90016 127324
rect 89952 127264 90016 127268
rect 90032 127324 90096 127328
rect 90032 127268 90036 127324
rect 90036 127268 90092 127324
rect 90092 127268 90096 127324
rect 90032 127264 90096 127268
rect 90112 127324 90176 127328
rect 90112 127268 90116 127324
rect 90116 127268 90172 127324
rect 90172 127268 90176 127324
rect 90112 127264 90176 127268
rect 90192 127324 90256 127328
rect 90192 127268 90196 127324
rect 90196 127268 90252 127324
rect 90252 127268 90256 127324
rect 90192 127264 90256 127268
rect 84516 126924 84580 126988
rect 3952 126780 4016 126784
rect 3952 126724 3956 126780
rect 3956 126724 4012 126780
rect 4012 126724 4016 126780
rect 3952 126720 4016 126724
rect 4032 126780 4096 126784
rect 4032 126724 4036 126780
rect 4036 126724 4092 126780
rect 4092 126724 4096 126780
rect 4032 126720 4096 126724
rect 4112 126780 4176 126784
rect 4112 126724 4116 126780
rect 4116 126724 4172 126780
rect 4172 126724 4176 126780
rect 4112 126720 4176 126724
rect 4192 126780 4256 126784
rect 4192 126724 4196 126780
rect 4196 126724 4252 126780
rect 4252 126724 4256 126780
rect 4192 126720 4256 126724
rect 87952 126780 88016 126784
rect 87952 126724 87956 126780
rect 87956 126724 88012 126780
rect 88012 126724 88016 126780
rect 87952 126720 88016 126724
rect 88032 126780 88096 126784
rect 88032 126724 88036 126780
rect 88036 126724 88092 126780
rect 88092 126724 88096 126780
rect 88032 126720 88096 126724
rect 88112 126780 88176 126784
rect 88112 126724 88116 126780
rect 88116 126724 88172 126780
rect 88172 126724 88176 126780
rect 88112 126720 88176 126724
rect 88192 126780 88256 126784
rect 88192 126724 88196 126780
rect 88196 126724 88252 126780
rect 88252 126724 88256 126780
rect 88192 126720 88256 126724
rect 1952 126236 2016 126240
rect 1952 126180 1956 126236
rect 1956 126180 2012 126236
rect 2012 126180 2016 126236
rect 1952 126176 2016 126180
rect 2032 126236 2096 126240
rect 2032 126180 2036 126236
rect 2036 126180 2092 126236
rect 2092 126180 2096 126236
rect 2032 126176 2096 126180
rect 2112 126236 2176 126240
rect 2112 126180 2116 126236
rect 2116 126180 2172 126236
rect 2172 126180 2176 126236
rect 2112 126176 2176 126180
rect 2192 126236 2256 126240
rect 2192 126180 2196 126236
rect 2196 126180 2252 126236
rect 2252 126180 2256 126236
rect 2192 126176 2256 126180
rect 85952 126236 86016 126240
rect 85952 126180 85956 126236
rect 85956 126180 86012 126236
rect 86012 126180 86016 126236
rect 85952 126176 86016 126180
rect 86032 126236 86096 126240
rect 86032 126180 86036 126236
rect 86036 126180 86092 126236
rect 86092 126180 86096 126236
rect 86032 126176 86096 126180
rect 86112 126236 86176 126240
rect 86112 126180 86116 126236
rect 86116 126180 86172 126236
rect 86172 126180 86176 126236
rect 86112 126176 86176 126180
rect 86192 126236 86256 126240
rect 86192 126180 86196 126236
rect 86196 126180 86252 126236
rect 86252 126180 86256 126236
rect 86192 126176 86256 126180
rect 89952 126236 90016 126240
rect 89952 126180 89956 126236
rect 89956 126180 90012 126236
rect 90012 126180 90016 126236
rect 89952 126176 90016 126180
rect 90032 126236 90096 126240
rect 90032 126180 90036 126236
rect 90036 126180 90092 126236
rect 90092 126180 90096 126236
rect 90032 126176 90096 126180
rect 90112 126236 90176 126240
rect 90112 126180 90116 126236
rect 90116 126180 90172 126236
rect 90172 126180 90176 126236
rect 90112 126176 90176 126180
rect 90192 126236 90256 126240
rect 90192 126180 90196 126236
rect 90196 126180 90252 126236
rect 90252 126180 90256 126236
rect 90192 126176 90256 126180
rect 84700 125700 84764 125764
rect 3952 125692 4016 125696
rect 3952 125636 3956 125692
rect 3956 125636 4012 125692
rect 4012 125636 4016 125692
rect 3952 125632 4016 125636
rect 4032 125692 4096 125696
rect 4032 125636 4036 125692
rect 4036 125636 4092 125692
rect 4092 125636 4096 125692
rect 4032 125632 4096 125636
rect 4112 125692 4176 125696
rect 4112 125636 4116 125692
rect 4116 125636 4172 125692
rect 4172 125636 4176 125692
rect 4112 125632 4176 125636
rect 4192 125692 4256 125696
rect 4192 125636 4196 125692
rect 4196 125636 4252 125692
rect 4252 125636 4256 125692
rect 4192 125632 4256 125636
rect 87952 125692 88016 125696
rect 87952 125636 87956 125692
rect 87956 125636 88012 125692
rect 88012 125636 88016 125692
rect 87952 125632 88016 125636
rect 88032 125692 88096 125696
rect 88032 125636 88036 125692
rect 88036 125636 88092 125692
rect 88092 125636 88096 125692
rect 88032 125632 88096 125636
rect 88112 125692 88176 125696
rect 88112 125636 88116 125692
rect 88116 125636 88172 125692
rect 88172 125636 88176 125692
rect 88112 125632 88176 125636
rect 88192 125692 88256 125696
rect 88192 125636 88196 125692
rect 88196 125636 88252 125692
rect 88252 125636 88256 125692
rect 88192 125632 88256 125636
rect 1952 125148 2016 125152
rect 1952 125092 1956 125148
rect 1956 125092 2012 125148
rect 2012 125092 2016 125148
rect 1952 125088 2016 125092
rect 2032 125148 2096 125152
rect 2032 125092 2036 125148
rect 2036 125092 2092 125148
rect 2092 125092 2096 125148
rect 2032 125088 2096 125092
rect 2112 125148 2176 125152
rect 2112 125092 2116 125148
rect 2116 125092 2172 125148
rect 2172 125092 2176 125148
rect 2112 125088 2176 125092
rect 2192 125148 2256 125152
rect 2192 125092 2196 125148
rect 2196 125092 2252 125148
rect 2252 125092 2256 125148
rect 2192 125088 2256 125092
rect 85952 125148 86016 125152
rect 85952 125092 85956 125148
rect 85956 125092 86012 125148
rect 86012 125092 86016 125148
rect 85952 125088 86016 125092
rect 86032 125148 86096 125152
rect 86032 125092 86036 125148
rect 86036 125092 86092 125148
rect 86092 125092 86096 125148
rect 86032 125088 86096 125092
rect 86112 125148 86176 125152
rect 86112 125092 86116 125148
rect 86116 125092 86172 125148
rect 86172 125092 86176 125148
rect 86112 125088 86176 125092
rect 86192 125148 86256 125152
rect 86192 125092 86196 125148
rect 86196 125092 86252 125148
rect 86252 125092 86256 125148
rect 86192 125088 86256 125092
rect 89952 125148 90016 125152
rect 89952 125092 89956 125148
rect 89956 125092 90012 125148
rect 90012 125092 90016 125148
rect 89952 125088 90016 125092
rect 90032 125148 90096 125152
rect 90032 125092 90036 125148
rect 90036 125092 90092 125148
rect 90092 125092 90096 125148
rect 90032 125088 90096 125092
rect 90112 125148 90176 125152
rect 90112 125092 90116 125148
rect 90116 125092 90172 125148
rect 90172 125092 90176 125148
rect 90112 125088 90176 125092
rect 90192 125148 90256 125152
rect 90192 125092 90196 125148
rect 90196 125092 90252 125148
rect 90252 125092 90256 125148
rect 90192 125088 90256 125092
rect 3952 124604 4016 124608
rect 3952 124548 3956 124604
rect 3956 124548 4012 124604
rect 4012 124548 4016 124604
rect 3952 124544 4016 124548
rect 4032 124604 4096 124608
rect 4032 124548 4036 124604
rect 4036 124548 4092 124604
rect 4092 124548 4096 124604
rect 4032 124544 4096 124548
rect 4112 124604 4176 124608
rect 4112 124548 4116 124604
rect 4116 124548 4172 124604
rect 4172 124548 4176 124604
rect 4112 124544 4176 124548
rect 4192 124604 4256 124608
rect 4192 124548 4196 124604
rect 4196 124548 4252 124604
rect 4252 124548 4256 124604
rect 4192 124544 4256 124548
rect 87952 124604 88016 124608
rect 87952 124548 87956 124604
rect 87956 124548 88012 124604
rect 88012 124548 88016 124604
rect 87952 124544 88016 124548
rect 88032 124604 88096 124608
rect 88032 124548 88036 124604
rect 88036 124548 88092 124604
rect 88092 124548 88096 124604
rect 88032 124544 88096 124548
rect 88112 124604 88176 124608
rect 88112 124548 88116 124604
rect 88116 124548 88172 124604
rect 88172 124548 88176 124604
rect 88112 124544 88176 124548
rect 88192 124604 88256 124608
rect 88192 124548 88196 124604
rect 88196 124548 88252 124604
rect 88252 124548 88256 124604
rect 88192 124544 88256 124548
rect 1952 124060 2016 124064
rect 1952 124004 1956 124060
rect 1956 124004 2012 124060
rect 2012 124004 2016 124060
rect 1952 124000 2016 124004
rect 2032 124060 2096 124064
rect 2032 124004 2036 124060
rect 2036 124004 2092 124060
rect 2092 124004 2096 124060
rect 2032 124000 2096 124004
rect 2112 124060 2176 124064
rect 2112 124004 2116 124060
rect 2116 124004 2172 124060
rect 2172 124004 2176 124060
rect 2112 124000 2176 124004
rect 2192 124060 2256 124064
rect 2192 124004 2196 124060
rect 2196 124004 2252 124060
rect 2252 124004 2256 124060
rect 2192 124000 2256 124004
rect 85952 124060 86016 124064
rect 85952 124004 85956 124060
rect 85956 124004 86012 124060
rect 86012 124004 86016 124060
rect 85952 124000 86016 124004
rect 86032 124060 86096 124064
rect 86032 124004 86036 124060
rect 86036 124004 86092 124060
rect 86092 124004 86096 124060
rect 86032 124000 86096 124004
rect 86112 124060 86176 124064
rect 86112 124004 86116 124060
rect 86116 124004 86172 124060
rect 86172 124004 86176 124060
rect 86112 124000 86176 124004
rect 86192 124060 86256 124064
rect 86192 124004 86196 124060
rect 86196 124004 86252 124060
rect 86252 124004 86256 124060
rect 86192 124000 86256 124004
rect 89952 124060 90016 124064
rect 89952 124004 89956 124060
rect 89956 124004 90012 124060
rect 90012 124004 90016 124060
rect 89952 124000 90016 124004
rect 90032 124060 90096 124064
rect 90032 124004 90036 124060
rect 90036 124004 90092 124060
rect 90092 124004 90096 124060
rect 90032 124000 90096 124004
rect 90112 124060 90176 124064
rect 90112 124004 90116 124060
rect 90116 124004 90172 124060
rect 90172 124004 90176 124060
rect 90112 124000 90176 124004
rect 90192 124060 90256 124064
rect 90192 124004 90196 124060
rect 90196 124004 90252 124060
rect 90252 124004 90256 124060
rect 90192 124000 90256 124004
rect 3952 123516 4016 123520
rect 3952 123460 3956 123516
rect 3956 123460 4012 123516
rect 4012 123460 4016 123516
rect 3952 123456 4016 123460
rect 4032 123516 4096 123520
rect 4032 123460 4036 123516
rect 4036 123460 4092 123516
rect 4092 123460 4096 123516
rect 4032 123456 4096 123460
rect 4112 123516 4176 123520
rect 4112 123460 4116 123516
rect 4116 123460 4172 123516
rect 4172 123460 4176 123516
rect 4112 123456 4176 123460
rect 4192 123516 4256 123520
rect 4192 123460 4196 123516
rect 4196 123460 4252 123516
rect 4252 123460 4256 123516
rect 4192 123456 4256 123460
rect 87952 123516 88016 123520
rect 87952 123460 87956 123516
rect 87956 123460 88012 123516
rect 88012 123460 88016 123516
rect 87952 123456 88016 123460
rect 88032 123516 88096 123520
rect 88032 123460 88036 123516
rect 88036 123460 88092 123516
rect 88092 123460 88096 123516
rect 88032 123456 88096 123460
rect 88112 123516 88176 123520
rect 88112 123460 88116 123516
rect 88116 123460 88172 123516
rect 88172 123460 88176 123516
rect 88112 123456 88176 123460
rect 88192 123516 88256 123520
rect 88192 123460 88196 123516
rect 88196 123460 88252 123516
rect 88252 123460 88256 123516
rect 88192 123456 88256 123460
rect 1952 122972 2016 122976
rect 1952 122916 1956 122972
rect 1956 122916 2012 122972
rect 2012 122916 2016 122972
rect 1952 122912 2016 122916
rect 2032 122972 2096 122976
rect 2032 122916 2036 122972
rect 2036 122916 2092 122972
rect 2092 122916 2096 122972
rect 2032 122912 2096 122916
rect 2112 122972 2176 122976
rect 2112 122916 2116 122972
rect 2116 122916 2172 122972
rect 2172 122916 2176 122972
rect 2112 122912 2176 122916
rect 2192 122972 2256 122976
rect 2192 122916 2196 122972
rect 2196 122916 2252 122972
rect 2252 122916 2256 122972
rect 2192 122912 2256 122916
rect 85952 122972 86016 122976
rect 85952 122916 85956 122972
rect 85956 122916 86012 122972
rect 86012 122916 86016 122972
rect 85952 122912 86016 122916
rect 86032 122972 86096 122976
rect 86032 122916 86036 122972
rect 86036 122916 86092 122972
rect 86092 122916 86096 122972
rect 86032 122912 86096 122916
rect 86112 122972 86176 122976
rect 86112 122916 86116 122972
rect 86116 122916 86172 122972
rect 86172 122916 86176 122972
rect 86112 122912 86176 122916
rect 86192 122972 86256 122976
rect 86192 122916 86196 122972
rect 86196 122916 86252 122972
rect 86252 122916 86256 122972
rect 86192 122912 86256 122916
rect 89952 122972 90016 122976
rect 89952 122916 89956 122972
rect 89956 122916 90012 122972
rect 90012 122916 90016 122972
rect 89952 122912 90016 122916
rect 90032 122972 90096 122976
rect 90032 122916 90036 122972
rect 90036 122916 90092 122972
rect 90092 122916 90096 122972
rect 90032 122912 90096 122916
rect 90112 122972 90176 122976
rect 90112 122916 90116 122972
rect 90116 122916 90172 122972
rect 90172 122916 90176 122972
rect 90112 122912 90176 122916
rect 90192 122972 90256 122976
rect 90192 122916 90196 122972
rect 90196 122916 90252 122972
rect 90252 122916 90256 122972
rect 90192 122912 90256 122916
rect 86908 122572 86972 122636
rect 90588 122572 90652 122636
rect 3952 122428 4016 122432
rect 3952 122372 3956 122428
rect 3956 122372 4012 122428
rect 4012 122372 4016 122428
rect 3952 122368 4016 122372
rect 4032 122428 4096 122432
rect 4032 122372 4036 122428
rect 4036 122372 4092 122428
rect 4092 122372 4096 122428
rect 4032 122368 4096 122372
rect 4112 122428 4176 122432
rect 4112 122372 4116 122428
rect 4116 122372 4172 122428
rect 4172 122372 4176 122428
rect 4112 122368 4176 122372
rect 4192 122428 4256 122432
rect 4192 122372 4196 122428
rect 4196 122372 4252 122428
rect 4252 122372 4256 122428
rect 4192 122368 4256 122372
rect 87952 122428 88016 122432
rect 87952 122372 87956 122428
rect 87956 122372 88012 122428
rect 88012 122372 88016 122428
rect 87952 122368 88016 122372
rect 88032 122428 88096 122432
rect 88032 122372 88036 122428
rect 88036 122372 88092 122428
rect 88092 122372 88096 122428
rect 88032 122368 88096 122372
rect 88112 122428 88176 122432
rect 88112 122372 88116 122428
rect 88116 122372 88172 122428
rect 88172 122372 88176 122428
rect 88112 122368 88176 122372
rect 88192 122428 88256 122432
rect 88192 122372 88196 122428
rect 88196 122372 88252 122428
rect 88252 122372 88256 122428
rect 88192 122368 88256 122372
rect 86908 122300 86972 122364
rect 1952 121884 2016 121888
rect 1952 121828 1956 121884
rect 1956 121828 2012 121884
rect 2012 121828 2016 121884
rect 1952 121824 2016 121828
rect 2032 121884 2096 121888
rect 2032 121828 2036 121884
rect 2036 121828 2092 121884
rect 2092 121828 2096 121884
rect 2032 121824 2096 121828
rect 2112 121884 2176 121888
rect 2112 121828 2116 121884
rect 2116 121828 2172 121884
rect 2172 121828 2176 121884
rect 2112 121824 2176 121828
rect 2192 121884 2256 121888
rect 2192 121828 2196 121884
rect 2196 121828 2252 121884
rect 2252 121828 2256 121884
rect 2192 121824 2256 121828
rect 85952 121884 86016 121888
rect 85952 121828 85956 121884
rect 85956 121828 86012 121884
rect 86012 121828 86016 121884
rect 85952 121824 86016 121828
rect 86032 121884 86096 121888
rect 86032 121828 86036 121884
rect 86036 121828 86092 121884
rect 86092 121828 86096 121884
rect 86032 121824 86096 121828
rect 86112 121884 86176 121888
rect 86112 121828 86116 121884
rect 86116 121828 86172 121884
rect 86172 121828 86176 121884
rect 86112 121824 86176 121828
rect 86192 121884 86256 121888
rect 86192 121828 86196 121884
rect 86196 121828 86252 121884
rect 86252 121828 86256 121884
rect 86192 121824 86256 121828
rect 89952 121884 90016 121888
rect 89952 121828 89956 121884
rect 89956 121828 90012 121884
rect 90012 121828 90016 121884
rect 89952 121824 90016 121828
rect 90032 121884 90096 121888
rect 90032 121828 90036 121884
rect 90036 121828 90092 121884
rect 90092 121828 90096 121884
rect 90032 121824 90096 121828
rect 90112 121884 90176 121888
rect 90112 121828 90116 121884
rect 90116 121828 90172 121884
rect 90172 121828 90176 121884
rect 90112 121824 90176 121828
rect 90192 121884 90256 121888
rect 90192 121828 90196 121884
rect 90196 121828 90252 121884
rect 90252 121828 90256 121884
rect 90192 121824 90256 121828
rect 6132 121484 6196 121548
rect 3952 121340 4016 121344
rect 3952 121284 3956 121340
rect 3956 121284 4012 121340
rect 4012 121284 4016 121340
rect 3952 121280 4016 121284
rect 4032 121340 4096 121344
rect 4032 121284 4036 121340
rect 4036 121284 4092 121340
rect 4092 121284 4096 121340
rect 4032 121280 4096 121284
rect 4112 121340 4176 121344
rect 4112 121284 4116 121340
rect 4116 121284 4172 121340
rect 4172 121284 4176 121340
rect 4112 121280 4176 121284
rect 4192 121340 4256 121344
rect 4192 121284 4196 121340
rect 4196 121284 4252 121340
rect 4252 121284 4256 121340
rect 4192 121280 4256 121284
rect 87952 121340 88016 121344
rect 87952 121284 87956 121340
rect 87956 121284 88012 121340
rect 88012 121284 88016 121340
rect 87952 121280 88016 121284
rect 88032 121340 88096 121344
rect 88032 121284 88036 121340
rect 88036 121284 88092 121340
rect 88092 121284 88096 121340
rect 88032 121280 88096 121284
rect 88112 121340 88176 121344
rect 88112 121284 88116 121340
rect 88116 121284 88172 121340
rect 88172 121284 88176 121340
rect 88112 121280 88176 121284
rect 88192 121340 88256 121344
rect 88192 121284 88196 121340
rect 88196 121284 88252 121340
rect 88252 121284 88256 121340
rect 88192 121280 88256 121284
rect 1952 120796 2016 120800
rect 1952 120740 1956 120796
rect 1956 120740 2012 120796
rect 2012 120740 2016 120796
rect 1952 120736 2016 120740
rect 2032 120796 2096 120800
rect 2032 120740 2036 120796
rect 2036 120740 2092 120796
rect 2092 120740 2096 120796
rect 2032 120736 2096 120740
rect 2112 120796 2176 120800
rect 2112 120740 2116 120796
rect 2116 120740 2172 120796
rect 2172 120740 2176 120796
rect 2112 120736 2176 120740
rect 2192 120796 2256 120800
rect 2192 120740 2196 120796
rect 2196 120740 2252 120796
rect 2252 120740 2256 120796
rect 2192 120736 2256 120740
rect 85952 120796 86016 120800
rect 85952 120740 85956 120796
rect 85956 120740 86012 120796
rect 86012 120740 86016 120796
rect 85952 120736 86016 120740
rect 86032 120796 86096 120800
rect 86032 120740 86036 120796
rect 86036 120740 86092 120796
rect 86092 120740 86096 120796
rect 86032 120736 86096 120740
rect 86112 120796 86176 120800
rect 86112 120740 86116 120796
rect 86116 120740 86172 120796
rect 86172 120740 86176 120796
rect 86112 120736 86176 120740
rect 86192 120796 86256 120800
rect 86192 120740 86196 120796
rect 86196 120740 86252 120796
rect 86252 120740 86256 120796
rect 86192 120736 86256 120740
rect 89952 120796 90016 120800
rect 89952 120740 89956 120796
rect 89956 120740 90012 120796
rect 90012 120740 90016 120796
rect 89952 120736 90016 120740
rect 90032 120796 90096 120800
rect 90032 120740 90036 120796
rect 90036 120740 90092 120796
rect 90092 120740 90096 120796
rect 90032 120736 90096 120740
rect 90112 120796 90176 120800
rect 90112 120740 90116 120796
rect 90116 120740 90172 120796
rect 90172 120740 90176 120796
rect 90112 120736 90176 120740
rect 90192 120796 90256 120800
rect 90192 120740 90196 120796
rect 90196 120740 90252 120796
rect 90252 120740 90256 120796
rect 90192 120736 90256 120740
rect 3952 120252 4016 120256
rect 3952 120196 3956 120252
rect 3956 120196 4012 120252
rect 4012 120196 4016 120252
rect 3952 120192 4016 120196
rect 4032 120252 4096 120256
rect 4032 120196 4036 120252
rect 4036 120196 4092 120252
rect 4092 120196 4096 120252
rect 4032 120192 4096 120196
rect 4112 120252 4176 120256
rect 4112 120196 4116 120252
rect 4116 120196 4172 120252
rect 4172 120196 4176 120252
rect 4112 120192 4176 120196
rect 4192 120252 4256 120256
rect 4192 120196 4196 120252
rect 4196 120196 4252 120252
rect 4252 120196 4256 120252
rect 4192 120192 4256 120196
rect 87952 120252 88016 120256
rect 87952 120196 87956 120252
rect 87956 120196 88012 120252
rect 88012 120196 88016 120252
rect 87952 120192 88016 120196
rect 88032 120252 88096 120256
rect 88032 120196 88036 120252
rect 88036 120196 88092 120252
rect 88092 120196 88096 120252
rect 88032 120192 88096 120196
rect 88112 120252 88176 120256
rect 88112 120196 88116 120252
rect 88116 120196 88172 120252
rect 88172 120196 88176 120252
rect 88112 120192 88176 120196
rect 88192 120252 88256 120256
rect 88192 120196 88196 120252
rect 88196 120196 88252 120252
rect 88252 120196 88256 120252
rect 88192 120192 88256 120196
rect 84332 120124 84396 120188
rect 1952 119708 2016 119712
rect 1952 119652 1956 119708
rect 1956 119652 2012 119708
rect 2012 119652 2016 119708
rect 1952 119648 2016 119652
rect 2032 119708 2096 119712
rect 2032 119652 2036 119708
rect 2036 119652 2092 119708
rect 2092 119652 2096 119708
rect 2032 119648 2096 119652
rect 2112 119708 2176 119712
rect 2112 119652 2116 119708
rect 2116 119652 2172 119708
rect 2172 119652 2176 119708
rect 2112 119648 2176 119652
rect 2192 119708 2256 119712
rect 2192 119652 2196 119708
rect 2196 119652 2252 119708
rect 2252 119652 2256 119708
rect 2192 119648 2256 119652
rect 85952 119708 86016 119712
rect 85952 119652 85956 119708
rect 85956 119652 86012 119708
rect 86012 119652 86016 119708
rect 85952 119648 86016 119652
rect 86032 119708 86096 119712
rect 86032 119652 86036 119708
rect 86036 119652 86092 119708
rect 86092 119652 86096 119708
rect 86032 119648 86096 119652
rect 86112 119708 86176 119712
rect 86112 119652 86116 119708
rect 86116 119652 86172 119708
rect 86172 119652 86176 119708
rect 86112 119648 86176 119652
rect 86192 119708 86256 119712
rect 86192 119652 86196 119708
rect 86196 119652 86252 119708
rect 86252 119652 86256 119708
rect 86192 119648 86256 119652
rect 89952 119708 90016 119712
rect 89952 119652 89956 119708
rect 89956 119652 90012 119708
rect 90012 119652 90016 119708
rect 89952 119648 90016 119652
rect 90032 119708 90096 119712
rect 90032 119652 90036 119708
rect 90036 119652 90092 119708
rect 90092 119652 90096 119708
rect 90032 119648 90096 119652
rect 90112 119708 90176 119712
rect 90112 119652 90116 119708
rect 90116 119652 90172 119708
rect 90172 119652 90176 119708
rect 90112 119648 90176 119652
rect 90192 119708 90256 119712
rect 90192 119652 90196 119708
rect 90196 119652 90252 119708
rect 90252 119652 90256 119708
rect 90192 119648 90256 119652
rect 3952 119164 4016 119168
rect 3952 119108 3956 119164
rect 3956 119108 4012 119164
rect 4012 119108 4016 119164
rect 3952 119104 4016 119108
rect 4032 119164 4096 119168
rect 4032 119108 4036 119164
rect 4036 119108 4092 119164
rect 4092 119108 4096 119164
rect 4032 119104 4096 119108
rect 4112 119164 4176 119168
rect 4112 119108 4116 119164
rect 4116 119108 4172 119164
rect 4172 119108 4176 119164
rect 4112 119104 4176 119108
rect 4192 119164 4256 119168
rect 4192 119108 4196 119164
rect 4196 119108 4252 119164
rect 4252 119108 4256 119164
rect 4192 119104 4256 119108
rect 87952 119164 88016 119168
rect 87952 119108 87956 119164
rect 87956 119108 88012 119164
rect 88012 119108 88016 119164
rect 87952 119104 88016 119108
rect 88032 119164 88096 119168
rect 88032 119108 88036 119164
rect 88036 119108 88092 119164
rect 88092 119108 88096 119164
rect 88032 119104 88096 119108
rect 88112 119164 88176 119168
rect 88112 119108 88116 119164
rect 88116 119108 88172 119164
rect 88172 119108 88176 119164
rect 88112 119104 88176 119108
rect 88192 119164 88256 119168
rect 88192 119108 88196 119164
rect 88196 119108 88252 119164
rect 88252 119108 88256 119164
rect 88192 119104 88256 119108
rect 1952 118620 2016 118624
rect 1952 118564 1956 118620
rect 1956 118564 2012 118620
rect 2012 118564 2016 118620
rect 1952 118560 2016 118564
rect 2032 118620 2096 118624
rect 2032 118564 2036 118620
rect 2036 118564 2092 118620
rect 2092 118564 2096 118620
rect 2032 118560 2096 118564
rect 2112 118620 2176 118624
rect 2112 118564 2116 118620
rect 2116 118564 2172 118620
rect 2172 118564 2176 118620
rect 2112 118560 2176 118564
rect 2192 118620 2256 118624
rect 2192 118564 2196 118620
rect 2196 118564 2252 118620
rect 2252 118564 2256 118620
rect 2192 118560 2256 118564
rect 85952 118620 86016 118624
rect 85952 118564 85956 118620
rect 85956 118564 86012 118620
rect 86012 118564 86016 118620
rect 85952 118560 86016 118564
rect 86032 118620 86096 118624
rect 86032 118564 86036 118620
rect 86036 118564 86092 118620
rect 86092 118564 86096 118620
rect 86032 118560 86096 118564
rect 86112 118620 86176 118624
rect 86112 118564 86116 118620
rect 86116 118564 86172 118620
rect 86172 118564 86176 118620
rect 86112 118560 86176 118564
rect 86192 118620 86256 118624
rect 86192 118564 86196 118620
rect 86196 118564 86252 118620
rect 86252 118564 86256 118620
rect 86192 118560 86256 118564
rect 89952 118620 90016 118624
rect 89952 118564 89956 118620
rect 89956 118564 90012 118620
rect 90012 118564 90016 118620
rect 89952 118560 90016 118564
rect 90032 118620 90096 118624
rect 90032 118564 90036 118620
rect 90036 118564 90092 118620
rect 90092 118564 90096 118620
rect 90032 118560 90096 118564
rect 90112 118620 90176 118624
rect 90112 118564 90116 118620
rect 90116 118564 90172 118620
rect 90172 118564 90176 118620
rect 90112 118560 90176 118564
rect 90192 118620 90256 118624
rect 90192 118564 90196 118620
rect 90196 118564 90252 118620
rect 90252 118564 90256 118620
rect 90192 118560 90256 118564
rect 86908 118492 86972 118556
rect 3952 118076 4016 118080
rect 3952 118020 3956 118076
rect 3956 118020 4012 118076
rect 4012 118020 4016 118076
rect 3952 118016 4016 118020
rect 4032 118076 4096 118080
rect 4032 118020 4036 118076
rect 4036 118020 4092 118076
rect 4092 118020 4096 118076
rect 4032 118016 4096 118020
rect 4112 118076 4176 118080
rect 4112 118020 4116 118076
rect 4116 118020 4172 118076
rect 4172 118020 4176 118076
rect 4112 118016 4176 118020
rect 4192 118076 4256 118080
rect 4192 118020 4196 118076
rect 4196 118020 4252 118076
rect 4252 118020 4256 118076
rect 4192 118016 4256 118020
rect 87952 118076 88016 118080
rect 87952 118020 87956 118076
rect 87956 118020 88012 118076
rect 88012 118020 88016 118076
rect 87952 118016 88016 118020
rect 88032 118076 88096 118080
rect 88032 118020 88036 118076
rect 88036 118020 88092 118076
rect 88092 118020 88096 118076
rect 88032 118016 88096 118020
rect 88112 118076 88176 118080
rect 88112 118020 88116 118076
rect 88116 118020 88172 118076
rect 88172 118020 88176 118076
rect 88112 118016 88176 118020
rect 88192 118076 88256 118080
rect 88192 118020 88196 118076
rect 88196 118020 88252 118076
rect 88252 118020 88256 118076
rect 88192 118016 88256 118020
rect 1952 117532 2016 117536
rect 1952 117476 1956 117532
rect 1956 117476 2012 117532
rect 2012 117476 2016 117532
rect 1952 117472 2016 117476
rect 2032 117532 2096 117536
rect 2032 117476 2036 117532
rect 2036 117476 2092 117532
rect 2092 117476 2096 117532
rect 2032 117472 2096 117476
rect 2112 117532 2176 117536
rect 2112 117476 2116 117532
rect 2116 117476 2172 117532
rect 2172 117476 2176 117532
rect 2112 117472 2176 117476
rect 2192 117532 2256 117536
rect 2192 117476 2196 117532
rect 2196 117476 2252 117532
rect 2252 117476 2256 117532
rect 2192 117472 2256 117476
rect 85952 117532 86016 117536
rect 85952 117476 85956 117532
rect 85956 117476 86012 117532
rect 86012 117476 86016 117532
rect 85952 117472 86016 117476
rect 86032 117532 86096 117536
rect 86032 117476 86036 117532
rect 86036 117476 86092 117532
rect 86092 117476 86096 117532
rect 86032 117472 86096 117476
rect 86112 117532 86176 117536
rect 86112 117476 86116 117532
rect 86116 117476 86172 117532
rect 86172 117476 86176 117532
rect 86112 117472 86176 117476
rect 86192 117532 86256 117536
rect 86192 117476 86196 117532
rect 86196 117476 86252 117532
rect 86252 117476 86256 117532
rect 86192 117472 86256 117476
rect 89952 117532 90016 117536
rect 89952 117476 89956 117532
rect 89956 117476 90012 117532
rect 90012 117476 90016 117532
rect 89952 117472 90016 117476
rect 90032 117532 90096 117536
rect 90032 117476 90036 117532
rect 90036 117476 90092 117532
rect 90092 117476 90096 117532
rect 90032 117472 90096 117476
rect 90112 117532 90176 117536
rect 90112 117476 90116 117532
rect 90116 117476 90172 117532
rect 90172 117476 90176 117532
rect 90112 117472 90176 117476
rect 90192 117532 90256 117536
rect 90192 117476 90196 117532
rect 90196 117476 90252 117532
rect 90252 117476 90256 117532
rect 90192 117472 90256 117476
rect 3952 116988 4016 116992
rect 3952 116932 3956 116988
rect 3956 116932 4012 116988
rect 4012 116932 4016 116988
rect 3952 116928 4016 116932
rect 4032 116988 4096 116992
rect 4032 116932 4036 116988
rect 4036 116932 4092 116988
rect 4092 116932 4096 116988
rect 4032 116928 4096 116932
rect 4112 116988 4176 116992
rect 4112 116932 4116 116988
rect 4116 116932 4172 116988
rect 4172 116932 4176 116988
rect 4112 116928 4176 116932
rect 4192 116988 4256 116992
rect 4192 116932 4196 116988
rect 4196 116932 4252 116988
rect 4252 116932 4256 116988
rect 4192 116928 4256 116932
rect 87952 116988 88016 116992
rect 87952 116932 87956 116988
rect 87956 116932 88012 116988
rect 88012 116932 88016 116988
rect 87952 116928 88016 116932
rect 88032 116988 88096 116992
rect 88032 116932 88036 116988
rect 88036 116932 88092 116988
rect 88092 116932 88096 116988
rect 88032 116928 88096 116932
rect 88112 116988 88176 116992
rect 88112 116932 88116 116988
rect 88116 116932 88172 116988
rect 88172 116932 88176 116988
rect 88112 116928 88176 116932
rect 88192 116988 88256 116992
rect 88192 116932 88196 116988
rect 88196 116932 88252 116988
rect 88252 116932 88256 116988
rect 88192 116928 88256 116932
rect 5396 116648 5460 116652
rect 5396 116592 5410 116648
rect 5410 116592 5460 116648
rect 5396 116588 5460 116592
rect 1952 116444 2016 116448
rect 1952 116388 1956 116444
rect 1956 116388 2012 116444
rect 2012 116388 2016 116444
rect 1952 116384 2016 116388
rect 2032 116444 2096 116448
rect 2032 116388 2036 116444
rect 2036 116388 2092 116444
rect 2092 116388 2096 116444
rect 2032 116384 2096 116388
rect 2112 116444 2176 116448
rect 2112 116388 2116 116444
rect 2116 116388 2172 116444
rect 2172 116388 2176 116444
rect 2112 116384 2176 116388
rect 2192 116444 2256 116448
rect 2192 116388 2196 116444
rect 2196 116388 2252 116444
rect 2252 116388 2256 116444
rect 2192 116384 2256 116388
rect 85952 116444 86016 116448
rect 85952 116388 85956 116444
rect 85956 116388 86012 116444
rect 86012 116388 86016 116444
rect 85952 116384 86016 116388
rect 86032 116444 86096 116448
rect 86032 116388 86036 116444
rect 86036 116388 86092 116444
rect 86092 116388 86096 116444
rect 86032 116384 86096 116388
rect 86112 116444 86176 116448
rect 86112 116388 86116 116444
rect 86116 116388 86172 116444
rect 86172 116388 86176 116444
rect 86112 116384 86176 116388
rect 86192 116444 86256 116448
rect 86192 116388 86196 116444
rect 86196 116388 86252 116444
rect 86252 116388 86256 116444
rect 86192 116384 86256 116388
rect 89952 116444 90016 116448
rect 89952 116388 89956 116444
rect 89956 116388 90012 116444
rect 90012 116388 90016 116444
rect 89952 116384 90016 116388
rect 90032 116444 90096 116448
rect 90032 116388 90036 116444
rect 90036 116388 90092 116444
rect 90092 116388 90096 116444
rect 90032 116384 90096 116388
rect 90112 116444 90176 116448
rect 90112 116388 90116 116444
rect 90116 116388 90172 116444
rect 90172 116388 90176 116444
rect 90112 116384 90176 116388
rect 90192 116444 90256 116448
rect 90192 116388 90196 116444
rect 90196 116388 90252 116444
rect 90252 116388 90256 116444
rect 90192 116384 90256 116388
rect 3952 115900 4016 115904
rect 3952 115844 3956 115900
rect 3956 115844 4012 115900
rect 4012 115844 4016 115900
rect 3952 115840 4016 115844
rect 4032 115900 4096 115904
rect 4032 115844 4036 115900
rect 4036 115844 4092 115900
rect 4092 115844 4096 115900
rect 4032 115840 4096 115844
rect 4112 115900 4176 115904
rect 4112 115844 4116 115900
rect 4116 115844 4172 115900
rect 4172 115844 4176 115900
rect 4112 115840 4176 115844
rect 4192 115900 4256 115904
rect 4192 115844 4196 115900
rect 4196 115844 4252 115900
rect 4252 115844 4256 115900
rect 4192 115840 4256 115844
rect 87952 115900 88016 115904
rect 87952 115844 87956 115900
rect 87956 115844 88012 115900
rect 88012 115844 88016 115900
rect 87952 115840 88016 115844
rect 88032 115900 88096 115904
rect 88032 115844 88036 115900
rect 88036 115844 88092 115900
rect 88092 115844 88096 115900
rect 88032 115840 88096 115844
rect 88112 115900 88176 115904
rect 88112 115844 88116 115900
rect 88116 115844 88172 115900
rect 88172 115844 88176 115900
rect 88112 115840 88176 115844
rect 88192 115900 88256 115904
rect 88192 115844 88196 115900
rect 88196 115844 88252 115900
rect 88252 115844 88256 115900
rect 88192 115840 88256 115844
rect 1952 115356 2016 115360
rect 1952 115300 1956 115356
rect 1956 115300 2012 115356
rect 2012 115300 2016 115356
rect 1952 115296 2016 115300
rect 2032 115356 2096 115360
rect 2032 115300 2036 115356
rect 2036 115300 2092 115356
rect 2092 115300 2096 115356
rect 2032 115296 2096 115300
rect 2112 115356 2176 115360
rect 2112 115300 2116 115356
rect 2116 115300 2172 115356
rect 2172 115300 2176 115356
rect 2112 115296 2176 115300
rect 2192 115356 2256 115360
rect 2192 115300 2196 115356
rect 2196 115300 2252 115356
rect 2252 115300 2256 115356
rect 2192 115296 2256 115300
rect 85952 115356 86016 115360
rect 85952 115300 85956 115356
rect 85956 115300 86012 115356
rect 86012 115300 86016 115356
rect 85952 115296 86016 115300
rect 86032 115356 86096 115360
rect 86032 115300 86036 115356
rect 86036 115300 86092 115356
rect 86092 115300 86096 115356
rect 86032 115296 86096 115300
rect 86112 115356 86176 115360
rect 86112 115300 86116 115356
rect 86116 115300 86172 115356
rect 86172 115300 86176 115356
rect 86112 115296 86176 115300
rect 86192 115356 86256 115360
rect 86192 115300 86196 115356
rect 86196 115300 86252 115356
rect 86252 115300 86256 115356
rect 86192 115296 86256 115300
rect 89952 115356 90016 115360
rect 89952 115300 89956 115356
rect 89956 115300 90012 115356
rect 90012 115300 90016 115356
rect 89952 115296 90016 115300
rect 90032 115356 90096 115360
rect 90032 115300 90036 115356
rect 90036 115300 90092 115356
rect 90092 115300 90096 115356
rect 90032 115296 90096 115300
rect 90112 115356 90176 115360
rect 90112 115300 90116 115356
rect 90116 115300 90172 115356
rect 90172 115300 90176 115356
rect 90112 115296 90176 115300
rect 90192 115356 90256 115360
rect 90192 115300 90196 115356
rect 90196 115300 90252 115356
rect 90252 115300 90256 115356
rect 90192 115296 90256 115300
rect 3952 114812 4016 114816
rect 3952 114756 3956 114812
rect 3956 114756 4012 114812
rect 4012 114756 4016 114812
rect 3952 114752 4016 114756
rect 4032 114812 4096 114816
rect 4032 114756 4036 114812
rect 4036 114756 4092 114812
rect 4092 114756 4096 114812
rect 4032 114752 4096 114756
rect 4112 114812 4176 114816
rect 4112 114756 4116 114812
rect 4116 114756 4172 114812
rect 4172 114756 4176 114812
rect 4112 114752 4176 114756
rect 4192 114812 4256 114816
rect 4192 114756 4196 114812
rect 4196 114756 4252 114812
rect 4252 114756 4256 114812
rect 4192 114752 4256 114756
rect 87952 114812 88016 114816
rect 87952 114756 87956 114812
rect 87956 114756 88012 114812
rect 88012 114756 88016 114812
rect 87952 114752 88016 114756
rect 88032 114812 88096 114816
rect 88032 114756 88036 114812
rect 88036 114756 88092 114812
rect 88092 114756 88096 114812
rect 88032 114752 88096 114756
rect 88112 114812 88176 114816
rect 88112 114756 88116 114812
rect 88116 114756 88172 114812
rect 88172 114756 88176 114812
rect 88112 114752 88176 114756
rect 88192 114812 88256 114816
rect 88192 114756 88196 114812
rect 88196 114756 88252 114812
rect 88252 114756 88256 114812
rect 88192 114752 88256 114756
rect 83412 114276 83476 114340
rect 1952 114268 2016 114272
rect 1952 114212 1956 114268
rect 1956 114212 2012 114268
rect 2012 114212 2016 114268
rect 1952 114208 2016 114212
rect 2032 114268 2096 114272
rect 2032 114212 2036 114268
rect 2036 114212 2092 114268
rect 2092 114212 2096 114268
rect 2032 114208 2096 114212
rect 2112 114268 2176 114272
rect 2112 114212 2116 114268
rect 2116 114212 2172 114268
rect 2172 114212 2176 114268
rect 2112 114208 2176 114212
rect 2192 114268 2256 114272
rect 2192 114212 2196 114268
rect 2196 114212 2252 114268
rect 2252 114212 2256 114268
rect 2192 114208 2256 114212
rect 85952 114268 86016 114272
rect 85952 114212 85956 114268
rect 85956 114212 86012 114268
rect 86012 114212 86016 114268
rect 85952 114208 86016 114212
rect 86032 114268 86096 114272
rect 86032 114212 86036 114268
rect 86036 114212 86092 114268
rect 86092 114212 86096 114268
rect 86032 114208 86096 114212
rect 86112 114268 86176 114272
rect 86112 114212 86116 114268
rect 86116 114212 86172 114268
rect 86172 114212 86176 114268
rect 86112 114208 86176 114212
rect 86192 114268 86256 114272
rect 86192 114212 86196 114268
rect 86196 114212 86252 114268
rect 86252 114212 86256 114268
rect 86192 114208 86256 114212
rect 89952 114268 90016 114272
rect 89952 114212 89956 114268
rect 89956 114212 90012 114268
rect 90012 114212 90016 114268
rect 89952 114208 90016 114212
rect 90032 114268 90096 114272
rect 90032 114212 90036 114268
rect 90036 114212 90092 114268
rect 90092 114212 90096 114268
rect 90032 114208 90096 114212
rect 90112 114268 90176 114272
rect 90112 114212 90116 114268
rect 90116 114212 90172 114268
rect 90172 114212 90176 114268
rect 90112 114208 90176 114212
rect 90192 114268 90256 114272
rect 90192 114212 90196 114268
rect 90196 114212 90252 114268
rect 90252 114212 90256 114268
rect 90192 114208 90256 114212
rect 83412 113868 83476 113932
rect 83964 113868 84028 113932
rect 3952 113724 4016 113728
rect 3952 113668 3956 113724
rect 3956 113668 4012 113724
rect 4012 113668 4016 113724
rect 3952 113664 4016 113668
rect 4032 113724 4096 113728
rect 4032 113668 4036 113724
rect 4036 113668 4092 113724
rect 4092 113668 4096 113724
rect 4032 113664 4096 113668
rect 4112 113724 4176 113728
rect 4112 113668 4116 113724
rect 4116 113668 4172 113724
rect 4172 113668 4176 113724
rect 4112 113664 4176 113668
rect 4192 113724 4256 113728
rect 4192 113668 4196 113724
rect 4196 113668 4252 113724
rect 4252 113668 4256 113724
rect 4192 113664 4256 113668
rect 87952 113724 88016 113728
rect 87952 113668 87956 113724
rect 87956 113668 88012 113724
rect 88012 113668 88016 113724
rect 87952 113664 88016 113668
rect 88032 113724 88096 113728
rect 88032 113668 88036 113724
rect 88036 113668 88092 113724
rect 88092 113668 88096 113724
rect 88032 113664 88096 113668
rect 88112 113724 88176 113728
rect 88112 113668 88116 113724
rect 88116 113668 88172 113724
rect 88172 113668 88176 113724
rect 88112 113664 88176 113668
rect 88192 113724 88256 113728
rect 88192 113668 88196 113724
rect 88196 113668 88252 113724
rect 88252 113668 88256 113724
rect 88192 113664 88256 113668
rect 1952 113180 2016 113184
rect 1952 113124 1956 113180
rect 1956 113124 2012 113180
rect 2012 113124 2016 113180
rect 1952 113120 2016 113124
rect 2032 113180 2096 113184
rect 2032 113124 2036 113180
rect 2036 113124 2092 113180
rect 2092 113124 2096 113180
rect 2032 113120 2096 113124
rect 2112 113180 2176 113184
rect 2112 113124 2116 113180
rect 2116 113124 2172 113180
rect 2172 113124 2176 113180
rect 2112 113120 2176 113124
rect 2192 113180 2256 113184
rect 2192 113124 2196 113180
rect 2196 113124 2252 113180
rect 2252 113124 2256 113180
rect 2192 113120 2256 113124
rect 85952 113180 86016 113184
rect 85952 113124 85956 113180
rect 85956 113124 86012 113180
rect 86012 113124 86016 113180
rect 85952 113120 86016 113124
rect 86032 113180 86096 113184
rect 86032 113124 86036 113180
rect 86036 113124 86092 113180
rect 86092 113124 86096 113180
rect 86032 113120 86096 113124
rect 86112 113180 86176 113184
rect 86112 113124 86116 113180
rect 86116 113124 86172 113180
rect 86172 113124 86176 113180
rect 86112 113120 86176 113124
rect 86192 113180 86256 113184
rect 86192 113124 86196 113180
rect 86196 113124 86252 113180
rect 86252 113124 86256 113180
rect 86192 113120 86256 113124
rect 89952 113180 90016 113184
rect 89952 113124 89956 113180
rect 89956 113124 90012 113180
rect 90012 113124 90016 113180
rect 89952 113120 90016 113124
rect 90032 113180 90096 113184
rect 90032 113124 90036 113180
rect 90036 113124 90092 113180
rect 90092 113124 90096 113180
rect 90032 113120 90096 113124
rect 90112 113180 90176 113184
rect 90112 113124 90116 113180
rect 90116 113124 90172 113180
rect 90172 113124 90176 113180
rect 90112 113120 90176 113124
rect 90192 113180 90256 113184
rect 90192 113124 90196 113180
rect 90196 113124 90252 113180
rect 90252 113124 90256 113180
rect 90192 113120 90256 113124
rect 3952 112636 4016 112640
rect 3952 112580 3956 112636
rect 3956 112580 4012 112636
rect 4012 112580 4016 112636
rect 3952 112576 4016 112580
rect 4032 112636 4096 112640
rect 4032 112580 4036 112636
rect 4036 112580 4092 112636
rect 4092 112580 4096 112636
rect 4032 112576 4096 112580
rect 4112 112636 4176 112640
rect 4112 112580 4116 112636
rect 4116 112580 4172 112636
rect 4172 112580 4176 112636
rect 4112 112576 4176 112580
rect 4192 112636 4256 112640
rect 4192 112580 4196 112636
rect 4196 112580 4252 112636
rect 4252 112580 4256 112636
rect 4192 112576 4256 112580
rect 87952 112636 88016 112640
rect 87952 112580 87956 112636
rect 87956 112580 88012 112636
rect 88012 112580 88016 112636
rect 87952 112576 88016 112580
rect 88032 112636 88096 112640
rect 88032 112580 88036 112636
rect 88036 112580 88092 112636
rect 88092 112580 88096 112636
rect 88032 112576 88096 112580
rect 88112 112636 88176 112640
rect 88112 112580 88116 112636
rect 88116 112580 88172 112636
rect 88172 112580 88176 112636
rect 88112 112576 88176 112580
rect 88192 112636 88256 112640
rect 88192 112580 88196 112636
rect 88196 112580 88252 112636
rect 88252 112580 88256 112636
rect 88192 112576 88256 112580
rect 1952 112092 2016 112096
rect 1952 112036 1956 112092
rect 1956 112036 2012 112092
rect 2012 112036 2016 112092
rect 1952 112032 2016 112036
rect 2032 112092 2096 112096
rect 2032 112036 2036 112092
rect 2036 112036 2092 112092
rect 2092 112036 2096 112092
rect 2032 112032 2096 112036
rect 2112 112092 2176 112096
rect 2112 112036 2116 112092
rect 2116 112036 2172 112092
rect 2172 112036 2176 112092
rect 2112 112032 2176 112036
rect 2192 112092 2256 112096
rect 2192 112036 2196 112092
rect 2196 112036 2252 112092
rect 2252 112036 2256 112092
rect 2192 112032 2256 112036
rect 85952 112092 86016 112096
rect 85952 112036 85956 112092
rect 85956 112036 86012 112092
rect 86012 112036 86016 112092
rect 85952 112032 86016 112036
rect 86032 112092 86096 112096
rect 86032 112036 86036 112092
rect 86036 112036 86092 112092
rect 86092 112036 86096 112092
rect 86032 112032 86096 112036
rect 86112 112092 86176 112096
rect 86112 112036 86116 112092
rect 86116 112036 86172 112092
rect 86172 112036 86176 112092
rect 86112 112032 86176 112036
rect 86192 112092 86256 112096
rect 86192 112036 86196 112092
rect 86196 112036 86252 112092
rect 86252 112036 86256 112092
rect 86192 112032 86256 112036
rect 89952 112092 90016 112096
rect 89952 112036 89956 112092
rect 89956 112036 90012 112092
rect 90012 112036 90016 112092
rect 89952 112032 90016 112036
rect 90032 112092 90096 112096
rect 90032 112036 90036 112092
rect 90036 112036 90092 112092
rect 90092 112036 90096 112092
rect 90032 112032 90096 112036
rect 90112 112092 90176 112096
rect 90112 112036 90116 112092
rect 90116 112036 90172 112092
rect 90172 112036 90176 112092
rect 90112 112032 90176 112036
rect 90192 112092 90256 112096
rect 90192 112036 90196 112092
rect 90196 112036 90252 112092
rect 90252 112036 90256 112092
rect 90192 112032 90256 112036
rect 3952 111548 4016 111552
rect 3952 111492 3956 111548
rect 3956 111492 4012 111548
rect 4012 111492 4016 111548
rect 3952 111488 4016 111492
rect 4032 111548 4096 111552
rect 4032 111492 4036 111548
rect 4036 111492 4092 111548
rect 4092 111492 4096 111548
rect 4032 111488 4096 111492
rect 4112 111548 4176 111552
rect 4112 111492 4116 111548
rect 4116 111492 4172 111548
rect 4172 111492 4176 111548
rect 4112 111488 4176 111492
rect 4192 111548 4256 111552
rect 4192 111492 4196 111548
rect 4196 111492 4252 111548
rect 4252 111492 4256 111548
rect 4192 111488 4256 111492
rect 87952 111548 88016 111552
rect 87952 111492 87956 111548
rect 87956 111492 88012 111548
rect 88012 111492 88016 111548
rect 87952 111488 88016 111492
rect 88032 111548 88096 111552
rect 88032 111492 88036 111548
rect 88036 111492 88092 111548
rect 88092 111492 88096 111548
rect 88032 111488 88096 111492
rect 88112 111548 88176 111552
rect 88112 111492 88116 111548
rect 88116 111492 88172 111548
rect 88172 111492 88176 111548
rect 88112 111488 88176 111492
rect 88192 111548 88256 111552
rect 88192 111492 88196 111548
rect 88196 111492 88252 111548
rect 88252 111492 88256 111548
rect 88192 111488 88256 111492
rect 1952 111004 2016 111008
rect 1952 110948 1956 111004
rect 1956 110948 2012 111004
rect 2012 110948 2016 111004
rect 1952 110944 2016 110948
rect 2032 111004 2096 111008
rect 2032 110948 2036 111004
rect 2036 110948 2092 111004
rect 2092 110948 2096 111004
rect 2032 110944 2096 110948
rect 2112 111004 2176 111008
rect 2112 110948 2116 111004
rect 2116 110948 2172 111004
rect 2172 110948 2176 111004
rect 2112 110944 2176 110948
rect 2192 111004 2256 111008
rect 2192 110948 2196 111004
rect 2196 110948 2252 111004
rect 2252 110948 2256 111004
rect 2192 110944 2256 110948
rect 85952 111004 86016 111008
rect 85952 110948 85956 111004
rect 85956 110948 86012 111004
rect 86012 110948 86016 111004
rect 85952 110944 86016 110948
rect 86032 111004 86096 111008
rect 86032 110948 86036 111004
rect 86036 110948 86092 111004
rect 86092 110948 86096 111004
rect 86032 110944 86096 110948
rect 86112 111004 86176 111008
rect 86112 110948 86116 111004
rect 86116 110948 86172 111004
rect 86172 110948 86176 111004
rect 86112 110944 86176 110948
rect 86192 111004 86256 111008
rect 86192 110948 86196 111004
rect 86196 110948 86252 111004
rect 86252 110948 86256 111004
rect 86192 110944 86256 110948
rect 89952 111004 90016 111008
rect 89952 110948 89956 111004
rect 89956 110948 90012 111004
rect 90012 110948 90016 111004
rect 89952 110944 90016 110948
rect 90032 111004 90096 111008
rect 90032 110948 90036 111004
rect 90036 110948 90092 111004
rect 90092 110948 90096 111004
rect 90032 110944 90096 110948
rect 90112 111004 90176 111008
rect 90112 110948 90116 111004
rect 90116 110948 90172 111004
rect 90172 110948 90176 111004
rect 90112 110944 90176 110948
rect 90192 111004 90256 111008
rect 90192 110948 90196 111004
rect 90196 110948 90252 111004
rect 90252 110948 90256 111004
rect 90192 110944 90256 110948
rect 3952 110460 4016 110464
rect 3952 110404 3956 110460
rect 3956 110404 4012 110460
rect 4012 110404 4016 110460
rect 3952 110400 4016 110404
rect 4032 110460 4096 110464
rect 4032 110404 4036 110460
rect 4036 110404 4092 110460
rect 4092 110404 4096 110460
rect 4032 110400 4096 110404
rect 4112 110460 4176 110464
rect 4112 110404 4116 110460
rect 4116 110404 4172 110460
rect 4172 110404 4176 110460
rect 4112 110400 4176 110404
rect 4192 110460 4256 110464
rect 4192 110404 4196 110460
rect 4196 110404 4252 110460
rect 4252 110404 4256 110460
rect 4192 110400 4256 110404
rect 87952 110460 88016 110464
rect 87952 110404 87956 110460
rect 87956 110404 88012 110460
rect 88012 110404 88016 110460
rect 87952 110400 88016 110404
rect 88032 110460 88096 110464
rect 88032 110404 88036 110460
rect 88036 110404 88092 110460
rect 88092 110404 88096 110460
rect 88032 110400 88096 110404
rect 88112 110460 88176 110464
rect 88112 110404 88116 110460
rect 88116 110404 88172 110460
rect 88172 110404 88176 110460
rect 88112 110400 88176 110404
rect 88192 110460 88256 110464
rect 88192 110404 88196 110460
rect 88196 110404 88252 110460
rect 88252 110404 88256 110460
rect 88192 110400 88256 110404
rect 1952 109916 2016 109920
rect 1952 109860 1956 109916
rect 1956 109860 2012 109916
rect 2012 109860 2016 109916
rect 1952 109856 2016 109860
rect 2032 109916 2096 109920
rect 2032 109860 2036 109916
rect 2036 109860 2092 109916
rect 2092 109860 2096 109916
rect 2032 109856 2096 109860
rect 2112 109916 2176 109920
rect 2112 109860 2116 109916
rect 2116 109860 2172 109916
rect 2172 109860 2176 109916
rect 2112 109856 2176 109860
rect 2192 109916 2256 109920
rect 2192 109860 2196 109916
rect 2196 109860 2252 109916
rect 2252 109860 2256 109916
rect 2192 109856 2256 109860
rect 85952 109916 86016 109920
rect 85952 109860 85956 109916
rect 85956 109860 86012 109916
rect 86012 109860 86016 109916
rect 85952 109856 86016 109860
rect 86032 109916 86096 109920
rect 86032 109860 86036 109916
rect 86036 109860 86092 109916
rect 86092 109860 86096 109916
rect 86032 109856 86096 109860
rect 86112 109916 86176 109920
rect 86112 109860 86116 109916
rect 86116 109860 86172 109916
rect 86172 109860 86176 109916
rect 86112 109856 86176 109860
rect 86192 109916 86256 109920
rect 86192 109860 86196 109916
rect 86196 109860 86252 109916
rect 86252 109860 86256 109916
rect 86192 109856 86256 109860
rect 89952 109916 90016 109920
rect 89952 109860 89956 109916
rect 89956 109860 90012 109916
rect 90012 109860 90016 109916
rect 89952 109856 90016 109860
rect 90032 109916 90096 109920
rect 90032 109860 90036 109916
rect 90036 109860 90092 109916
rect 90092 109860 90096 109916
rect 90032 109856 90096 109860
rect 90112 109916 90176 109920
rect 90112 109860 90116 109916
rect 90116 109860 90172 109916
rect 90172 109860 90176 109916
rect 90112 109856 90176 109860
rect 90192 109916 90256 109920
rect 90192 109860 90196 109916
rect 90196 109860 90252 109916
rect 90252 109860 90256 109916
rect 90192 109856 90256 109860
rect 3952 109372 4016 109376
rect 3952 109316 3956 109372
rect 3956 109316 4012 109372
rect 4012 109316 4016 109372
rect 3952 109312 4016 109316
rect 4032 109372 4096 109376
rect 4032 109316 4036 109372
rect 4036 109316 4092 109372
rect 4092 109316 4096 109372
rect 4032 109312 4096 109316
rect 4112 109372 4176 109376
rect 4112 109316 4116 109372
rect 4116 109316 4172 109372
rect 4172 109316 4176 109372
rect 4112 109312 4176 109316
rect 4192 109372 4256 109376
rect 4192 109316 4196 109372
rect 4196 109316 4252 109372
rect 4252 109316 4256 109372
rect 4192 109312 4256 109316
rect 87952 109372 88016 109376
rect 87952 109316 87956 109372
rect 87956 109316 88012 109372
rect 88012 109316 88016 109372
rect 87952 109312 88016 109316
rect 88032 109372 88096 109376
rect 88032 109316 88036 109372
rect 88036 109316 88092 109372
rect 88092 109316 88096 109372
rect 88032 109312 88096 109316
rect 88112 109372 88176 109376
rect 88112 109316 88116 109372
rect 88116 109316 88172 109372
rect 88172 109316 88176 109372
rect 88112 109312 88176 109316
rect 88192 109372 88256 109376
rect 88192 109316 88196 109372
rect 88196 109316 88252 109372
rect 88252 109316 88256 109372
rect 88192 109312 88256 109316
rect 86908 109108 86972 109172
rect 1952 108828 2016 108832
rect 1952 108772 1956 108828
rect 1956 108772 2012 108828
rect 2012 108772 2016 108828
rect 1952 108768 2016 108772
rect 2032 108828 2096 108832
rect 2032 108772 2036 108828
rect 2036 108772 2092 108828
rect 2092 108772 2096 108828
rect 2032 108768 2096 108772
rect 2112 108828 2176 108832
rect 2112 108772 2116 108828
rect 2116 108772 2172 108828
rect 2172 108772 2176 108828
rect 2112 108768 2176 108772
rect 2192 108828 2256 108832
rect 2192 108772 2196 108828
rect 2196 108772 2252 108828
rect 2252 108772 2256 108828
rect 2192 108768 2256 108772
rect 85952 108828 86016 108832
rect 85952 108772 85956 108828
rect 85956 108772 86012 108828
rect 86012 108772 86016 108828
rect 85952 108768 86016 108772
rect 86032 108828 86096 108832
rect 86032 108772 86036 108828
rect 86036 108772 86092 108828
rect 86092 108772 86096 108828
rect 86032 108768 86096 108772
rect 86112 108828 86176 108832
rect 86112 108772 86116 108828
rect 86116 108772 86172 108828
rect 86172 108772 86176 108828
rect 86112 108768 86176 108772
rect 86192 108828 86256 108832
rect 86192 108772 86196 108828
rect 86196 108772 86252 108828
rect 86252 108772 86256 108828
rect 86192 108768 86256 108772
rect 89952 108828 90016 108832
rect 89952 108772 89956 108828
rect 89956 108772 90012 108828
rect 90012 108772 90016 108828
rect 89952 108768 90016 108772
rect 90032 108828 90096 108832
rect 90032 108772 90036 108828
rect 90036 108772 90092 108828
rect 90092 108772 90096 108828
rect 90032 108768 90096 108772
rect 90112 108828 90176 108832
rect 90112 108772 90116 108828
rect 90116 108772 90172 108828
rect 90172 108772 90176 108828
rect 90112 108768 90176 108772
rect 90192 108828 90256 108832
rect 90192 108772 90196 108828
rect 90196 108772 90252 108828
rect 90252 108772 90256 108828
rect 90192 108768 90256 108772
rect 86908 108700 86972 108764
rect 85620 108564 85684 108628
rect 3952 108284 4016 108288
rect 3952 108228 3956 108284
rect 3956 108228 4012 108284
rect 4012 108228 4016 108284
rect 3952 108224 4016 108228
rect 4032 108284 4096 108288
rect 4032 108228 4036 108284
rect 4036 108228 4092 108284
rect 4092 108228 4096 108284
rect 4032 108224 4096 108228
rect 4112 108284 4176 108288
rect 4112 108228 4116 108284
rect 4116 108228 4172 108284
rect 4172 108228 4176 108284
rect 4112 108224 4176 108228
rect 4192 108284 4256 108288
rect 4192 108228 4196 108284
rect 4196 108228 4252 108284
rect 4252 108228 4256 108284
rect 4192 108224 4256 108228
rect 87952 108284 88016 108288
rect 87952 108228 87956 108284
rect 87956 108228 88012 108284
rect 88012 108228 88016 108284
rect 87952 108224 88016 108228
rect 88032 108284 88096 108288
rect 88032 108228 88036 108284
rect 88036 108228 88092 108284
rect 88092 108228 88096 108284
rect 88032 108224 88096 108228
rect 88112 108284 88176 108288
rect 88112 108228 88116 108284
rect 88116 108228 88172 108284
rect 88172 108228 88176 108284
rect 88112 108224 88176 108228
rect 88192 108284 88256 108288
rect 88192 108228 88196 108284
rect 88196 108228 88252 108284
rect 88252 108228 88256 108284
rect 88192 108224 88256 108228
rect 1952 107740 2016 107744
rect 1952 107684 1956 107740
rect 1956 107684 2012 107740
rect 2012 107684 2016 107740
rect 1952 107680 2016 107684
rect 2032 107740 2096 107744
rect 2032 107684 2036 107740
rect 2036 107684 2092 107740
rect 2092 107684 2096 107740
rect 2032 107680 2096 107684
rect 2112 107740 2176 107744
rect 2112 107684 2116 107740
rect 2116 107684 2172 107740
rect 2172 107684 2176 107740
rect 2112 107680 2176 107684
rect 2192 107740 2256 107744
rect 2192 107684 2196 107740
rect 2196 107684 2252 107740
rect 2252 107684 2256 107740
rect 2192 107680 2256 107684
rect 85952 107740 86016 107744
rect 85952 107684 85956 107740
rect 85956 107684 86012 107740
rect 86012 107684 86016 107740
rect 85952 107680 86016 107684
rect 86032 107740 86096 107744
rect 86032 107684 86036 107740
rect 86036 107684 86092 107740
rect 86092 107684 86096 107740
rect 86032 107680 86096 107684
rect 86112 107740 86176 107744
rect 86112 107684 86116 107740
rect 86116 107684 86172 107740
rect 86172 107684 86176 107740
rect 86112 107680 86176 107684
rect 86192 107740 86256 107744
rect 86192 107684 86196 107740
rect 86196 107684 86252 107740
rect 86252 107684 86256 107740
rect 86192 107680 86256 107684
rect 89952 107740 90016 107744
rect 89952 107684 89956 107740
rect 89956 107684 90012 107740
rect 90012 107684 90016 107740
rect 89952 107680 90016 107684
rect 90032 107740 90096 107744
rect 90032 107684 90036 107740
rect 90036 107684 90092 107740
rect 90092 107684 90096 107740
rect 90032 107680 90096 107684
rect 90112 107740 90176 107744
rect 90112 107684 90116 107740
rect 90116 107684 90172 107740
rect 90172 107684 90176 107740
rect 90112 107680 90176 107684
rect 90192 107740 90256 107744
rect 90192 107684 90196 107740
rect 90196 107684 90252 107740
rect 90252 107684 90256 107740
rect 90192 107680 90256 107684
rect 3952 107196 4016 107200
rect 3952 107140 3956 107196
rect 3956 107140 4012 107196
rect 4012 107140 4016 107196
rect 3952 107136 4016 107140
rect 4032 107196 4096 107200
rect 4032 107140 4036 107196
rect 4036 107140 4092 107196
rect 4092 107140 4096 107196
rect 4032 107136 4096 107140
rect 4112 107196 4176 107200
rect 4112 107140 4116 107196
rect 4116 107140 4172 107196
rect 4172 107140 4176 107196
rect 4112 107136 4176 107140
rect 4192 107196 4256 107200
rect 4192 107140 4196 107196
rect 4196 107140 4252 107196
rect 4252 107140 4256 107196
rect 4192 107136 4256 107140
rect 87952 107196 88016 107200
rect 87952 107140 87956 107196
rect 87956 107140 88012 107196
rect 88012 107140 88016 107196
rect 87952 107136 88016 107140
rect 88032 107196 88096 107200
rect 88032 107140 88036 107196
rect 88036 107140 88092 107196
rect 88092 107140 88096 107196
rect 88032 107136 88096 107140
rect 88112 107196 88176 107200
rect 88112 107140 88116 107196
rect 88116 107140 88172 107196
rect 88172 107140 88176 107196
rect 88112 107136 88176 107140
rect 88192 107196 88256 107200
rect 88192 107140 88196 107196
rect 88196 107140 88252 107196
rect 88252 107140 88256 107196
rect 88192 107136 88256 107140
rect 1952 106652 2016 106656
rect 1952 106596 1956 106652
rect 1956 106596 2012 106652
rect 2012 106596 2016 106652
rect 1952 106592 2016 106596
rect 2032 106652 2096 106656
rect 2032 106596 2036 106652
rect 2036 106596 2092 106652
rect 2092 106596 2096 106652
rect 2032 106592 2096 106596
rect 2112 106652 2176 106656
rect 2112 106596 2116 106652
rect 2116 106596 2172 106652
rect 2172 106596 2176 106652
rect 2112 106592 2176 106596
rect 2192 106652 2256 106656
rect 2192 106596 2196 106652
rect 2196 106596 2252 106652
rect 2252 106596 2256 106652
rect 2192 106592 2256 106596
rect 85952 106652 86016 106656
rect 85952 106596 85956 106652
rect 85956 106596 86012 106652
rect 86012 106596 86016 106652
rect 85952 106592 86016 106596
rect 86032 106652 86096 106656
rect 86032 106596 86036 106652
rect 86036 106596 86092 106652
rect 86092 106596 86096 106652
rect 86032 106592 86096 106596
rect 86112 106652 86176 106656
rect 86112 106596 86116 106652
rect 86116 106596 86172 106652
rect 86172 106596 86176 106652
rect 86112 106592 86176 106596
rect 86192 106652 86256 106656
rect 86192 106596 86196 106652
rect 86196 106596 86252 106652
rect 86252 106596 86256 106652
rect 86192 106592 86256 106596
rect 89952 106652 90016 106656
rect 89952 106596 89956 106652
rect 89956 106596 90012 106652
rect 90012 106596 90016 106652
rect 89952 106592 90016 106596
rect 90032 106652 90096 106656
rect 90032 106596 90036 106652
rect 90036 106596 90092 106652
rect 90092 106596 90096 106652
rect 90032 106592 90096 106596
rect 90112 106652 90176 106656
rect 90112 106596 90116 106652
rect 90116 106596 90172 106652
rect 90172 106596 90176 106652
rect 90112 106592 90176 106596
rect 90192 106652 90256 106656
rect 90192 106596 90196 106652
rect 90196 106596 90252 106652
rect 90252 106596 90256 106652
rect 90192 106592 90256 106596
rect 3952 106108 4016 106112
rect 3952 106052 3956 106108
rect 3956 106052 4012 106108
rect 4012 106052 4016 106108
rect 3952 106048 4016 106052
rect 4032 106108 4096 106112
rect 4032 106052 4036 106108
rect 4036 106052 4092 106108
rect 4092 106052 4096 106108
rect 4032 106048 4096 106052
rect 4112 106108 4176 106112
rect 4112 106052 4116 106108
rect 4116 106052 4172 106108
rect 4172 106052 4176 106108
rect 4112 106048 4176 106052
rect 4192 106108 4256 106112
rect 4192 106052 4196 106108
rect 4196 106052 4252 106108
rect 4252 106052 4256 106108
rect 4192 106048 4256 106052
rect 87952 106108 88016 106112
rect 87952 106052 87956 106108
rect 87956 106052 88012 106108
rect 88012 106052 88016 106108
rect 87952 106048 88016 106052
rect 88032 106108 88096 106112
rect 88032 106052 88036 106108
rect 88036 106052 88092 106108
rect 88092 106052 88096 106108
rect 88032 106048 88096 106052
rect 88112 106108 88176 106112
rect 88112 106052 88116 106108
rect 88116 106052 88172 106108
rect 88172 106052 88176 106108
rect 88112 106048 88176 106052
rect 88192 106108 88256 106112
rect 88192 106052 88196 106108
rect 88196 106052 88252 106108
rect 88252 106052 88256 106108
rect 88192 106048 88256 106052
rect 1952 105564 2016 105568
rect 1952 105508 1956 105564
rect 1956 105508 2012 105564
rect 2012 105508 2016 105564
rect 1952 105504 2016 105508
rect 2032 105564 2096 105568
rect 2032 105508 2036 105564
rect 2036 105508 2092 105564
rect 2092 105508 2096 105564
rect 2032 105504 2096 105508
rect 2112 105564 2176 105568
rect 2112 105508 2116 105564
rect 2116 105508 2172 105564
rect 2172 105508 2176 105564
rect 2112 105504 2176 105508
rect 2192 105564 2256 105568
rect 2192 105508 2196 105564
rect 2196 105508 2252 105564
rect 2252 105508 2256 105564
rect 2192 105504 2256 105508
rect 85952 105564 86016 105568
rect 85952 105508 85956 105564
rect 85956 105508 86012 105564
rect 86012 105508 86016 105564
rect 85952 105504 86016 105508
rect 86032 105564 86096 105568
rect 86032 105508 86036 105564
rect 86036 105508 86092 105564
rect 86092 105508 86096 105564
rect 86032 105504 86096 105508
rect 86112 105564 86176 105568
rect 86112 105508 86116 105564
rect 86116 105508 86172 105564
rect 86172 105508 86176 105564
rect 86112 105504 86176 105508
rect 86192 105564 86256 105568
rect 86192 105508 86196 105564
rect 86196 105508 86252 105564
rect 86252 105508 86256 105564
rect 86192 105504 86256 105508
rect 89952 105564 90016 105568
rect 89952 105508 89956 105564
rect 89956 105508 90012 105564
rect 90012 105508 90016 105564
rect 89952 105504 90016 105508
rect 90032 105564 90096 105568
rect 90032 105508 90036 105564
rect 90036 105508 90092 105564
rect 90092 105508 90096 105564
rect 90032 105504 90096 105508
rect 90112 105564 90176 105568
rect 90112 105508 90116 105564
rect 90116 105508 90172 105564
rect 90172 105508 90176 105564
rect 90112 105504 90176 105508
rect 90192 105564 90256 105568
rect 90192 105508 90196 105564
rect 90196 105508 90252 105564
rect 90252 105508 90256 105564
rect 90192 105504 90256 105508
rect 3952 105020 4016 105024
rect 3952 104964 3956 105020
rect 3956 104964 4012 105020
rect 4012 104964 4016 105020
rect 3952 104960 4016 104964
rect 4032 105020 4096 105024
rect 4032 104964 4036 105020
rect 4036 104964 4092 105020
rect 4092 104964 4096 105020
rect 4032 104960 4096 104964
rect 4112 105020 4176 105024
rect 4112 104964 4116 105020
rect 4116 104964 4172 105020
rect 4172 104964 4176 105020
rect 4112 104960 4176 104964
rect 4192 105020 4256 105024
rect 4192 104964 4196 105020
rect 4196 104964 4252 105020
rect 4252 104964 4256 105020
rect 4192 104960 4256 104964
rect 87952 105020 88016 105024
rect 87952 104964 87956 105020
rect 87956 104964 88012 105020
rect 88012 104964 88016 105020
rect 87952 104960 88016 104964
rect 88032 105020 88096 105024
rect 88032 104964 88036 105020
rect 88036 104964 88092 105020
rect 88092 104964 88096 105020
rect 88032 104960 88096 104964
rect 88112 105020 88176 105024
rect 88112 104964 88116 105020
rect 88116 104964 88172 105020
rect 88172 104964 88176 105020
rect 88112 104960 88176 104964
rect 88192 105020 88256 105024
rect 88192 104964 88196 105020
rect 88196 104964 88252 105020
rect 88252 104964 88256 105020
rect 88192 104960 88256 104964
rect 1952 104476 2016 104480
rect 1952 104420 1956 104476
rect 1956 104420 2012 104476
rect 2012 104420 2016 104476
rect 1952 104416 2016 104420
rect 2032 104476 2096 104480
rect 2032 104420 2036 104476
rect 2036 104420 2092 104476
rect 2092 104420 2096 104476
rect 2032 104416 2096 104420
rect 2112 104476 2176 104480
rect 2112 104420 2116 104476
rect 2116 104420 2172 104476
rect 2172 104420 2176 104476
rect 2112 104416 2176 104420
rect 2192 104476 2256 104480
rect 2192 104420 2196 104476
rect 2196 104420 2252 104476
rect 2252 104420 2256 104476
rect 2192 104416 2256 104420
rect 85952 104476 86016 104480
rect 85952 104420 85956 104476
rect 85956 104420 86012 104476
rect 86012 104420 86016 104476
rect 85952 104416 86016 104420
rect 86032 104476 86096 104480
rect 86032 104420 86036 104476
rect 86036 104420 86092 104476
rect 86092 104420 86096 104476
rect 86032 104416 86096 104420
rect 86112 104476 86176 104480
rect 86112 104420 86116 104476
rect 86116 104420 86172 104476
rect 86172 104420 86176 104476
rect 86112 104416 86176 104420
rect 86192 104476 86256 104480
rect 86192 104420 86196 104476
rect 86196 104420 86252 104476
rect 86252 104420 86256 104476
rect 86192 104416 86256 104420
rect 89952 104476 90016 104480
rect 89952 104420 89956 104476
rect 89956 104420 90012 104476
rect 90012 104420 90016 104476
rect 89952 104416 90016 104420
rect 90032 104476 90096 104480
rect 90032 104420 90036 104476
rect 90036 104420 90092 104476
rect 90092 104420 90096 104476
rect 90032 104416 90096 104420
rect 90112 104476 90176 104480
rect 90112 104420 90116 104476
rect 90116 104420 90172 104476
rect 90172 104420 90176 104476
rect 90112 104416 90176 104420
rect 90192 104476 90256 104480
rect 90192 104420 90196 104476
rect 90196 104420 90252 104476
rect 90252 104420 90256 104476
rect 90192 104416 90256 104420
rect 3952 103932 4016 103936
rect 3952 103876 3956 103932
rect 3956 103876 4012 103932
rect 4012 103876 4016 103932
rect 3952 103872 4016 103876
rect 4032 103932 4096 103936
rect 4032 103876 4036 103932
rect 4036 103876 4092 103932
rect 4092 103876 4096 103932
rect 4032 103872 4096 103876
rect 4112 103932 4176 103936
rect 4112 103876 4116 103932
rect 4116 103876 4172 103932
rect 4172 103876 4176 103932
rect 4112 103872 4176 103876
rect 4192 103932 4256 103936
rect 4192 103876 4196 103932
rect 4196 103876 4252 103932
rect 4252 103876 4256 103932
rect 4192 103872 4256 103876
rect 87952 103932 88016 103936
rect 87952 103876 87956 103932
rect 87956 103876 88012 103932
rect 88012 103876 88016 103932
rect 87952 103872 88016 103876
rect 88032 103932 88096 103936
rect 88032 103876 88036 103932
rect 88036 103876 88092 103932
rect 88092 103876 88096 103932
rect 88032 103872 88096 103876
rect 88112 103932 88176 103936
rect 88112 103876 88116 103932
rect 88116 103876 88172 103932
rect 88172 103876 88176 103932
rect 88112 103872 88176 103876
rect 88192 103932 88256 103936
rect 88192 103876 88196 103932
rect 88196 103876 88252 103932
rect 88252 103876 88256 103932
rect 88192 103872 88256 103876
rect 86724 103668 86788 103732
rect 1952 103388 2016 103392
rect 1952 103332 1956 103388
rect 1956 103332 2012 103388
rect 2012 103332 2016 103388
rect 1952 103328 2016 103332
rect 2032 103388 2096 103392
rect 2032 103332 2036 103388
rect 2036 103332 2092 103388
rect 2092 103332 2096 103388
rect 2032 103328 2096 103332
rect 2112 103388 2176 103392
rect 2112 103332 2116 103388
rect 2116 103332 2172 103388
rect 2172 103332 2176 103388
rect 2112 103328 2176 103332
rect 2192 103388 2256 103392
rect 2192 103332 2196 103388
rect 2196 103332 2252 103388
rect 2252 103332 2256 103388
rect 2192 103328 2256 103332
rect 85952 103388 86016 103392
rect 85952 103332 85956 103388
rect 85956 103332 86012 103388
rect 86012 103332 86016 103388
rect 85952 103328 86016 103332
rect 86032 103388 86096 103392
rect 86032 103332 86036 103388
rect 86036 103332 86092 103388
rect 86092 103332 86096 103388
rect 86032 103328 86096 103332
rect 86112 103388 86176 103392
rect 86112 103332 86116 103388
rect 86116 103332 86172 103388
rect 86172 103332 86176 103388
rect 86112 103328 86176 103332
rect 86192 103388 86256 103392
rect 86192 103332 86196 103388
rect 86196 103332 86252 103388
rect 86252 103332 86256 103388
rect 86192 103328 86256 103332
rect 89952 103388 90016 103392
rect 89952 103332 89956 103388
rect 89956 103332 90012 103388
rect 90012 103332 90016 103388
rect 89952 103328 90016 103332
rect 90032 103388 90096 103392
rect 90032 103332 90036 103388
rect 90036 103332 90092 103388
rect 90092 103332 90096 103388
rect 90032 103328 90096 103332
rect 90112 103388 90176 103392
rect 90112 103332 90116 103388
rect 90116 103332 90172 103388
rect 90172 103332 90176 103388
rect 90112 103328 90176 103332
rect 90192 103388 90256 103392
rect 90192 103332 90196 103388
rect 90196 103332 90252 103388
rect 90252 103332 90256 103388
rect 90192 103328 90256 103332
rect 3952 102844 4016 102848
rect 3952 102788 3956 102844
rect 3956 102788 4012 102844
rect 4012 102788 4016 102844
rect 3952 102784 4016 102788
rect 4032 102844 4096 102848
rect 4032 102788 4036 102844
rect 4036 102788 4092 102844
rect 4092 102788 4096 102844
rect 4032 102784 4096 102788
rect 4112 102844 4176 102848
rect 4112 102788 4116 102844
rect 4116 102788 4172 102844
rect 4172 102788 4176 102844
rect 4112 102784 4176 102788
rect 4192 102844 4256 102848
rect 4192 102788 4196 102844
rect 4196 102788 4252 102844
rect 4252 102788 4256 102844
rect 4192 102784 4256 102788
rect 87952 102844 88016 102848
rect 87952 102788 87956 102844
rect 87956 102788 88012 102844
rect 88012 102788 88016 102844
rect 87952 102784 88016 102788
rect 88032 102844 88096 102848
rect 88032 102788 88036 102844
rect 88036 102788 88092 102844
rect 88092 102788 88096 102844
rect 88032 102784 88096 102788
rect 88112 102844 88176 102848
rect 88112 102788 88116 102844
rect 88116 102788 88172 102844
rect 88172 102788 88176 102844
rect 88112 102784 88176 102788
rect 88192 102844 88256 102848
rect 88192 102788 88196 102844
rect 88196 102788 88252 102844
rect 88252 102788 88256 102844
rect 88192 102784 88256 102788
rect 86908 102580 86972 102644
rect 1952 102300 2016 102304
rect 1952 102244 1956 102300
rect 1956 102244 2012 102300
rect 2012 102244 2016 102300
rect 1952 102240 2016 102244
rect 2032 102300 2096 102304
rect 2032 102244 2036 102300
rect 2036 102244 2092 102300
rect 2092 102244 2096 102300
rect 2032 102240 2096 102244
rect 2112 102300 2176 102304
rect 2112 102244 2116 102300
rect 2116 102244 2172 102300
rect 2172 102244 2176 102300
rect 2112 102240 2176 102244
rect 2192 102300 2256 102304
rect 2192 102244 2196 102300
rect 2196 102244 2252 102300
rect 2252 102244 2256 102300
rect 2192 102240 2256 102244
rect 85952 102300 86016 102304
rect 85952 102244 85956 102300
rect 85956 102244 86012 102300
rect 86012 102244 86016 102300
rect 85952 102240 86016 102244
rect 86032 102300 86096 102304
rect 86032 102244 86036 102300
rect 86036 102244 86092 102300
rect 86092 102244 86096 102300
rect 86032 102240 86096 102244
rect 86112 102300 86176 102304
rect 86112 102244 86116 102300
rect 86116 102244 86172 102300
rect 86172 102244 86176 102300
rect 86112 102240 86176 102244
rect 86192 102300 86256 102304
rect 86192 102244 86196 102300
rect 86196 102244 86252 102300
rect 86252 102244 86256 102300
rect 86192 102240 86256 102244
rect 89952 102300 90016 102304
rect 89952 102244 89956 102300
rect 89956 102244 90012 102300
rect 90012 102244 90016 102300
rect 89952 102240 90016 102244
rect 90032 102300 90096 102304
rect 90032 102244 90036 102300
rect 90036 102244 90092 102300
rect 90092 102244 90096 102300
rect 90032 102240 90096 102244
rect 90112 102300 90176 102304
rect 90112 102244 90116 102300
rect 90116 102244 90172 102300
rect 90172 102244 90176 102300
rect 90112 102240 90176 102244
rect 90192 102300 90256 102304
rect 90192 102244 90196 102300
rect 90196 102244 90252 102300
rect 90252 102244 90256 102300
rect 90192 102240 90256 102244
rect 3952 101756 4016 101760
rect 3952 101700 3956 101756
rect 3956 101700 4012 101756
rect 4012 101700 4016 101756
rect 3952 101696 4016 101700
rect 4032 101756 4096 101760
rect 4032 101700 4036 101756
rect 4036 101700 4092 101756
rect 4092 101700 4096 101756
rect 4032 101696 4096 101700
rect 4112 101756 4176 101760
rect 4112 101700 4116 101756
rect 4116 101700 4172 101756
rect 4172 101700 4176 101756
rect 4112 101696 4176 101700
rect 4192 101756 4256 101760
rect 4192 101700 4196 101756
rect 4196 101700 4252 101756
rect 4252 101700 4256 101756
rect 4192 101696 4256 101700
rect 87952 101756 88016 101760
rect 87952 101700 87956 101756
rect 87956 101700 88012 101756
rect 88012 101700 88016 101756
rect 87952 101696 88016 101700
rect 88032 101756 88096 101760
rect 88032 101700 88036 101756
rect 88036 101700 88092 101756
rect 88092 101700 88096 101756
rect 88032 101696 88096 101700
rect 88112 101756 88176 101760
rect 88112 101700 88116 101756
rect 88116 101700 88172 101756
rect 88172 101700 88176 101756
rect 88112 101696 88176 101700
rect 88192 101756 88256 101760
rect 88192 101700 88196 101756
rect 88196 101700 88252 101756
rect 88252 101700 88256 101756
rect 88192 101696 88256 101700
rect 1952 101212 2016 101216
rect 1952 101156 1956 101212
rect 1956 101156 2012 101212
rect 2012 101156 2016 101212
rect 1952 101152 2016 101156
rect 2032 101212 2096 101216
rect 2032 101156 2036 101212
rect 2036 101156 2092 101212
rect 2092 101156 2096 101212
rect 2032 101152 2096 101156
rect 2112 101212 2176 101216
rect 2112 101156 2116 101212
rect 2116 101156 2172 101212
rect 2172 101156 2176 101212
rect 2112 101152 2176 101156
rect 2192 101212 2256 101216
rect 2192 101156 2196 101212
rect 2196 101156 2252 101212
rect 2252 101156 2256 101212
rect 2192 101152 2256 101156
rect 85952 101212 86016 101216
rect 85952 101156 85956 101212
rect 85956 101156 86012 101212
rect 86012 101156 86016 101212
rect 85952 101152 86016 101156
rect 86032 101212 86096 101216
rect 86032 101156 86036 101212
rect 86036 101156 86092 101212
rect 86092 101156 86096 101212
rect 86032 101152 86096 101156
rect 86112 101212 86176 101216
rect 86112 101156 86116 101212
rect 86116 101156 86172 101212
rect 86172 101156 86176 101212
rect 86112 101152 86176 101156
rect 86192 101212 86256 101216
rect 86192 101156 86196 101212
rect 86196 101156 86252 101212
rect 86252 101156 86256 101212
rect 86192 101152 86256 101156
rect 89952 101212 90016 101216
rect 89952 101156 89956 101212
rect 89956 101156 90012 101212
rect 90012 101156 90016 101212
rect 89952 101152 90016 101156
rect 90032 101212 90096 101216
rect 90032 101156 90036 101212
rect 90036 101156 90092 101212
rect 90092 101156 90096 101212
rect 90032 101152 90096 101156
rect 90112 101212 90176 101216
rect 90112 101156 90116 101212
rect 90116 101156 90172 101212
rect 90172 101156 90176 101212
rect 90112 101152 90176 101156
rect 90192 101212 90256 101216
rect 90192 101156 90196 101212
rect 90196 101156 90252 101212
rect 90252 101156 90256 101212
rect 90192 101152 90256 101156
rect 3952 100668 4016 100672
rect 3952 100612 3956 100668
rect 3956 100612 4012 100668
rect 4012 100612 4016 100668
rect 3952 100608 4016 100612
rect 4032 100668 4096 100672
rect 4032 100612 4036 100668
rect 4036 100612 4092 100668
rect 4092 100612 4096 100668
rect 4032 100608 4096 100612
rect 4112 100668 4176 100672
rect 4112 100612 4116 100668
rect 4116 100612 4172 100668
rect 4172 100612 4176 100668
rect 4112 100608 4176 100612
rect 4192 100668 4256 100672
rect 4192 100612 4196 100668
rect 4196 100612 4252 100668
rect 4252 100612 4256 100668
rect 4192 100608 4256 100612
rect 87952 100668 88016 100672
rect 87952 100612 87956 100668
rect 87956 100612 88012 100668
rect 88012 100612 88016 100668
rect 87952 100608 88016 100612
rect 88032 100668 88096 100672
rect 88032 100612 88036 100668
rect 88036 100612 88092 100668
rect 88092 100612 88096 100668
rect 88032 100608 88096 100612
rect 88112 100668 88176 100672
rect 88112 100612 88116 100668
rect 88116 100612 88172 100668
rect 88172 100612 88176 100668
rect 88112 100608 88176 100612
rect 88192 100668 88256 100672
rect 88192 100612 88196 100668
rect 88196 100612 88252 100668
rect 88252 100612 88256 100668
rect 88192 100608 88256 100612
rect 1952 100124 2016 100128
rect 1952 100068 1956 100124
rect 1956 100068 2012 100124
rect 2012 100068 2016 100124
rect 1952 100064 2016 100068
rect 2032 100124 2096 100128
rect 2032 100068 2036 100124
rect 2036 100068 2092 100124
rect 2092 100068 2096 100124
rect 2032 100064 2096 100068
rect 2112 100124 2176 100128
rect 2112 100068 2116 100124
rect 2116 100068 2172 100124
rect 2172 100068 2176 100124
rect 2112 100064 2176 100068
rect 2192 100124 2256 100128
rect 2192 100068 2196 100124
rect 2196 100068 2252 100124
rect 2252 100068 2256 100124
rect 2192 100064 2256 100068
rect 85952 100124 86016 100128
rect 85952 100068 85956 100124
rect 85956 100068 86012 100124
rect 86012 100068 86016 100124
rect 85952 100064 86016 100068
rect 86032 100124 86096 100128
rect 86032 100068 86036 100124
rect 86036 100068 86092 100124
rect 86092 100068 86096 100124
rect 86032 100064 86096 100068
rect 86112 100124 86176 100128
rect 86112 100068 86116 100124
rect 86116 100068 86172 100124
rect 86172 100068 86176 100124
rect 86112 100064 86176 100068
rect 86192 100124 86256 100128
rect 86192 100068 86196 100124
rect 86196 100068 86252 100124
rect 86252 100068 86256 100124
rect 86192 100064 86256 100068
rect 89952 100124 90016 100128
rect 89952 100068 89956 100124
rect 89956 100068 90012 100124
rect 90012 100068 90016 100124
rect 89952 100064 90016 100068
rect 90032 100124 90096 100128
rect 90032 100068 90036 100124
rect 90036 100068 90092 100124
rect 90092 100068 90096 100124
rect 90032 100064 90096 100068
rect 90112 100124 90176 100128
rect 90112 100068 90116 100124
rect 90116 100068 90172 100124
rect 90172 100068 90176 100124
rect 90112 100064 90176 100068
rect 90192 100124 90256 100128
rect 90192 100068 90196 100124
rect 90196 100068 90252 100124
rect 90252 100068 90256 100124
rect 90192 100064 90256 100068
rect 3952 99580 4016 99584
rect 3952 99524 3956 99580
rect 3956 99524 4012 99580
rect 4012 99524 4016 99580
rect 3952 99520 4016 99524
rect 4032 99580 4096 99584
rect 4032 99524 4036 99580
rect 4036 99524 4092 99580
rect 4092 99524 4096 99580
rect 4032 99520 4096 99524
rect 4112 99580 4176 99584
rect 4112 99524 4116 99580
rect 4116 99524 4172 99580
rect 4172 99524 4176 99580
rect 4112 99520 4176 99524
rect 4192 99580 4256 99584
rect 4192 99524 4196 99580
rect 4196 99524 4252 99580
rect 4252 99524 4256 99580
rect 4192 99520 4256 99524
rect 84516 99452 84580 99516
rect 85436 99452 85500 99516
rect 86908 99452 86972 99516
rect 87952 99580 88016 99584
rect 87952 99524 87956 99580
rect 87956 99524 88012 99580
rect 88012 99524 88016 99580
rect 87952 99520 88016 99524
rect 88032 99580 88096 99584
rect 88032 99524 88036 99580
rect 88036 99524 88092 99580
rect 88092 99524 88096 99580
rect 88032 99520 88096 99524
rect 88112 99580 88176 99584
rect 88112 99524 88116 99580
rect 88116 99524 88172 99580
rect 88172 99524 88176 99580
rect 88112 99520 88176 99524
rect 88192 99580 88256 99584
rect 88192 99524 88196 99580
rect 88196 99524 88252 99580
rect 88252 99524 88256 99580
rect 88192 99520 88256 99524
rect 84516 99316 84580 99380
rect 86724 99316 86788 99380
rect 85436 99104 85500 99108
rect 85436 99048 85450 99104
rect 85450 99048 85500 99104
rect 85436 99044 85500 99048
rect 1952 99036 2016 99040
rect 1952 98980 1956 99036
rect 1956 98980 2012 99036
rect 2012 98980 2016 99036
rect 1952 98976 2016 98980
rect 2032 99036 2096 99040
rect 2032 98980 2036 99036
rect 2036 98980 2092 99036
rect 2092 98980 2096 99036
rect 2032 98976 2096 98980
rect 2112 99036 2176 99040
rect 2112 98980 2116 99036
rect 2116 98980 2172 99036
rect 2172 98980 2176 99036
rect 2112 98976 2176 98980
rect 2192 99036 2256 99040
rect 2192 98980 2196 99036
rect 2196 98980 2252 99036
rect 2252 98980 2256 99036
rect 2192 98976 2256 98980
rect 85952 99036 86016 99040
rect 85952 98980 85956 99036
rect 85956 98980 86012 99036
rect 86012 98980 86016 99036
rect 85952 98976 86016 98980
rect 86032 99036 86096 99040
rect 86032 98980 86036 99036
rect 86036 98980 86092 99036
rect 86092 98980 86096 99036
rect 86032 98976 86096 98980
rect 86112 99036 86176 99040
rect 86112 98980 86116 99036
rect 86116 98980 86172 99036
rect 86172 98980 86176 99036
rect 86112 98976 86176 98980
rect 86192 99036 86256 99040
rect 86192 98980 86196 99036
rect 86196 98980 86252 99036
rect 86252 98980 86256 99036
rect 86192 98976 86256 98980
rect 89952 99036 90016 99040
rect 89952 98980 89956 99036
rect 89956 98980 90012 99036
rect 90012 98980 90016 99036
rect 89952 98976 90016 98980
rect 90032 99036 90096 99040
rect 90032 98980 90036 99036
rect 90036 98980 90092 99036
rect 90092 98980 90096 99036
rect 90032 98976 90096 98980
rect 90112 99036 90176 99040
rect 90112 98980 90116 99036
rect 90116 98980 90172 99036
rect 90172 98980 90176 99036
rect 90112 98976 90176 98980
rect 90192 99036 90256 99040
rect 90192 98980 90196 99036
rect 90196 98980 90252 99036
rect 90252 98980 90256 99036
rect 90192 98976 90256 98980
rect 3952 98492 4016 98496
rect 3952 98436 3956 98492
rect 3956 98436 4012 98492
rect 4012 98436 4016 98492
rect 3952 98432 4016 98436
rect 4032 98492 4096 98496
rect 4032 98436 4036 98492
rect 4036 98436 4092 98492
rect 4092 98436 4096 98492
rect 4032 98432 4096 98436
rect 4112 98492 4176 98496
rect 4112 98436 4116 98492
rect 4116 98436 4172 98492
rect 4172 98436 4176 98492
rect 4112 98432 4176 98436
rect 4192 98492 4256 98496
rect 4192 98436 4196 98492
rect 4196 98436 4252 98492
rect 4252 98436 4256 98492
rect 4192 98432 4256 98436
rect 87952 98492 88016 98496
rect 87952 98436 87956 98492
rect 87956 98436 88012 98492
rect 88012 98436 88016 98492
rect 87952 98432 88016 98436
rect 88032 98492 88096 98496
rect 88032 98436 88036 98492
rect 88036 98436 88092 98492
rect 88092 98436 88096 98492
rect 88032 98432 88096 98436
rect 88112 98492 88176 98496
rect 88112 98436 88116 98492
rect 88116 98436 88172 98492
rect 88172 98436 88176 98492
rect 88112 98432 88176 98436
rect 88192 98492 88256 98496
rect 88192 98436 88196 98492
rect 88196 98436 88252 98492
rect 88252 98436 88256 98492
rect 88192 98432 88256 98436
rect 89116 98092 89180 98156
rect 90588 98092 90652 98156
rect 1952 97948 2016 97952
rect 1952 97892 1956 97948
rect 1956 97892 2012 97948
rect 2012 97892 2016 97948
rect 1952 97888 2016 97892
rect 2032 97948 2096 97952
rect 2032 97892 2036 97948
rect 2036 97892 2092 97948
rect 2092 97892 2096 97948
rect 2032 97888 2096 97892
rect 2112 97948 2176 97952
rect 2112 97892 2116 97948
rect 2116 97892 2172 97948
rect 2172 97892 2176 97948
rect 2112 97888 2176 97892
rect 2192 97948 2256 97952
rect 2192 97892 2196 97948
rect 2196 97892 2252 97948
rect 2252 97892 2256 97948
rect 2192 97888 2256 97892
rect 85952 97948 86016 97952
rect 85952 97892 85956 97948
rect 85956 97892 86012 97948
rect 86012 97892 86016 97948
rect 85952 97888 86016 97892
rect 86032 97948 86096 97952
rect 86032 97892 86036 97948
rect 86036 97892 86092 97948
rect 86092 97892 86096 97948
rect 86032 97888 86096 97892
rect 86112 97948 86176 97952
rect 86112 97892 86116 97948
rect 86116 97892 86172 97948
rect 86172 97892 86176 97948
rect 86112 97888 86176 97892
rect 86192 97948 86256 97952
rect 86192 97892 86196 97948
rect 86196 97892 86252 97948
rect 86252 97892 86256 97948
rect 86192 97888 86256 97892
rect 89952 97948 90016 97952
rect 89952 97892 89956 97948
rect 89956 97892 90012 97948
rect 90012 97892 90016 97948
rect 89952 97888 90016 97892
rect 90032 97948 90096 97952
rect 90032 97892 90036 97948
rect 90036 97892 90092 97948
rect 90092 97892 90096 97948
rect 90032 97888 90096 97892
rect 90112 97948 90176 97952
rect 90112 97892 90116 97948
rect 90116 97892 90172 97948
rect 90172 97892 90176 97948
rect 90112 97888 90176 97892
rect 90192 97948 90256 97952
rect 90192 97892 90196 97948
rect 90196 97892 90252 97948
rect 90252 97892 90256 97948
rect 90192 97888 90256 97892
rect 89300 97820 89364 97884
rect 3952 97404 4016 97408
rect 3952 97348 3956 97404
rect 3956 97348 4012 97404
rect 4012 97348 4016 97404
rect 3952 97344 4016 97348
rect 4032 97404 4096 97408
rect 4032 97348 4036 97404
rect 4036 97348 4092 97404
rect 4092 97348 4096 97404
rect 4032 97344 4096 97348
rect 4112 97404 4176 97408
rect 4112 97348 4116 97404
rect 4116 97348 4172 97404
rect 4172 97348 4176 97404
rect 4112 97344 4176 97348
rect 4192 97404 4256 97408
rect 4192 97348 4196 97404
rect 4196 97348 4252 97404
rect 4252 97348 4256 97404
rect 4192 97344 4256 97348
rect 87952 97404 88016 97408
rect 87952 97348 87956 97404
rect 87956 97348 88012 97404
rect 88012 97348 88016 97404
rect 87952 97344 88016 97348
rect 88032 97404 88096 97408
rect 88032 97348 88036 97404
rect 88036 97348 88092 97404
rect 88092 97348 88096 97404
rect 88032 97344 88096 97348
rect 88112 97404 88176 97408
rect 88112 97348 88116 97404
rect 88116 97348 88172 97404
rect 88172 97348 88176 97404
rect 88112 97344 88176 97348
rect 88192 97404 88256 97408
rect 88192 97348 88196 97404
rect 88196 97348 88252 97404
rect 88252 97348 88256 97404
rect 88192 97344 88256 97348
rect 85252 97276 85316 97340
rect 22692 97200 22756 97204
rect 22692 97144 22706 97200
rect 22706 97144 22756 97200
rect 22692 97140 22756 97144
rect 40356 97140 40420 97204
rect 14596 97064 14660 97068
rect 14596 97008 14646 97064
rect 14646 97008 14660 97064
rect 14596 97004 14660 97008
rect 17172 97064 17236 97068
rect 17172 97008 17186 97064
rect 17186 97008 17236 97064
rect 17172 97004 17236 97008
rect 18092 97064 18156 97068
rect 18092 97008 18106 97064
rect 18106 97008 18156 97064
rect 18092 97004 18156 97008
rect 24348 97064 24412 97068
rect 24348 97008 24362 97064
rect 24362 97008 24412 97064
rect 24348 97004 24412 97008
rect 25452 97064 25516 97068
rect 25452 97008 25466 97064
rect 25466 97008 25516 97064
rect 25452 97004 25516 97008
rect 30052 97064 30116 97068
rect 30052 97008 30102 97064
rect 30102 97008 30116 97064
rect 30052 97004 30116 97008
rect 32076 97064 32140 97068
rect 32076 97008 32090 97064
rect 32090 97008 32140 97064
rect 32076 97004 32140 97008
rect 33180 97064 33244 97068
rect 33180 97008 33194 97064
rect 33194 97008 33244 97064
rect 33180 97004 33244 97008
rect 35940 96868 36004 96932
rect 42932 97004 42996 97068
rect 1952 96860 2016 96864
rect 1952 96804 1956 96860
rect 1956 96804 2012 96860
rect 2012 96804 2016 96860
rect 1952 96800 2016 96804
rect 2032 96860 2096 96864
rect 2032 96804 2036 96860
rect 2036 96804 2092 96860
rect 2092 96804 2096 96860
rect 2032 96800 2096 96804
rect 2112 96860 2176 96864
rect 2112 96804 2116 96860
rect 2116 96804 2172 96860
rect 2172 96804 2176 96860
rect 2112 96800 2176 96804
rect 2192 96860 2256 96864
rect 2192 96804 2196 96860
rect 2196 96804 2252 96860
rect 2252 96804 2256 96860
rect 2192 96800 2256 96804
rect 40540 96732 40604 96796
rect 47164 96732 47228 96796
rect 54156 96868 54220 96932
rect 79916 97140 79980 97204
rect 87276 97140 87340 97204
rect 84884 96868 84948 96932
rect 52132 96732 52196 96796
rect 60596 96732 60660 96796
rect 61516 96792 61580 96796
rect 61516 96736 61566 96792
rect 61566 96736 61580 96792
rect 61516 96732 61580 96736
rect 61700 96792 61764 96796
rect 61700 96736 61750 96792
rect 61750 96736 61764 96792
rect 61700 96732 61764 96736
rect 42748 96596 42812 96660
rect 57836 96656 57900 96660
rect 57836 96600 57886 96656
rect 57886 96600 57900 96656
rect 57836 96596 57900 96600
rect 58020 96656 58084 96660
rect 58020 96600 58070 96656
rect 58070 96600 58084 96656
rect 58020 96596 58084 96600
rect 58388 96596 58452 96660
rect 59676 96656 59740 96660
rect 59676 96600 59726 96656
rect 59726 96600 59740 96656
rect 59676 96596 59740 96600
rect 60228 96596 60292 96660
rect 82492 96732 82556 96796
rect 87460 97004 87524 97068
rect 85952 96860 86016 96864
rect 85952 96804 85956 96860
rect 85956 96804 86012 96860
rect 86012 96804 86016 96860
rect 85952 96800 86016 96804
rect 86032 96860 86096 96864
rect 86032 96804 86036 96860
rect 86036 96804 86092 96860
rect 86092 96804 86096 96860
rect 86032 96800 86096 96804
rect 86112 96860 86176 96864
rect 86112 96804 86116 96860
rect 86116 96804 86172 96860
rect 86172 96804 86176 96860
rect 86112 96800 86176 96804
rect 86192 96860 86256 96864
rect 86192 96804 86196 96860
rect 86196 96804 86252 96860
rect 86252 96804 86256 96860
rect 86192 96800 86256 96804
rect 89952 96860 90016 96864
rect 89952 96804 89956 96860
rect 89956 96804 90012 96860
rect 90012 96804 90016 96860
rect 89952 96800 90016 96804
rect 90032 96860 90096 96864
rect 90032 96804 90036 96860
rect 90036 96804 90092 96860
rect 90092 96804 90096 96860
rect 90032 96800 90096 96804
rect 90112 96860 90176 96864
rect 90112 96804 90116 96860
rect 90116 96804 90172 96860
rect 90172 96804 90176 96860
rect 90112 96800 90176 96804
rect 90192 96860 90256 96864
rect 90192 96804 90196 96860
rect 90196 96804 90252 96860
rect 90252 96804 90256 96860
rect 90192 96800 90256 96804
rect 87644 96732 87708 96796
rect 16436 96520 16500 96524
rect 16436 96464 16486 96520
rect 16486 96464 16500 96520
rect 16436 96460 16500 96464
rect 15700 96384 15764 96388
rect 15700 96328 15750 96384
rect 15750 96328 15764 96384
rect 15700 96324 15764 96328
rect 21220 96324 21284 96388
rect 85804 96460 85868 96524
rect 50476 96324 50540 96388
rect 51028 96324 51092 96388
rect 3952 96316 4016 96320
rect 3952 96260 3956 96316
rect 3956 96260 4012 96316
rect 4012 96260 4016 96316
rect 3952 96256 4016 96260
rect 4032 96316 4096 96320
rect 4032 96260 4036 96316
rect 4036 96260 4092 96316
rect 4092 96260 4096 96316
rect 4032 96256 4096 96260
rect 4112 96316 4176 96320
rect 4112 96260 4116 96316
rect 4116 96260 4172 96316
rect 4172 96260 4176 96316
rect 4112 96256 4176 96260
rect 4192 96316 4256 96320
rect 4192 96260 4196 96316
rect 4196 96260 4252 96316
rect 4252 96260 4256 96316
rect 4192 96256 4256 96260
rect 9628 96248 9692 96252
rect 9628 96192 9642 96248
rect 9642 96192 9692 96248
rect 9628 96188 9692 96192
rect 22140 96248 22204 96252
rect 22140 96192 22154 96248
rect 22154 96192 22204 96248
rect 22140 96188 22204 96192
rect 27984 96248 28048 96252
rect 27984 96192 27986 96248
rect 27986 96192 28042 96248
rect 28042 96192 28048 96248
rect 27984 96188 28048 96192
rect 29152 96248 29216 96252
rect 29152 96192 29182 96248
rect 29182 96192 29216 96248
rect 29152 96188 29216 96192
rect 42000 96248 42064 96252
rect 87952 96316 88016 96320
rect 87952 96260 87956 96316
rect 87956 96260 88012 96316
rect 88012 96260 88016 96316
rect 87952 96256 88016 96260
rect 88032 96316 88096 96320
rect 88032 96260 88036 96316
rect 88036 96260 88092 96316
rect 88092 96260 88096 96316
rect 88032 96256 88096 96260
rect 88112 96316 88176 96320
rect 88112 96260 88116 96316
rect 88116 96260 88172 96316
rect 88172 96260 88176 96316
rect 88112 96256 88176 96260
rect 88192 96316 88256 96320
rect 88192 96260 88196 96316
rect 88196 96260 88252 96316
rect 88252 96260 88256 96316
rect 88192 96256 88256 96260
rect 42000 96192 42026 96248
rect 42026 96192 42064 96248
rect 42000 96188 42064 96192
rect 20976 96112 21040 96116
rect 20976 96056 20994 96112
rect 20994 96056 21040 96112
rect 20976 96052 21040 96056
rect 26816 96112 26880 96116
rect 26816 96056 26846 96112
rect 26846 96056 26880 96112
rect 26816 96052 26880 96056
rect 31488 96112 31552 96116
rect 31488 96056 31538 96112
rect 31538 96056 31552 96112
rect 31488 96052 31552 96056
rect 34992 96112 35056 96116
rect 34992 96056 35034 96112
rect 35034 96056 35056 96112
rect 34992 96052 35056 96056
rect 39620 95976 39684 95980
rect 39620 95920 39634 95976
rect 39634 95920 39684 95976
rect 39620 95916 39684 95920
rect 38516 95840 38580 95844
rect 38516 95784 38530 95840
rect 38530 95784 38580 95840
rect 38516 95780 38580 95784
rect 1952 95772 2016 95776
rect 1952 95716 1956 95772
rect 1956 95716 2012 95772
rect 2012 95716 2016 95772
rect 1952 95712 2016 95716
rect 2032 95772 2096 95776
rect 2032 95716 2036 95772
rect 2036 95716 2092 95772
rect 2092 95716 2096 95772
rect 2032 95712 2096 95716
rect 2112 95772 2176 95776
rect 2112 95716 2116 95772
rect 2116 95716 2172 95772
rect 2172 95716 2176 95772
rect 2112 95712 2176 95716
rect 2192 95772 2256 95776
rect 2192 95716 2196 95772
rect 2196 95716 2252 95772
rect 2252 95716 2256 95772
rect 2192 95712 2256 95716
rect 85952 95772 86016 95776
rect 85952 95716 85956 95772
rect 85956 95716 86012 95772
rect 86012 95716 86016 95772
rect 85952 95712 86016 95716
rect 86032 95772 86096 95776
rect 86032 95716 86036 95772
rect 86036 95716 86092 95772
rect 86092 95716 86096 95772
rect 86032 95712 86096 95716
rect 86112 95772 86176 95776
rect 86112 95716 86116 95772
rect 86116 95716 86172 95772
rect 86172 95716 86176 95772
rect 86112 95712 86176 95716
rect 86192 95772 86256 95776
rect 86192 95716 86196 95772
rect 86196 95716 86252 95772
rect 86252 95716 86256 95772
rect 86192 95712 86256 95716
rect 89952 95772 90016 95776
rect 89952 95716 89956 95772
rect 89956 95716 90012 95772
rect 90012 95716 90016 95772
rect 89952 95712 90016 95716
rect 90032 95772 90096 95776
rect 90032 95716 90036 95772
rect 90036 95716 90092 95772
rect 90092 95716 90096 95772
rect 90032 95712 90096 95716
rect 90112 95772 90176 95776
rect 90112 95716 90116 95772
rect 90116 95716 90172 95772
rect 90172 95716 90176 95772
rect 90112 95712 90176 95716
rect 90192 95772 90256 95776
rect 90192 95716 90196 95772
rect 90196 95716 90252 95772
rect 90252 95716 90256 95772
rect 90192 95712 90256 95716
rect 32996 95644 33060 95708
rect 28764 95508 28828 95572
rect 75132 95568 75196 95572
rect 75132 95512 75182 95568
rect 75182 95512 75196 95568
rect 75132 95508 75196 95512
rect 79180 95508 79244 95572
rect 23980 95372 24044 95436
rect 24532 95296 24596 95300
rect 24532 95240 24582 95296
rect 24582 95240 24596 95296
rect 24532 95236 24596 95240
rect 37780 95296 37844 95300
rect 37780 95240 37830 95296
rect 37830 95240 37844 95296
rect 37780 95236 37844 95240
rect 41092 95296 41156 95300
rect 41092 95240 41142 95296
rect 41142 95240 41156 95296
rect 41092 95236 41156 95240
rect 45324 95296 45388 95300
rect 45324 95240 45374 95296
rect 45374 95240 45388 95296
rect 45324 95236 45388 95240
rect 47900 95296 47964 95300
rect 47900 95240 47950 95296
rect 47950 95240 47964 95296
rect 47900 95236 47964 95240
rect 64092 95296 64156 95300
rect 64092 95240 64142 95296
rect 64142 95240 64156 95296
rect 64092 95236 64156 95240
rect 85620 95236 85684 95300
rect 3952 95228 4016 95232
rect 3952 95172 3956 95228
rect 3956 95172 4012 95228
rect 4012 95172 4016 95228
rect 3952 95168 4016 95172
rect 4032 95228 4096 95232
rect 4032 95172 4036 95228
rect 4036 95172 4092 95228
rect 4092 95172 4096 95228
rect 4032 95168 4096 95172
rect 4112 95228 4176 95232
rect 4112 95172 4116 95228
rect 4116 95172 4172 95228
rect 4172 95172 4176 95228
rect 4112 95168 4176 95172
rect 4192 95228 4256 95232
rect 4192 95172 4196 95228
rect 4196 95172 4252 95228
rect 4252 95172 4256 95228
rect 4192 95168 4256 95172
rect 87952 95228 88016 95232
rect 87952 95172 87956 95228
rect 87956 95172 88012 95228
rect 88012 95172 88016 95228
rect 87952 95168 88016 95172
rect 88032 95228 88096 95232
rect 88032 95172 88036 95228
rect 88036 95172 88092 95228
rect 88092 95172 88096 95228
rect 88032 95168 88096 95172
rect 88112 95228 88176 95232
rect 88112 95172 88116 95228
rect 88116 95172 88172 95228
rect 88172 95172 88176 95228
rect 88112 95168 88176 95172
rect 88192 95228 88256 95232
rect 88192 95172 88196 95228
rect 88196 95172 88252 95228
rect 88252 95172 88256 95228
rect 88192 95168 88256 95172
rect 12756 95160 12820 95164
rect 12756 95104 12806 95160
rect 12806 95104 12820 95160
rect 12756 95100 12820 95104
rect 19380 95160 19444 95164
rect 19380 95104 19394 95160
rect 19394 95104 19444 95160
rect 19380 95100 19444 95104
rect 24716 95160 24780 95164
rect 24716 95104 24766 95160
rect 24766 95104 24780 95160
rect 24716 95100 24780 95104
rect 25820 95100 25884 95164
rect 27476 95100 27540 95164
rect 22876 94964 22940 95028
rect 29868 94964 29932 95028
rect 30972 94964 31036 95028
rect 37964 95100 38028 95164
rect 43852 95100 43916 95164
rect 44404 95100 44468 95164
rect 45508 95160 45572 95164
rect 45508 95104 45558 95160
rect 45558 95104 45572 95160
rect 45508 95100 45572 95104
rect 46612 95160 46676 95164
rect 46612 95104 46662 95160
rect 46662 95104 46676 95160
rect 46612 95100 46676 95104
rect 48084 95160 48148 95164
rect 48084 95104 48134 95160
rect 48134 95104 48148 95160
rect 48084 95100 48148 95104
rect 79732 94964 79796 95028
rect 80468 95024 80532 95028
rect 80468 94968 80518 95024
rect 80518 94968 80532 95024
rect 80468 94964 80532 94968
rect 19932 94828 19996 94892
rect 31708 94828 31772 94892
rect 83780 94828 83844 94892
rect 34468 94692 34532 94756
rect 1952 94684 2016 94688
rect 1952 94628 1956 94684
rect 1956 94628 2012 94684
rect 2012 94628 2016 94684
rect 1952 94624 2016 94628
rect 2032 94684 2096 94688
rect 2032 94628 2036 94684
rect 2036 94628 2092 94684
rect 2092 94628 2096 94684
rect 2032 94624 2096 94628
rect 2112 94684 2176 94688
rect 2112 94628 2116 94684
rect 2116 94628 2172 94684
rect 2172 94628 2176 94684
rect 2112 94624 2176 94628
rect 2192 94684 2256 94688
rect 2192 94628 2196 94684
rect 2196 94628 2252 94684
rect 2252 94628 2256 94684
rect 2192 94624 2256 94628
rect 85952 94684 86016 94688
rect 85952 94628 85956 94684
rect 85956 94628 86012 94684
rect 86012 94628 86016 94684
rect 85952 94624 86016 94628
rect 86032 94684 86096 94688
rect 86032 94628 86036 94684
rect 86036 94628 86092 94684
rect 86092 94628 86096 94684
rect 86032 94624 86096 94628
rect 86112 94684 86176 94688
rect 86112 94628 86116 94684
rect 86116 94628 86172 94684
rect 86172 94628 86176 94684
rect 86112 94624 86176 94628
rect 86192 94684 86256 94688
rect 86192 94628 86196 94684
rect 86196 94628 86252 94684
rect 86252 94628 86256 94684
rect 86192 94624 86256 94628
rect 89952 94684 90016 94688
rect 89952 94628 89956 94684
rect 89956 94628 90012 94684
rect 90012 94628 90016 94684
rect 89952 94624 90016 94628
rect 90032 94684 90096 94688
rect 90032 94628 90036 94684
rect 90036 94628 90092 94684
rect 90092 94628 90096 94684
rect 90032 94624 90096 94628
rect 90112 94684 90176 94688
rect 90112 94628 90116 94684
rect 90116 94628 90172 94684
rect 90172 94628 90176 94684
rect 90112 94624 90176 94628
rect 90192 94684 90256 94688
rect 90192 94628 90196 94684
rect 90196 94628 90252 94684
rect 90252 94628 90256 94684
rect 90192 94624 90256 94628
rect 37228 94616 37292 94620
rect 37228 94560 37278 94616
rect 37278 94560 37292 94616
rect 37228 94556 37292 94560
rect 36860 94420 36924 94484
rect 42564 94420 42628 94484
rect 44956 94420 45020 94484
rect 46244 94420 46308 94484
rect 84148 94420 84212 94484
rect 39988 94284 40052 94348
rect 83596 94284 83660 94348
rect 39252 94148 39316 94212
rect 3952 94140 4016 94144
rect 3952 94084 3956 94140
rect 3956 94084 4012 94140
rect 4012 94084 4016 94140
rect 3952 94080 4016 94084
rect 4032 94140 4096 94144
rect 4032 94084 4036 94140
rect 4036 94084 4092 94140
rect 4092 94084 4096 94140
rect 4032 94080 4096 94084
rect 4112 94140 4176 94144
rect 4112 94084 4116 94140
rect 4116 94084 4172 94140
rect 4172 94084 4176 94140
rect 4112 94080 4176 94084
rect 4192 94140 4256 94144
rect 4192 94084 4196 94140
rect 4196 94084 4252 94140
rect 4252 94084 4256 94140
rect 4192 94080 4256 94084
rect 41276 94012 41340 94076
rect 83412 94148 83476 94212
rect 87952 94140 88016 94144
rect 87952 94084 87956 94140
rect 87956 94084 88012 94140
rect 88012 94084 88016 94140
rect 87952 94080 88016 94084
rect 88032 94140 88096 94144
rect 88032 94084 88036 94140
rect 88036 94084 88092 94140
rect 88092 94084 88096 94140
rect 88032 94080 88096 94084
rect 88112 94140 88176 94144
rect 88112 94084 88116 94140
rect 88116 94084 88172 94140
rect 88172 94084 88176 94140
rect 88112 94080 88176 94084
rect 88192 94140 88256 94144
rect 88192 94084 88196 94140
rect 88196 94084 88252 94140
rect 88252 94084 88256 94140
rect 88192 94080 88256 94084
rect 19196 93876 19260 93940
rect 86540 94012 86604 94076
rect 86356 93876 86420 93940
rect 35756 93740 35820 93804
rect 82492 93740 82556 93804
rect 83412 93740 83476 93804
rect 31708 93604 31772 93668
rect 42564 93664 42628 93668
rect 42564 93608 42614 93664
rect 42614 93608 42628 93664
rect 42564 93604 42628 93608
rect 44036 93664 44100 93668
rect 44036 93608 44086 93664
rect 44086 93608 44100 93664
rect 44036 93604 44100 93608
rect 46612 93664 46676 93668
rect 46612 93608 46662 93664
rect 46662 93608 46676 93664
rect 46612 93604 46676 93608
rect 47900 93664 47964 93668
rect 47900 93608 47950 93664
rect 47950 93608 47964 93664
rect 47900 93604 47964 93608
rect 48268 93604 48332 93668
rect 49004 93664 49068 93668
rect 49004 93608 49054 93664
rect 49054 93608 49068 93664
rect 49004 93604 49068 93608
rect 49188 93604 49252 93668
rect 49924 93664 49988 93668
rect 49924 93608 49974 93664
rect 49974 93608 49988 93664
rect 49924 93604 49988 93608
rect 50292 93604 50356 93668
rect 51212 93664 51276 93668
rect 51212 93608 51262 93664
rect 51262 93608 51276 93664
rect 51212 93604 51276 93608
rect 51396 93664 51460 93668
rect 51396 93608 51446 93664
rect 51446 93608 51460 93664
rect 51396 93604 51460 93608
rect 52132 93664 52196 93668
rect 52132 93608 52182 93664
rect 52182 93608 52196 93664
rect 52132 93604 52196 93608
rect 52500 93664 52564 93668
rect 52500 93608 52550 93664
rect 52550 93608 52564 93664
rect 52500 93604 52564 93608
rect 53236 93664 53300 93668
rect 53236 93608 53286 93664
rect 53286 93608 53300 93664
rect 53236 93604 53300 93608
rect 53788 93664 53852 93668
rect 53788 93608 53802 93664
rect 53802 93608 53852 93664
rect 53788 93604 53852 93608
rect 53972 93664 54036 93668
rect 53972 93608 54022 93664
rect 54022 93608 54036 93664
rect 53972 93604 54036 93608
rect 54340 93604 54404 93668
rect 54524 93664 54588 93668
rect 54524 93608 54574 93664
rect 54574 93608 54588 93664
rect 54524 93604 54588 93608
rect 54892 93664 54956 93668
rect 54892 93608 54942 93664
rect 54942 93608 54956 93664
rect 54892 93604 54956 93608
rect 55260 93604 55324 93668
rect 1952 93596 2016 93600
rect 1952 93540 1956 93596
rect 1956 93540 2012 93596
rect 2012 93540 2016 93596
rect 1952 93536 2016 93540
rect 2032 93596 2096 93600
rect 2032 93540 2036 93596
rect 2036 93540 2092 93596
rect 2092 93540 2096 93596
rect 2032 93536 2096 93540
rect 2112 93596 2176 93600
rect 2112 93540 2116 93596
rect 2116 93540 2172 93596
rect 2172 93540 2176 93596
rect 2112 93536 2176 93540
rect 2192 93596 2256 93600
rect 2192 93540 2196 93596
rect 2196 93540 2252 93596
rect 2252 93540 2256 93596
rect 2192 93536 2256 93540
rect 84332 93604 84396 93668
rect 85068 93664 85132 93668
rect 85068 93608 85118 93664
rect 85118 93608 85132 93664
rect 85068 93604 85132 93608
rect 85952 93596 86016 93600
rect 85952 93540 85956 93596
rect 85956 93540 86012 93596
rect 86012 93540 86016 93596
rect 85952 93536 86016 93540
rect 86032 93596 86096 93600
rect 86032 93540 86036 93596
rect 86036 93540 86092 93596
rect 86092 93540 86096 93596
rect 86032 93536 86096 93540
rect 86112 93596 86176 93600
rect 86112 93540 86116 93596
rect 86116 93540 86172 93596
rect 86172 93540 86176 93596
rect 86112 93536 86176 93540
rect 86192 93596 86256 93600
rect 86192 93540 86196 93596
rect 86196 93540 86252 93596
rect 86252 93540 86256 93596
rect 86192 93536 86256 93540
rect 89952 93596 90016 93600
rect 89952 93540 89956 93596
rect 89956 93540 90012 93596
rect 90012 93540 90016 93596
rect 89952 93536 90016 93540
rect 90032 93596 90096 93600
rect 90032 93540 90036 93596
rect 90036 93540 90092 93596
rect 90092 93540 90096 93596
rect 90032 93536 90096 93540
rect 90112 93596 90176 93600
rect 90112 93540 90116 93596
rect 90116 93540 90172 93596
rect 90172 93540 90176 93596
rect 90112 93536 90176 93540
rect 90192 93596 90256 93600
rect 90192 93540 90196 93596
rect 90196 93540 90252 93596
rect 90252 93540 90256 93596
rect 90192 93536 90256 93540
rect 30236 93332 30300 93396
rect 27476 93196 27540 93260
rect 83780 93332 83844 93396
rect 28948 93060 29012 93124
rect 83596 93060 83660 93124
rect 3952 93052 4016 93056
rect 3952 92996 3956 93052
rect 3956 92996 4012 93052
rect 4012 92996 4016 93052
rect 3952 92992 4016 92996
rect 4032 93052 4096 93056
rect 4032 92996 4036 93052
rect 4036 92996 4092 93052
rect 4092 92996 4096 93052
rect 4032 92992 4096 92996
rect 4112 93052 4176 93056
rect 4112 92996 4116 93052
rect 4116 92996 4172 93052
rect 4172 92996 4176 93052
rect 4112 92992 4176 92996
rect 4192 93052 4256 93056
rect 4192 92996 4196 93052
rect 4196 92996 4252 93052
rect 4252 92996 4256 93052
rect 4192 92992 4256 92996
rect 87952 93052 88016 93056
rect 87952 92996 87956 93052
rect 87956 92996 88012 93052
rect 88012 92996 88016 93052
rect 87952 92992 88016 92996
rect 88032 93052 88096 93056
rect 88032 92996 88036 93052
rect 88036 92996 88092 93052
rect 88092 92996 88096 93052
rect 88032 92992 88096 92996
rect 88112 93052 88176 93056
rect 88112 92996 88116 93052
rect 88116 92996 88172 93052
rect 88172 92996 88176 93052
rect 88112 92992 88176 92996
rect 88192 93052 88256 93056
rect 88192 92996 88196 93052
rect 88196 92996 88252 93052
rect 88252 92996 88256 93052
rect 88192 92992 88256 92996
rect 26188 92924 26252 92988
rect 32812 92848 32876 92852
rect 32812 92792 32862 92848
rect 32862 92792 32876 92848
rect 32812 92788 32876 92792
rect 34100 92848 34164 92852
rect 34100 92792 34150 92848
rect 34150 92792 34164 92848
rect 34100 92788 34164 92792
rect 35204 92848 35268 92852
rect 35204 92792 35254 92848
rect 35254 92792 35268 92848
rect 35204 92788 35268 92792
rect 36676 92848 36740 92852
rect 36676 92792 36726 92848
rect 36726 92792 36740 92848
rect 36676 92788 36740 92792
rect 38332 92848 38396 92852
rect 38332 92792 38382 92848
rect 38382 92792 38396 92848
rect 38332 92788 38396 92792
rect 39988 92848 40052 92852
rect 39988 92792 40002 92848
rect 40002 92792 40052 92848
rect 39988 92788 40052 92792
rect 80100 92788 80164 92852
rect 87276 92788 87340 92852
rect 1952 92508 2016 92512
rect 1952 92452 1956 92508
rect 1956 92452 2012 92508
rect 2012 92452 2016 92508
rect 1952 92448 2016 92452
rect 2032 92508 2096 92512
rect 2032 92452 2036 92508
rect 2036 92452 2092 92508
rect 2092 92452 2096 92508
rect 2032 92448 2096 92452
rect 2112 92508 2176 92512
rect 2112 92452 2116 92508
rect 2116 92452 2172 92508
rect 2172 92452 2176 92508
rect 2112 92448 2176 92452
rect 2192 92508 2256 92512
rect 2192 92452 2196 92508
rect 2196 92452 2252 92508
rect 2252 92452 2256 92508
rect 2192 92448 2256 92452
rect 85952 92508 86016 92512
rect 85952 92452 85956 92508
rect 85956 92452 86012 92508
rect 86012 92452 86016 92508
rect 85952 92448 86016 92452
rect 86032 92508 86096 92512
rect 86032 92452 86036 92508
rect 86036 92452 86092 92508
rect 86092 92452 86096 92508
rect 86032 92448 86096 92452
rect 86112 92508 86176 92512
rect 86112 92452 86116 92508
rect 86116 92452 86172 92508
rect 86172 92452 86176 92508
rect 86112 92448 86176 92452
rect 86192 92508 86256 92512
rect 86192 92452 86196 92508
rect 86196 92452 86252 92508
rect 86252 92452 86256 92508
rect 86192 92448 86256 92452
rect 89952 92508 90016 92512
rect 89952 92452 89956 92508
rect 89956 92452 90012 92508
rect 90012 92452 90016 92508
rect 89952 92448 90016 92452
rect 90032 92508 90096 92512
rect 90032 92452 90036 92508
rect 90036 92452 90092 92508
rect 90092 92452 90096 92508
rect 90032 92448 90096 92452
rect 90112 92508 90176 92512
rect 90112 92452 90116 92508
rect 90116 92452 90172 92508
rect 90172 92452 90176 92508
rect 90112 92448 90176 92452
rect 90192 92508 90256 92512
rect 90192 92452 90196 92508
rect 90196 92452 90252 92508
rect 90252 92452 90256 92508
rect 90192 92448 90256 92452
rect 4844 92380 4908 92444
rect 3952 91964 4016 91968
rect 3952 91908 3956 91964
rect 3956 91908 4012 91964
rect 4012 91908 4016 91964
rect 3952 91904 4016 91908
rect 4032 91964 4096 91968
rect 4032 91908 4036 91964
rect 4036 91908 4092 91964
rect 4092 91908 4096 91964
rect 4032 91904 4096 91908
rect 4112 91964 4176 91968
rect 4112 91908 4116 91964
rect 4116 91908 4172 91964
rect 4172 91908 4176 91964
rect 4112 91904 4176 91908
rect 4192 91964 4256 91968
rect 4192 91908 4196 91964
rect 4196 91908 4252 91964
rect 4252 91908 4256 91964
rect 4192 91904 4256 91908
rect 87952 91964 88016 91968
rect 87952 91908 87956 91964
rect 87956 91908 88012 91964
rect 88012 91908 88016 91964
rect 87952 91904 88016 91908
rect 88032 91964 88096 91968
rect 88032 91908 88036 91964
rect 88036 91908 88092 91964
rect 88092 91908 88096 91964
rect 88032 91904 88096 91908
rect 88112 91964 88176 91968
rect 88112 91908 88116 91964
rect 88116 91908 88172 91964
rect 88172 91908 88176 91964
rect 88112 91904 88176 91908
rect 88192 91964 88256 91968
rect 88192 91908 88196 91964
rect 88196 91908 88252 91964
rect 88252 91908 88256 91964
rect 88192 91904 88256 91908
rect 86908 91700 86972 91764
rect 1952 91420 2016 91424
rect 1952 91364 1956 91420
rect 1956 91364 2012 91420
rect 2012 91364 2016 91420
rect 1952 91360 2016 91364
rect 2032 91420 2096 91424
rect 2032 91364 2036 91420
rect 2036 91364 2092 91420
rect 2092 91364 2096 91420
rect 2032 91360 2096 91364
rect 2112 91420 2176 91424
rect 2112 91364 2116 91420
rect 2116 91364 2172 91420
rect 2172 91364 2176 91420
rect 2112 91360 2176 91364
rect 2192 91420 2256 91424
rect 2192 91364 2196 91420
rect 2196 91364 2252 91420
rect 2252 91364 2256 91420
rect 2192 91360 2256 91364
rect 85952 91420 86016 91424
rect 85952 91364 85956 91420
rect 85956 91364 86012 91420
rect 86012 91364 86016 91420
rect 85952 91360 86016 91364
rect 86032 91420 86096 91424
rect 86032 91364 86036 91420
rect 86036 91364 86092 91420
rect 86092 91364 86096 91420
rect 86032 91360 86096 91364
rect 86112 91420 86176 91424
rect 86112 91364 86116 91420
rect 86116 91364 86172 91420
rect 86172 91364 86176 91420
rect 86112 91360 86176 91364
rect 86192 91420 86256 91424
rect 86192 91364 86196 91420
rect 86196 91364 86252 91420
rect 86252 91364 86256 91420
rect 86192 91360 86256 91364
rect 89952 91420 90016 91424
rect 89952 91364 89956 91420
rect 89956 91364 90012 91420
rect 90012 91364 90016 91420
rect 89952 91360 90016 91364
rect 90032 91420 90096 91424
rect 90032 91364 90036 91420
rect 90036 91364 90092 91420
rect 90092 91364 90096 91420
rect 90032 91360 90096 91364
rect 90112 91420 90176 91424
rect 90112 91364 90116 91420
rect 90116 91364 90172 91420
rect 90172 91364 90176 91420
rect 90112 91360 90176 91364
rect 90192 91420 90256 91424
rect 90192 91364 90196 91420
rect 90196 91364 90252 91420
rect 90252 91364 90256 91420
rect 90192 91360 90256 91364
rect 3952 90876 4016 90880
rect 3952 90820 3956 90876
rect 3956 90820 4012 90876
rect 4012 90820 4016 90876
rect 3952 90816 4016 90820
rect 4032 90876 4096 90880
rect 4032 90820 4036 90876
rect 4036 90820 4092 90876
rect 4092 90820 4096 90876
rect 4032 90816 4096 90820
rect 4112 90876 4176 90880
rect 4112 90820 4116 90876
rect 4116 90820 4172 90876
rect 4172 90820 4176 90876
rect 4112 90816 4176 90820
rect 4192 90876 4256 90880
rect 4192 90820 4196 90876
rect 4196 90820 4252 90876
rect 4252 90820 4256 90876
rect 4192 90816 4256 90820
rect 87952 90876 88016 90880
rect 87952 90820 87956 90876
rect 87956 90820 88012 90876
rect 88012 90820 88016 90876
rect 87952 90816 88016 90820
rect 88032 90876 88096 90880
rect 88032 90820 88036 90876
rect 88036 90820 88092 90876
rect 88092 90820 88096 90876
rect 88032 90816 88096 90820
rect 88112 90876 88176 90880
rect 88112 90820 88116 90876
rect 88116 90820 88172 90876
rect 88172 90820 88176 90876
rect 88112 90816 88176 90820
rect 88192 90876 88256 90880
rect 88192 90820 88196 90876
rect 88196 90820 88252 90876
rect 88252 90820 88256 90876
rect 88192 90816 88256 90820
rect 86908 90476 86972 90540
rect 1952 90332 2016 90336
rect 1952 90276 1956 90332
rect 1956 90276 2012 90332
rect 2012 90276 2016 90332
rect 1952 90272 2016 90276
rect 2032 90332 2096 90336
rect 2032 90276 2036 90332
rect 2036 90276 2092 90332
rect 2092 90276 2096 90332
rect 2032 90272 2096 90276
rect 2112 90332 2176 90336
rect 2112 90276 2116 90332
rect 2116 90276 2172 90332
rect 2172 90276 2176 90332
rect 2112 90272 2176 90276
rect 2192 90332 2256 90336
rect 2192 90276 2196 90332
rect 2196 90276 2252 90332
rect 2252 90276 2256 90332
rect 2192 90272 2256 90276
rect 85952 90332 86016 90336
rect 85952 90276 85956 90332
rect 85956 90276 86012 90332
rect 86012 90276 86016 90332
rect 85952 90272 86016 90276
rect 86032 90332 86096 90336
rect 86032 90276 86036 90332
rect 86036 90276 86092 90332
rect 86092 90276 86096 90332
rect 86032 90272 86096 90276
rect 86112 90332 86176 90336
rect 86112 90276 86116 90332
rect 86116 90276 86172 90332
rect 86172 90276 86176 90332
rect 86112 90272 86176 90276
rect 86192 90332 86256 90336
rect 86192 90276 86196 90332
rect 86196 90276 86252 90332
rect 86252 90276 86256 90332
rect 86192 90272 86256 90276
rect 89952 90332 90016 90336
rect 89952 90276 89956 90332
rect 89956 90276 90012 90332
rect 90012 90276 90016 90332
rect 89952 90272 90016 90276
rect 90032 90332 90096 90336
rect 90032 90276 90036 90332
rect 90036 90276 90092 90332
rect 90092 90276 90096 90332
rect 90032 90272 90096 90276
rect 90112 90332 90176 90336
rect 90112 90276 90116 90332
rect 90116 90276 90172 90332
rect 90172 90276 90176 90332
rect 90112 90272 90176 90276
rect 90192 90332 90256 90336
rect 90192 90276 90196 90332
rect 90196 90276 90252 90332
rect 90252 90276 90256 90332
rect 90192 90272 90256 90276
rect 3952 89788 4016 89792
rect 3952 89732 3956 89788
rect 3956 89732 4012 89788
rect 4012 89732 4016 89788
rect 3952 89728 4016 89732
rect 4032 89788 4096 89792
rect 4032 89732 4036 89788
rect 4036 89732 4092 89788
rect 4092 89732 4096 89788
rect 4032 89728 4096 89732
rect 4112 89788 4176 89792
rect 4112 89732 4116 89788
rect 4116 89732 4172 89788
rect 4172 89732 4176 89788
rect 4112 89728 4176 89732
rect 4192 89788 4256 89792
rect 4192 89732 4196 89788
rect 4196 89732 4252 89788
rect 4252 89732 4256 89788
rect 4192 89728 4256 89732
rect 87952 89788 88016 89792
rect 87952 89732 87956 89788
rect 87956 89732 88012 89788
rect 88012 89732 88016 89788
rect 87952 89728 88016 89732
rect 88032 89788 88096 89792
rect 88032 89732 88036 89788
rect 88036 89732 88092 89788
rect 88092 89732 88096 89788
rect 88032 89728 88096 89732
rect 88112 89788 88176 89792
rect 88112 89732 88116 89788
rect 88116 89732 88172 89788
rect 88172 89732 88176 89788
rect 88112 89728 88176 89732
rect 88192 89788 88256 89792
rect 88192 89732 88196 89788
rect 88196 89732 88252 89788
rect 88252 89732 88256 89788
rect 88192 89728 88256 89732
rect 5212 89448 5276 89452
rect 5212 89392 5226 89448
rect 5226 89392 5276 89448
rect 5212 89388 5276 89392
rect 1952 89244 2016 89248
rect 1952 89188 1956 89244
rect 1956 89188 2012 89244
rect 2012 89188 2016 89244
rect 1952 89184 2016 89188
rect 2032 89244 2096 89248
rect 2032 89188 2036 89244
rect 2036 89188 2092 89244
rect 2092 89188 2096 89244
rect 2032 89184 2096 89188
rect 2112 89244 2176 89248
rect 2112 89188 2116 89244
rect 2116 89188 2172 89244
rect 2172 89188 2176 89244
rect 2112 89184 2176 89188
rect 2192 89244 2256 89248
rect 2192 89188 2196 89244
rect 2196 89188 2252 89244
rect 2252 89188 2256 89244
rect 2192 89184 2256 89188
rect 85952 89244 86016 89248
rect 85952 89188 85956 89244
rect 85956 89188 86012 89244
rect 86012 89188 86016 89244
rect 85952 89184 86016 89188
rect 86032 89244 86096 89248
rect 86032 89188 86036 89244
rect 86036 89188 86092 89244
rect 86092 89188 86096 89244
rect 86032 89184 86096 89188
rect 86112 89244 86176 89248
rect 86112 89188 86116 89244
rect 86116 89188 86172 89244
rect 86172 89188 86176 89244
rect 86112 89184 86176 89188
rect 86192 89244 86256 89248
rect 86192 89188 86196 89244
rect 86196 89188 86252 89244
rect 86252 89188 86256 89244
rect 86192 89184 86256 89188
rect 89952 89244 90016 89248
rect 89952 89188 89956 89244
rect 89956 89188 90012 89244
rect 90012 89188 90016 89244
rect 89952 89184 90016 89188
rect 90032 89244 90096 89248
rect 90032 89188 90036 89244
rect 90036 89188 90092 89244
rect 90092 89188 90096 89244
rect 90032 89184 90096 89188
rect 90112 89244 90176 89248
rect 90112 89188 90116 89244
rect 90116 89188 90172 89244
rect 90172 89188 90176 89244
rect 90112 89184 90176 89188
rect 90192 89244 90256 89248
rect 90192 89188 90196 89244
rect 90196 89188 90252 89244
rect 90252 89188 90256 89244
rect 90192 89184 90256 89188
rect 5580 89116 5644 89180
rect 86908 88980 86972 89044
rect 4844 88904 4908 88908
rect 4844 88848 4858 88904
rect 4858 88848 4908 88904
rect 4844 88844 4908 88848
rect 5212 88768 5276 88772
rect 5212 88712 5262 88768
rect 5262 88712 5276 88768
rect 5212 88708 5276 88712
rect 3952 88700 4016 88704
rect 3952 88644 3956 88700
rect 3956 88644 4012 88700
rect 4012 88644 4016 88700
rect 3952 88640 4016 88644
rect 4032 88700 4096 88704
rect 4032 88644 4036 88700
rect 4036 88644 4092 88700
rect 4092 88644 4096 88700
rect 4032 88640 4096 88644
rect 4112 88700 4176 88704
rect 4112 88644 4116 88700
rect 4116 88644 4172 88700
rect 4172 88644 4176 88700
rect 4112 88640 4176 88644
rect 4192 88700 4256 88704
rect 4192 88644 4196 88700
rect 4196 88644 4252 88700
rect 4252 88644 4256 88700
rect 4192 88640 4256 88644
rect 87952 88700 88016 88704
rect 87952 88644 87956 88700
rect 87956 88644 88012 88700
rect 88012 88644 88016 88700
rect 87952 88640 88016 88644
rect 88032 88700 88096 88704
rect 88032 88644 88036 88700
rect 88036 88644 88092 88700
rect 88092 88644 88096 88700
rect 88032 88640 88096 88644
rect 88112 88700 88176 88704
rect 88112 88644 88116 88700
rect 88116 88644 88172 88700
rect 88172 88644 88176 88700
rect 88112 88640 88176 88644
rect 88192 88700 88256 88704
rect 88192 88644 88196 88700
rect 88196 88644 88252 88700
rect 88252 88644 88256 88700
rect 88192 88640 88256 88644
rect 1952 88156 2016 88160
rect 1952 88100 1956 88156
rect 1956 88100 2012 88156
rect 2012 88100 2016 88156
rect 1952 88096 2016 88100
rect 2032 88156 2096 88160
rect 2032 88100 2036 88156
rect 2036 88100 2092 88156
rect 2092 88100 2096 88156
rect 2032 88096 2096 88100
rect 2112 88156 2176 88160
rect 2112 88100 2116 88156
rect 2116 88100 2172 88156
rect 2172 88100 2176 88156
rect 2112 88096 2176 88100
rect 2192 88156 2256 88160
rect 2192 88100 2196 88156
rect 2196 88100 2252 88156
rect 2252 88100 2256 88156
rect 2192 88096 2256 88100
rect 85952 88156 86016 88160
rect 85952 88100 85956 88156
rect 85956 88100 86012 88156
rect 86012 88100 86016 88156
rect 85952 88096 86016 88100
rect 86032 88156 86096 88160
rect 86032 88100 86036 88156
rect 86036 88100 86092 88156
rect 86092 88100 86096 88156
rect 86032 88096 86096 88100
rect 86112 88156 86176 88160
rect 86112 88100 86116 88156
rect 86116 88100 86172 88156
rect 86172 88100 86176 88156
rect 86112 88096 86176 88100
rect 86192 88156 86256 88160
rect 86192 88100 86196 88156
rect 86196 88100 86252 88156
rect 86252 88100 86256 88156
rect 86192 88096 86256 88100
rect 89952 88156 90016 88160
rect 89952 88100 89956 88156
rect 89956 88100 90012 88156
rect 90012 88100 90016 88156
rect 89952 88096 90016 88100
rect 90032 88156 90096 88160
rect 90032 88100 90036 88156
rect 90036 88100 90092 88156
rect 90092 88100 90096 88156
rect 90032 88096 90096 88100
rect 90112 88156 90176 88160
rect 90112 88100 90116 88156
rect 90116 88100 90172 88156
rect 90172 88100 90176 88156
rect 90112 88096 90176 88100
rect 90192 88156 90256 88160
rect 90192 88100 90196 88156
rect 90196 88100 90252 88156
rect 90252 88100 90256 88156
rect 90192 88096 90256 88100
rect 3952 87612 4016 87616
rect 3952 87556 3956 87612
rect 3956 87556 4012 87612
rect 4012 87556 4016 87612
rect 3952 87552 4016 87556
rect 4032 87612 4096 87616
rect 4032 87556 4036 87612
rect 4036 87556 4092 87612
rect 4092 87556 4096 87612
rect 4032 87552 4096 87556
rect 4112 87612 4176 87616
rect 4112 87556 4116 87612
rect 4116 87556 4172 87612
rect 4172 87556 4176 87612
rect 4112 87552 4176 87556
rect 4192 87612 4256 87616
rect 4192 87556 4196 87612
rect 4196 87556 4252 87612
rect 4252 87556 4256 87612
rect 4192 87552 4256 87556
rect 87952 87612 88016 87616
rect 87952 87556 87956 87612
rect 87956 87556 88012 87612
rect 88012 87556 88016 87612
rect 87952 87552 88016 87556
rect 88032 87612 88096 87616
rect 88032 87556 88036 87612
rect 88036 87556 88092 87612
rect 88092 87556 88096 87612
rect 88032 87552 88096 87556
rect 88112 87612 88176 87616
rect 88112 87556 88116 87612
rect 88116 87556 88172 87612
rect 88172 87556 88176 87612
rect 88112 87552 88176 87556
rect 88192 87612 88256 87616
rect 88192 87556 88196 87612
rect 88196 87556 88252 87612
rect 88252 87556 88256 87612
rect 88192 87552 88256 87556
rect 1952 87068 2016 87072
rect 1952 87012 1956 87068
rect 1956 87012 2012 87068
rect 2012 87012 2016 87068
rect 1952 87008 2016 87012
rect 2032 87068 2096 87072
rect 2032 87012 2036 87068
rect 2036 87012 2092 87068
rect 2092 87012 2096 87068
rect 2032 87008 2096 87012
rect 2112 87068 2176 87072
rect 2112 87012 2116 87068
rect 2116 87012 2172 87068
rect 2172 87012 2176 87068
rect 2112 87008 2176 87012
rect 2192 87068 2256 87072
rect 2192 87012 2196 87068
rect 2196 87012 2252 87068
rect 2252 87012 2256 87068
rect 2192 87008 2256 87012
rect 85952 87068 86016 87072
rect 85952 87012 85956 87068
rect 85956 87012 86012 87068
rect 86012 87012 86016 87068
rect 85952 87008 86016 87012
rect 86032 87068 86096 87072
rect 86032 87012 86036 87068
rect 86036 87012 86092 87068
rect 86092 87012 86096 87068
rect 86032 87008 86096 87012
rect 86112 87068 86176 87072
rect 86112 87012 86116 87068
rect 86116 87012 86172 87068
rect 86172 87012 86176 87068
rect 86112 87008 86176 87012
rect 86192 87068 86256 87072
rect 86192 87012 86196 87068
rect 86196 87012 86252 87068
rect 86252 87012 86256 87068
rect 86192 87008 86256 87012
rect 89952 87068 90016 87072
rect 89952 87012 89956 87068
rect 89956 87012 90012 87068
rect 90012 87012 90016 87068
rect 89952 87008 90016 87012
rect 90032 87068 90096 87072
rect 90032 87012 90036 87068
rect 90036 87012 90092 87068
rect 90092 87012 90096 87068
rect 90032 87008 90096 87012
rect 90112 87068 90176 87072
rect 90112 87012 90116 87068
rect 90116 87012 90172 87068
rect 90172 87012 90176 87068
rect 90112 87008 90176 87012
rect 90192 87068 90256 87072
rect 90192 87012 90196 87068
rect 90196 87012 90252 87068
rect 90252 87012 90256 87068
rect 90192 87008 90256 87012
rect 5396 86668 5460 86732
rect 3952 86524 4016 86528
rect 3952 86468 3956 86524
rect 3956 86468 4012 86524
rect 4012 86468 4016 86524
rect 3952 86464 4016 86468
rect 4032 86524 4096 86528
rect 4032 86468 4036 86524
rect 4036 86468 4092 86524
rect 4092 86468 4096 86524
rect 4032 86464 4096 86468
rect 4112 86524 4176 86528
rect 4112 86468 4116 86524
rect 4116 86468 4172 86524
rect 4172 86468 4176 86524
rect 4112 86464 4176 86468
rect 4192 86524 4256 86528
rect 4192 86468 4196 86524
rect 4196 86468 4252 86524
rect 4252 86468 4256 86524
rect 4192 86464 4256 86468
rect 87952 86524 88016 86528
rect 87952 86468 87956 86524
rect 87956 86468 88012 86524
rect 88012 86468 88016 86524
rect 87952 86464 88016 86468
rect 88032 86524 88096 86528
rect 88032 86468 88036 86524
rect 88036 86468 88092 86524
rect 88092 86468 88096 86524
rect 88032 86464 88096 86468
rect 88112 86524 88176 86528
rect 88112 86468 88116 86524
rect 88116 86468 88172 86524
rect 88172 86468 88176 86524
rect 88112 86464 88176 86468
rect 88192 86524 88256 86528
rect 88192 86468 88196 86524
rect 88196 86468 88252 86524
rect 88252 86468 88256 86524
rect 88192 86464 88256 86468
rect 1952 85980 2016 85984
rect 1952 85924 1956 85980
rect 1956 85924 2012 85980
rect 2012 85924 2016 85980
rect 1952 85920 2016 85924
rect 2032 85980 2096 85984
rect 2032 85924 2036 85980
rect 2036 85924 2092 85980
rect 2092 85924 2096 85980
rect 2032 85920 2096 85924
rect 2112 85980 2176 85984
rect 2112 85924 2116 85980
rect 2116 85924 2172 85980
rect 2172 85924 2176 85980
rect 2112 85920 2176 85924
rect 2192 85980 2256 85984
rect 2192 85924 2196 85980
rect 2196 85924 2252 85980
rect 2252 85924 2256 85980
rect 2192 85920 2256 85924
rect 85952 85980 86016 85984
rect 85952 85924 85956 85980
rect 85956 85924 86012 85980
rect 86012 85924 86016 85980
rect 85952 85920 86016 85924
rect 86032 85980 86096 85984
rect 86032 85924 86036 85980
rect 86036 85924 86092 85980
rect 86092 85924 86096 85980
rect 86032 85920 86096 85924
rect 86112 85980 86176 85984
rect 86112 85924 86116 85980
rect 86116 85924 86172 85980
rect 86172 85924 86176 85980
rect 86112 85920 86176 85924
rect 86192 85980 86256 85984
rect 86192 85924 86196 85980
rect 86196 85924 86252 85980
rect 86252 85924 86256 85980
rect 86192 85920 86256 85924
rect 89952 85980 90016 85984
rect 89952 85924 89956 85980
rect 89956 85924 90012 85980
rect 90012 85924 90016 85980
rect 89952 85920 90016 85924
rect 90032 85980 90096 85984
rect 90032 85924 90036 85980
rect 90036 85924 90092 85980
rect 90092 85924 90096 85980
rect 90032 85920 90096 85924
rect 90112 85980 90176 85984
rect 90112 85924 90116 85980
rect 90116 85924 90172 85980
rect 90172 85924 90176 85980
rect 90112 85920 90176 85924
rect 90192 85980 90256 85984
rect 90192 85924 90196 85980
rect 90196 85924 90252 85980
rect 90252 85924 90256 85980
rect 90192 85920 90256 85924
rect 3952 85436 4016 85440
rect 3952 85380 3956 85436
rect 3956 85380 4012 85436
rect 4012 85380 4016 85436
rect 3952 85376 4016 85380
rect 4032 85436 4096 85440
rect 4032 85380 4036 85436
rect 4036 85380 4092 85436
rect 4092 85380 4096 85436
rect 4032 85376 4096 85380
rect 4112 85436 4176 85440
rect 4112 85380 4116 85436
rect 4116 85380 4172 85436
rect 4172 85380 4176 85436
rect 4112 85376 4176 85380
rect 4192 85436 4256 85440
rect 4192 85380 4196 85436
rect 4196 85380 4252 85436
rect 4252 85380 4256 85436
rect 4192 85376 4256 85380
rect 87952 85436 88016 85440
rect 87952 85380 87956 85436
rect 87956 85380 88012 85436
rect 88012 85380 88016 85436
rect 87952 85376 88016 85380
rect 88032 85436 88096 85440
rect 88032 85380 88036 85436
rect 88036 85380 88092 85436
rect 88092 85380 88096 85436
rect 88032 85376 88096 85380
rect 88112 85436 88176 85440
rect 88112 85380 88116 85436
rect 88116 85380 88172 85436
rect 88172 85380 88176 85436
rect 88112 85376 88176 85380
rect 88192 85436 88256 85440
rect 88192 85380 88196 85436
rect 88196 85380 88252 85436
rect 88252 85380 88256 85436
rect 88192 85376 88256 85380
rect 1952 84892 2016 84896
rect 1952 84836 1956 84892
rect 1956 84836 2012 84892
rect 2012 84836 2016 84892
rect 1952 84832 2016 84836
rect 2032 84892 2096 84896
rect 2032 84836 2036 84892
rect 2036 84836 2092 84892
rect 2092 84836 2096 84892
rect 2032 84832 2096 84836
rect 2112 84892 2176 84896
rect 2112 84836 2116 84892
rect 2116 84836 2172 84892
rect 2172 84836 2176 84892
rect 2112 84832 2176 84836
rect 2192 84892 2256 84896
rect 2192 84836 2196 84892
rect 2196 84836 2252 84892
rect 2252 84836 2256 84892
rect 2192 84832 2256 84836
rect 85952 84892 86016 84896
rect 85952 84836 85956 84892
rect 85956 84836 86012 84892
rect 86012 84836 86016 84892
rect 85952 84832 86016 84836
rect 86032 84892 86096 84896
rect 86032 84836 86036 84892
rect 86036 84836 86092 84892
rect 86092 84836 86096 84892
rect 86032 84832 86096 84836
rect 86112 84892 86176 84896
rect 86112 84836 86116 84892
rect 86116 84836 86172 84892
rect 86172 84836 86176 84892
rect 86112 84832 86176 84836
rect 86192 84892 86256 84896
rect 86192 84836 86196 84892
rect 86196 84836 86252 84892
rect 86252 84836 86256 84892
rect 86192 84832 86256 84836
rect 89952 84892 90016 84896
rect 89952 84836 89956 84892
rect 89956 84836 90012 84892
rect 90012 84836 90016 84892
rect 89952 84832 90016 84836
rect 90032 84892 90096 84896
rect 90032 84836 90036 84892
rect 90036 84836 90092 84892
rect 90092 84836 90096 84892
rect 90032 84832 90096 84836
rect 90112 84892 90176 84896
rect 90112 84836 90116 84892
rect 90116 84836 90172 84892
rect 90172 84836 90176 84892
rect 90112 84832 90176 84836
rect 90192 84892 90256 84896
rect 90192 84836 90196 84892
rect 90196 84836 90252 84892
rect 90252 84836 90256 84892
rect 90192 84832 90256 84836
rect 3952 84348 4016 84352
rect 3952 84292 3956 84348
rect 3956 84292 4012 84348
rect 4012 84292 4016 84348
rect 3952 84288 4016 84292
rect 4032 84348 4096 84352
rect 4032 84292 4036 84348
rect 4036 84292 4092 84348
rect 4092 84292 4096 84348
rect 4032 84288 4096 84292
rect 4112 84348 4176 84352
rect 4112 84292 4116 84348
rect 4116 84292 4172 84348
rect 4172 84292 4176 84348
rect 4112 84288 4176 84292
rect 4192 84348 4256 84352
rect 4192 84292 4196 84348
rect 4196 84292 4252 84348
rect 4252 84292 4256 84348
rect 4192 84288 4256 84292
rect 87952 84348 88016 84352
rect 87952 84292 87956 84348
rect 87956 84292 88012 84348
rect 88012 84292 88016 84348
rect 87952 84288 88016 84292
rect 88032 84348 88096 84352
rect 88032 84292 88036 84348
rect 88036 84292 88092 84348
rect 88092 84292 88096 84348
rect 88032 84288 88096 84292
rect 88112 84348 88176 84352
rect 88112 84292 88116 84348
rect 88116 84292 88172 84348
rect 88172 84292 88176 84348
rect 88112 84288 88176 84292
rect 88192 84348 88256 84352
rect 88192 84292 88196 84348
rect 88196 84292 88252 84348
rect 88252 84292 88256 84348
rect 88192 84288 88256 84292
rect 1952 83804 2016 83808
rect 1952 83748 1956 83804
rect 1956 83748 2012 83804
rect 2012 83748 2016 83804
rect 1952 83744 2016 83748
rect 2032 83804 2096 83808
rect 2032 83748 2036 83804
rect 2036 83748 2092 83804
rect 2092 83748 2096 83804
rect 2032 83744 2096 83748
rect 2112 83804 2176 83808
rect 2112 83748 2116 83804
rect 2116 83748 2172 83804
rect 2172 83748 2176 83804
rect 2112 83744 2176 83748
rect 2192 83804 2256 83808
rect 2192 83748 2196 83804
rect 2196 83748 2252 83804
rect 2252 83748 2256 83804
rect 2192 83744 2256 83748
rect 85952 83804 86016 83808
rect 85952 83748 85956 83804
rect 85956 83748 86012 83804
rect 86012 83748 86016 83804
rect 85952 83744 86016 83748
rect 86032 83804 86096 83808
rect 86032 83748 86036 83804
rect 86036 83748 86092 83804
rect 86092 83748 86096 83804
rect 86032 83744 86096 83748
rect 86112 83804 86176 83808
rect 86112 83748 86116 83804
rect 86116 83748 86172 83804
rect 86172 83748 86176 83804
rect 86112 83744 86176 83748
rect 86192 83804 86256 83808
rect 86192 83748 86196 83804
rect 86196 83748 86252 83804
rect 86252 83748 86256 83804
rect 86192 83744 86256 83748
rect 89952 83804 90016 83808
rect 89952 83748 89956 83804
rect 89956 83748 90012 83804
rect 90012 83748 90016 83804
rect 89952 83744 90016 83748
rect 90032 83804 90096 83808
rect 90032 83748 90036 83804
rect 90036 83748 90092 83804
rect 90092 83748 90096 83804
rect 90032 83744 90096 83748
rect 90112 83804 90176 83808
rect 90112 83748 90116 83804
rect 90116 83748 90172 83804
rect 90172 83748 90176 83804
rect 90112 83744 90176 83748
rect 90192 83804 90256 83808
rect 90192 83748 90196 83804
rect 90196 83748 90252 83804
rect 90252 83748 90256 83804
rect 90192 83744 90256 83748
rect 3952 83260 4016 83264
rect 3952 83204 3956 83260
rect 3956 83204 4012 83260
rect 4012 83204 4016 83260
rect 3952 83200 4016 83204
rect 4032 83260 4096 83264
rect 4032 83204 4036 83260
rect 4036 83204 4092 83260
rect 4092 83204 4096 83260
rect 4032 83200 4096 83204
rect 4112 83260 4176 83264
rect 4112 83204 4116 83260
rect 4116 83204 4172 83260
rect 4172 83204 4176 83260
rect 4112 83200 4176 83204
rect 4192 83260 4256 83264
rect 4192 83204 4196 83260
rect 4196 83204 4252 83260
rect 4252 83204 4256 83260
rect 4192 83200 4256 83204
rect 87952 83260 88016 83264
rect 87952 83204 87956 83260
rect 87956 83204 88012 83260
rect 88012 83204 88016 83260
rect 87952 83200 88016 83204
rect 88032 83260 88096 83264
rect 88032 83204 88036 83260
rect 88036 83204 88092 83260
rect 88092 83204 88096 83260
rect 88032 83200 88096 83204
rect 88112 83260 88176 83264
rect 88112 83204 88116 83260
rect 88116 83204 88172 83260
rect 88172 83204 88176 83260
rect 88112 83200 88176 83204
rect 88192 83260 88256 83264
rect 88192 83204 88196 83260
rect 88196 83204 88252 83260
rect 88252 83204 88256 83260
rect 88192 83200 88256 83204
rect 1952 82716 2016 82720
rect 1952 82660 1956 82716
rect 1956 82660 2012 82716
rect 2012 82660 2016 82716
rect 1952 82656 2016 82660
rect 2032 82716 2096 82720
rect 2032 82660 2036 82716
rect 2036 82660 2092 82716
rect 2092 82660 2096 82716
rect 2032 82656 2096 82660
rect 2112 82716 2176 82720
rect 2112 82660 2116 82716
rect 2116 82660 2172 82716
rect 2172 82660 2176 82716
rect 2112 82656 2176 82660
rect 2192 82716 2256 82720
rect 2192 82660 2196 82716
rect 2196 82660 2252 82716
rect 2252 82660 2256 82716
rect 2192 82656 2256 82660
rect 85952 82716 86016 82720
rect 85952 82660 85956 82716
rect 85956 82660 86012 82716
rect 86012 82660 86016 82716
rect 85952 82656 86016 82660
rect 86032 82716 86096 82720
rect 86032 82660 86036 82716
rect 86036 82660 86092 82716
rect 86092 82660 86096 82716
rect 86032 82656 86096 82660
rect 86112 82716 86176 82720
rect 86112 82660 86116 82716
rect 86116 82660 86172 82716
rect 86172 82660 86176 82716
rect 86112 82656 86176 82660
rect 86192 82716 86256 82720
rect 86192 82660 86196 82716
rect 86196 82660 86252 82716
rect 86252 82660 86256 82716
rect 86192 82656 86256 82660
rect 89952 82716 90016 82720
rect 89952 82660 89956 82716
rect 89956 82660 90012 82716
rect 90012 82660 90016 82716
rect 89952 82656 90016 82660
rect 90032 82716 90096 82720
rect 90032 82660 90036 82716
rect 90036 82660 90092 82716
rect 90092 82660 90096 82716
rect 90032 82656 90096 82660
rect 90112 82716 90176 82720
rect 90112 82660 90116 82716
rect 90116 82660 90172 82716
rect 90172 82660 90176 82716
rect 90112 82656 90176 82660
rect 90192 82716 90256 82720
rect 90192 82660 90196 82716
rect 90196 82660 90252 82716
rect 90252 82660 90256 82716
rect 90192 82656 90256 82660
rect 3952 82172 4016 82176
rect 3952 82116 3956 82172
rect 3956 82116 4012 82172
rect 4012 82116 4016 82172
rect 3952 82112 4016 82116
rect 4032 82172 4096 82176
rect 4032 82116 4036 82172
rect 4036 82116 4092 82172
rect 4092 82116 4096 82172
rect 4032 82112 4096 82116
rect 4112 82172 4176 82176
rect 4112 82116 4116 82172
rect 4116 82116 4172 82172
rect 4172 82116 4176 82172
rect 4112 82112 4176 82116
rect 4192 82172 4256 82176
rect 4192 82116 4196 82172
rect 4196 82116 4252 82172
rect 4252 82116 4256 82172
rect 4192 82112 4256 82116
rect 87952 82172 88016 82176
rect 87952 82116 87956 82172
rect 87956 82116 88012 82172
rect 88012 82116 88016 82172
rect 87952 82112 88016 82116
rect 88032 82172 88096 82176
rect 88032 82116 88036 82172
rect 88036 82116 88092 82172
rect 88092 82116 88096 82172
rect 88032 82112 88096 82116
rect 88112 82172 88176 82176
rect 88112 82116 88116 82172
rect 88116 82116 88172 82172
rect 88172 82116 88176 82172
rect 88112 82112 88176 82116
rect 88192 82172 88256 82176
rect 88192 82116 88196 82172
rect 88196 82116 88252 82172
rect 88252 82116 88256 82172
rect 88192 82112 88256 82116
rect 1952 81628 2016 81632
rect 1952 81572 1956 81628
rect 1956 81572 2012 81628
rect 2012 81572 2016 81628
rect 1952 81568 2016 81572
rect 2032 81628 2096 81632
rect 2032 81572 2036 81628
rect 2036 81572 2092 81628
rect 2092 81572 2096 81628
rect 2032 81568 2096 81572
rect 2112 81628 2176 81632
rect 2112 81572 2116 81628
rect 2116 81572 2172 81628
rect 2172 81572 2176 81628
rect 2112 81568 2176 81572
rect 2192 81628 2256 81632
rect 2192 81572 2196 81628
rect 2196 81572 2252 81628
rect 2252 81572 2256 81628
rect 2192 81568 2256 81572
rect 85952 81628 86016 81632
rect 85952 81572 85956 81628
rect 85956 81572 86012 81628
rect 86012 81572 86016 81628
rect 85952 81568 86016 81572
rect 86032 81628 86096 81632
rect 86032 81572 86036 81628
rect 86036 81572 86092 81628
rect 86092 81572 86096 81628
rect 86032 81568 86096 81572
rect 86112 81628 86176 81632
rect 86112 81572 86116 81628
rect 86116 81572 86172 81628
rect 86172 81572 86176 81628
rect 86112 81568 86176 81572
rect 86192 81628 86256 81632
rect 86192 81572 86196 81628
rect 86196 81572 86252 81628
rect 86252 81572 86256 81628
rect 86192 81568 86256 81572
rect 89952 81628 90016 81632
rect 89952 81572 89956 81628
rect 89956 81572 90012 81628
rect 90012 81572 90016 81628
rect 89952 81568 90016 81572
rect 90032 81628 90096 81632
rect 90032 81572 90036 81628
rect 90036 81572 90092 81628
rect 90092 81572 90096 81628
rect 90032 81568 90096 81572
rect 90112 81628 90176 81632
rect 90112 81572 90116 81628
rect 90116 81572 90172 81628
rect 90172 81572 90176 81628
rect 90112 81568 90176 81572
rect 90192 81628 90256 81632
rect 90192 81572 90196 81628
rect 90196 81572 90252 81628
rect 90252 81572 90256 81628
rect 90192 81568 90256 81572
rect 3952 81084 4016 81088
rect 3952 81028 3956 81084
rect 3956 81028 4012 81084
rect 4012 81028 4016 81084
rect 3952 81024 4016 81028
rect 4032 81084 4096 81088
rect 4032 81028 4036 81084
rect 4036 81028 4092 81084
rect 4092 81028 4096 81084
rect 4032 81024 4096 81028
rect 4112 81084 4176 81088
rect 4112 81028 4116 81084
rect 4116 81028 4172 81084
rect 4172 81028 4176 81084
rect 4112 81024 4176 81028
rect 4192 81084 4256 81088
rect 4192 81028 4196 81084
rect 4196 81028 4252 81084
rect 4252 81028 4256 81084
rect 4192 81024 4256 81028
rect 87952 81084 88016 81088
rect 87952 81028 87956 81084
rect 87956 81028 88012 81084
rect 88012 81028 88016 81084
rect 87952 81024 88016 81028
rect 88032 81084 88096 81088
rect 88032 81028 88036 81084
rect 88036 81028 88092 81084
rect 88092 81028 88096 81084
rect 88032 81024 88096 81028
rect 88112 81084 88176 81088
rect 88112 81028 88116 81084
rect 88116 81028 88172 81084
rect 88172 81028 88176 81084
rect 88112 81024 88176 81028
rect 88192 81084 88256 81088
rect 88192 81028 88196 81084
rect 88196 81028 88252 81084
rect 88252 81028 88256 81084
rect 88192 81024 88256 81028
rect 1952 80540 2016 80544
rect 1952 80484 1956 80540
rect 1956 80484 2012 80540
rect 2012 80484 2016 80540
rect 1952 80480 2016 80484
rect 2032 80540 2096 80544
rect 2032 80484 2036 80540
rect 2036 80484 2092 80540
rect 2092 80484 2096 80540
rect 2032 80480 2096 80484
rect 2112 80540 2176 80544
rect 2112 80484 2116 80540
rect 2116 80484 2172 80540
rect 2172 80484 2176 80540
rect 2112 80480 2176 80484
rect 2192 80540 2256 80544
rect 2192 80484 2196 80540
rect 2196 80484 2252 80540
rect 2252 80484 2256 80540
rect 2192 80480 2256 80484
rect 85952 80540 86016 80544
rect 85952 80484 85956 80540
rect 85956 80484 86012 80540
rect 86012 80484 86016 80540
rect 85952 80480 86016 80484
rect 86032 80540 86096 80544
rect 86032 80484 86036 80540
rect 86036 80484 86092 80540
rect 86092 80484 86096 80540
rect 86032 80480 86096 80484
rect 86112 80540 86176 80544
rect 86112 80484 86116 80540
rect 86116 80484 86172 80540
rect 86172 80484 86176 80540
rect 86112 80480 86176 80484
rect 86192 80540 86256 80544
rect 86192 80484 86196 80540
rect 86196 80484 86252 80540
rect 86252 80484 86256 80540
rect 86192 80480 86256 80484
rect 89952 80540 90016 80544
rect 89952 80484 89956 80540
rect 89956 80484 90012 80540
rect 90012 80484 90016 80540
rect 89952 80480 90016 80484
rect 90032 80540 90096 80544
rect 90032 80484 90036 80540
rect 90036 80484 90092 80540
rect 90092 80484 90096 80540
rect 90032 80480 90096 80484
rect 90112 80540 90176 80544
rect 90112 80484 90116 80540
rect 90116 80484 90172 80540
rect 90172 80484 90176 80540
rect 90112 80480 90176 80484
rect 90192 80540 90256 80544
rect 90192 80484 90196 80540
rect 90196 80484 90252 80540
rect 90252 80484 90256 80540
rect 90192 80480 90256 80484
rect 3952 79996 4016 80000
rect 3952 79940 3956 79996
rect 3956 79940 4012 79996
rect 4012 79940 4016 79996
rect 3952 79936 4016 79940
rect 4032 79996 4096 80000
rect 4032 79940 4036 79996
rect 4036 79940 4092 79996
rect 4092 79940 4096 79996
rect 4032 79936 4096 79940
rect 4112 79996 4176 80000
rect 4112 79940 4116 79996
rect 4116 79940 4172 79996
rect 4172 79940 4176 79996
rect 4112 79936 4176 79940
rect 4192 79996 4256 80000
rect 4192 79940 4196 79996
rect 4196 79940 4252 79996
rect 4252 79940 4256 79996
rect 4192 79936 4256 79940
rect 87952 79996 88016 80000
rect 87952 79940 87956 79996
rect 87956 79940 88012 79996
rect 88012 79940 88016 79996
rect 87952 79936 88016 79940
rect 88032 79996 88096 80000
rect 88032 79940 88036 79996
rect 88036 79940 88092 79996
rect 88092 79940 88096 79996
rect 88032 79936 88096 79940
rect 88112 79996 88176 80000
rect 88112 79940 88116 79996
rect 88116 79940 88172 79996
rect 88172 79940 88176 79996
rect 88112 79936 88176 79940
rect 88192 79996 88256 80000
rect 88192 79940 88196 79996
rect 88196 79940 88252 79996
rect 88252 79940 88256 79996
rect 88192 79936 88256 79940
rect 1952 79452 2016 79456
rect 1952 79396 1956 79452
rect 1956 79396 2012 79452
rect 2012 79396 2016 79452
rect 1952 79392 2016 79396
rect 2032 79452 2096 79456
rect 2032 79396 2036 79452
rect 2036 79396 2092 79452
rect 2092 79396 2096 79452
rect 2032 79392 2096 79396
rect 2112 79452 2176 79456
rect 2112 79396 2116 79452
rect 2116 79396 2172 79452
rect 2172 79396 2176 79452
rect 2112 79392 2176 79396
rect 2192 79452 2256 79456
rect 2192 79396 2196 79452
rect 2196 79396 2252 79452
rect 2252 79396 2256 79452
rect 2192 79392 2256 79396
rect 85952 79452 86016 79456
rect 85952 79396 85956 79452
rect 85956 79396 86012 79452
rect 86012 79396 86016 79452
rect 85952 79392 86016 79396
rect 86032 79452 86096 79456
rect 86032 79396 86036 79452
rect 86036 79396 86092 79452
rect 86092 79396 86096 79452
rect 86032 79392 86096 79396
rect 86112 79452 86176 79456
rect 86112 79396 86116 79452
rect 86116 79396 86172 79452
rect 86172 79396 86176 79452
rect 86112 79392 86176 79396
rect 86192 79452 86256 79456
rect 86192 79396 86196 79452
rect 86196 79396 86252 79452
rect 86252 79396 86256 79452
rect 86192 79392 86256 79396
rect 89952 79452 90016 79456
rect 89952 79396 89956 79452
rect 89956 79396 90012 79452
rect 90012 79396 90016 79452
rect 89952 79392 90016 79396
rect 90032 79452 90096 79456
rect 90032 79396 90036 79452
rect 90036 79396 90092 79452
rect 90092 79396 90096 79452
rect 90032 79392 90096 79396
rect 90112 79452 90176 79456
rect 90112 79396 90116 79452
rect 90116 79396 90172 79452
rect 90172 79396 90176 79452
rect 90112 79392 90176 79396
rect 90192 79452 90256 79456
rect 90192 79396 90196 79452
rect 90196 79396 90252 79452
rect 90252 79396 90256 79452
rect 90192 79392 90256 79396
rect 3952 78908 4016 78912
rect 3952 78852 3956 78908
rect 3956 78852 4012 78908
rect 4012 78852 4016 78908
rect 3952 78848 4016 78852
rect 4032 78908 4096 78912
rect 4032 78852 4036 78908
rect 4036 78852 4092 78908
rect 4092 78852 4096 78908
rect 4032 78848 4096 78852
rect 4112 78908 4176 78912
rect 4112 78852 4116 78908
rect 4116 78852 4172 78908
rect 4172 78852 4176 78908
rect 4112 78848 4176 78852
rect 4192 78908 4256 78912
rect 4192 78852 4196 78908
rect 4196 78852 4252 78908
rect 4252 78852 4256 78908
rect 4192 78848 4256 78852
rect 87952 78908 88016 78912
rect 87952 78852 87956 78908
rect 87956 78852 88012 78908
rect 88012 78852 88016 78908
rect 87952 78848 88016 78852
rect 88032 78908 88096 78912
rect 88032 78852 88036 78908
rect 88036 78852 88092 78908
rect 88092 78852 88096 78908
rect 88032 78848 88096 78852
rect 88112 78908 88176 78912
rect 88112 78852 88116 78908
rect 88116 78852 88172 78908
rect 88172 78852 88176 78908
rect 88112 78848 88176 78852
rect 88192 78908 88256 78912
rect 88192 78852 88196 78908
rect 88196 78852 88252 78908
rect 88252 78852 88256 78908
rect 88192 78848 88256 78852
rect 1952 78364 2016 78368
rect 1952 78308 1956 78364
rect 1956 78308 2012 78364
rect 2012 78308 2016 78364
rect 1952 78304 2016 78308
rect 2032 78364 2096 78368
rect 2032 78308 2036 78364
rect 2036 78308 2092 78364
rect 2092 78308 2096 78364
rect 2032 78304 2096 78308
rect 2112 78364 2176 78368
rect 2112 78308 2116 78364
rect 2116 78308 2172 78364
rect 2172 78308 2176 78364
rect 2112 78304 2176 78308
rect 2192 78364 2256 78368
rect 2192 78308 2196 78364
rect 2196 78308 2252 78364
rect 2252 78308 2256 78364
rect 2192 78304 2256 78308
rect 85952 78364 86016 78368
rect 85952 78308 85956 78364
rect 85956 78308 86012 78364
rect 86012 78308 86016 78364
rect 85952 78304 86016 78308
rect 86032 78364 86096 78368
rect 86032 78308 86036 78364
rect 86036 78308 86092 78364
rect 86092 78308 86096 78364
rect 86032 78304 86096 78308
rect 86112 78364 86176 78368
rect 86112 78308 86116 78364
rect 86116 78308 86172 78364
rect 86172 78308 86176 78364
rect 86112 78304 86176 78308
rect 86192 78364 86256 78368
rect 86192 78308 86196 78364
rect 86196 78308 86252 78364
rect 86252 78308 86256 78364
rect 86192 78304 86256 78308
rect 89952 78364 90016 78368
rect 89952 78308 89956 78364
rect 89956 78308 90012 78364
rect 90012 78308 90016 78364
rect 89952 78304 90016 78308
rect 90032 78364 90096 78368
rect 90032 78308 90036 78364
rect 90036 78308 90092 78364
rect 90092 78308 90096 78364
rect 90032 78304 90096 78308
rect 90112 78364 90176 78368
rect 90112 78308 90116 78364
rect 90116 78308 90172 78364
rect 90172 78308 90176 78364
rect 90112 78304 90176 78308
rect 90192 78364 90256 78368
rect 90192 78308 90196 78364
rect 90196 78308 90252 78364
rect 90252 78308 90256 78364
rect 90192 78304 90256 78308
rect 3952 77820 4016 77824
rect 3952 77764 3956 77820
rect 3956 77764 4012 77820
rect 4012 77764 4016 77820
rect 3952 77760 4016 77764
rect 4032 77820 4096 77824
rect 4032 77764 4036 77820
rect 4036 77764 4092 77820
rect 4092 77764 4096 77820
rect 4032 77760 4096 77764
rect 4112 77820 4176 77824
rect 4112 77764 4116 77820
rect 4116 77764 4172 77820
rect 4172 77764 4176 77820
rect 4112 77760 4176 77764
rect 4192 77820 4256 77824
rect 4192 77764 4196 77820
rect 4196 77764 4252 77820
rect 4252 77764 4256 77820
rect 4192 77760 4256 77764
rect 87952 77820 88016 77824
rect 87952 77764 87956 77820
rect 87956 77764 88012 77820
rect 88012 77764 88016 77820
rect 87952 77760 88016 77764
rect 88032 77820 88096 77824
rect 88032 77764 88036 77820
rect 88036 77764 88092 77820
rect 88092 77764 88096 77820
rect 88032 77760 88096 77764
rect 88112 77820 88176 77824
rect 88112 77764 88116 77820
rect 88116 77764 88172 77820
rect 88172 77764 88176 77820
rect 88112 77760 88176 77764
rect 88192 77820 88256 77824
rect 88192 77764 88196 77820
rect 88196 77764 88252 77820
rect 88252 77764 88256 77820
rect 88192 77760 88256 77764
rect 1952 77276 2016 77280
rect 1952 77220 1956 77276
rect 1956 77220 2012 77276
rect 2012 77220 2016 77276
rect 1952 77216 2016 77220
rect 2032 77276 2096 77280
rect 2032 77220 2036 77276
rect 2036 77220 2092 77276
rect 2092 77220 2096 77276
rect 2032 77216 2096 77220
rect 2112 77276 2176 77280
rect 2112 77220 2116 77276
rect 2116 77220 2172 77276
rect 2172 77220 2176 77276
rect 2112 77216 2176 77220
rect 2192 77276 2256 77280
rect 2192 77220 2196 77276
rect 2196 77220 2252 77276
rect 2252 77220 2256 77276
rect 2192 77216 2256 77220
rect 85952 77276 86016 77280
rect 85952 77220 85956 77276
rect 85956 77220 86012 77276
rect 86012 77220 86016 77276
rect 85952 77216 86016 77220
rect 86032 77276 86096 77280
rect 86032 77220 86036 77276
rect 86036 77220 86092 77276
rect 86092 77220 86096 77276
rect 86032 77216 86096 77220
rect 86112 77276 86176 77280
rect 86112 77220 86116 77276
rect 86116 77220 86172 77276
rect 86172 77220 86176 77276
rect 86112 77216 86176 77220
rect 86192 77276 86256 77280
rect 86192 77220 86196 77276
rect 86196 77220 86252 77276
rect 86252 77220 86256 77276
rect 86192 77216 86256 77220
rect 89952 77276 90016 77280
rect 89952 77220 89956 77276
rect 89956 77220 90012 77276
rect 90012 77220 90016 77276
rect 89952 77216 90016 77220
rect 90032 77276 90096 77280
rect 90032 77220 90036 77276
rect 90036 77220 90092 77276
rect 90092 77220 90096 77276
rect 90032 77216 90096 77220
rect 90112 77276 90176 77280
rect 90112 77220 90116 77276
rect 90116 77220 90172 77276
rect 90172 77220 90176 77276
rect 90112 77216 90176 77220
rect 90192 77276 90256 77280
rect 90192 77220 90196 77276
rect 90196 77220 90252 77276
rect 90252 77220 90256 77276
rect 90192 77216 90256 77220
rect 3952 76732 4016 76736
rect 3952 76676 3956 76732
rect 3956 76676 4012 76732
rect 4012 76676 4016 76732
rect 3952 76672 4016 76676
rect 4032 76732 4096 76736
rect 4032 76676 4036 76732
rect 4036 76676 4092 76732
rect 4092 76676 4096 76732
rect 4032 76672 4096 76676
rect 4112 76732 4176 76736
rect 4112 76676 4116 76732
rect 4116 76676 4172 76732
rect 4172 76676 4176 76732
rect 4112 76672 4176 76676
rect 4192 76732 4256 76736
rect 4192 76676 4196 76732
rect 4196 76676 4252 76732
rect 4252 76676 4256 76732
rect 4192 76672 4256 76676
rect 87952 76732 88016 76736
rect 87952 76676 87956 76732
rect 87956 76676 88012 76732
rect 88012 76676 88016 76732
rect 87952 76672 88016 76676
rect 88032 76732 88096 76736
rect 88032 76676 88036 76732
rect 88036 76676 88092 76732
rect 88092 76676 88096 76732
rect 88032 76672 88096 76676
rect 88112 76732 88176 76736
rect 88112 76676 88116 76732
rect 88116 76676 88172 76732
rect 88172 76676 88176 76732
rect 88112 76672 88176 76676
rect 88192 76732 88256 76736
rect 88192 76676 88196 76732
rect 88196 76676 88252 76732
rect 88252 76676 88256 76732
rect 88192 76672 88256 76676
rect 1952 76188 2016 76192
rect 1952 76132 1956 76188
rect 1956 76132 2012 76188
rect 2012 76132 2016 76188
rect 1952 76128 2016 76132
rect 2032 76188 2096 76192
rect 2032 76132 2036 76188
rect 2036 76132 2092 76188
rect 2092 76132 2096 76188
rect 2032 76128 2096 76132
rect 2112 76188 2176 76192
rect 2112 76132 2116 76188
rect 2116 76132 2172 76188
rect 2172 76132 2176 76188
rect 2112 76128 2176 76132
rect 2192 76188 2256 76192
rect 2192 76132 2196 76188
rect 2196 76132 2252 76188
rect 2252 76132 2256 76188
rect 2192 76128 2256 76132
rect 85952 76188 86016 76192
rect 85952 76132 85956 76188
rect 85956 76132 86012 76188
rect 86012 76132 86016 76188
rect 85952 76128 86016 76132
rect 86032 76188 86096 76192
rect 86032 76132 86036 76188
rect 86036 76132 86092 76188
rect 86092 76132 86096 76188
rect 86032 76128 86096 76132
rect 86112 76188 86176 76192
rect 86112 76132 86116 76188
rect 86116 76132 86172 76188
rect 86172 76132 86176 76188
rect 86112 76128 86176 76132
rect 86192 76188 86256 76192
rect 86192 76132 86196 76188
rect 86196 76132 86252 76188
rect 86252 76132 86256 76188
rect 86192 76128 86256 76132
rect 89952 76188 90016 76192
rect 89952 76132 89956 76188
rect 89956 76132 90012 76188
rect 90012 76132 90016 76188
rect 89952 76128 90016 76132
rect 90032 76188 90096 76192
rect 90032 76132 90036 76188
rect 90036 76132 90092 76188
rect 90092 76132 90096 76188
rect 90032 76128 90096 76132
rect 90112 76188 90176 76192
rect 90112 76132 90116 76188
rect 90116 76132 90172 76188
rect 90172 76132 90176 76188
rect 90112 76128 90176 76132
rect 90192 76188 90256 76192
rect 90192 76132 90196 76188
rect 90196 76132 90252 76188
rect 90252 76132 90256 76188
rect 90192 76128 90256 76132
rect 3952 75644 4016 75648
rect 3952 75588 3956 75644
rect 3956 75588 4012 75644
rect 4012 75588 4016 75644
rect 3952 75584 4016 75588
rect 4032 75644 4096 75648
rect 4032 75588 4036 75644
rect 4036 75588 4092 75644
rect 4092 75588 4096 75644
rect 4032 75584 4096 75588
rect 4112 75644 4176 75648
rect 4112 75588 4116 75644
rect 4116 75588 4172 75644
rect 4172 75588 4176 75644
rect 4112 75584 4176 75588
rect 4192 75644 4256 75648
rect 4192 75588 4196 75644
rect 4196 75588 4252 75644
rect 4252 75588 4256 75644
rect 4192 75584 4256 75588
rect 87952 75644 88016 75648
rect 87952 75588 87956 75644
rect 87956 75588 88012 75644
rect 88012 75588 88016 75644
rect 87952 75584 88016 75588
rect 88032 75644 88096 75648
rect 88032 75588 88036 75644
rect 88036 75588 88092 75644
rect 88092 75588 88096 75644
rect 88032 75584 88096 75588
rect 88112 75644 88176 75648
rect 88112 75588 88116 75644
rect 88116 75588 88172 75644
rect 88172 75588 88176 75644
rect 88112 75584 88176 75588
rect 88192 75644 88256 75648
rect 88192 75588 88196 75644
rect 88196 75588 88252 75644
rect 88252 75588 88256 75644
rect 88192 75584 88256 75588
rect 1952 75100 2016 75104
rect 1952 75044 1956 75100
rect 1956 75044 2012 75100
rect 2012 75044 2016 75100
rect 1952 75040 2016 75044
rect 2032 75100 2096 75104
rect 2032 75044 2036 75100
rect 2036 75044 2092 75100
rect 2092 75044 2096 75100
rect 2032 75040 2096 75044
rect 2112 75100 2176 75104
rect 2112 75044 2116 75100
rect 2116 75044 2172 75100
rect 2172 75044 2176 75100
rect 2112 75040 2176 75044
rect 2192 75100 2256 75104
rect 2192 75044 2196 75100
rect 2196 75044 2252 75100
rect 2252 75044 2256 75100
rect 2192 75040 2256 75044
rect 85952 75100 86016 75104
rect 85952 75044 85956 75100
rect 85956 75044 86012 75100
rect 86012 75044 86016 75100
rect 85952 75040 86016 75044
rect 86032 75100 86096 75104
rect 86032 75044 86036 75100
rect 86036 75044 86092 75100
rect 86092 75044 86096 75100
rect 86032 75040 86096 75044
rect 86112 75100 86176 75104
rect 86112 75044 86116 75100
rect 86116 75044 86172 75100
rect 86172 75044 86176 75100
rect 86112 75040 86176 75044
rect 86192 75100 86256 75104
rect 86192 75044 86196 75100
rect 86196 75044 86252 75100
rect 86252 75044 86256 75100
rect 86192 75040 86256 75044
rect 89952 75100 90016 75104
rect 89952 75044 89956 75100
rect 89956 75044 90012 75100
rect 90012 75044 90016 75100
rect 89952 75040 90016 75044
rect 90032 75100 90096 75104
rect 90032 75044 90036 75100
rect 90036 75044 90092 75100
rect 90092 75044 90096 75100
rect 90032 75040 90096 75044
rect 90112 75100 90176 75104
rect 90112 75044 90116 75100
rect 90116 75044 90172 75100
rect 90172 75044 90176 75100
rect 90112 75040 90176 75044
rect 90192 75100 90256 75104
rect 90192 75044 90196 75100
rect 90196 75044 90252 75100
rect 90252 75044 90256 75100
rect 90192 75040 90256 75044
rect 3952 74556 4016 74560
rect 3952 74500 3956 74556
rect 3956 74500 4012 74556
rect 4012 74500 4016 74556
rect 3952 74496 4016 74500
rect 4032 74556 4096 74560
rect 4032 74500 4036 74556
rect 4036 74500 4092 74556
rect 4092 74500 4096 74556
rect 4032 74496 4096 74500
rect 4112 74556 4176 74560
rect 4112 74500 4116 74556
rect 4116 74500 4172 74556
rect 4172 74500 4176 74556
rect 4112 74496 4176 74500
rect 4192 74556 4256 74560
rect 4192 74500 4196 74556
rect 4196 74500 4252 74556
rect 4252 74500 4256 74556
rect 4192 74496 4256 74500
rect 87952 74556 88016 74560
rect 87952 74500 87956 74556
rect 87956 74500 88012 74556
rect 88012 74500 88016 74556
rect 87952 74496 88016 74500
rect 88032 74556 88096 74560
rect 88032 74500 88036 74556
rect 88036 74500 88092 74556
rect 88092 74500 88096 74556
rect 88032 74496 88096 74500
rect 88112 74556 88176 74560
rect 88112 74500 88116 74556
rect 88116 74500 88172 74556
rect 88172 74500 88176 74556
rect 88112 74496 88176 74500
rect 88192 74556 88256 74560
rect 88192 74500 88196 74556
rect 88196 74500 88252 74556
rect 88252 74500 88256 74556
rect 88192 74496 88256 74500
rect 1952 74012 2016 74016
rect 1952 73956 1956 74012
rect 1956 73956 2012 74012
rect 2012 73956 2016 74012
rect 1952 73952 2016 73956
rect 2032 74012 2096 74016
rect 2032 73956 2036 74012
rect 2036 73956 2092 74012
rect 2092 73956 2096 74012
rect 2032 73952 2096 73956
rect 2112 74012 2176 74016
rect 2112 73956 2116 74012
rect 2116 73956 2172 74012
rect 2172 73956 2176 74012
rect 2112 73952 2176 73956
rect 2192 74012 2256 74016
rect 2192 73956 2196 74012
rect 2196 73956 2252 74012
rect 2252 73956 2256 74012
rect 2192 73952 2256 73956
rect 85952 74012 86016 74016
rect 85952 73956 85956 74012
rect 85956 73956 86012 74012
rect 86012 73956 86016 74012
rect 85952 73952 86016 73956
rect 86032 74012 86096 74016
rect 86032 73956 86036 74012
rect 86036 73956 86092 74012
rect 86092 73956 86096 74012
rect 86032 73952 86096 73956
rect 86112 74012 86176 74016
rect 86112 73956 86116 74012
rect 86116 73956 86172 74012
rect 86172 73956 86176 74012
rect 86112 73952 86176 73956
rect 86192 74012 86256 74016
rect 86192 73956 86196 74012
rect 86196 73956 86252 74012
rect 86252 73956 86256 74012
rect 86192 73952 86256 73956
rect 89952 74012 90016 74016
rect 89952 73956 89956 74012
rect 89956 73956 90012 74012
rect 90012 73956 90016 74012
rect 89952 73952 90016 73956
rect 90032 74012 90096 74016
rect 90032 73956 90036 74012
rect 90036 73956 90092 74012
rect 90092 73956 90096 74012
rect 90032 73952 90096 73956
rect 90112 74012 90176 74016
rect 90112 73956 90116 74012
rect 90116 73956 90172 74012
rect 90172 73956 90176 74012
rect 90112 73952 90176 73956
rect 90192 74012 90256 74016
rect 90192 73956 90196 74012
rect 90196 73956 90252 74012
rect 90252 73956 90256 74012
rect 90192 73952 90256 73956
rect 3952 73468 4016 73472
rect 3952 73412 3956 73468
rect 3956 73412 4012 73468
rect 4012 73412 4016 73468
rect 3952 73408 4016 73412
rect 4032 73468 4096 73472
rect 4032 73412 4036 73468
rect 4036 73412 4092 73468
rect 4092 73412 4096 73468
rect 4032 73408 4096 73412
rect 4112 73468 4176 73472
rect 4112 73412 4116 73468
rect 4116 73412 4172 73468
rect 4172 73412 4176 73468
rect 4112 73408 4176 73412
rect 4192 73468 4256 73472
rect 4192 73412 4196 73468
rect 4196 73412 4252 73468
rect 4252 73412 4256 73468
rect 4192 73408 4256 73412
rect 87952 73468 88016 73472
rect 87952 73412 87956 73468
rect 87956 73412 88012 73468
rect 88012 73412 88016 73468
rect 87952 73408 88016 73412
rect 88032 73468 88096 73472
rect 88032 73412 88036 73468
rect 88036 73412 88092 73468
rect 88092 73412 88096 73468
rect 88032 73408 88096 73412
rect 88112 73468 88176 73472
rect 88112 73412 88116 73468
rect 88116 73412 88172 73468
rect 88172 73412 88176 73468
rect 88112 73408 88176 73412
rect 88192 73468 88256 73472
rect 88192 73412 88196 73468
rect 88196 73412 88252 73468
rect 88252 73412 88256 73468
rect 88192 73408 88256 73412
rect 1952 72924 2016 72928
rect 1952 72868 1956 72924
rect 1956 72868 2012 72924
rect 2012 72868 2016 72924
rect 1952 72864 2016 72868
rect 2032 72924 2096 72928
rect 2032 72868 2036 72924
rect 2036 72868 2092 72924
rect 2092 72868 2096 72924
rect 2032 72864 2096 72868
rect 2112 72924 2176 72928
rect 2112 72868 2116 72924
rect 2116 72868 2172 72924
rect 2172 72868 2176 72924
rect 2112 72864 2176 72868
rect 2192 72924 2256 72928
rect 2192 72868 2196 72924
rect 2196 72868 2252 72924
rect 2252 72868 2256 72924
rect 2192 72864 2256 72868
rect 85952 72924 86016 72928
rect 85952 72868 85956 72924
rect 85956 72868 86012 72924
rect 86012 72868 86016 72924
rect 85952 72864 86016 72868
rect 86032 72924 86096 72928
rect 86032 72868 86036 72924
rect 86036 72868 86092 72924
rect 86092 72868 86096 72924
rect 86032 72864 86096 72868
rect 86112 72924 86176 72928
rect 86112 72868 86116 72924
rect 86116 72868 86172 72924
rect 86172 72868 86176 72924
rect 86112 72864 86176 72868
rect 86192 72924 86256 72928
rect 86192 72868 86196 72924
rect 86196 72868 86252 72924
rect 86252 72868 86256 72924
rect 86192 72864 86256 72868
rect 89952 72924 90016 72928
rect 89952 72868 89956 72924
rect 89956 72868 90012 72924
rect 90012 72868 90016 72924
rect 89952 72864 90016 72868
rect 90032 72924 90096 72928
rect 90032 72868 90036 72924
rect 90036 72868 90092 72924
rect 90092 72868 90096 72924
rect 90032 72864 90096 72868
rect 90112 72924 90176 72928
rect 90112 72868 90116 72924
rect 90116 72868 90172 72924
rect 90172 72868 90176 72924
rect 90112 72864 90176 72868
rect 90192 72924 90256 72928
rect 90192 72868 90196 72924
rect 90196 72868 90252 72924
rect 90252 72868 90256 72924
rect 90192 72864 90256 72868
rect 3952 72380 4016 72384
rect 3952 72324 3956 72380
rect 3956 72324 4012 72380
rect 4012 72324 4016 72380
rect 3952 72320 4016 72324
rect 4032 72380 4096 72384
rect 4032 72324 4036 72380
rect 4036 72324 4092 72380
rect 4092 72324 4096 72380
rect 4032 72320 4096 72324
rect 4112 72380 4176 72384
rect 4112 72324 4116 72380
rect 4116 72324 4172 72380
rect 4172 72324 4176 72380
rect 4112 72320 4176 72324
rect 4192 72380 4256 72384
rect 4192 72324 4196 72380
rect 4196 72324 4252 72380
rect 4252 72324 4256 72380
rect 4192 72320 4256 72324
rect 87952 72380 88016 72384
rect 87952 72324 87956 72380
rect 87956 72324 88012 72380
rect 88012 72324 88016 72380
rect 87952 72320 88016 72324
rect 88032 72380 88096 72384
rect 88032 72324 88036 72380
rect 88036 72324 88092 72380
rect 88092 72324 88096 72380
rect 88032 72320 88096 72324
rect 88112 72380 88176 72384
rect 88112 72324 88116 72380
rect 88116 72324 88172 72380
rect 88172 72324 88176 72380
rect 88112 72320 88176 72324
rect 88192 72380 88256 72384
rect 88192 72324 88196 72380
rect 88196 72324 88252 72380
rect 88252 72324 88256 72380
rect 88192 72320 88256 72324
rect 1952 71836 2016 71840
rect 1952 71780 1956 71836
rect 1956 71780 2012 71836
rect 2012 71780 2016 71836
rect 1952 71776 2016 71780
rect 2032 71836 2096 71840
rect 2032 71780 2036 71836
rect 2036 71780 2092 71836
rect 2092 71780 2096 71836
rect 2032 71776 2096 71780
rect 2112 71836 2176 71840
rect 2112 71780 2116 71836
rect 2116 71780 2172 71836
rect 2172 71780 2176 71836
rect 2112 71776 2176 71780
rect 2192 71836 2256 71840
rect 2192 71780 2196 71836
rect 2196 71780 2252 71836
rect 2252 71780 2256 71836
rect 2192 71776 2256 71780
rect 85952 71836 86016 71840
rect 85952 71780 85956 71836
rect 85956 71780 86012 71836
rect 86012 71780 86016 71836
rect 85952 71776 86016 71780
rect 86032 71836 86096 71840
rect 86032 71780 86036 71836
rect 86036 71780 86092 71836
rect 86092 71780 86096 71836
rect 86032 71776 86096 71780
rect 86112 71836 86176 71840
rect 86112 71780 86116 71836
rect 86116 71780 86172 71836
rect 86172 71780 86176 71836
rect 86112 71776 86176 71780
rect 86192 71836 86256 71840
rect 86192 71780 86196 71836
rect 86196 71780 86252 71836
rect 86252 71780 86256 71836
rect 86192 71776 86256 71780
rect 89952 71836 90016 71840
rect 89952 71780 89956 71836
rect 89956 71780 90012 71836
rect 90012 71780 90016 71836
rect 89952 71776 90016 71780
rect 90032 71836 90096 71840
rect 90032 71780 90036 71836
rect 90036 71780 90092 71836
rect 90092 71780 90096 71836
rect 90032 71776 90096 71780
rect 90112 71836 90176 71840
rect 90112 71780 90116 71836
rect 90116 71780 90172 71836
rect 90172 71780 90176 71836
rect 90112 71776 90176 71780
rect 90192 71836 90256 71840
rect 90192 71780 90196 71836
rect 90196 71780 90252 71836
rect 90252 71780 90256 71836
rect 90192 71776 90256 71780
rect 3952 71292 4016 71296
rect 3952 71236 3956 71292
rect 3956 71236 4012 71292
rect 4012 71236 4016 71292
rect 3952 71232 4016 71236
rect 4032 71292 4096 71296
rect 4032 71236 4036 71292
rect 4036 71236 4092 71292
rect 4092 71236 4096 71292
rect 4032 71232 4096 71236
rect 4112 71292 4176 71296
rect 4112 71236 4116 71292
rect 4116 71236 4172 71292
rect 4172 71236 4176 71292
rect 4112 71232 4176 71236
rect 4192 71292 4256 71296
rect 4192 71236 4196 71292
rect 4196 71236 4252 71292
rect 4252 71236 4256 71292
rect 4192 71232 4256 71236
rect 87952 71292 88016 71296
rect 87952 71236 87956 71292
rect 87956 71236 88012 71292
rect 88012 71236 88016 71292
rect 87952 71232 88016 71236
rect 88032 71292 88096 71296
rect 88032 71236 88036 71292
rect 88036 71236 88092 71292
rect 88092 71236 88096 71292
rect 88032 71232 88096 71236
rect 88112 71292 88176 71296
rect 88112 71236 88116 71292
rect 88116 71236 88172 71292
rect 88172 71236 88176 71292
rect 88112 71232 88176 71236
rect 88192 71292 88256 71296
rect 88192 71236 88196 71292
rect 88196 71236 88252 71292
rect 88252 71236 88256 71292
rect 88192 71232 88256 71236
rect 1952 70748 2016 70752
rect 1952 70692 1956 70748
rect 1956 70692 2012 70748
rect 2012 70692 2016 70748
rect 1952 70688 2016 70692
rect 2032 70748 2096 70752
rect 2032 70692 2036 70748
rect 2036 70692 2092 70748
rect 2092 70692 2096 70748
rect 2032 70688 2096 70692
rect 2112 70748 2176 70752
rect 2112 70692 2116 70748
rect 2116 70692 2172 70748
rect 2172 70692 2176 70748
rect 2112 70688 2176 70692
rect 2192 70748 2256 70752
rect 2192 70692 2196 70748
rect 2196 70692 2252 70748
rect 2252 70692 2256 70748
rect 2192 70688 2256 70692
rect 85952 70748 86016 70752
rect 85952 70692 85956 70748
rect 85956 70692 86012 70748
rect 86012 70692 86016 70748
rect 85952 70688 86016 70692
rect 86032 70748 86096 70752
rect 86032 70692 86036 70748
rect 86036 70692 86092 70748
rect 86092 70692 86096 70748
rect 86032 70688 86096 70692
rect 86112 70748 86176 70752
rect 86112 70692 86116 70748
rect 86116 70692 86172 70748
rect 86172 70692 86176 70748
rect 86112 70688 86176 70692
rect 86192 70748 86256 70752
rect 86192 70692 86196 70748
rect 86196 70692 86252 70748
rect 86252 70692 86256 70748
rect 86192 70688 86256 70692
rect 89952 70748 90016 70752
rect 89952 70692 89956 70748
rect 89956 70692 90012 70748
rect 90012 70692 90016 70748
rect 89952 70688 90016 70692
rect 90032 70748 90096 70752
rect 90032 70692 90036 70748
rect 90036 70692 90092 70748
rect 90092 70692 90096 70748
rect 90032 70688 90096 70692
rect 90112 70748 90176 70752
rect 90112 70692 90116 70748
rect 90116 70692 90172 70748
rect 90172 70692 90176 70748
rect 90112 70688 90176 70692
rect 90192 70748 90256 70752
rect 90192 70692 90196 70748
rect 90196 70692 90252 70748
rect 90252 70692 90256 70748
rect 90192 70688 90256 70692
rect 3952 70204 4016 70208
rect 3952 70148 3956 70204
rect 3956 70148 4012 70204
rect 4012 70148 4016 70204
rect 3952 70144 4016 70148
rect 4032 70204 4096 70208
rect 4032 70148 4036 70204
rect 4036 70148 4092 70204
rect 4092 70148 4096 70204
rect 4032 70144 4096 70148
rect 4112 70204 4176 70208
rect 4112 70148 4116 70204
rect 4116 70148 4172 70204
rect 4172 70148 4176 70204
rect 4112 70144 4176 70148
rect 4192 70204 4256 70208
rect 4192 70148 4196 70204
rect 4196 70148 4252 70204
rect 4252 70148 4256 70204
rect 4192 70144 4256 70148
rect 87952 70204 88016 70208
rect 87952 70148 87956 70204
rect 87956 70148 88012 70204
rect 88012 70148 88016 70204
rect 87952 70144 88016 70148
rect 88032 70204 88096 70208
rect 88032 70148 88036 70204
rect 88036 70148 88092 70204
rect 88092 70148 88096 70204
rect 88032 70144 88096 70148
rect 88112 70204 88176 70208
rect 88112 70148 88116 70204
rect 88116 70148 88172 70204
rect 88172 70148 88176 70204
rect 88112 70144 88176 70148
rect 88192 70204 88256 70208
rect 88192 70148 88196 70204
rect 88196 70148 88252 70204
rect 88252 70148 88256 70204
rect 88192 70144 88256 70148
rect 1952 69660 2016 69664
rect 1952 69604 1956 69660
rect 1956 69604 2012 69660
rect 2012 69604 2016 69660
rect 1952 69600 2016 69604
rect 2032 69660 2096 69664
rect 2032 69604 2036 69660
rect 2036 69604 2092 69660
rect 2092 69604 2096 69660
rect 2032 69600 2096 69604
rect 2112 69660 2176 69664
rect 2112 69604 2116 69660
rect 2116 69604 2172 69660
rect 2172 69604 2176 69660
rect 2112 69600 2176 69604
rect 2192 69660 2256 69664
rect 2192 69604 2196 69660
rect 2196 69604 2252 69660
rect 2252 69604 2256 69660
rect 2192 69600 2256 69604
rect 85952 69660 86016 69664
rect 85952 69604 85956 69660
rect 85956 69604 86012 69660
rect 86012 69604 86016 69660
rect 85952 69600 86016 69604
rect 86032 69660 86096 69664
rect 86032 69604 86036 69660
rect 86036 69604 86092 69660
rect 86092 69604 86096 69660
rect 86032 69600 86096 69604
rect 86112 69660 86176 69664
rect 86112 69604 86116 69660
rect 86116 69604 86172 69660
rect 86172 69604 86176 69660
rect 86112 69600 86176 69604
rect 86192 69660 86256 69664
rect 86192 69604 86196 69660
rect 86196 69604 86252 69660
rect 86252 69604 86256 69660
rect 86192 69600 86256 69604
rect 89952 69660 90016 69664
rect 89952 69604 89956 69660
rect 89956 69604 90012 69660
rect 90012 69604 90016 69660
rect 89952 69600 90016 69604
rect 90032 69660 90096 69664
rect 90032 69604 90036 69660
rect 90036 69604 90092 69660
rect 90092 69604 90096 69660
rect 90032 69600 90096 69604
rect 90112 69660 90176 69664
rect 90112 69604 90116 69660
rect 90116 69604 90172 69660
rect 90172 69604 90176 69660
rect 90112 69600 90176 69604
rect 90192 69660 90256 69664
rect 90192 69604 90196 69660
rect 90196 69604 90252 69660
rect 90252 69604 90256 69660
rect 90192 69600 90256 69604
rect 3952 69116 4016 69120
rect 3952 69060 3956 69116
rect 3956 69060 4012 69116
rect 4012 69060 4016 69116
rect 3952 69056 4016 69060
rect 4032 69116 4096 69120
rect 4032 69060 4036 69116
rect 4036 69060 4092 69116
rect 4092 69060 4096 69116
rect 4032 69056 4096 69060
rect 4112 69116 4176 69120
rect 4112 69060 4116 69116
rect 4116 69060 4172 69116
rect 4172 69060 4176 69116
rect 4112 69056 4176 69060
rect 4192 69116 4256 69120
rect 4192 69060 4196 69116
rect 4196 69060 4252 69116
rect 4252 69060 4256 69116
rect 4192 69056 4256 69060
rect 87952 69116 88016 69120
rect 87952 69060 87956 69116
rect 87956 69060 88012 69116
rect 88012 69060 88016 69116
rect 87952 69056 88016 69060
rect 88032 69116 88096 69120
rect 88032 69060 88036 69116
rect 88036 69060 88092 69116
rect 88092 69060 88096 69116
rect 88032 69056 88096 69060
rect 88112 69116 88176 69120
rect 88112 69060 88116 69116
rect 88116 69060 88172 69116
rect 88172 69060 88176 69116
rect 88112 69056 88176 69060
rect 88192 69116 88256 69120
rect 88192 69060 88196 69116
rect 88196 69060 88252 69116
rect 88252 69060 88256 69116
rect 88192 69056 88256 69060
rect 1952 68572 2016 68576
rect 1952 68516 1956 68572
rect 1956 68516 2012 68572
rect 2012 68516 2016 68572
rect 1952 68512 2016 68516
rect 2032 68572 2096 68576
rect 2032 68516 2036 68572
rect 2036 68516 2092 68572
rect 2092 68516 2096 68572
rect 2032 68512 2096 68516
rect 2112 68572 2176 68576
rect 2112 68516 2116 68572
rect 2116 68516 2172 68572
rect 2172 68516 2176 68572
rect 2112 68512 2176 68516
rect 2192 68572 2256 68576
rect 2192 68516 2196 68572
rect 2196 68516 2252 68572
rect 2252 68516 2256 68572
rect 2192 68512 2256 68516
rect 85952 68572 86016 68576
rect 85952 68516 85956 68572
rect 85956 68516 86012 68572
rect 86012 68516 86016 68572
rect 85952 68512 86016 68516
rect 86032 68572 86096 68576
rect 86032 68516 86036 68572
rect 86036 68516 86092 68572
rect 86092 68516 86096 68572
rect 86032 68512 86096 68516
rect 86112 68572 86176 68576
rect 86112 68516 86116 68572
rect 86116 68516 86172 68572
rect 86172 68516 86176 68572
rect 86112 68512 86176 68516
rect 86192 68572 86256 68576
rect 86192 68516 86196 68572
rect 86196 68516 86252 68572
rect 86252 68516 86256 68572
rect 86192 68512 86256 68516
rect 89952 68572 90016 68576
rect 89952 68516 89956 68572
rect 89956 68516 90012 68572
rect 90012 68516 90016 68572
rect 89952 68512 90016 68516
rect 90032 68572 90096 68576
rect 90032 68516 90036 68572
rect 90036 68516 90092 68572
rect 90092 68516 90096 68572
rect 90032 68512 90096 68516
rect 90112 68572 90176 68576
rect 90112 68516 90116 68572
rect 90116 68516 90172 68572
rect 90172 68516 90176 68572
rect 90112 68512 90176 68516
rect 90192 68572 90256 68576
rect 90192 68516 90196 68572
rect 90196 68516 90252 68572
rect 90252 68516 90256 68572
rect 90192 68512 90256 68516
rect 3952 68028 4016 68032
rect 3952 67972 3956 68028
rect 3956 67972 4012 68028
rect 4012 67972 4016 68028
rect 3952 67968 4016 67972
rect 4032 68028 4096 68032
rect 4032 67972 4036 68028
rect 4036 67972 4092 68028
rect 4092 67972 4096 68028
rect 4032 67968 4096 67972
rect 4112 68028 4176 68032
rect 4112 67972 4116 68028
rect 4116 67972 4172 68028
rect 4172 67972 4176 68028
rect 4112 67968 4176 67972
rect 4192 68028 4256 68032
rect 4192 67972 4196 68028
rect 4196 67972 4252 68028
rect 4252 67972 4256 68028
rect 4192 67968 4256 67972
rect 87952 68028 88016 68032
rect 87952 67972 87956 68028
rect 87956 67972 88012 68028
rect 88012 67972 88016 68028
rect 87952 67968 88016 67972
rect 88032 68028 88096 68032
rect 88032 67972 88036 68028
rect 88036 67972 88092 68028
rect 88092 67972 88096 68028
rect 88032 67968 88096 67972
rect 88112 68028 88176 68032
rect 88112 67972 88116 68028
rect 88116 67972 88172 68028
rect 88172 67972 88176 68028
rect 88112 67968 88176 67972
rect 88192 68028 88256 68032
rect 88192 67972 88196 68028
rect 88196 67972 88252 68028
rect 88252 67972 88256 68028
rect 88192 67968 88256 67972
rect 1952 67484 2016 67488
rect 1952 67428 1956 67484
rect 1956 67428 2012 67484
rect 2012 67428 2016 67484
rect 1952 67424 2016 67428
rect 2032 67484 2096 67488
rect 2032 67428 2036 67484
rect 2036 67428 2092 67484
rect 2092 67428 2096 67484
rect 2032 67424 2096 67428
rect 2112 67484 2176 67488
rect 2112 67428 2116 67484
rect 2116 67428 2172 67484
rect 2172 67428 2176 67484
rect 2112 67424 2176 67428
rect 2192 67484 2256 67488
rect 2192 67428 2196 67484
rect 2196 67428 2252 67484
rect 2252 67428 2256 67484
rect 2192 67424 2256 67428
rect 85952 67484 86016 67488
rect 85952 67428 85956 67484
rect 85956 67428 86012 67484
rect 86012 67428 86016 67484
rect 85952 67424 86016 67428
rect 86032 67484 86096 67488
rect 86032 67428 86036 67484
rect 86036 67428 86092 67484
rect 86092 67428 86096 67484
rect 86032 67424 86096 67428
rect 86112 67484 86176 67488
rect 86112 67428 86116 67484
rect 86116 67428 86172 67484
rect 86172 67428 86176 67484
rect 86112 67424 86176 67428
rect 86192 67484 86256 67488
rect 86192 67428 86196 67484
rect 86196 67428 86252 67484
rect 86252 67428 86256 67484
rect 86192 67424 86256 67428
rect 89952 67484 90016 67488
rect 89952 67428 89956 67484
rect 89956 67428 90012 67484
rect 90012 67428 90016 67484
rect 89952 67424 90016 67428
rect 90032 67484 90096 67488
rect 90032 67428 90036 67484
rect 90036 67428 90092 67484
rect 90092 67428 90096 67484
rect 90032 67424 90096 67428
rect 90112 67484 90176 67488
rect 90112 67428 90116 67484
rect 90116 67428 90172 67484
rect 90172 67428 90176 67484
rect 90112 67424 90176 67428
rect 90192 67484 90256 67488
rect 90192 67428 90196 67484
rect 90196 67428 90252 67484
rect 90252 67428 90256 67484
rect 90192 67424 90256 67428
rect 3952 66940 4016 66944
rect 3952 66884 3956 66940
rect 3956 66884 4012 66940
rect 4012 66884 4016 66940
rect 3952 66880 4016 66884
rect 4032 66940 4096 66944
rect 4032 66884 4036 66940
rect 4036 66884 4092 66940
rect 4092 66884 4096 66940
rect 4032 66880 4096 66884
rect 4112 66940 4176 66944
rect 4112 66884 4116 66940
rect 4116 66884 4172 66940
rect 4172 66884 4176 66940
rect 4112 66880 4176 66884
rect 4192 66940 4256 66944
rect 4192 66884 4196 66940
rect 4196 66884 4252 66940
rect 4252 66884 4256 66940
rect 4192 66880 4256 66884
rect 87952 66940 88016 66944
rect 87952 66884 87956 66940
rect 87956 66884 88012 66940
rect 88012 66884 88016 66940
rect 87952 66880 88016 66884
rect 88032 66940 88096 66944
rect 88032 66884 88036 66940
rect 88036 66884 88092 66940
rect 88092 66884 88096 66940
rect 88032 66880 88096 66884
rect 88112 66940 88176 66944
rect 88112 66884 88116 66940
rect 88116 66884 88172 66940
rect 88172 66884 88176 66940
rect 88112 66880 88176 66884
rect 88192 66940 88256 66944
rect 88192 66884 88196 66940
rect 88196 66884 88252 66940
rect 88252 66884 88256 66940
rect 88192 66880 88256 66884
rect 1952 66396 2016 66400
rect 1952 66340 1956 66396
rect 1956 66340 2012 66396
rect 2012 66340 2016 66396
rect 1952 66336 2016 66340
rect 2032 66396 2096 66400
rect 2032 66340 2036 66396
rect 2036 66340 2092 66396
rect 2092 66340 2096 66396
rect 2032 66336 2096 66340
rect 2112 66396 2176 66400
rect 2112 66340 2116 66396
rect 2116 66340 2172 66396
rect 2172 66340 2176 66396
rect 2112 66336 2176 66340
rect 2192 66396 2256 66400
rect 2192 66340 2196 66396
rect 2196 66340 2252 66396
rect 2252 66340 2256 66396
rect 2192 66336 2256 66340
rect 85952 66396 86016 66400
rect 85952 66340 85956 66396
rect 85956 66340 86012 66396
rect 86012 66340 86016 66396
rect 85952 66336 86016 66340
rect 86032 66396 86096 66400
rect 86032 66340 86036 66396
rect 86036 66340 86092 66396
rect 86092 66340 86096 66396
rect 86032 66336 86096 66340
rect 86112 66396 86176 66400
rect 86112 66340 86116 66396
rect 86116 66340 86172 66396
rect 86172 66340 86176 66396
rect 86112 66336 86176 66340
rect 86192 66396 86256 66400
rect 86192 66340 86196 66396
rect 86196 66340 86252 66396
rect 86252 66340 86256 66396
rect 86192 66336 86256 66340
rect 89952 66396 90016 66400
rect 89952 66340 89956 66396
rect 89956 66340 90012 66396
rect 90012 66340 90016 66396
rect 89952 66336 90016 66340
rect 90032 66396 90096 66400
rect 90032 66340 90036 66396
rect 90036 66340 90092 66396
rect 90092 66340 90096 66396
rect 90032 66336 90096 66340
rect 90112 66396 90176 66400
rect 90112 66340 90116 66396
rect 90116 66340 90172 66396
rect 90172 66340 90176 66396
rect 90112 66336 90176 66340
rect 90192 66396 90256 66400
rect 90192 66340 90196 66396
rect 90196 66340 90252 66396
rect 90252 66340 90256 66396
rect 90192 66336 90256 66340
rect 3952 65852 4016 65856
rect 3952 65796 3956 65852
rect 3956 65796 4012 65852
rect 4012 65796 4016 65852
rect 3952 65792 4016 65796
rect 4032 65852 4096 65856
rect 4032 65796 4036 65852
rect 4036 65796 4092 65852
rect 4092 65796 4096 65852
rect 4032 65792 4096 65796
rect 4112 65852 4176 65856
rect 4112 65796 4116 65852
rect 4116 65796 4172 65852
rect 4172 65796 4176 65852
rect 4112 65792 4176 65796
rect 4192 65852 4256 65856
rect 4192 65796 4196 65852
rect 4196 65796 4252 65852
rect 4252 65796 4256 65852
rect 4192 65792 4256 65796
rect 87952 65852 88016 65856
rect 87952 65796 87956 65852
rect 87956 65796 88012 65852
rect 88012 65796 88016 65852
rect 87952 65792 88016 65796
rect 88032 65852 88096 65856
rect 88032 65796 88036 65852
rect 88036 65796 88092 65852
rect 88092 65796 88096 65852
rect 88032 65792 88096 65796
rect 88112 65852 88176 65856
rect 88112 65796 88116 65852
rect 88116 65796 88172 65852
rect 88172 65796 88176 65852
rect 88112 65792 88176 65796
rect 88192 65852 88256 65856
rect 88192 65796 88196 65852
rect 88196 65796 88252 65852
rect 88252 65796 88256 65852
rect 88192 65792 88256 65796
rect 1952 65308 2016 65312
rect 1952 65252 1956 65308
rect 1956 65252 2012 65308
rect 2012 65252 2016 65308
rect 1952 65248 2016 65252
rect 2032 65308 2096 65312
rect 2032 65252 2036 65308
rect 2036 65252 2092 65308
rect 2092 65252 2096 65308
rect 2032 65248 2096 65252
rect 2112 65308 2176 65312
rect 2112 65252 2116 65308
rect 2116 65252 2172 65308
rect 2172 65252 2176 65308
rect 2112 65248 2176 65252
rect 2192 65308 2256 65312
rect 2192 65252 2196 65308
rect 2196 65252 2252 65308
rect 2252 65252 2256 65308
rect 2192 65248 2256 65252
rect 85952 65308 86016 65312
rect 85952 65252 85956 65308
rect 85956 65252 86012 65308
rect 86012 65252 86016 65308
rect 85952 65248 86016 65252
rect 86032 65308 86096 65312
rect 86032 65252 86036 65308
rect 86036 65252 86092 65308
rect 86092 65252 86096 65308
rect 86032 65248 86096 65252
rect 86112 65308 86176 65312
rect 86112 65252 86116 65308
rect 86116 65252 86172 65308
rect 86172 65252 86176 65308
rect 86112 65248 86176 65252
rect 86192 65308 86256 65312
rect 86192 65252 86196 65308
rect 86196 65252 86252 65308
rect 86252 65252 86256 65308
rect 86192 65248 86256 65252
rect 89952 65308 90016 65312
rect 89952 65252 89956 65308
rect 89956 65252 90012 65308
rect 90012 65252 90016 65308
rect 89952 65248 90016 65252
rect 90032 65308 90096 65312
rect 90032 65252 90036 65308
rect 90036 65252 90092 65308
rect 90092 65252 90096 65308
rect 90032 65248 90096 65252
rect 90112 65308 90176 65312
rect 90112 65252 90116 65308
rect 90116 65252 90172 65308
rect 90172 65252 90176 65308
rect 90112 65248 90176 65252
rect 90192 65308 90256 65312
rect 90192 65252 90196 65308
rect 90196 65252 90252 65308
rect 90252 65252 90256 65308
rect 90192 65248 90256 65252
rect 3952 64764 4016 64768
rect 3952 64708 3956 64764
rect 3956 64708 4012 64764
rect 4012 64708 4016 64764
rect 3952 64704 4016 64708
rect 4032 64764 4096 64768
rect 4032 64708 4036 64764
rect 4036 64708 4092 64764
rect 4092 64708 4096 64764
rect 4032 64704 4096 64708
rect 4112 64764 4176 64768
rect 4112 64708 4116 64764
rect 4116 64708 4172 64764
rect 4172 64708 4176 64764
rect 4112 64704 4176 64708
rect 4192 64764 4256 64768
rect 4192 64708 4196 64764
rect 4196 64708 4252 64764
rect 4252 64708 4256 64764
rect 4192 64704 4256 64708
rect 87952 64764 88016 64768
rect 87952 64708 87956 64764
rect 87956 64708 88012 64764
rect 88012 64708 88016 64764
rect 87952 64704 88016 64708
rect 88032 64764 88096 64768
rect 88032 64708 88036 64764
rect 88036 64708 88092 64764
rect 88092 64708 88096 64764
rect 88032 64704 88096 64708
rect 88112 64764 88176 64768
rect 88112 64708 88116 64764
rect 88116 64708 88172 64764
rect 88172 64708 88176 64764
rect 88112 64704 88176 64708
rect 88192 64764 88256 64768
rect 88192 64708 88196 64764
rect 88196 64708 88252 64764
rect 88252 64708 88256 64764
rect 88192 64704 88256 64708
rect 1952 64220 2016 64224
rect 1952 64164 1956 64220
rect 1956 64164 2012 64220
rect 2012 64164 2016 64220
rect 1952 64160 2016 64164
rect 2032 64220 2096 64224
rect 2032 64164 2036 64220
rect 2036 64164 2092 64220
rect 2092 64164 2096 64220
rect 2032 64160 2096 64164
rect 2112 64220 2176 64224
rect 2112 64164 2116 64220
rect 2116 64164 2172 64220
rect 2172 64164 2176 64220
rect 2112 64160 2176 64164
rect 2192 64220 2256 64224
rect 2192 64164 2196 64220
rect 2196 64164 2252 64220
rect 2252 64164 2256 64220
rect 2192 64160 2256 64164
rect 85952 64220 86016 64224
rect 85952 64164 85956 64220
rect 85956 64164 86012 64220
rect 86012 64164 86016 64220
rect 85952 64160 86016 64164
rect 86032 64220 86096 64224
rect 86032 64164 86036 64220
rect 86036 64164 86092 64220
rect 86092 64164 86096 64220
rect 86032 64160 86096 64164
rect 86112 64220 86176 64224
rect 86112 64164 86116 64220
rect 86116 64164 86172 64220
rect 86172 64164 86176 64220
rect 86112 64160 86176 64164
rect 86192 64220 86256 64224
rect 86192 64164 86196 64220
rect 86196 64164 86252 64220
rect 86252 64164 86256 64220
rect 86192 64160 86256 64164
rect 89952 64220 90016 64224
rect 89952 64164 89956 64220
rect 89956 64164 90012 64220
rect 90012 64164 90016 64220
rect 89952 64160 90016 64164
rect 90032 64220 90096 64224
rect 90032 64164 90036 64220
rect 90036 64164 90092 64220
rect 90092 64164 90096 64220
rect 90032 64160 90096 64164
rect 90112 64220 90176 64224
rect 90112 64164 90116 64220
rect 90116 64164 90172 64220
rect 90172 64164 90176 64220
rect 90112 64160 90176 64164
rect 90192 64220 90256 64224
rect 90192 64164 90196 64220
rect 90196 64164 90252 64220
rect 90252 64164 90256 64220
rect 90192 64160 90256 64164
rect 3952 63676 4016 63680
rect 3952 63620 3956 63676
rect 3956 63620 4012 63676
rect 4012 63620 4016 63676
rect 3952 63616 4016 63620
rect 4032 63676 4096 63680
rect 4032 63620 4036 63676
rect 4036 63620 4092 63676
rect 4092 63620 4096 63676
rect 4032 63616 4096 63620
rect 4112 63676 4176 63680
rect 4112 63620 4116 63676
rect 4116 63620 4172 63676
rect 4172 63620 4176 63676
rect 4112 63616 4176 63620
rect 4192 63676 4256 63680
rect 4192 63620 4196 63676
rect 4196 63620 4252 63676
rect 4252 63620 4256 63676
rect 4192 63616 4256 63620
rect 87952 63676 88016 63680
rect 87952 63620 87956 63676
rect 87956 63620 88012 63676
rect 88012 63620 88016 63676
rect 87952 63616 88016 63620
rect 88032 63676 88096 63680
rect 88032 63620 88036 63676
rect 88036 63620 88092 63676
rect 88092 63620 88096 63676
rect 88032 63616 88096 63620
rect 88112 63676 88176 63680
rect 88112 63620 88116 63676
rect 88116 63620 88172 63676
rect 88172 63620 88176 63676
rect 88112 63616 88176 63620
rect 88192 63676 88256 63680
rect 88192 63620 88196 63676
rect 88196 63620 88252 63676
rect 88252 63620 88256 63676
rect 88192 63616 88256 63620
rect 1952 63132 2016 63136
rect 1952 63076 1956 63132
rect 1956 63076 2012 63132
rect 2012 63076 2016 63132
rect 1952 63072 2016 63076
rect 2032 63132 2096 63136
rect 2032 63076 2036 63132
rect 2036 63076 2092 63132
rect 2092 63076 2096 63132
rect 2032 63072 2096 63076
rect 2112 63132 2176 63136
rect 2112 63076 2116 63132
rect 2116 63076 2172 63132
rect 2172 63076 2176 63132
rect 2112 63072 2176 63076
rect 2192 63132 2256 63136
rect 2192 63076 2196 63132
rect 2196 63076 2252 63132
rect 2252 63076 2256 63132
rect 2192 63072 2256 63076
rect 85952 63132 86016 63136
rect 85952 63076 85956 63132
rect 85956 63076 86012 63132
rect 86012 63076 86016 63132
rect 85952 63072 86016 63076
rect 86032 63132 86096 63136
rect 86032 63076 86036 63132
rect 86036 63076 86092 63132
rect 86092 63076 86096 63132
rect 86032 63072 86096 63076
rect 86112 63132 86176 63136
rect 86112 63076 86116 63132
rect 86116 63076 86172 63132
rect 86172 63076 86176 63132
rect 86112 63072 86176 63076
rect 86192 63132 86256 63136
rect 86192 63076 86196 63132
rect 86196 63076 86252 63132
rect 86252 63076 86256 63132
rect 86192 63072 86256 63076
rect 89952 63132 90016 63136
rect 89952 63076 89956 63132
rect 89956 63076 90012 63132
rect 90012 63076 90016 63132
rect 89952 63072 90016 63076
rect 90032 63132 90096 63136
rect 90032 63076 90036 63132
rect 90036 63076 90092 63132
rect 90092 63076 90096 63132
rect 90032 63072 90096 63076
rect 90112 63132 90176 63136
rect 90112 63076 90116 63132
rect 90116 63076 90172 63132
rect 90172 63076 90176 63132
rect 90112 63072 90176 63076
rect 90192 63132 90256 63136
rect 90192 63076 90196 63132
rect 90196 63076 90252 63132
rect 90252 63076 90256 63132
rect 90192 63072 90256 63076
rect 3952 62588 4016 62592
rect 3952 62532 3956 62588
rect 3956 62532 4012 62588
rect 4012 62532 4016 62588
rect 3952 62528 4016 62532
rect 4032 62588 4096 62592
rect 4032 62532 4036 62588
rect 4036 62532 4092 62588
rect 4092 62532 4096 62588
rect 4032 62528 4096 62532
rect 4112 62588 4176 62592
rect 4112 62532 4116 62588
rect 4116 62532 4172 62588
rect 4172 62532 4176 62588
rect 4112 62528 4176 62532
rect 4192 62588 4256 62592
rect 4192 62532 4196 62588
rect 4196 62532 4252 62588
rect 4252 62532 4256 62588
rect 4192 62528 4256 62532
rect 87952 62588 88016 62592
rect 87952 62532 87956 62588
rect 87956 62532 88012 62588
rect 88012 62532 88016 62588
rect 87952 62528 88016 62532
rect 88032 62588 88096 62592
rect 88032 62532 88036 62588
rect 88036 62532 88092 62588
rect 88092 62532 88096 62588
rect 88032 62528 88096 62532
rect 88112 62588 88176 62592
rect 88112 62532 88116 62588
rect 88116 62532 88172 62588
rect 88172 62532 88176 62588
rect 88112 62528 88176 62532
rect 88192 62588 88256 62592
rect 88192 62532 88196 62588
rect 88196 62532 88252 62588
rect 88252 62532 88256 62588
rect 88192 62528 88256 62532
rect 1952 62044 2016 62048
rect 1952 61988 1956 62044
rect 1956 61988 2012 62044
rect 2012 61988 2016 62044
rect 1952 61984 2016 61988
rect 2032 62044 2096 62048
rect 2032 61988 2036 62044
rect 2036 61988 2092 62044
rect 2092 61988 2096 62044
rect 2032 61984 2096 61988
rect 2112 62044 2176 62048
rect 2112 61988 2116 62044
rect 2116 61988 2172 62044
rect 2172 61988 2176 62044
rect 2112 61984 2176 61988
rect 2192 62044 2256 62048
rect 2192 61988 2196 62044
rect 2196 61988 2252 62044
rect 2252 61988 2256 62044
rect 2192 61984 2256 61988
rect 85952 62044 86016 62048
rect 85952 61988 85956 62044
rect 85956 61988 86012 62044
rect 86012 61988 86016 62044
rect 85952 61984 86016 61988
rect 86032 62044 86096 62048
rect 86032 61988 86036 62044
rect 86036 61988 86092 62044
rect 86092 61988 86096 62044
rect 86032 61984 86096 61988
rect 86112 62044 86176 62048
rect 86112 61988 86116 62044
rect 86116 61988 86172 62044
rect 86172 61988 86176 62044
rect 86112 61984 86176 61988
rect 86192 62044 86256 62048
rect 86192 61988 86196 62044
rect 86196 61988 86252 62044
rect 86252 61988 86256 62044
rect 86192 61984 86256 61988
rect 89952 62044 90016 62048
rect 89952 61988 89956 62044
rect 89956 61988 90012 62044
rect 90012 61988 90016 62044
rect 89952 61984 90016 61988
rect 90032 62044 90096 62048
rect 90032 61988 90036 62044
rect 90036 61988 90092 62044
rect 90092 61988 90096 62044
rect 90032 61984 90096 61988
rect 90112 62044 90176 62048
rect 90112 61988 90116 62044
rect 90116 61988 90172 62044
rect 90172 61988 90176 62044
rect 90112 61984 90176 61988
rect 90192 62044 90256 62048
rect 90192 61988 90196 62044
rect 90196 61988 90252 62044
rect 90252 61988 90256 62044
rect 90192 61984 90256 61988
rect 3952 61500 4016 61504
rect 3952 61444 3956 61500
rect 3956 61444 4012 61500
rect 4012 61444 4016 61500
rect 3952 61440 4016 61444
rect 4032 61500 4096 61504
rect 4032 61444 4036 61500
rect 4036 61444 4092 61500
rect 4092 61444 4096 61500
rect 4032 61440 4096 61444
rect 4112 61500 4176 61504
rect 4112 61444 4116 61500
rect 4116 61444 4172 61500
rect 4172 61444 4176 61500
rect 4112 61440 4176 61444
rect 4192 61500 4256 61504
rect 4192 61444 4196 61500
rect 4196 61444 4252 61500
rect 4252 61444 4256 61500
rect 4192 61440 4256 61444
rect 87952 61500 88016 61504
rect 87952 61444 87956 61500
rect 87956 61444 88012 61500
rect 88012 61444 88016 61500
rect 87952 61440 88016 61444
rect 88032 61500 88096 61504
rect 88032 61444 88036 61500
rect 88036 61444 88092 61500
rect 88092 61444 88096 61500
rect 88032 61440 88096 61444
rect 88112 61500 88176 61504
rect 88112 61444 88116 61500
rect 88116 61444 88172 61500
rect 88172 61444 88176 61500
rect 88112 61440 88176 61444
rect 88192 61500 88256 61504
rect 88192 61444 88196 61500
rect 88196 61444 88252 61500
rect 88252 61444 88256 61500
rect 88192 61440 88256 61444
rect 1952 60956 2016 60960
rect 1952 60900 1956 60956
rect 1956 60900 2012 60956
rect 2012 60900 2016 60956
rect 1952 60896 2016 60900
rect 2032 60956 2096 60960
rect 2032 60900 2036 60956
rect 2036 60900 2092 60956
rect 2092 60900 2096 60956
rect 2032 60896 2096 60900
rect 2112 60956 2176 60960
rect 2112 60900 2116 60956
rect 2116 60900 2172 60956
rect 2172 60900 2176 60956
rect 2112 60896 2176 60900
rect 2192 60956 2256 60960
rect 2192 60900 2196 60956
rect 2196 60900 2252 60956
rect 2252 60900 2256 60956
rect 2192 60896 2256 60900
rect 85952 60956 86016 60960
rect 85952 60900 85956 60956
rect 85956 60900 86012 60956
rect 86012 60900 86016 60956
rect 85952 60896 86016 60900
rect 86032 60956 86096 60960
rect 86032 60900 86036 60956
rect 86036 60900 86092 60956
rect 86092 60900 86096 60956
rect 86032 60896 86096 60900
rect 86112 60956 86176 60960
rect 86112 60900 86116 60956
rect 86116 60900 86172 60956
rect 86172 60900 86176 60956
rect 86112 60896 86176 60900
rect 86192 60956 86256 60960
rect 86192 60900 86196 60956
rect 86196 60900 86252 60956
rect 86252 60900 86256 60956
rect 86192 60896 86256 60900
rect 89952 60956 90016 60960
rect 89952 60900 89956 60956
rect 89956 60900 90012 60956
rect 90012 60900 90016 60956
rect 89952 60896 90016 60900
rect 90032 60956 90096 60960
rect 90032 60900 90036 60956
rect 90036 60900 90092 60956
rect 90092 60900 90096 60956
rect 90032 60896 90096 60900
rect 90112 60956 90176 60960
rect 90112 60900 90116 60956
rect 90116 60900 90172 60956
rect 90172 60900 90176 60956
rect 90112 60896 90176 60900
rect 90192 60956 90256 60960
rect 90192 60900 90196 60956
rect 90196 60900 90252 60956
rect 90252 60900 90256 60956
rect 90192 60896 90256 60900
rect 3952 60412 4016 60416
rect 3952 60356 3956 60412
rect 3956 60356 4012 60412
rect 4012 60356 4016 60412
rect 3952 60352 4016 60356
rect 4032 60412 4096 60416
rect 4032 60356 4036 60412
rect 4036 60356 4092 60412
rect 4092 60356 4096 60412
rect 4032 60352 4096 60356
rect 4112 60412 4176 60416
rect 4112 60356 4116 60412
rect 4116 60356 4172 60412
rect 4172 60356 4176 60412
rect 4112 60352 4176 60356
rect 4192 60412 4256 60416
rect 4192 60356 4196 60412
rect 4196 60356 4252 60412
rect 4252 60356 4256 60412
rect 4192 60352 4256 60356
rect 87952 60412 88016 60416
rect 87952 60356 87956 60412
rect 87956 60356 88012 60412
rect 88012 60356 88016 60412
rect 87952 60352 88016 60356
rect 88032 60412 88096 60416
rect 88032 60356 88036 60412
rect 88036 60356 88092 60412
rect 88092 60356 88096 60412
rect 88032 60352 88096 60356
rect 88112 60412 88176 60416
rect 88112 60356 88116 60412
rect 88116 60356 88172 60412
rect 88172 60356 88176 60412
rect 88112 60352 88176 60356
rect 88192 60412 88256 60416
rect 88192 60356 88196 60412
rect 88196 60356 88252 60412
rect 88252 60356 88256 60412
rect 88192 60352 88256 60356
rect 1952 59868 2016 59872
rect 1952 59812 1956 59868
rect 1956 59812 2012 59868
rect 2012 59812 2016 59868
rect 1952 59808 2016 59812
rect 2032 59868 2096 59872
rect 2032 59812 2036 59868
rect 2036 59812 2092 59868
rect 2092 59812 2096 59868
rect 2032 59808 2096 59812
rect 2112 59868 2176 59872
rect 2112 59812 2116 59868
rect 2116 59812 2172 59868
rect 2172 59812 2176 59868
rect 2112 59808 2176 59812
rect 2192 59868 2256 59872
rect 2192 59812 2196 59868
rect 2196 59812 2252 59868
rect 2252 59812 2256 59868
rect 2192 59808 2256 59812
rect 85952 59868 86016 59872
rect 85952 59812 85956 59868
rect 85956 59812 86012 59868
rect 86012 59812 86016 59868
rect 85952 59808 86016 59812
rect 86032 59868 86096 59872
rect 86032 59812 86036 59868
rect 86036 59812 86092 59868
rect 86092 59812 86096 59868
rect 86032 59808 86096 59812
rect 86112 59868 86176 59872
rect 86112 59812 86116 59868
rect 86116 59812 86172 59868
rect 86172 59812 86176 59868
rect 86112 59808 86176 59812
rect 86192 59868 86256 59872
rect 86192 59812 86196 59868
rect 86196 59812 86252 59868
rect 86252 59812 86256 59868
rect 86192 59808 86256 59812
rect 89952 59868 90016 59872
rect 89952 59812 89956 59868
rect 89956 59812 90012 59868
rect 90012 59812 90016 59868
rect 89952 59808 90016 59812
rect 90032 59868 90096 59872
rect 90032 59812 90036 59868
rect 90036 59812 90092 59868
rect 90092 59812 90096 59868
rect 90032 59808 90096 59812
rect 90112 59868 90176 59872
rect 90112 59812 90116 59868
rect 90116 59812 90172 59868
rect 90172 59812 90176 59868
rect 90112 59808 90176 59812
rect 90192 59868 90256 59872
rect 90192 59812 90196 59868
rect 90196 59812 90252 59868
rect 90252 59812 90256 59868
rect 90192 59808 90256 59812
rect 3952 59324 4016 59328
rect 3952 59268 3956 59324
rect 3956 59268 4012 59324
rect 4012 59268 4016 59324
rect 3952 59264 4016 59268
rect 4032 59324 4096 59328
rect 4032 59268 4036 59324
rect 4036 59268 4092 59324
rect 4092 59268 4096 59324
rect 4032 59264 4096 59268
rect 4112 59324 4176 59328
rect 4112 59268 4116 59324
rect 4116 59268 4172 59324
rect 4172 59268 4176 59324
rect 4112 59264 4176 59268
rect 4192 59324 4256 59328
rect 4192 59268 4196 59324
rect 4196 59268 4252 59324
rect 4252 59268 4256 59324
rect 4192 59264 4256 59268
rect 87952 59324 88016 59328
rect 87952 59268 87956 59324
rect 87956 59268 88012 59324
rect 88012 59268 88016 59324
rect 87952 59264 88016 59268
rect 88032 59324 88096 59328
rect 88032 59268 88036 59324
rect 88036 59268 88092 59324
rect 88092 59268 88096 59324
rect 88032 59264 88096 59268
rect 88112 59324 88176 59328
rect 88112 59268 88116 59324
rect 88116 59268 88172 59324
rect 88172 59268 88176 59324
rect 88112 59264 88176 59268
rect 88192 59324 88256 59328
rect 88192 59268 88196 59324
rect 88196 59268 88252 59324
rect 88252 59268 88256 59324
rect 88192 59264 88256 59268
rect 1952 58780 2016 58784
rect 1952 58724 1956 58780
rect 1956 58724 2012 58780
rect 2012 58724 2016 58780
rect 1952 58720 2016 58724
rect 2032 58780 2096 58784
rect 2032 58724 2036 58780
rect 2036 58724 2092 58780
rect 2092 58724 2096 58780
rect 2032 58720 2096 58724
rect 2112 58780 2176 58784
rect 2112 58724 2116 58780
rect 2116 58724 2172 58780
rect 2172 58724 2176 58780
rect 2112 58720 2176 58724
rect 2192 58780 2256 58784
rect 2192 58724 2196 58780
rect 2196 58724 2252 58780
rect 2252 58724 2256 58780
rect 2192 58720 2256 58724
rect 85952 58780 86016 58784
rect 85952 58724 85956 58780
rect 85956 58724 86012 58780
rect 86012 58724 86016 58780
rect 85952 58720 86016 58724
rect 86032 58780 86096 58784
rect 86032 58724 86036 58780
rect 86036 58724 86092 58780
rect 86092 58724 86096 58780
rect 86032 58720 86096 58724
rect 86112 58780 86176 58784
rect 86112 58724 86116 58780
rect 86116 58724 86172 58780
rect 86172 58724 86176 58780
rect 86112 58720 86176 58724
rect 86192 58780 86256 58784
rect 86192 58724 86196 58780
rect 86196 58724 86252 58780
rect 86252 58724 86256 58780
rect 86192 58720 86256 58724
rect 89952 58780 90016 58784
rect 89952 58724 89956 58780
rect 89956 58724 90012 58780
rect 90012 58724 90016 58780
rect 89952 58720 90016 58724
rect 90032 58780 90096 58784
rect 90032 58724 90036 58780
rect 90036 58724 90092 58780
rect 90092 58724 90096 58780
rect 90032 58720 90096 58724
rect 90112 58780 90176 58784
rect 90112 58724 90116 58780
rect 90116 58724 90172 58780
rect 90172 58724 90176 58780
rect 90112 58720 90176 58724
rect 90192 58780 90256 58784
rect 90192 58724 90196 58780
rect 90196 58724 90252 58780
rect 90252 58724 90256 58780
rect 90192 58720 90256 58724
rect 3952 58236 4016 58240
rect 3952 58180 3956 58236
rect 3956 58180 4012 58236
rect 4012 58180 4016 58236
rect 3952 58176 4016 58180
rect 4032 58236 4096 58240
rect 4032 58180 4036 58236
rect 4036 58180 4092 58236
rect 4092 58180 4096 58236
rect 4032 58176 4096 58180
rect 4112 58236 4176 58240
rect 4112 58180 4116 58236
rect 4116 58180 4172 58236
rect 4172 58180 4176 58236
rect 4112 58176 4176 58180
rect 4192 58236 4256 58240
rect 4192 58180 4196 58236
rect 4196 58180 4252 58236
rect 4252 58180 4256 58236
rect 4192 58176 4256 58180
rect 87952 58236 88016 58240
rect 87952 58180 87956 58236
rect 87956 58180 88012 58236
rect 88012 58180 88016 58236
rect 87952 58176 88016 58180
rect 88032 58236 88096 58240
rect 88032 58180 88036 58236
rect 88036 58180 88092 58236
rect 88092 58180 88096 58236
rect 88032 58176 88096 58180
rect 88112 58236 88176 58240
rect 88112 58180 88116 58236
rect 88116 58180 88172 58236
rect 88172 58180 88176 58236
rect 88112 58176 88176 58180
rect 88192 58236 88256 58240
rect 88192 58180 88196 58236
rect 88196 58180 88252 58236
rect 88252 58180 88256 58236
rect 88192 58176 88256 58180
rect 1952 57692 2016 57696
rect 1952 57636 1956 57692
rect 1956 57636 2012 57692
rect 2012 57636 2016 57692
rect 1952 57632 2016 57636
rect 2032 57692 2096 57696
rect 2032 57636 2036 57692
rect 2036 57636 2092 57692
rect 2092 57636 2096 57692
rect 2032 57632 2096 57636
rect 2112 57692 2176 57696
rect 2112 57636 2116 57692
rect 2116 57636 2172 57692
rect 2172 57636 2176 57692
rect 2112 57632 2176 57636
rect 2192 57692 2256 57696
rect 2192 57636 2196 57692
rect 2196 57636 2252 57692
rect 2252 57636 2256 57692
rect 2192 57632 2256 57636
rect 85952 57692 86016 57696
rect 85952 57636 85956 57692
rect 85956 57636 86012 57692
rect 86012 57636 86016 57692
rect 85952 57632 86016 57636
rect 86032 57692 86096 57696
rect 86032 57636 86036 57692
rect 86036 57636 86092 57692
rect 86092 57636 86096 57692
rect 86032 57632 86096 57636
rect 86112 57692 86176 57696
rect 86112 57636 86116 57692
rect 86116 57636 86172 57692
rect 86172 57636 86176 57692
rect 86112 57632 86176 57636
rect 86192 57692 86256 57696
rect 86192 57636 86196 57692
rect 86196 57636 86252 57692
rect 86252 57636 86256 57692
rect 86192 57632 86256 57636
rect 89952 57692 90016 57696
rect 89952 57636 89956 57692
rect 89956 57636 90012 57692
rect 90012 57636 90016 57692
rect 89952 57632 90016 57636
rect 90032 57692 90096 57696
rect 90032 57636 90036 57692
rect 90036 57636 90092 57692
rect 90092 57636 90096 57692
rect 90032 57632 90096 57636
rect 90112 57692 90176 57696
rect 90112 57636 90116 57692
rect 90116 57636 90172 57692
rect 90172 57636 90176 57692
rect 90112 57632 90176 57636
rect 90192 57692 90256 57696
rect 90192 57636 90196 57692
rect 90196 57636 90252 57692
rect 90252 57636 90256 57692
rect 90192 57632 90256 57636
rect 3952 57148 4016 57152
rect 3952 57092 3956 57148
rect 3956 57092 4012 57148
rect 4012 57092 4016 57148
rect 3952 57088 4016 57092
rect 4032 57148 4096 57152
rect 4032 57092 4036 57148
rect 4036 57092 4092 57148
rect 4092 57092 4096 57148
rect 4032 57088 4096 57092
rect 4112 57148 4176 57152
rect 4112 57092 4116 57148
rect 4116 57092 4172 57148
rect 4172 57092 4176 57148
rect 4112 57088 4176 57092
rect 4192 57148 4256 57152
rect 4192 57092 4196 57148
rect 4196 57092 4252 57148
rect 4252 57092 4256 57148
rect 4192 57088 4256 57092
rect 87952 57148 88016 57152
rect 87952 57092 87956 57148
rect 87956 57092 88012 57148
rect 88012 57092 88016 57148
rect 87952 57088 88016 57092
rect 88032 57148 88096 57152
rect 88032 57092 88036 57148
rect 88036 57092 88092 57148
rect 88092 57092 88096 57148
rect 88032 57088 88096 57092
rect 88112 57148 88176 57152
rect 88112 57092 88116 57148
rect 88116 57092 88172 57148
rect 88172 57092 88176 57148
rect 88112 57088 88176 57092
rect 88192 57148 88256 57152
rect 88192 57092 88196 57148
rect 88196 57092 88252 57148
rect 88252 57092 88256 57148
rect 88192 57088 88256 57092
rect 1952 56604 2016 56608
rect 1952 56548 1956 56604
rect 1956 56548 2012 56604
rect 2012 56548 2016 56604
rect 1952 56544 2016 56548
rect 2032 56604 2096 56608
rect 2032 56548 2036 56604
rect 2036 56548 2092 56604
rect 2092 56548 2096 56604
rect 2032 56544 2096 56548
rect 2112 56604 2176 56608
rect 2112 56548 2116 56604
rect 2116 56548 2172 56604
rect 2172 56548 2176 56604
rect 2112 56544 2176 56548
rect 2192 56604 2256 56608
rect 2192 56548 2196 56604
rect 2196 56548 2252 56604
rect 2252 56548 2256 56604
rect 2192 56544 2256 56548
rect 85952 56604 86016 56608
rect 85952 56548 85956 56604
rect 85956 56548 86012 56604
rect 86012 56548 86016 56604
rect 85952 56544 86016 56548
rect 86032 56604 86096 56608
rect 86032 56548 86036 56604
rect 86036 56548 86092 56604
rect 86092 56548 86096 56604
rect 86032 56544 86096 56548
rect 86112 56604 86176 56608
rect 86112 56548 86116 56604
rect 86116 56548 86172 56604
rect 86172 56548 86176 56604
rect 86112 56544 86176 56548
rect 86192 56604 86256 56608
rect 86192 56548 86196 56604
rect 86196 56548 86252 56604
rect 86252 56548 86256 56604
rect 86192 56544 86256 56548
rect 89952 56604 90016 56608
rect 89952 56548 89956 56604
rect 89956 56548 90012 56604
rect 90012 56548 90016 56604
rect 89952 56544 90016 56548
rect 90032 56604 90096 56608
rect 90032 56548 90036 56604
rect 90036 56548 90092 56604
rect 90092 56548 90096 56604
rect 90032 56544 90096 56548
rect 90112 56604 90176 56608
rect 90112 56548 90116 56604
rect 90116 56548 90172 56604
rect 90172 56548 90176 56604
rect 90112 56544 90176 56548
rect 90192 56604 90256 56608
rect 90192 56548 90196 56604
rect 90196 56548 90252 56604
rect 90252 56548 90256 56604
rect 90192 56544 90256 56548
rect 3952 56060 4016 56064
rect 3952 56004 3956 56060
rect 3956 56004 4012 56060
rect 4012 56004 4016 56060
rect 3952 56000 4016 56004
rect 4032 56060 4096 56064
rect 4032 56004 4036 56060
rect 4036 56004 4092 56060
rect 4092 56004 4096 56060
rect 4032 56000 4096 56004
rect 4112 56060 4176 56064
rect 4112 56004 4116 56060
rect 4116 56004 4172 56060
rect 4172 56004 4176 56060
rect 4112 56000 4176 56004
rect 4192 56060 4256 56064
rect 4192 56004 4196 56060
rect 4196 56004 4252 56060
rect 4252 56004 4256 56060
rect 4192 56000 4256 56004
rect 87952 56060 88016 56064
rect 87952 56004 87956 56060
rect 87956 56004 88012 56060
rect 88012 56004 88016 56060
rect 87952 56000 88016 56004
rect 88032 56060 88096 56064
rect 88032 56004 88036 56060
rect 88036 56004 88092 56060
rect 88092 56004 88096 56060
rect 88032 56000 88096 56004
rect 88112 56060 88176 56064
rect 88112 56004 88116 56060
rect 88116 56004 88172 56060
rect 88172 56004 88176 56060
rect 88112 56000 88176 56004
rect 88192 56060 88256 56064
rect 88192 56004 88196 56060
rect 88196 56004 88252 56060
rect 88252 56004 88256 56060
rect 88192 56000 88256 56004
rect 1952 55516 2016 55520
rect 1952 55460 1956 55516
rect 1956 55460 2012 55516
rect 2012 55460 2016 55516
rect 1952 55456 2016 55460
rect 2032 55516 2096 55520
rect 2032 55460 2036 55516
rect 2036 55460 2092 55516
rect 2092 55460 2096 55516
rect 2032 55456 2096 55460
rect 2112 55516 2176 55520
rect 2112 55460 2116 55516
rect 2116 55460 2172 55516
rect 2172 55460 2176 55516
rect 2112 55456 2176 55460
rect 2192 55516 2256 55520
rect 2192 55460 2196 55516
rect 2196 55460 2252 55516
rect 2252 55460 2256 55516
rect 2192 55456 2256 55460
rect 85952 55516 86016 55520
rect 85952 55460 85956 55516
rect 85956 55460 86012 55516
rect 86012 55460 86016 55516
rect 85952 55456 86016 55460
rect 86032 55516 86096 55520
rect 86032 55460 86036 55516
rect 86036 55460 86092 55516
rect 86092 55460 86096 55516
rect 86032 55456 86096 55460
rect 86112 55516 86176 55520
rect 86112 55460 86116 55516
rect 86116 55460 86172 55516
rect 86172 55460 86176 55516
rect 86112 55456 86176 55460
rect 86192 55516 86256 55520
rect 86192 55460 86196 55516
rect 86196 55460 86252 55516
rect 86252 55460 86256 55516
rect 86192 55456 86256 55460
rect 89952 55516 90016 55520
rect 89952 55460 89956 55516
rect 89956 55460 90012 55516
rect 90012 55460 90016 55516
rect 89952 55456 90016 55460
rect 90032 55516 90096 55520
rect 90032 55460 90036 55516
rect 90036 55460 90092 55516
rect 90092 55460 90096 55516
rect 90032 55456 90096 55460
rect 90112 55516 90176 55520
rect 90112 55460 90116 55516
rect 90116 55460 90172 55516
rect 90172 55460 90176 55516
rect 90112 55456 90176 55460
rect 90192 55516 90256 55520
rect 90192 55460 90196 55516
rect 90196 55460 90252 55516
rect 90252 55460 90256 55516
rect 90192 55456 90256 55460
rect 84148 55252 84212 55316
rect 3952 54972 4016 54976
rect 3952 54916 3956 54972
rect 3956 54916 4012 54972
rect 4012 54916 4016 54972
rect 3952 54912 4016 54916
rect 4032 54972 4096 54976
rect 4032 54916 4036 54972
rect 4036 54916 4092 54972
rect 4092 54916 4096 54972
rect 4032 54912 4096 54916
rect 4112 54972 4176 54976
rect 4112 54916 4116 54972
rect 4116 54916 4172 54972
rect 4172 54916 4176 54972
rect 4112 54912 4176 54916
rect 4192 54972 4256 54976
rect 4192 54916 4196 54972
rect 4196 54916 4252 54972
rect 4252 54916 4256 54972
rect 4192 54912 4256 54916
rect 87952 54972 88016 54976
rect 87952 54916 87956 54972
rect 87956 54916 88012 54972
rect 88012 54916 88016 54972
rect 87952 54912 88016 54916
rect 88032 54972 88096 54976
rect 88032 54916 88036 54972
rect 88036 54916 88092 54972
rect 88092 54916 88096 54972
rect 88032 54912 88096 54916
rect 88112 54972 88176 54976
rect 88112 54916 88116 54972
rect 88116 54916 88172 54972
rect 88172 54916 88176 54972
rect 88112 54912 88176 54916
rect 88192 54972 88256 54976
rect 88192 54916 88196 54972
rect 88196 54916 88252 54972
rect 88252 54916 88256 54972
rect 88192 54912 88256 54916
rect 1952 54428 2016 54432
rect 1952 54372 1956 54428
rect 1956 54372 2012 54428
rect 2012 54372 2016 54428
rect 1952 54368 2016 54372
rect 2032 54428 2096 54432
rect 2032 54372 2036 54428
rect 2036 54372 2092 54428
rect 2092 54372 2096 54428
rect 2032 54368 2096 54372
rect 2112 54428 2176 54432
rect 2112 54372 2116 54428
rect 2116 54372 2172 54428
rect 2172 54372 2176 54428
rect 2112 54368 2176 54372
rect 2192 54428 2256 54432
rect 2192 54372 2196 54428
rect 2196 54372 2252 54428
rect 2252 54372 2256 54428
rect 2192 54368 2256 54372
rect 85952 54428 86016 54432
rect 85952 54372 85956 54428
rect 85956 54372 86012 54428
rect 86012 54372 86016 54428
rect 85952 54368 86016 54372
rect 86032 54428 86096 54432
rect 86032 54372 86036 54428
rect 86036 54372 86092 54428
rect 86092 54372 86096 54428
rect 86032 54368 86096 54372
rect 86112 54428 86176 54432
rect 86112 54372 86116 54428
rect 86116 54372 86172 54428
rect 86172 54372 86176 54428
rect 86112 54368 86176 54372
rect 86192 54428 86256 54432
rect 86192 54372 86196 54428
rect 86196 54372 86252 54428
rect 86252 54372 86256 54428
rect 86192 54368 86256 54372
rect 89952 54428 90016 54432
rect 89952 54372 89956 54428
rect 89956 54372 90012 54428
rect 90012 54372 90016 54428
rect 89952 54368 90016 54372
rect 90032 54428 90096 54432
rect 90032 54372 90036 54428
rect 90036 54372 90092 54428
rect 90092 54372 90096 54428
rect 90032 54368 90096 54372
rect 90112 54428 90176 54432
rect 90112 54372 90116 54428
rect 90116 54372 90172 54428
rect 90172 54372 90176 54428
rect 90112 54368 90176 54372
rect 90192 54428 90256 54432
rect 90192 54372 90196 54428
rect 90196 54372 90252 54428
rect 90252 54372 90256 54428
rect 90192 54368 90256 54372
rect 3952 53884 4016 53888
rect 3952 53828 3956 53884
rect 3956 53828 4012 53884
rect 4012 53828 4016 53884
rect 3952 53824 4016 53828
rect 4032 53884 4096 53888
rect 4032 53828 4036 53884
rect 4036 53828 4092 53884
rect 4092 53828 4096 53884
rect 4032 53824 4096 53828
rect 4112 53884 4176 53888
rect 4112 53828 4116 53884
rect 4116 53828 4172 53884
rect 4172 53828 4176 53884
rect 4112 53824 4176 53828
rect 4192 53884 4256 53888
rect 4192 53828 4196 53884
rect 4196 53828 4252 53884
rect 4252 53828 4256 53884
rect 4192 53824 4256 53828
rect 87952 53884 88016 53888
rect 87952 53828 87956 53884
rect 87956 53828 88012 53884
rect 88012 53828 88016 53884
rect 87952 53824 88016 53828
rect 88032 53884 88096 53888
rect 88032 53828 88036 53884
rect 88036 53828 88092 53884
rect 88092 53828 88096 53884
rect 88032 53824 88096 53828
rect 88112 53884 88176 53888
rect 88112 53828 88116 53884
rect 88116 53828 88172 53884
rect 88172 53828 88176 53884
rect 88112 53824 88176 53828
rect 88192 53884 88256 53888
rect 88192 53828 88196 53884
rect 88196 53828 88252 53884
rect 88252 53828 88256 53884
rect 88192 53824 88256 53828
rect 1952 53340 2016 53344
rect 1952 53284 1956 53340
rect 1956 53284 2012 53340
rect 2012 53284 2016 53340
rect 1952 53280 2016 53284
rect 2032 53340 2096 53344
rect 2032 53284 2036 53340
rect 2036 53284 2092 53340
rect 2092 53284 2096 53340
rect 2032 53280 2096 53284
rect 2112 53340 2176 53344
rect 2112 53284 2116 53340
rect 2116 53284 2172 53340
rect 2172 53284 2176 53340
rect 2112 53280 2176 53284
rect 2192 53340 2256 53344
rect 2192 53284 2196 53340
rect 2196 53284 2252 53340
rect 2252 53284 2256 53340
rect 2192 53280 2256 53284
rect 85952 53340 86016 53344
rect 85952 53284 85956 53340
rect 85956 53284 86012 53340
rect 86012 53284 86016 53340
rect 85952 53280 86016 53284
rect 86032 53340 86096 53344
rect 86032 53284 86036 53340
rect 86036 53284 86092 53340
rect 86092 53284 86096 53340
rect 86032 53280 86096 53284
rect 86112 53340 86176 53344
rect 86112 53284 86116 53340
rect 86116 53284 86172 53340
rect 86172 53284 86176 53340
rect 86112 53280 86176 53284
rect 86192 53340 86256 53344
rect 86192 53284 86196 53340
rect 86196 53284 86252 53340
rect 86252 53284 86256 53340
rect 86192 53280 86256 53284
rect 89952 53340 90016 53344
rect 89952 53284 89956 53340
rect 89956 53284 90012 53340
rect 90012 53284 90016 53340
rect 89952 53280 90016 53284
rect 90032 53340 90096 53344
rect 90032 53284 90036 53340
rect 90036 53284 90092 53340
rect 90092 53284 90096 53340
rect 90032 53280 90096 53284
rect 90112 53340 90176 53344
rect 90112 53284 90116 53340
rect 90116 53284 90172 53340
rect 90172 53284 90176 53340
rect 90112 53280 90176 53284
rect 90192 53340 90256 53344
rect 90192 53284 90196 53340
rect 90196 53284 90252 53340
rect 90252 53284 90256 53340
rect 90192 53280 90256 53284
rect 3952 52796 4016 52800
rect 3952 52740 3956 52796
rect 3956 52740 4012 52796
rect 4012 52740 4016 52796
rect 3952 52736 4016 52740
rect 4032 52796 4096 52800
rect 4032 52740 4036 52796
rect 4036 52740 4092 52796
rect 4092 52740 4096 52796
rect 4032 52736 4096 52740
rect 4112 52796 4176 52800
rect 4112 52740 4116 52796
rect 4116 52740 4172 52796
rect 4172 52740 4176 52796
rect 4112 52736 4176 52740
rect 4192 52796 4256 52800
rect 4192 52740 4196 52796
rect 4196 52740 4252 52796
rect 4252 52740 4256 52796
rect 4192 52736 4256 52740
rect 87952 52796 88016 52800
rect 87952 52740 87956 52796
rect 87956 52740 88012 52796
rect 88012 52740 88016 52796
rect 87952 52736 88016 52740
rect 88032 52796 88096 52800
rect 88032 52740 88036 52796
rect 88036 52740 88092 52796
rect 88092 52740 88096 52796
rect 88032 52736 88096 52740
rect 88112 52796 88176 52800
rect 88112 52740 88116 52796
rect 88116 52740 88172 52796
rect 88172 52740 88176 52796
rect 88112 52736 88176 52740
rect 88192 52796 88256 52800
rect 88192 52740 88196 52796
rect 88196 52740 88252 52796
rect 88252 52740 88256 52796
rect 88192 52736 88256 52740
rect 1952 52252 2016 52256
rect 1952 52196 1956 52252
rect 1956 52196 2012 52252
rect 2012 52196 2016 52252
rect 1952 52192 2016 52196
rect 2032 52252 2096 52256
rect 2032 52196 2036 52252
rect 2036 52196 2092 52252
rect 2092 52196 2096 52252
rect 2032 52192 2096 52196
rect 2112 52252 2176 52256
rect 2112 52196 2116 52252
rect 2116 52196 2172 52252
rect 2172 52196 2176 52252
rect 2112 52192 2176 52196
rect 2192 52252 2256 52256
rect 2192 52196 2196 52252
rect 2196 52196 2252 52252
rect 2252 52196 2256 52252
rect 2192 52192 2256 52196
rect 85952 52252 86016 52256
rect 85952 52196 85956 52252
rect 85956 52196 86012 52252
rect 86012 52196 86016 52252
rect 85952 52192 86016 52196
rect 86032 52252 86096 52256
rect 86032 52196 86036 52252
rect 86036 52196 86092 52252
rect 86092 52196 86096 52252
rect 86032 52192 86096 52196
rect 86112 52252 86176 52256
rect 86112 52196 86116 52252
rect 86116 52196 86172 52252
rect 86172 52196 86176 52252
rect 86112 52192 86176 52196
rect 86192 52252 86256 52256
rect 86192 52196 86196 52252
rect 86196 52196 86252 52252
rect 86252 52196 86256 52252
rect 86192 52192 86256 52196
rect 89952 52252 90016 52256
rect 89952 52196 89956 52252
rect 89956 52196 90012 52252
rect 90012 52196 90016 52252
rect 89952 52192 90016 52196
rect 90032 52252 90096 52256
rect 90032 52196 90036 52252
rect 90036 52196 90092 52252
rect 90092 52196 90096 52252
rect 90032 52192 90096 52196
rect 90112 52252 90176 52256
rect 90112 52196 90116 52252
rect 90116 52196 90172 52252
rect 90172 52196 90176 52252
rect 90112 52192 90176 52196
rect 90192 52252 90256 52256
rect 90192 52196 90196 52252
rect 90196 52196 90252 52252
rect 90252 52196 90256 52252
rect 90192 52192 90256 52196
rect 3952 51708 4016 51712
rect 3952 51652 3956 51708
rect 3956 51652 4012 51708
rect 4012 51652 4016 51708
rect 3952 51648 4016 51652
rect 4032 51708 4096 51712
rect 4032 51652 4036 51708
rect 4036 51652 4092 51708
rect 4092 51652 4096 51708
rect 4032 51648 4096 51652
rect 4112 51708 4176 51712
rect 4112 51652 4116 51708
rect 4116 51652 4172 51708
rect 4172 51652 4176 51708
rect 4112 51648 4176 51652
rect 4192 51708 4256 51712
rect 4192 51652 4196 51708
rect 4196 51652 4252 51708
rect 4252 51652 4256 51708
rect 4192 51648 4256 51652
rect 87952 51708 88016 51712
rect 87952 51652 87956 51708
rect 87956 51652 88012 51708
rect 88012 51652 88016 51708
rect 87952 51648 88016 51652
rect 88032 51708 88096 51712
rect 88032 51652 88036 51708
rect 88036 51652 88092 51708
rect 88092 51652 88096 51708
rect 88032 51648 88096 51652
rect 88112 51708 88176 51712
rect 88112 51652 88116 51708
rect 88116 51652 88172 51708
rect 88172 51652 88176 51708
rect 88112 51648 88176 51652
rect 88192 51708 88256 51712
rect 88192 51652 88196 51708
rect 88196 51652 88252 51708
rect 88252 51652 88256 51708
rect 88192 51648 88256 51652
rect 83780 51308 83844 51372
rect 1952 51164 2016 51168
rect 1952 51108 1956 51164
rect 1956 51108 2012 51164
rect 2012 51108 2016 51164
rect 1952 51104 2016 51108
rect 2032 51164 2096 51168
rect 2032 51108 2036 51164
rect 2036 51108 2092 51164
rect 2092 51108 2096 51164
rect 2032 51104 2096 51108
rect 2112 51164 2176 51168
rect 2112 51108 2116 51164
rect 2116 51108 2172 51164
rect 2172 51108 2176 51164
rect 2112 51104 2176 51108
rect 2192 51164 2256 51168
rect 2192 51108 2196 51164
rect 2196 51108 2252 51164
rect 2252 51108 2256 51164
rect 2192 51104 2256 51108
rect 85952 51164 86016 51168
rect 85952 51108 85956 51164
rect 85956 51108 86012 51164
rect 86012 51108 86016 51164
rect 85952 51104 86016 51108
rect 86032 51164 86096 51168
rect 86032 51108 86036 51164
rect 86036 51108 86092 51164
rect 86092 51108 86096 51164
rect 86032 51104 86096 51108
rect 86112 51164 86176 51168
rect 86112 51108 86116 51164
rect 86116 51108 86172 51164
rect 86172 51108 86176 51164
rect 86112 51104 86176 51108
rect 86192 51164 86256 51168
rect 86192 51108 86196 51164
rect 86196 51108 86252 51164
rect 86252 51108 86256 51164
rect 86192 51104 86256 51108
rect 89952 51164 90016 51168
rect 89952 51108 89956 51164
rect 89956 51108 90012 51164
rect 90012 51108 90016 51164
rect 89952 51104 90016 51108
rect 90032 51164 90096 51168
rect 90032 51108 90036 51164
rect 90036 51108 90092 51164
rect 90092 51108 90096 51164
rect 90032 51104 90096 51108
rect 90112 51164 90176 51168
rect 90112 51108 90116 51164
rect 90116 51108 90172 51164
rect 90172 51108 90176 51164
rect 90112 51104 90176 51108
rect 90192 51164 90256 51168
rect 90192 51108 90196 51164
rect 90196 51108 90252 51164
rect 90252 51108 90256 51164
rect 90192 51104 90256 51108
rect 3952 50620 4016 50624
rect 3952 50564 3956 50620
rect 3956 50564 4012 50620
rect 4012 50564 4016 50620
rect 3952 50560 4016 50564
rect 4032 50620 4096 50624
rect 4032 50564 4036 50620
rect 4036 50564 4092 50620
rect 4092 50564 4096 50620
rect 4032 50560 4096 50564
rect 4112 50620 4176 50624
rect 4112 50564 4116 50620
rect 4116 50564 4172 50620
rect 4172 50564 4176 50620
rect 4112 50560 4176 50564
rect 4192 50620 4256 50624
rect 4192 50564 4196 50620
rect 4196 50564 4252 50620
rect 4252 50564 4256 50620
rect 4192 50560 4256 50564
rect 87952 50620 88016 50624
rect 87952 50564 87956 50620
rect 87956 50564 88012 50620
rect 88012 50564 88016 50620
rect 87952 50560 88016 50564
rect 88032 50620 88096 50624
rect 88032 50564 88036 50620
rect 88036 50564 88092 50620
rect 88092 50564 88096 50620
rect 88032 50560 88096 50564
rect 88112 50620 88176 50624
rect 88112 50564 88116 50620
rect 88116 50564 88172 50620
rect 88172 50564 88176 50620
rect 88112 50560 88176 50564
rect 88192 50620 88256 50624
rect 88192 50564 88196 50620
rect 88196 50564 88252 50620
rect 88252 50564 88256 50620
rect 88192 50560 88256 50564
rect 1952 50076 2016 50080
rect 1952 50020 1956 50076
rect 1956 50020 2012 50076
rect 2012 50020 2016 50076
rect 1952 50016 2016 50020
rect 2032 50076 2096 50080
rect 2032 50020 2036 50076
rect 2036 50020 2092 50076
rect 2092 50020 2096 50076
rect 2032 50016 2096 50020
rect 2112 50076 2176 50080
rect 2112 50020 2116 50076
rect 2116 50020 2172 50076
rect 2172 50020 2176 50076
rect 2112 50016 2176 50020
rect 2192 50076 2256 50080
rect 2192 50020 2196 50076
rect 2196 50020 2252 50076
rect 2252 50020 2256 50076
rect 2192 50016 2256 50020
rect 83596 49676 83660 49740
rect 85952 50076 86016 50080
rect 85952 50020 85956 50076
rect 85956 50020 86012 50076
rect 86012 50020 86016 50076
rect 85952 50016 86016 50020
rect 86032 50076 86096 50080
rect 86032 50020 86036 50076
rect 86036 50020 86092 50076
rect 86092 50020 86096 50076
rect 86032 50016 86096 50020
rect 86112 50076 86176 50080
rect 86112 50020 86116 50076
rect 86116 50020 86172 50076
rect 86172 50020 86176 50076
rect 86112 50016 86176 50020
rect 86192 50076 86256 50080
rect 86192 50020 86196 50076
rect 86196 50020 86252 50076
rect 86252 50020 86256 50076
rect 86192 50016 86256 50020
rect 89952 50076 90016 50080
rect 89952 50020 89956 50076
rect 89956 50020 90012 50076
rect 90012 50020 90016 50076
rect 89952 50016 90016 50020
rect 90032 50076 90096 50080
rect 90032 50020 90036 50076
rect 90036 50020 90092 50076
rect 90092 50020 90096 50076
rect 90032 50016 90096 50020
rect 90112 50076 90176 50080
rect 90112 50020 90116 50076
rect 90116 50020 90172 50076
rect 90172 50020 90176 50076
rect 90112 50016 90176 50020
rect 90192 50076 90256 50080
rect 90192 50020 90196 50076
rect 90196 50020 90252 50076
rect 90252 50020 90256 50076
rect 90192 50016 90256 50020
rect 3952 49532 4016 49536
rect 3952 49476 3956 49532
rect 3956 49476 4012 49532
rect 4012 49476 4016 49532
rect 3952 49472 4016 49476
rect 4032 49532 4096 49536
rect 4032 49476 4036 49532
rect 4036 49476 4092 49532
rect 4092 49476 4096 49532
rect 4032 49472 4096 49476
rect 4112 49532 4176 49536
rect 4112 49476 4116 49532
rect 4116 49476 4172 49532
rect 4172 49476 4176 49532
rect 4112 49472 4176 49476
rect 4192 49532 4256 49536
rect 4192 49476 4196 49532
rect 4196 49476 4252 49532
rect 4252 49476 4256 49532
rect 4192 49472 4256 49476
rect 87952 49532 88016 49536
rect 87952 49476 87956 49532
rect 87956 49476 88012 49532
rect 88012 49476 88016 49532
rect 87952 49472 88016 49476
rect 88032 49532 88096 49536
rect 88032 49476 88036 49532
rect 88036 49476 88092 49532
rect 88092 49476 88096 49532
rect 88032 49472 88096 49476
rect 88112 49532 88176 49536
rect 88112 49476 88116 49532
rect 88116 49476 88172 49532
rect 88172 49476 88176 49532
rect 88112 49472 88176 49476
rect 88192 49532 88256 49536
rect 88192 49476 88196 49532
rect 88196 49476 88252 49532
rect 88252 49476 88256 49532
rect 88192 49472 88256 49476
rect 1952 48988 2016 48992
rect 1952 48932 1956 48988
rect 1956 48932 2012 48988
rect 2012 48932 2016 48988
rect 1952 48928 2016 48932
rect 2032 48988 2096 48992
rect 2032 48932 2036 48988
rect 2036 48932 2092 48988
rect 2092 48932 2096 48988
rect 2032 48928 2096 48932
rect 2112 48988 2176 48992
rect 2112 48932 2116 48988
rect 2116 48932 2172 48988
rect 2172 48932 2176 48988
rect 2112 48928 2176 48932
rect 2192 48988 2256 48992
rect 2192 48932 2196 48988
rect 2196 48932 2252 48988
rect 2252 48932 2256 48988
rect 2192 48928 2256 48932
rect 85952 48988 86016 48992
rect 85952 48932 85956 48988
rect 85956 48932 86012 48988
rect 86012 48932 86016 48988
rect 85952 48928 86016 48932
rect 86032 48988 86096 48992
rect 86032 48932 86036 48988
rect 86036 48932 86092 48988
rect 86092 48932 86096 48988
rect 86032 48928 86096 48932
rect 86112 48988 86176 48992
rect 86112 48932 86116 48988
rect 86116 48932 86172 48988
rect 86172 48932 86176 48988
rect 86112 48928 86176 48932
rect 86192 48988 86256 48992
rect 86192 48932 86196 48988
rect 86196 48932 86252 48988
rect 86252 48932 86256 48988
rect 86192 48928 86256 48932
rect 89952 48988 90016 48992
rect 89952 48932 89956 48988
rect 89956 48932 90012 48988
rect 90012 48932 90016 48988
rect 89952 48928 90016 48932
rect 90032 48988 90096 48992
rect 90032 48932 90036 48988
rect 90036 48932 90092 48988
rect 90092 48932 90096 48988
rect 90032 48928 90096 48932
rect 90112 48988 90176 48992
rect 90112 48932 90116 48988
rect 90116 48932 90172 48988
rect 90172 48932 90176 48988
rect 90112 48928 90176 48932
rect 90192 48988 90256 48992
rect 90192 48932 90196 48988
rect 90196 48932 90252 48988
rect 90252 48932 90256 48988
rect 90192 48928 90256 48932
rect 3952 48444 4016 48448
rect 3952 48388 3956 48444
rect 3956 48388 4012 48444
rect 4012 48388 4016 48444
rect 3952 48384 4016 48388
rect 4032 48444 4096 48448
rect 4032 48388 4036 48444
rect 4036 48388 4092 48444
rect 4092 48388 4096 48444
rect 4032 48384 4096 48388
rect 4112 48444 4176 48448
rect 4112 48388 4116 48444
rect 4116 48388 4172 48444
rect 4172 48388 4176 48444
rect 4112 48384 4176 48388
rect 4192 48444 4256 48448
rect 4192 48388 4196 48444
rect 4196 48388 4252 48444
rect 4252 48388 4256 48444
rect 4192 48384 4256 48388
rect 87952 48444 88016 48448
rect 87952 48388 87956 48444
rect 87956 48388 88012 48444
rect 88012 48388 88016 48444
rect 87952 48384 88016 48388
rect 88032 48444 88096 48448
rect 88032 48388 88036 48444
rect 88036 48388 88092 48444
rect 88092 48388 88096 48444
rect 88032 48384 88096 48388
rect 88112 48444 88176 48448
rect 88112 48388 88116 48444
rect 88116 48388 88172 48444
rect 88172 48388 88176 48444
rect 88112 48384 88176 48388
rect 88192 48444 88256 48448
rect 88192 48388 88196 48444
rect 88196 48388 88252 48444
rect 88252 48388 88256 48444
rect 88192 48384 88256 48388
rect 1952 47900 2016 47904
rect 1952 47844 1956 47900
rect 1956 47844 2012 47900
rect 2012 47844 2016 47900
rect 1952 47840 2016 47844
rect 2032 47900 2096 47904
rect 2032 47844 2036 47900
rect 2036 47844 2092 47900
rect 2092 47844 2096 47900
rect 2032 47840 2096 47844
rect 2112 47900 2176 47904
rect 2112 47844 2116 47900
rect 2116 47844 2172 47900
rect 2172 47844 2176 47900
rect 2112 47840 2176 47844
rect 2192 47900 2256 47904
rect 2192 47844 2196 47900
rect 2196 47844 2252 47900
rect 2252 47844 2256 47900
rect 2192 47840 2256 47844
rect 85952 47900 86016 47904
rect 85952 47844 85956 47900
rect 85956 47844 86012 47900
rect 86012 47844 86016 47900
rect 85952 47840 86016 47844
rect 86032 47900 86096 47904
rect 86032 47844 86036 47900
rect 86036 47844 86092 47900
rect 86092 47844 86096 47900
rect 86032 47840 86096 47844
rect 86112 47900 86176 47904
rect 86112 47844 86116 47900
rect 86116 47844 86172 47900
rect 86172 47844 86176 47900
rect 86112 47840 86176 47844
rect 86192 47900 86256 47904
rect 86192 47844 86196 47900
rect 86196 47844 86252 47900
rect 86252 47844 86256 47900
rect 86192 47840 86256 47844
rect 89952 47900 90016 47904
rect 89952 47844 89956 47900
rect 89956 47844 90012 47900
rect 90012 47844 90016 47900
rect 89952 47840 90016 47844
rect 90032 47900 90096 47904
rect 90032 47844 90036 47900
rect 90036 47844 90092 47900
rect 90092 47844 90096 47900
rect 90032 47840 90096 47844
rect 90112 47900 90176 47904
rect 90112 47844 90116 47900
rect 90116 47844 90172 47900
rect 90172 47844 90176 47900
rect 90112 47840 90176 47844
rect 90192 47900 90256 47904
rect 90192 47844 90196 47900
rect 90196 47844 90252 47900
rect 90252 47844 90256 47900
rect 90192 47840 90256 47844
rect 3952 47356 4016 47360
rect 3952 47300 3956 47356
rect 3956 47300 4012 47356
rect 4012 47300 4016 47356
rect 3952 47296 4016 47300
rect 4032 47356 4096 47360
rect 4032 47300 4036 47356
rect 4036 47300 4092 47356
rect 4092 47300 4096 47356
rect 4032 47296 4096 47300
rect 4112 47356 4176 47360
rect 4112 47300 4116 47356
rect 4116 47300 4172 47356
rect 4172 47300 4176 47356
rect 4112 47296 4176 47300
rect 4192 47356 4256 47360
rect 4192 47300 4196 47356
rect 4196 47300 4252 47356
rect 4252 47300 4256 47356
rect 4192 47296 4256 47300
rect 87952 47356 88016 47360
rect 87952 47300 87956 47356
rect 87956 47300 88012 47356
rect 88012 47300 88016 47356
rect 87952 47296 88016 47300
rect 88032 47356 88096 47360
rect 88032 47300 88036 47356
rect 88036 47300 88092 47356
rect 88092 47300 88096 47356
rect 88032 47296 88096 47300
rect 88112 47356 88176 47360
rect 88112 47300 88116 47356
rect 88116 47300 88172 47356
rect 88172 47300 88176 47356
rect 88112 47296 88176 47300
rect 88192 47356 88256 47360
rect 88192 47300 88196 47356
rect 88196 47300 88252 47356
rect 88252 47300 88256 47356
rect 88192 47296 88256 47300
rect 1952 46812 2016 46816
rect 1952 46756 1956 46812
rect 1956 46756 2012 46812
rect 2012 46756 2016 46812
rect 1952 46752 2016 46756
rect 2032 46812 2096 46816
rect 2032 46756 2036 46812
rect 2036 46756 2092 46812
rect 2092 46756 2096 46812
rect 2032 46752 2096 46756
rect 2112 46812 2176 46816
rect 2112 46756 2116 46812
rect 2116 46756 2172 46812
rect 2172 46756 2176 46812
rect 2112 46752 2176 46756
rect 2192 46812 2256 46816
rect 2192 46756 2196 46812
rect 2196 46756 2252 46812
rect 2252 46756 2256 46812
rect 2192 46752 2256 46756
rect 85952 46812 86016 46816
rect 85952 46756 85956 46812
rect 85956 46756 86012 46812
rect 86012 46756 86016 46812
rect 85952 46752 86016 46756
rect 86032 46812 86096 46816
rect 86032 46756 86036 46812
rect 86036 46756 86092 46812
rect 86092 46756 86096 46812
rect 86032 46752 86096 46756
rect 86112 46812 86176 46816
rect 86112 46756 86116 46812
rect 86116 46756 86172 46812
rect 86172 46756 86176 46812
rect 86112 46752 86176 46756
rect 86192 46812 86256 46816
rect 86192 46756 86196 46812
rect 86196 46756 86252 46812
rect 86252 46756 86256 46812
rect 86192 46752 86256 46756
rect 89952 46812 90016 46816
rect 89952 46756 89956 46812
rect 89956 46756 90012 46812
rect 90012 46756 90016 46812
rect 89952 46752 90016 46756
rect 90032 46812 90096 46816
rect 90032 46756 90036 46812
rect 90036 46756 90092 46812
rect 90092 46756 90096 46812
rect 90032 46752 90096 46756
rect 90112 46812 90176 46816
rect 90112 46756 90116 46812
rect 90116 46756 90172 46812
rect 90172 46756 90176 46812
rect 90112 46752 90176 46756
rect 90192 46812 90256 46816
rect 90192 46756 90196 46812
rect 90196 46756 90252 46812
rect 90252 46756 90256 46812
rect 90192 46752 90256 46756
rect 3952 46268 4016 46272
rect 3952 46212 3956 46268
rect 3956 46212 4012 46268
rect 4012 46212 4016 46268
rect 3952 46208 4016 46212
rect 4032 46268 4096 46272
rect 4032 46212 4036 46268
rect 4036 46212 4092 46268
rect 4092 46212 4096 46268
rect 4032 46208 4096 46212
rect 4112 46268 4176 46272
rect 4112 46212 4116 46268
rect 4116 46212 4172 46268
rect 4172 46212 4176 46268
rect 4112 46208 4176 46212
rect 4192 46268 4256 46272
rect 4192 46212 4196 46268
rect 4196 46212 4252 46268
rect 4252 46212 4256 46268
rect 4192 46208 4256 46212
rect 87952 46268 88016 46272
rect 87952 46212 87956 46268
rect 87956 46212 88012 46268
rect 88012 46212 88016 46268
rect 87952 46208 88016 46212
rect 88032 46268 88096 46272
rect 88032 46212 88036 46268
rect 88036 46212 88092 46268
rect 88092 46212 88096 46268
rect 88032 46208 88096 46212
rect 88112 46268 88176 46272
rect 88112 46212 88116 46268
rect 88116 46212 88172 46268
rect 88172 46212 88176 46268
rect 88112 46208 88176 46212
rect 88192 46268 88256 46272
rect 88192 46212 88196 46268
rect 88196 46212 88252 46268
rect 88252 46212 88256 46268
rect 88192 46208 88256 46212
rect 1952 45724 2016 45728
rect 1952 45668 1956 45724
rect 1956 45668 2012 45724
rect 2012 45668 2016 45724
rect 1952 45664 2016 45668
rect 2032 45724 2096 45728
rect 2032 45668 2036 45724
rect 2036 45668 2092 45724
rect 2092 45668 2096 45724
rect 2032 45664 2096 45668
rect 2112 45724 2176 45728
rect 2112 45668 2116 45724
rect 2116 45668 2172 45724
rect 2172 45668 2176 45724
rect 2112 45664 2176 45668
rect 2192 45724 2256 45728
rect 2192 45668 2196 45724
rect 2196 45668 2252 45724
rect 2252 45668 2256 45724
rect 2192 45664 2256 45668
rect 85952 45724 86016 45728
rect 85952 45668 85956 45724
rect 85956 45668 86012 45724
rect 86012 45668 86016 45724
rect 85952 45664 86016 45668
rect 86032 45724 86096 45728
rect 86032 45668 86036 45724
rect 86036 45668 86092 45724
rect 86092 45668 86096 45724
rect 86032 45664 86096 45668
rect 86112 45724 86176 45728
rect 86112 45668 86116 45724
rect 86116 45668 86172 45724
rect 86172 45668 86176 45724
rect 86112 45664 86176 45668
rect 86192 45724 86256 45728
rect 86192 45668 86196 45724
rect 86196 45668 86252 45724
rect 86252 45668 86256 45724
rect 86192 45664 86256 45668
rect 89952 45724 90016 45728
rect 89952 45668 89956 45724
rect 89956 45668 90012 45724
rect 90012 45668 90016 45724
rect 89952 45664 90016 45668
rect 90032 45724 90096 45728
rect 90032 45668 90036 45724
rect 90036 45668 90092 45724
rect 90092 45668 90096 45724
rect 90032 45664 90096 45668
rect 90112 45724 90176 45728
rect 90112 45668 90116 45724
rect 90116 45668 90172 45724
rect 90172 45668 90176 45724
rect 90112 45664 90176 45668
rect 90192 45724 90256 45728
rect 90192 45668 90196 45724
rect 90196 45668 90252 45724
rect 90252 45668 90256 45724
rect 90192 45664 90256 45668
rect 83412 45460 83476 45524
rect 3952 45180 4016 45184
rect 3952 45124 3956 45180
rect 3956 45124 4012 45180
rect 4012 45124 4016 45180
rect 3952 45120 4016 45124
rect 4032 45180 4096 45184
rect 4032 45124 4036 45180
rect 4036 45124 4092 45180
rect 4092 45124 4096 45180
rect 4032 45120 4096 45124
rect 4112 45180 4176 45184
rect 4112 45124 4116 45180
rect 4116 45124 4172 45180
rect 4172 45124 4176 45180
rect 4112 45120 4176 45124
rect 4192 45180 4256 45184
rect 4192 45124 4196 45180
rect 4196 45124 4252 45180
rect 4252 45124 4256 45180
rect 4192 45120 4256 45124
rect 87952 45180 88016 45184
rect 87952 45124 87956 45180
rect 87956 45124 88012 45180
rect 88012 45124 88016 45180
rect 87952 45120 88016 45124
rect 88032 45180 88096 45184
rect 88032 45124 88036 45180
rect 88036 45124 88092 45180
rect 88092 45124 88096 45180
rect 88032 45120 88096 45124
rect 88112 45180 88176 45184
rect 88112 45124 88116 45180
rect 88116 45124 88172 45180
rect 88172 45124 88176 45180
rect 88112 45120 88176 45124
rect 88192 45180 88256 45184
rect 88192 45124 88196 45180
rect 88196 45124 88252 45180
rect 88252 45124 88256 45180
rect 88192 45120 88256 45124
rect 1952 44636 2016 44640
rect 1952 44580 1956 44636
rect 1956 44580 2012 44636
rect 2012 44580 2016 44636
rect 1952 44576 2016 44580
rect 2032 44636 2096 44640
rect 2032 44580 2036 44636
rect 2036 44580 2092 44636
rect 2092 44580 2096 44636
rect 2032 44576 2096 44580
rect 2112 44636 2176 44640
rect 2112 44580 2116 44636
rect 2116 44580 2172 44636
rect 2172 44580 2176 44636
rect 2112 44576 2176 44580
rect 2192 44636 2256 44640
rect 2192 44580 2196 44636
rect 2196 44580 2252 44636
rect 2252 44580 2256 44636
rect 2192 44576 2256 44580
rect 85952 44636 86016 44640
rect 85952 44580 85956 44636
rect 85956 44580 86012 44636
rect 86012 44580 86016 44636
rect 85952 44576 86016 44580
rect 86032 44636 86096 44640
rect 86032 44580 86036 44636
rect 86036 44580 86092 44636
rect 86092 44580 86096 44636
rect 86032 44576 86096 44580
rect 86112 44636 86176 44640
rect 86112 44580 86116 44636
rect 86116 44580 86172 44636
rect 86172 44580 86176 44636
rect 86112 44576 86176 44580
rect 86192 44636 86256 44640
rect 86192 44580 86196 44636
rect 86196 44580 86252 44636
rect 86252 44580 86256 44636
rect 86192 44576 86256 44580
rect 89952 44636 90016 44640
rect 89952 44580 89956 44636
rect 89956 44580 90012 44636
rect 90012 44580 90016 44636
rect 89952 44576 90016 44580
rect 90032 44636 90096 44640
rect 90032 44580 90036 44636
rect 90036 44580 90092 44636
rect 90092 44580 90096 44636
rect 90032 44576 90096 44580
rect 90112 44636 90176 44640
rect 90112 44580 90116 44636
rect 90116 44580 90172 44636
rect 90172 44580 90176 44636
rect 90112 44576 90176 44580
rect 90192 44636 90256 44640
rect 90192 44580 90196 44636
rect 90196 44580 90252 44636
rect 90252 44580 90256 44636
rect 90192 44576 90256 44580
rect 3952 44092 4016 44096
rect 3952 44036 3956 44092
rect 3956 44036 4012 44092
rect 4012 44036 4016 44092
rect 3952 44032 4016 44036
rect 4032 44092 4096 44096
rect 4032 44036 4036 44092
rect 4036 44036 4092 44092
rect 4092 44036 4096 44092
rect 4032 44032 4096 44036
rect 4112 44092 4176 44096
rect 4112 44036 4116 44092
rect 4116 44036 4172 44092
rect 4172 44036 4176 44092
rect 4112 44032 4176 44036
rect 4192 44092 4256 44096
rect 4192 44036 4196 44092
rect 4196 44036 4252 44092
rect 4252 44036 4256 44092
rect 4192 44032 4256 44036
rect 87952 44092 88016 44096
rect 87952 44036 87956 44092
rect 87956 44036 88012 44092
rect 88012 44036 88016 44092
rect 87952 44032 88016 44036
rect 88032 44092 88096 44096
rect 88032 44036 88036 44092
rect 88036 44036 88092 44092
rect 88092 44036 88096 44092
rect 88032 44032 88096 44036
rect 88112 44092 88176 44096
rect 88112 44036 88116 44092
rect 88116 44036 88172 44092
rect 88172 44036 88176 44092
rect 88112 44032 88176 44036
rect 88192 44092 88256 44096
rect 88192 44036 88196 44092
rect 88196 44036 88252 44092
rect 88252 44036 88256 44092
rect 88192 44032 88256 44036
rect 1952 43548 2016 43552
rect 1952 43492 1956 43548
rect 1956 43492 2012 43548
rect 2012 43492 2016 43548
rect 1952 43488 2016 43492
rect 2032 43548 2096 43552
rect 2032 43492 2036 43548
rect 2036 43492 2092 43548
rect 2092 43492 2096 43548
rect 2032 43488 2096 43492
rect 2112 43548 2176 43552
rect 2112 43492 2116 43548
rect 2116 43492 2172 43548
rect 2172 43492 2176 43548
rect 2112 43488 2176 43492
rect 2192 43548 2256 43552
rect 2192 43492 2196 43548
rect 2196 43492 2252 43548
rect 2252 43492 2256 43548
rect 2192 43488 2256 43492
rect 85952 43548 86016 43552
rect 85952 43492 85956 43548
rect 85956 43492 86012 43548
rect 86012 43492 86016 43548
rect 85952 43488 86016 43492
rect 86032 43548 86096 43552
rect 86032 43492 86036 43548
rect 86036 43492 86092 43548
rect 86092 43492 86096 43548
rect 86032 43488 86096 43492
rect 86112 43548 86176 43552
rect 86112 43492 86116 43548
rect 86116 43492 86172 43548
rect 86172 43492 86176 43548
rect 86112 43488 86176 43492
rect 86192 43548 86256 43552
rect 86192 43492 86196 43548
rect 86196 43492 86252 43548
rect 86252 43492 86256 43548
rect 86192 43488 86256 43492
rect 89952 43548 90016 43552
rect 89952 43492 89956 43548
rect 89956 43492 90012 43548
rect 90012 43492 90016 43548
rect 89952 43488 90016 43492
rect 90032 43548 90096 43552
rect 90032 43492 90036 43548
rect 90036 43492 90092 43548
rect 90092 43492 90096 43548
rect 90032 43488 90096 43492
rect 90112 43548 90176 43552
rect 90112 43492 90116 43548
rect 90116 43492 90172 43548
rect 90172 43492 90176 43548
rect 90112 43488 90176 43492
rect 90192 43548 90256 43552
rect 90192 43492 90196 43548
rect 90196 43492 90252 43548
rect 90252 43492 90256 43548
rect 90192 43488 90256 43492
rect 3952 43004 4016 43008
rect 3952 42948 3956 43004
rect 3956 42948 4012 43004
rect 4012 42948 4016 43004
rect 3952 42944 4016 42948
rect 4032 43004 4096 43008
rect 4032 42948 4036 43004
rect 4036 42948 4092 43004
rect 4092 42948 4096 43004
rect 4032 42944 4096 42948
rect 4112 43004 4176 43008
rect 4112 42948 4116 43004
rect 4116 42948 4172 43004
rect 4172 42948 4176 43004
rect 4112 42944 4176 42948
rect 4192 43004 4256 43008
rect 4192 42948 4196 43004
rect 4196 42948 4252 43004
rect 4252 42948 4256 43004
rect 4192 42944 4256 42948
rect 87952 43004 88016 43008
rect 87952 42948 87956 43004
rect 87956 42948 88012 43004
rect 88012 42948 88016 43004
rect 87952 42944 88016 42948
rect 88032 43004 88096 43008
rect 88032 42948 88036 43004
rect 88036 42948 88092 43004
rect 88092 42948 88096 43004
rect 88032 42944 88096 42948
rect 88112 43004 88176 43008
rect 88112 42948 88116 43004
rect 88116 42948 88172 43004
rect 88172 42948 88176 43004
rect 88112 42944 88176 42948
rect 88192 43004 88256 43008
rect 88192 42948 88196 43004
rect 88196 42948 88252 43004
rect 88252 42948 88256 43004
rect 88192 42944 88256 42948
rect 1952 42460 2016 42464
rect 1952 42404 1956 42460
rect 1956 42404 2012 42460
rect 2012 42404 2016 42460
rect 1952 42400 2016 42404
rect 2032 42460 2096 42464
rect 2032 42404 2036 42460
rect 2036 42404 2092 42460
rect 2092 42404 2096 42460
rect 2032 42400 2096 42404
rect 2112 42460 2176 42464
rect 2112 42404 2116 42460
rect 2116 42404 2172 42460
rect 2172 42404 2176 42460
rect 2112 42400 2176 42404
rect 2192 42460 2256 42464
rect 2192 42404 2196 42460
rect 2196 42404 2252 42460
rect 2252 42404 2256 42460
rect 2192 42400 2256 42404
rect 85952 42460 86016 42464
rect 85952 42404 85956 42460
rect 85956 42404 86012 42460
rect 86012 42404 86016 42460
rect 85952 42400 86016 42404
rect 86032 42460 86096 42464
rect 86032 42404 86036 42460
rect 86036 42404 86092 42460
rect 86092 42404 86096 42460
rect 86032 42400 86096 42404
rect 86112 42460 86176 42464
rect 86112 42404 86116 42460
rect 86116 42404 86172 42460
rect 86172 42404 86176 42460
rect 86112 42400 86176 42404
rect 86192 42460 86256 42464
rect 86192 42404 86196 42460
rect 86196 42404 86252 42460
rect 86252 42404 86256 42460
rect 86192 42400 86256 42404
rect 89952 42460 90016 42464
rect 89952 42404 89956 42460
rect 89956 42404 90012 42460
rect 90012 42404 90016 42460
rect 89952 42400 90016 42404
rect 90032 42460 90096 42464
rect 90032 42404 90036 42460
rect 90036 42404 90092 42460
rect 90092 42404 90096 42460
rect 90032 42400 90096 42404
rect 90112 42460 90176 42464
rect 90112 42404 90116 42460
rect 90116 42404 90172 42460
rect 90172 42404 90176 42460
rect 90112 42400 90176 42404
rect 90192 42460 90256 42464
rect 90192 42404 90196 42460
rect 90196 42404 90252 42460
rect 90252 42404 90256 42460
rect 90192 42400 90256 42404
rect 3952 41916 4016 41920
rect 3952 41860 3956 41916
rect 3956 41860 4012 41916
rect 4012 41860 4016 41916
rect 3952 41856 4016 41860
rect 4032 41916 4096 41920
rect 4032 41860 4036 41916
rect 4036 41860 4092 41916
rect 4092 41860 4096 41916
rect 4032 41856 4096 41860
rect 4112 41916 4176 41920
rect 4112 41860 4116 41916
rect 4116 41860 4172 41916
rect 4172 41860 4176 41916
rect 4112 41856 4176 41860
rect 4192 41916 4256 41920
rect 4192 41860 4196 41916
rect 4196 41860 4252 41916
rect 4252 41860 4256 41916
rect 4192 41856 4256 41860
rect 87952 41916 88016 41920
rect 87952 41860 87956 41916
rect 87956 41860 88012 41916
rect 88012 41860 88016 41916
rect 87952 41856 88016 41860
rect 88032 41916 88096 41920
rect 88032 41860 88036 41916
rect 88036 41860 88092 41916
rect 88092 41860 88096 41916
rect 88032 41856 88096 41860
rect 88112 41916 88176 41920
rect 88112 41860 88116 41916
rect 88116 41860 88172 41916
rect 88172 41860 88176 41916
rect 88112 41856 88176 41860
rect 88192 41916 88256 41920
rect 88192 41860 88196 41916
rect 88196 41860 88252 41916
rect 88252 41860 88256 41916
rect 88192 41856 88256 41860
rect 1952 41372 2016 41376
rect 1952 41316 1956 41372
rect 1956 41316 2012 41372
rect 2012 41316 2016 41372
rect 1952 41312 2016 41316
rect 2032 41372 2096 41376
rect 2032 41316 2036 41372
rect 2036 41316 2092 41372
rect 2092 41316 2096 41372
rect 2032 41312 2096 41316
rect 2112 41372 2176 41376
rect 2112 41316 2116 41372
rect 2116 41316 2172 41372
rect 2172 41316 2176 41372
rect 2112 41312 2176 41316
rect 2192 41372 2256 41376
rect 2192 41316 2196 41372
rect 2196 41316 2252 41372
rect 2252 41316 2256 41372
rect 2192 41312 2256 41316
rect 85952 41372 86016 41376
rect 85952 41316 85956 41372
rect 85956 41316 86012 41372
rect 86012 41316 86016 41372
rect 85952 41312 86016 41316
rect 86032 41372 86096 41376
rect 86032 41316 86036 41372
rect 86036 41316 86092 41372
rect 86092 41316 86096 41372
rect 86032 41312 86096 41316
rect 86112 41372 86176 41376
rect 86112 41316 86116 41372
rect 86116 41316 86172 41372
rect 86172 41316 86176 41372
rect 86112 41312 86176 41316
rect 86192 41372 86256 41376
rect 86192 41316 86196 41372
rect 86196 41316 86252 41372
rect 86252 41316 86256 41372
rect 86192 41312 86256 41316
rect 89952 41372 90016 41376
rect 89952 41316 89956 41372
rect 89956 41316 90012 41372
rect 90012 41316 90016 41372
rect 89952 41312 90016 41316
rect 90032 41372 90096 41376
rect 90032 41316 90036 41372
rect 90036 41316 90092 41372
rect 90092 41316 90096 41372
rect 90032 41312 90096 41316
rect 90112 41372 90176 41376
rect 90112 41316 90116 41372
rect 90116 41316 90172 41372
rect 90172 41316 90176 41372
rect 90112 41312 90176 41316
rect 90192 41372 90256 41376
rect 90192 41316 90196 41372
rect 90196 41316 90252 41372
rect 90252 41316 90256 41372
rect 90192 41312 90256 41316
rect 3952 40828 4016 40832
rect 3952 40772 3956 40828
rect 3956 40772 4012 40828
rect 4012 40772 4016 40828
rect 3952 40768 4016 40772
rect 4032 40828 4096 40832
rect 4032 40772 4036 40828
rect 4036 40772 4092 40828
rect 4092 40772 4096 40828
rect 4032 40768 4096 40772
rect 4112 40828 4176 40832
rect 4112 40772 4116 40828
rect 4116 40772 4172 40828
rect 4172 40772 4176 40828
rect 4112 40768 4176 40772
rect 4192 40828 4256 40832
rect 4192 40772 4196 40828
rect 4196 40772 4252 40828
rect 4252 40772 4256 40828
rect 4192 40768 4256 40772
rect 87952 40828 88016 40832
rect 87952 40772 87956 40828
rect 87956 40772 88012 40828
rect 88012 40772 88016 40828
rect 87952 40768 88016 40772
rect 88032 40828 88096 40832
rect 88032 40772 88036 40828
rect 88036 40772 88092 40828
rect 88092 40772 88096 40828
rect 88032 40768 88096 40772
rect 88112 40828 88176 40832
rect 88112 40772 88116 40828
rect 88116 40772 88172 40828
rect 88172 40772 88176 40828
rect 88112 40768 88176 40772
rect 88192 40828 88256 40832
rect 88192 40772 88196 40828
rect 88196 40772 88252 40828
rect 88252 40772 88256 40828
rect 88192 40768 88256 40772
rect 1952 40284 2016 40288
rect 1952 40228 1956 40284
rect 1956 40228 2012 40284
rect 2012 40228 2016 40284
rect 1952 40224 2016 40228
rect 2032 40284 2096 40288
rect 2032 40228 2036 40284
rect 2036 40228 2092 40284
rect 2092 40228 2096 40284
rect 2032 40224 2096 40228
rect 2112 40284 2176 40288
rect 2112 40228 2116 40284
rect 2116 40228 2172 40284
rect 2172 40228 2176 40284
rect 2112 40224 2176 40228
rect 2192 40284 2256 40288
rect 2192 40228 2196 40284
rect 2196 40228 2252 40284
rect 2252 40228 2256 40284
rect 2192 40224 2256 40228
rect 85952 40284 86016 40288
rect 85952 40228 85956 40284
rect 85956 40228 86012 40284
rect 86012 40228 86016 40284
rect 85952 40224 86016 40228
rect 86032 40284 86096 40288
rect 86032 40228 86036 40284
rect 86036 40228 86092 40284
rect 86092 40228 86096 40284
rect 86032 40224 86096 40228
rect 86112 40284 86176 40288
rect 86112 40228 86116 40284
rect 86116 40228 86172 40284
rect 86172 40228 86176 40284
rect 86112 40224 86176 40228
rect 86192 40284 86256 40288
rect 86192 40228 86196 40284
rect 86196 40228 86252 40284
rect 86252 40228 86256 40284
rect 86192 40224 86256 40228
rect 89952 40284 90016 40288
rect 89952 40228 89956 40284
rect 89956 40228 90012 40284
rect 90012 40228 90016 40284
rect 89952 40224 90016 40228
rect 90032 40284 90096 40288
rect 90032 40228 90036 40284
rect 90036 40228 90092 40284
rect 90092 40228 90096 40284
rect 90032 40224 90096 40228
rect 90112 40284 90176 40288
rect 90112 40228 90116 40284
rect 90116 40228 90172 40284
rect 90172 40228 90176 40284
rect 90112 40224 90176 40228
rect 90192 40284 90256 40288
rect 90192 40228 90196 40284
rect 90196 40228 90252 40284
rect 90252 40228 90256 40284
rect 90192 40224 90256 40228
rect 3952 39740 4016 39744
rect 3952 39684 3956 39740
rect 3956 39684 4012 39740
rect 4012 39684 4016 39740
rect 3952 39680 4016 39684
rect 4032 39740 4096 39744
rect 4032 39684 4036 39740
rect 4036 39684 4092 39740
rect 4092 39684 4096 39740
rect 4032 39680 4096 39684
rect 4112 39740 4176 39744
rect 4112 39684 4116 39740
rect 4116 39684 4172 39740
rect 4172 39684 4176 39740
rect 4112 39680 4176 39684
rect 4192 39740 4256 39744
rect 4192 39684 4196 39740
rect 4196 39684 4252 39740
rect 4252 39684 4256 39740
rect 4192 39680 4256 39684
rect 87952 39740 88016 39744
rect 87952 39684 87956 39740
rect 87956 39684 88012 39740
rect 88012 39684 88016 39740
rect 87952 39680 88016 39684
rect 88032 39740 88096 39744
rect 88032 39684 88036 39740
rect 88036 39684 88092 39740
rect 88092 39684 88096 39740
rect 88032 39680 88096 39684
rect 88112 39740 88176 39744
rect 88112 39684 88116 39740
rect 88116 39684 88172 39740
rect 88172 39684 88176 39740
rect 88112 39680 88176 39684
rect 88192 39740 88256 39744
rect 88192 39684 88196 39740
rect 88196 39684 88252 39740
rect 88252 39684 88256 39740
rect 88192 39680 88256 39684
rect 1952 39196 2016 39200
rect 1952 39140 1956 39196
rect 1956 39140 2012 39196
rect 2012 39140 2016 39196
rect 1952 39136 2016 39140
rect 2032 39196 2096 39200
rect 2032 39140 2036 39196
rect 2036 39140 2092 39196
rect 2092 39140 2096 39196
rect 2032 39136 2096 39140
rect 2112 39196 2176 39200
rect 2112 39140 2116 39196
rect 2116 39140 2172 39196
rect 2172 39140 2176 39196
rect 2112 39136 2176 39140
rect 2192 39196 2256 39200
rect 2192 39140 2196 39196
rect 2196 39140 2252 39196
rect 2252 39140 2256 39196
rect 2192 39136 2256 39140
rect 85952 39196 86016 39200
rect 85952 39140 85956 39196
rect 85956 39140 86012 39196
rect 86012 39140 86016 39196
rect 85952 39136 86016 39140
rect 86032 39196 86096 39200
rect 86032 39140 86036 39196
rect 86036 39140 86092 39196
rect 86092 39140 86096 39196
rect 86032 39136 86096 39140
rect 86112 39196 86176 39200
rect 86112 39140 86116 39196
rect 86116 39140 86172 39196
rect 86172 39140 86176 39196
rect 86112 39136 86176 39140
rect 86192 39196 86256 39200
rect 86192 39140 86196 39196
rect 86196 39140 86252 39196
rect 86252 39140 86256 39196
rect 86192 39136 86256 39140
rect 89952 39196 90016 39200
rect 89952 39140 89956 39196
rect 89956 39140 90012 39196
rect 90012 39140 90016 39196
rect 89952 39136 90016 39140
rect 90032 39196 90096 39200
rect 90032 39140 90036 39196
rect 90036 39140 90092 39196
rect 90092 39140 90096 39196
rect 90032 39136 90096 39140
rect 90112 39196 90176 39200
rect 90112 39140 90116 39196
rect 90116 39140 90172 39196
rect 90172 39140 90176 39196
rect 90112 39136 90176 39140
rect 90192 39196 90256 39200
rect 90192 39140 90196 39196
rect 90196 39140 90252 39196
rect 90252 39140 90256 39196
rect 90192 39136 90256 39140
rect 3952 38652 4016 38656
rect 3952 38596 3956 38652
rect 3956 38596 4012 38652
rect 4012 38596 4016 38652
rect 3952 38592 4016 38596
rect 4032 38652 4096 38656
rect 4032 38596 4036 38652
rect 4036 38596 4092 38652
rect 4092 38596 4096 38652
rect 4032 38592 4096 38596
rect 4112 38652 4176 38656
rect 4112 38596 4116 38652
rect 4116 38596 4172 38652
rect 4172 38596 4176 38652
rect 4112 38592 4176 38596
rect 4192 38652 4256 38656
rect 4192 38596 4196 38652
rect 4196 38596 4252 38652
rect 4252 38596 4256 38652
rect 4192 38592 4256 38596
rect 87952 38652 88016 38656
rect 87952 38596 87956 38652
rect 87956 38596 88012 38652
rect 88012 38596 88016 38652
rect 87952 38592 88016 38596
rect 88032 38652 88096 38656
rect 88032 38596 88036 38652
rect 88036 38596 88092 38652
rect 88092 38596 88096 38652
rect 88032 38592 88096 38596
rect 88112 38652 88176 38656
rect 88112 38596 88116 38652
rect 88116 38596 88172 38652
rect 88172 38596 88176 38652
rect 88112 38592 88176 38596
rect 88192 38652 88256 38656
rect 88192 38596 88196 38652
rect 88196 38596 88252 38652
rect 88252 38596 88256 38652
rect 88192 38592 88256 38596
rect 1952 38108 2016 38112
rect 1952 38052 1956 38108
rect 1956 38052 2012 38108
rect 2012 38052 2016 38108
rect 1952 38048 2016 38052
rect 2032 38108 2096 38112
rect 2032 38052 2036 38108
rect 2036 38052 2092 38108
rect 2092 38052 2096 38108
rect 2032 38048 2096 38052
rect 2112 38108 2176 38112
rect 2112 38052 2116 38108
rect 2116 38052 2172 38108
rect 2172 38052 2176 38108
rect 2112 38048 2176 38052
rect 2192 38108 2256 38112
rect 2192 38052 2196 38108
rect 2196 38052 2252 38108
rect 2252 38052 2256 38108
rect 2192 38048 2256 38052
rect 85952 38108 86016 38112
rect 85952 38052 85956 38108
rect 85956 38052 86012 38108
rect 86012 38052 86016 38108
rect 85952 38048 86016 38052
rect 86032 38108 86096 38112
rect 86032 38052 86036 38108
rect 86036 38052 86092 38108
rect 86092 38052 86096 38108
rect 86032 38048 86096 38052
rect 86112 38108 86176 38112
rect 86112 38052 86116 38108
rect 86116 38052 86172 38108
rect 86172 38052 86176 38108
rect 86112 38048 86176 38052
rect 86192 38108 86256 38112
rect 86192 38052 86196 38108
rect 86196 38052 86252 38108
rect 86252 38052 86256 38108
rect 86192 38048 86256 38052
rect 89952 38108 90016 38112
rect 89952 38052 89956 38108
rect 89956 38052 90012 38108
rect 90012 38052 90016 38108
rect 89952 38048 90016 38052
rect 90032 38108 90096 38112
rect 90032 38052 90036 38108
rect 90036 38052 90092 38108
rect 90092 38052 90096 38108
rect 90032 38048 90096 38052
rect 90112 38108 90176 38112
rect 90112 38052 90116 38108
rect 90116 38052 90172 38108
rect 90172 38052 90176 38108
rect 90112 38048 90176 38052
rect 90192 38108 90256 38112
rect 90192 38052 90196 38108
rect 90196 38052 90252 38108
rect 90252 38052 90256 38108
rect 90192 38048 90256 38052
rect 3952 37564 4016 37568
rect 3952 37508 3956 37564
rect 3956 37508 4012 37564
rect 4012 37508 4016 37564
rect 3952 37504 4016 37508
rect 4032 37564 4096 37568
rect 4032 37508 4036 37564
rect 4036 37508 4092 37564
rect 4092 37508 4096 37564
rect 4032 37504 4096 37508
rect 4112 37564 4176 37568
rect 4112 37508 4116 37564
rect 4116 37508 4172 37564
rect 4172 37508 4176 37564
rect 4112 37504 4176 37508
rect 4192 37564 4256 37568
rect 4192 37508 4196 37564
rect 4196 37508 4252 37564
rect 4252 37508 4256 37564
rect 4192 37504 4256 37508
rect 87952 37564 88016 37568
rect 87952 37508 87956 37564
rect 87956 37508 88012 37564
rect 88012 37508 88016 37564
rect 87952 37504 88016 37508
rect 88032 37564 88096 37568
rect 88032 37508 88036 37564
rect 88036 37508 88092 37564
rect 88092 37508 88096 37564
rect 88032 37504 88096 37508
rect 88112 37564 88176 37568
rect 88112 37508 88116 37564
rect 88116 37508 88172 37564
rect 88172 37508 88176 37564
rect 88112 37504 88176 37508
rect 88192 37564 88256 37568
rect 88192 37508 88196 37564
rect 88196 37508 88252 37564
rect 88252 37508 88256 37564
rect 88192 37504 88256 37508
rect 1952 37020 2016 37024
rect 1952 36964 1956 37020
rect 1956 36964 2012 37020
rect 2012 36964 2016 37020
rect 1952 36960 2016 36964
rect 2032 37020 2096 37024
rect 2032 36964 2036 37020
rect 2036 36964 2092 37020
rect 2092 36964 2096 37020
rect 2032 36960 2096 36964
rect 2112 37020 2176 37024
rect 2112 36964 2116 37020
rect 2116 36964 2172 37020
rect 2172 36964 2176 37020
rect 2112 36960 2176 36964
rect 2192 37020 2256 37024
rect 2192 36964 2196 37020
rect 2196 36964 2252 37020
rect 2252 36964 2256 37020
rect 2192 36960 2256 36964
rect 85952 37020 86016 37024
rect 85952 36964 85956 37020
rect 85956 36964 86012 37020
rect 86012 36964 86016 37020
rect 85952 36960 86016 36964
rect 86032 37020 86096 37024
rect 86032 36964 86036 37020
rect 86036 36964 86092 37020
rect 86092 36964 86096 37020
rect 86032 36960 86096 36964
rect 86112 37020 86176 37024
rect 86112 36964 86116 37020
rect 86116 36964 86172 37020
rect 86172 36964 86176 37020
rect 86112 36960 86176 36964
rect 86192 37020 86256 37024
rect 86192 36964 86196 37020
rect 86196 36964 86252 37020
rect 86252 36964 86256 37020
rect 86192 36960 86256 36964
rect 89952 37020 90016 37024
rect 89952 36964 89956 37020
rect 89956 36964 90012 37020
rect 90012 36964 90016 37020
rect 89952 36960 90016 36964
rect 90032 37020 90096 37024
rect 90032 36964 90036 37020
rect 90036 36964 90092 37020
rect 90092 36964 90096 37020
rect 90032 36960 90096 36964
rect 90112 37020 90176 37024
rect 90112 36964 90116 37020
rect 90116 36964 90172 37020
rect 90172 36964 90176 37020
rect 90112 36960 90176 36964
rect 90192 37020 90256 37024
rect 90192 36964 90196 37020
rect 90196 36964 90252 37020
rect 90252 36964 90256 37020
rect 90192 36960 90256 36964
rect 3952 36476 4016 36480
rect 3952 36420 3956 36476
rect 3956 36420 4012 36476
rect 4012 36420 4016 36476
rect 3952 36416 4016 36420
rect 4032 36476 4096 36480
rect 4032 36420 4036 36476
rect 4036 36420 4092 36476
rect 4092 36420 4096 36476
rect 4032 36416 4096 36420
rect 4112 36476 4176 36480
rect 4112 36420 4116 36476
rect 4116 36420 4172 36476
rect 4172 36420 4176 36476
rect 4112 36416 4176 36420
rect 4192 36476 4256 36480
rect 4192 36420 4196 36476
rect 4196 36420 4252 36476
rect 4252 36420 4256 36476
rect 4192 36416 4256 36420
rect 87952 36476 88016 36480
rect 87952 36420 87956 36476
rect 87956 36420 88012 36476
rect 88012 36420 88016 36476
rect 87952 36416 88016 36420
rect 88032 36476 88096 36480
rect 88032 36420 88036 36476
rect 88036 36420 88092 36476
rect 88092 36420 88096 36476
rect 88032 36416 88096 36420
rect 88112 36476 88176 36480
rect 88112 36420 88116 36476
rect 88116 36420 88172 36476
rect 88172 36420 88176 36476
rect 88112 36416 88176 36420
rect 88192 36476 88256 36480
rect 88192 36420 88196 36476
rect 88196 36420 88252 36476
rect 88252 36420 88256 36476
rect 88192 36416 88256 36420
rect 1952 35932 2016 35936
rect 1952 35876 1956 35932
rect 1956 35876 2012 35932
rect 2012 35876 2016 35932
rect 1952 35872 2016 35876
rect 2032 35932 2096 35936
rect 2032 35876 2036 35932
rect 2036 35876 2092 35932
rect 2092 35876 2096 35932
rect 2032 35872 2096 35876
rect 2112 35932 2176 35936
rect 2112 35876 2116 35932
rect 2116 35876 2172 35932
rect 2172 35876 2176 35932
rect 2112 35872 2176 35876
rect 2192 35932 2256 35936
rect 2192 35876 2196 35932
rect 2196 35876 2252 35932
rect 2252 35876 2256 35932
rect 2192 35872 2256 35876
rect 85952 35932 86016 35936
rect 85952 35876 85956 35932
rect 85956 35876 86012 35932
rect 86012 35876 86016 35932
rect 85952 35872 86016 35876
rect 86032 35932 86096 35936
rect 86032 35876 86036 35932
rect 86036 35876 86092 35932
rect 86092 35876 86096 35932
rect 86032 35872 86096 35876
rect 86112 35932 86176 35936
rect 86112 35876 86116 35932
rect 86116 35876 86172 35932
rect 86172 35876 86176 35932
rect 86112 35872 86176 35876
rect 86192 35932 86256 35936
rect 86192 35876 86196 35932
rect 86196 35876 86252 35932
rect 86252 35876 86256 35932
rect 86192 35872 86256 35876
rect 89952 35932 90016 35936
rect 89952 35876 89956 35932
rect 89956 35876 90012 35932
rect 90012 35876 90016 35932
rect 89952 35872 90016 35876
rect 90032 35932 90096 35936
rect 90032 35876 90036 35932
rect 90036 35876 90092 35932
rect 90092 35876 90096 35932
rect 90032 35872 90096 35876
rect 90112 35932 90176 35936
rect 90112 35876 90116 35932
rect 90116 35876 90172 35932
rect 90172 35876 90176 35932
rect 90112 35872 90176 35876
rect 90192 35932 90256 35936
rect 90192 35876 90196 35932
rect 90196 35876 90252 35932
rect 90252 35876 90256 35932
rect 90192 35872 90256 35876
rect 3952 35388 4016 35392
rect 3952 35332 3956 35388
rect 3956 35332 4012 35388
rect 4012 35332 4016 35388
rect 3952 35328 4016 35332
rect 4032 35388 4096 35392
rect 4032 35332 4036 35388
rect 4036 35332 4092 35388
rect 4092 35332 4096 35388
rect 4032 35328 4096 35332
rect 4112 35388 4176 35392
rect 4112 35332 4116 35388
rect 4116 35332 4172 35388
rect 4172 35332 4176 35388
rect 4112 35328 4176 35332
rect 4192 35388 4256 35392
rect 4192 35332 4196 35388
rect 4196 35332 4252 35388
rect 4252 35332 4256 35388
rect 4192 35328 4256 35332
rect 87952 35388 88016 35392
rect 87952 35332 87956 35388
rect 87956 35332 88012 35388
rect 88012 35332 88016 35388
rect 87952 35328 88016 35332
rect 88032 35388 88096 35392
rect 88032 35332 88036 35388
rect 88036 35332 88092 35388
rect 88092 35332 88096 35388
rect 88032 35328 88096 35332
rect 88112 35388 88176 35392
rect 88112 35332 88116 35388
rect 88116 35332 88172 35388
rect 88172 35332 88176 35388
rect 88112 35328 88176 35332
rect 88192 35388 88256 35392
rect 88192 35332 88196 35388
rect 88196 35332 88252 35388
rect 88252 35332 88256 35388
rect 88192 35328 88256 35332
rect 1952 34844 2016 34848
rect 1952 34788 1956 34844
rect 1956 34788 2012 34844
rect 2012 34788 2016 34844
rect 1952 34784 2016 34788
rect 2032 34844 2096 34848
rect 2032 34788 2036 34844
rect 2036 34788 2092 34844
rect 2092 34788 2096 34844
rect 2032 34784 2096 34788
rect 2112 34844 2176 34848
rect 2112 34788 2116 34844
rect 2116 34788 2172 34844
rect 2172 34788 2176 34844
rect 2112 34784 2176 34788
rect 2192 34844 2256 34848
rect 2192 34788 2196 34844
rect 2196 34788 2252 34844
rect 2252 34788 2256 34844
rect 2192 34784 2256 34788
rect 85952 34844 86016 34848
rect 85952 34788 85956 34844
rect 85956 34788 86012 34844
rect 86012 34788 86016 34844
rect 85952 34784 86016 34788
rect 86032 34844 86096 34848
rect 86032 34788 86036 34844
rect 86036 34788 86092 34844
rect 86092 34788 86096 34844
rect 86032 34784 86096 34788
rect 86112 34844 86176 34848
rect 86112 34788 86116 34844
rect 86116 34788 86172 34844
rect 86172 34788 86176 34844
rect 86112 34784 86176 34788
rect 86192 34844 86256 34848
rect 86192 34788 86196 34844
rect 86196 34788 86252 34844
rect 86252 34788 86256 34844
rect 86192 34784 86256 34788
rect 89952 34844 90016 34848
rect 89952 34788 89956 34844
rect 89956 34788 90012 34844
rect 90012 34788 90016 34844
rect 89952 34784 90016 34788
rect 90032 34844 90096 34848
rect 90032 34788 90036 34844
rect 90036 34788 90092 34844
rect 90092 34788 90096 34844
rect 90032 34784 90096 34788
rect 90112 34844 90176 34848
rect 90112 34788 90116 34844
rect 90116 34788 90172 34844
rect 90172 34788 90176 34844
rect 90112 34784 90176 34788
rect 90192 34844 90256 34848
rect 90192 34788 90196 34844
rect 90196 34788 90252 34844
rect 90252 34788 90256 34844
rect 90192 34784 90256 34788
rect 3952 34300 4016 34304
rect 3952 34244 3956 34300
rect 3956 34244 4012 34300
rect 4012 34244 4016 34300
rect 3952 34240 4016 34244
rect 4032 34300 4096 34304
rect 4032 34244 4036 34300
rect 4036 34244 4092 34300
rect 4092 34244 4096 34300
rect 4032 34240 4096 34244
rect 4112 34300 4176 34304
rect 4112 34244 4116 34300
rect 4116 34244 4172 34300
rect 4172 34244 4176 34300
rect 4112 34240 4176 34244
rect 4192 34300 4256 34304
rect 4192 34244 4196 34300
rect 4196 34244 4252 34300
rect 4252 34244 4256 34300
rect 4192 34240 4256 34244
rect 87952 34300 88016 34304
rect 87952 34244 87956 34300
rect 87956 34244 88012 34300
rect 88012 34244 88016 34300
rect 87952 34240 88016 34244
rect 88032 34300 88096 34304
rect 88032 34244 88036 34300
rect 88036 34244 88092 34300
rect 88092 34244 88096 34300
rect 88032 34240 88096 34244
rect 88112 34300 88176 34304
rect 88112 34244 88116 34300
rect 88116 34244 88172 34300
rect 88172 34244 88176 34300
rect 88112 34240 88176 34244
rect 88192 34300 88256 34304
rect 88192 34244 88196 34300
rect 88196 34244 88252 34300
rect 88252 34244 88256 34300
rect 88192 34240 88256 34244
rect 83412 33764 83476 33828
rect 83964 33764 84028 33828
rect 1952 33756 2016 33760
rect 1952 33700 1956 33756
rect 1956 33700 2012 33756
rect 2012 33700 2016 33756
rect 1952 33696 2016 33700
rect 2032 33756 2096 33760
rect 2032 33700 2036 33756
rect 2036 33700 2092 33756
rect 2092 33700 2096 33756
rect 2032 33696 2096 33700
rect 2112 33756 2176 33760
rect 2112 33700 2116 33756
rect 2116 33700 2172 33756
rect 2172 33700 2176 33756
rect 2112 33696 2176 33700
rect 2192 33756 2256 33760
rect 2192 33700 2196 33756
rect 2196 33700 2252 33756
rect 2252 33700 2256 33756
rect 2192 33696 2256 33700
rect 85952 33756 86016 33760
rect 85952 33700 85956 33756
rect 85956 33700 86012 33756
rect 86012 33700 86016 33756
rect 85952 33696 86016 33700
rect 86032 33756 86096 33760
rect 86032 33700 86036 33756
rect 86036 33700 86092 33756
rect 86092 33700 86096 33756
rect 86032 33696 86096 33700
rect 86112 33756 86176 33760
rect 86112 33700 86116 33756
rect 86116 33700 86172 33756
rect 86172 33700 86176 33756
rect 86112 33696 86176 33700
rect 86192 33756 86256 33760
rect 86192 33700 86196 33756
rect 86196 33700 86252 33756
rect 86252 33700 86256 33756
rect 86192 33696 86256 33700
rect 89952 33756 90016 33760
rect 89952 33700 89956 33756
rect 89956 33700 90012 33756
rect 90012 33700 90016 33756
rect 89952 33696 90016 33700
rect 90032 33756 90096 33760
rect 90032 33700 90036 33756
rect 90036 33700 90092 33756
rect 90092 33700 90096 33756
rect 90032 33696 90096 33700
rect 90112 33756 90176 33760
rect 90112 33700 90116 33756
rect 90116 33700 90172 33756
rect 90172 33700 90176 33756
rect 90112 33696 90176 33700
rect 90192 33756 90256 33760
rect 90192 33700 90196 33756
rect 90196 33700 90252 33756
rect 90252 33700 90256 33756
rect 90192 33696 90256 33700
rect 3952 33212 4016 33216
rect 3952 33156 3956 33212
rect 3956 33156 4012 33212
rect 4012 33156 4016 33212
rect 3952 33152 4016 33156
rect 4032 33212 4096 33216
rect 4032 33156 4036 33212
rect 4036 33156 4092 33212
rect 4092 33156 4096 33212
rect 4032 33152 4096 33156
rect 4112 33212 4176 33216
rect 4112 33156 4116 33212
rect 4116 33156 4172 33212
rect 4172 33156 4176 33212
rect 4112 33152 4176 33156
rect 4192 33212 4256 33216
rect 4192 33156 4196 33212
rect 4196 33156 4252 33212
rect 4252 33156 4256 33212
rect 4192 33152 4256 33156
rect 87952 33212 88016 33216
rect 87952 33156 87956 33212
rect 87956 33156 88012 33212
rect 88012 33156 88016 33212
rect 87952 33152 88016 33156
rect 88032 33212 88096 33216
rect 88032 33156 88036 33212
rect 88036 33156 88092 33212
rect 88092 33156 88096 33212
rect 88032 33152 88096 33156
rect 88112 33212 88176 33216
rect 88112 33156 88116 33212
rect 88116 33156 88172 33212
rect 88172 33156 88176 33212
rect 88112 33152 88176 33156
rect 88192 33212 88256 33216
rect 88192 33156 88196 33212
rect 88196 33156 88252 33212
rect 88252 33156 88256 33212
rect 88192 33152 88256 33156
rect 1952 32668 2016 32672
rect 1952 32612 1956 32668
rect 1956 32612 2012 32668
rect 2012 32612 2016 32668
rect 1952 32608 2016 32612
rect 2032 32668 2096 32672
rect 2032 32612 2036 32668
rect 2036 32612 2092 32668
rect 2092 32612 2096 32668
rect 2032 32608 2096 32612
rect 2112 32668 2176 32672
rect 2112 32612 2116 32668
rect 2116 32612 2172 32668
rect 2172 32612 2176 32668
rect 2112 32608 2176 32612
rect 2192 32668 2256 32672
rect 2192 32612 2196 32668
rect 2196 32612 2252 32668
rect 2252 32612 2256 32668
rect 2192 32608 2256 32612
rect 85952 32668 86016 32672
rect 85952 32612 85956 32668
rect 85956 32612 86012 32668
rect 86012 32612 86016 32668
rect 85952 32608 86016 32612
rect 86032 32668 86096 32672
rect 86032 32612 86036 32668
rect 86036 32612 86092 32668
rect 86092 32612 86096 32668
rect 86032 32608 86096 32612
rect 86112 32668 86176 32672
rect 86112 32612 86116 32668
rect 86116 32612 86172 32668
rect 86172 32612 86176 32668
rect 86112 32608 86176 32612
rect 86192 32668 86256 32672
rect 86192 32612 86196 32668
rect 86196 32612 86252 32668
rect 86252 32612 86256 32668
rect 86192 32608 86256 32612
rect 89952 32668 90016 32672
rect 89952 32612 89956 32668
rect 89956 32612 90012 32668
rect 90012 32612 90016 32668
rect 89952 32608 90016 32612
rect 90032 32668 90096 32672
rect 90032 32612 90036 32668
rect 90036 32612 90092 32668
rect 90092 32612 90096 32668
rect 90032 32608 90096 32612
rect 90112 32668 90176 32672
rect 90112 32612 90116 32668
rect 90116 32612 90172 32668
rect 90172 32612 90176 32668
rect 90112 32608 90176 32612
rect 90192 32668 90256 32672
rect 90192 32612 90196 32668
rect 90196 32612 90252 32668
rect 90252 32612 90256 32668
rect 90192 32608 90256 32612
rect 3952 32124 4016 32128
rect 3952 32068 3956 32124
rect 3956 32068 4012 32124
rect 4012 32068 4016 32124
rect 3952 32064 4016 32068
rect 4032 32124 4096 32128
rect 4032 32068 4036 32124
rect 4036 32068 4092 32124
rect 4092 32068 4096 32124
rect 4032 32064 4096 32068
rect 4112 32124 4176 32128
rect 4112 32068 4116 32124
rect 4116 32068 4172 32124
rect 4172 32068 4176 32124
rect 4112 32064 4176 32068
rect 4192 32124 4256 32128
rect 4192 32068 4196 32124
rect 4196 32068 4252 32124
rect 4252 32068 4256 32124
rect 4192 32064 4256 32068
rect 87952 32124 88016 32128
rect 87952 32068 87956 32124
rect 87956 32068 88012 32124
rect 88012 32068 88016 32124
rect 87952 32064 88016 32068
rect 88032 32124 88096 32128
rect 88032 32068 88036 32124
rect 88036 32068 88092 32124
rect 88092 32068 88096 32124
rect 88032 32064 88096 32068
rect 88112 32124 88176 32128
rect 88112 32068 88116 32124
rect 88116 32068 88172 32124
rect 88172 32068 88176 32124
rect 88112 32064 88176 32068
rect 88192 32124 88256 32128
rect 88192 32068 88196 32124
rect 88196 32068 88252 32124
rect 88252 32068 88256 32124
rect 88192 32064 88256 32068
rect 1952 31580 2016 31584
rect 1952 31524 1956 31580
rect 1956 31524 2012 31580
rect 2012 31524 2016 31580
rect 1952 31520 2016 31524
rect 2032 31580 2096 31584
rect 2032 31524 2036 31580
rect 2036 31524 2092 31580
rect 2092 31524 2096 31580
rect 2032 31520 2096 31524
rect 2112 31580 2176 31584
rect 2112 31524 2116 31580
rect 2116 31524 2172 31580
rect 2172 31524 2176 31580
rect 2112 31520 2176 31524
rect 2192 31580 2256 31584
rect 2192 31524 2196 31580
rect 2196 31524 2252 31580
rect 2252 31524 2256 31580
rect 2192 31520 2256 31524
rect 85952 31580 86016 31584
rect 85952 31524 85956 31580
rect 85956 31524 86012 31580
rect 86012 31524 86016 31580
rect 85952 31520 86016 31524
rect 86032 31580 86096 31584
rect 86032 31524 86036 31580
rect 86036 31524 86092 31580
rect 86092 31524 86096 31580
rect 86032 31520 86096 31524
rect 86112 31580 86176 31584
rect 86112 31524 86116 31580
rect 86116 31524 86172 31580
rect 86172 31524 86176 31580
rect 86112 31520 86176 31524
rect 86192 31580 86256 31584
rect 86192 31524 86196 31580
rect 86196 31524 86252 31580
rect 86252 31524 86256 31580
rect 86192 31520 86256 31524
rect 89952 31580 90016 31584
rect 89952 31524 89956 31580
rect 89956 31524 90012 31580
rect 90012 31524 90016 31580
rect 89952 31520 90016 31524
rect 90032 31580 90096 31584
rect 90032 31524 90036 31580
rect 90036 31524 90092 31580
rect 90092 31524 90096 31580
rect 90032 31520 90096 31524
rect 90112 31580 90176 31584
rect 90112 31524 90116 31580
rect 90116 31524 90172 31580
rect 90172 31524 90176 31580
rect 90112 31520 90176 31524
rect 90192 31580 90256 31584
rect 90192 31524 90196 31580
rect 90196 31524 90252 31580
rect 90252 31524 90256 31580
rect 90192 31520 90256 31524
rect 3952 31036 4016 31040
rect 3952 30980 3956 31036
rect 3956 30980 4012 31036
rect 4012 30980 4016 31036
rect 3952 30976 4016 30980
rect 4032 31036 4096 31040
rect 4032 30980 4036 31036
rect 4036 30980 4092 31036
rect 4092 30980 4096 31036
rect 4032 30976 4096 30980
rect 4112 31036 4176 31040
rect 4112 30980 4116 31036
rect 4116 30980 4172 31036
rect 4172 30980 4176 31036
rect 4112 30976 4176 30980
rect 4192 31036 4256 31040
rect 4192 30980 4196 31036
rect 4196 30980 4252 31036
rect 4252 30980 4256 31036
rect 4192 30976 4256 30980
rect 87952 31036 88016 31040
rect 87952 30980 87956 31036
rect 87956 30980 88012 31036
rect 88012 30980 88016 31036
rect 87952 30976 88016 30980
rect 88032 31036 88096 31040
rect 88032 30980 88036 31036
rect 88036 30980 88092 31036
rect 88092 30980 88096 31036
rect 88032 30976 88096 30980
rect 88112 31036 88176 31040
rect 88112 30980 88116 31036
rect 88116 30980 88172 31036
rect 88172 30980 88176 31036
rect 88112 30976 88176 30980
rect 88192 31036 88256 31040
rect 88192 30980 88196 31036
rect 88196 30980 88252 31036
rect 88252 30980 88256 31036
rect 88192 30976 88256 30980
rect 1952 30492 2016 30496
rect 1952 30436 1956 30492
rect 1956 30436 2012 30492
rect 2012 30436 2016 30492
rect 1952 30432 2016 30436
rect 2032 30492 2096 30496
rect 2032 30436 2036 30492
rect 2036 30436 2092 30492
rect 2092 30436 2096 30492
rect 2032 30432 2096 30436
rect 2112 30492 2176 30496
rect 2112 30436 2116 30492
rect 2116 30436 2172 30492
rect 2172 30436 2176 30492
rect 2112 30432 2176 30436
rect 2192 30492 2256 30496
rect 2192 30436 2196 30492
rect 2196 30436 2252 30492
rect 2252 30436 2256 30492
rect 2192 30432 2256 30436
rect 85952 30492 86016 30496
rect 85952 30436 85956 30492
rect 85956 30436 86012 30492
rect 86012 30436 86016 30492
rect 85952 30432 86016 30436
rect 86032 30492 86096 30496
rect 86032 30436 86036 30492
rect 86036 30436 86092 30492
rect 86092 30436 86096 30492
rect 86032 30432 86096 30436
rect 86112 30492 86176 30496
rect 86112 30436 86116 30492
rect 86116 30436 86172 30492
rect 86172 30436 86176 30492
rect 86112 30432 86176 30436
rect 86192 30492 86256 30496
rect 86192 30436 86196 30492
rect 86196 30436 86252 30492
rect 86252 30436 86256 30492
rect 86192 30432 86256 30436
rect 89952 30492 90016 30496
rect 89952 30436 89956 30492
rect 89956 30436 90012 30492
rect 90012 30436 90016 30492
rect 89952 30432 90016 30436
rect 90032 30492 90096 30496
rect 90032 30436 90036 30492
rect 90036 30436 90092 30492
rect 90092 30436 90096 30492
rect 90032 30432 90096 30436
rect 90112 30492 90176 30496
rect 90112 30436 90116 30492
rect 90116 30436 90172 30492
rect 90172 30436 90176 30492
rect 90112 30432 90176 30436
rect 90192 30492 90256 30496
rect 90192 30436 90196 30492
rect 90196 30436 90252 30492
rect 90252 30436 90256 30492
rect 90192 30432 90256 30436
rect 3952 29948 4016 29952
rect 3952 29892 3956 29948
rect 3956 29892 4012 29948
rect 4012 29892 4016 29948
rect 3952 29888 4016 29892
rect 4032 29948 4096 29952
rect 4032 29892 4036 29948
rect 4036 29892 4092 29948
rect 4092 29892 4096 29948
rect 4032 29888 4096 29892
rect 4112 29948 4176 29952
rect 4112 29892 4116 29948
rect 4116 29892 4172 29948
rect 4172 29892 4176 29948
rect 4112 29888 4176 29892
rect 4192 29948 4256 29952
rect 4192 29892 4196 29948
rect 4196 29892 4252 29948
rect 4252 29892 4256 29948
rect 4192 29888 4256 29892
rect 87952 29948 88016 29952
rect 87952 29892 87956 29948
rect 87956 29892 88012 29948
rect 88012 29892 88016 29948
rect 87952 29888 88016 29892
rect 88032 29948 88096 29952
rect 88032 29892 88036 29948
rect 88036 29892 88092 29948
rect 88092 29892 88096 29948
rect 88032 29888 88096 29892
rect 88112 29948 88176 29952
rect 88112 29892 88116 29948
rect 88116 29892 88172 29948
rect 88172 29892 88176 29948
rect 88112 29888 88176 29892
rect 88192 29948 88256 29952
rect 88192 29892 88196 29948
rect 88196 29892 88252 29948
rect 88252 29892 88256 29948
rect 88192 29888 88256 29892
rect 1952 29404 2016 29408
rect 1952 29348 1956 29404
rect 1956 29348 2012 29404
rect 2012 29348 2016 29404
rect 1952 29344 2016 29348
rect 2032 29404 2096 29408
rect 2032 29348 2036 29404
rect 2036 29348 2092 29404
rect 2092 29348 2096 29404
rect 2032 29344 2096 29348
rect 2112 29404 2176 29408
rect 2112 29348 2116 29404
rect 2116 29348 2172 29404
rect 2172 29348 2176 29404
rect 2112 29344 2176 29348
rect 2192 29404 2256 29408
rect 2192 29348 2196 29404
rect 2196 29348 2252 29404
rect 2252 29348 2256 29404
rect 2192 29344 2256 29348
rect 85952 29404 86016 29408
rect 85952 29348 85956 29404
rect 85956 29348 86012 29404
rect 86012 29348 86016 29404
rect 85952 29344 86016 29348
rect 86032 29404 86096 29408
rect 86032 29348 86036 29404
rect 86036 29348 86092 29404
rect 86092 29348 86096 29404
rect 86032 29344 86096 29348
rect 86112 29404 86176 29408
rect 86112 29348 86116 29404
rect 86116 29348 86172 29404
rect 86172 29348 86176 29404
rect 86112 29344 86176 29348
rect 86192 29404 86256 29408
rect 86192 29348 86196 29404
rect 86196 29348 86252 29404
rect 86252 29348 86256 29404
rect 86192 29344 86256 29348
rect 89952 29404 90016 29408
rect 89952 29348 89956 29404
rect 89956 29348 90012 29404
rect 90012 29348 90016 29404
rect 89952 29344 90016 29348
rect 90032 29404 90096 29408
rect 90032 29348 90036 29404
rect 90036 29348 90092 29404
rect 90092 29348 90096 29404
rect 90032 29344 90096 29348
rect 90112 29404 90176 29408
rect 90112 29348 90116 29404
rect 90116 29348 90172 29404
rect 90172 29348 90176 29404
rect 90112 29344 90176 29348
rect 90192 29404 90256 29408
rect 90192 29348 90196 29404
rect 90196 29348 90252 29404
rect 90252 29348 90256 29404
rect 90192 29344 90256 29348
rect 3952 28860 4016 28864
rect 3952 28804 3956 28860
rect 3956 28804 4012 28860
rect 4012 28804 4016 28860
rect 3952 28800 4016 28804
rect 4032 28860 4096 28864
rect 4032 28804 4036 28860
rect 4036 28804 4092 28860
rect 4092 28804 4096 28860
rect 4032 28800 4096 28804
rect 4112 28860 4176 28864
rect 4112 28804 4116 28860
rect 4116 28804 4172 28860
rect 4172 28804 4176 28860
rect 4112 28800 4176 28804
rect 4192 28860 4256 28864
rect 4192 28804 4196 28860
rect 4196 28804 4252 28860
rect 4252 28804 4256 28860
rect 4192 28800 4256 28804
rect 87952 28860 88016 28864
rect 87952 28804 87956 28860
rect 87956 28804 88012 28860
rect 88012 28804 88016 28860
rect 87952 28800 88016 28804
rect 88032 28860 88096 28864
rect 88032 28804 88036 28860
rect 88036 28804 88092 28860
rect 88092 28804 88096 28860
rect 88032 28800 88096 28804
rect 88112 28860 88176 28864
rect 88112 28804 88116 28860
rect 88116 28804 88172 28860
rect 88172 28804 88176 28860
rect 88112 28800 88176 28804
rect 88192 28860 88256 28864
rect 88192 28804 88196 28860
rect 88196 28804 88252 28860
rect 88252 28804 88256 28860
rect 88192 28800 88256 28804
rect 1952 28316 2016 28320
rect 1952 28260 1956 28316
rect 1956 28260 2012 28316
rect 2012 28260 2016 28316
rect 1952 28256 2016 28260
rect 2032 28316 2096 28320
rect 2032 28260 2036 28316
rect 2036 28260 2092 28316
rect 2092 28260 2096 28316
rect 2032 28256 2096 28260
rect 2112 28316 2176 28320
rect 2112 28260 2116 28316
rect 2116 28260 2172 28316
rect 2172 28260 2176 28316
rect 2112 28256 2176 28260
rect 2192 28316 2256 28320
rect 2192 28260 2196 28316
rect 2196 28260 2252 28316
rect 2252 28260 2256 28316
rect 2192 28256 2256 28260
rect 85952 28316 86016 28320
rect 85952 28260 85956 28316
rect 85956 28260 86012 28316
rect 86012 28260 86016 28316
rect 85952 28256 86016 28260
rect 86032 28316 86096 28320
rect 86032 28260 86036 28316
rect 86036 28260 86092 28316
rect 86092 28260 86096 28316
rect 86032 28256 86096 28260
rect 86112 28316 86176 28320
rect 86112 28260 86116 28316
rect 86116 28260 86172 28316
rect 86172 28260 86176 28316
rect 86112 28256 86176 28260
rect 86192 28316 86256 28320
rect 86192 28260 86196 28316
rect 86196 28260 86252 28316
rect 86252 28260 86256 28316
rect 86192 28256 86256 28260
rect 89952 28316 90016 28320
rect 89952 28260 89956 28316
rect 89956 28260 90012 28316
rect 90012 28260 90016 28316
rect 89952 28256 90016 28260
rect 90032 28316 90096 28320
rect 90032 28260 90036 28316
rect 90036 28260 90092 28316
rect 90092 28260 90096 28316
rect 90032 28256 90096 28260
rect 90112 28316 90176 28320
rect 90112 28260 90116 28316
rect 90116 28260 90172 28316
rect 90172 28260 90176 28316
rect 90112 28256 90176 28260
rect 90192 28316 90256 28320
rect 90192 28260 90196 28316
rect 90196 28260 90252 28316
rect 90252 28260 90256 28316
rect 90192 28256 90256 28260
rect 3952 27772 4016 27776
rect 3952 27716 3956 27772
rect 3956 27716 4012 27772
rect 4012 27716 4016 27772
rect 3952 27712 4016 27716
rect 4032 27772 4096 27776
rect 4032 27716 4036 27772
rect 4036 27716 4092 27772
rect 4092 27716 4096 27772
rect 4032 27712 4096 27716
rect 4112 27772 4176 27776
rect 4112 27716 4116 27772
rect 4116 27716 4172 27772
rect 4172 27716 4176 27772
rect 4112 27712 4176 27716
rect 4192 27772 4256 27776
rect 4192 27716 4196 27772
rect 4196 27716 4252 27772
rect 4252 27716 4256 27772
rect 4192 27712 4256 27716
rect 87952 27772 88016 27776
rect 87952 27716 87956 27772
rect 87956 27716 88012 27772
rect 88012 27716 88016 27772
rect 87952 27712 88016 27716
rect 88032 27772 88096 27776
rect 88032 27716 88036 27772
rect 88036 27716 88092 27772
rect 88092 27716 88096 27772
rect 88032 27712 88096 27716
rect 88112 27772 88176 27776
rect 88112 27716 88116 27772
rect 88116 27716 88172 27772
rect 88172 27716 88176 27772
rect 88112 27712 88176 27716
rect 88192 27772 88256 27776
rect 88192 27716 88196 27772
rect 88196 27716 88252 27772
rect 88252 27716 88256 27772
rect 88192 27712 88256 27716
rect 1952 27228 2016 27232
rect 1952 27172 1956 27228
rect 1956 27172 2012 27228
rect 2012 27172 2016 27228
rect 1952 27168 2016 27172
rect 2032 27228 2096 27232
rect 2032 27172 2036 27228
rect 2036 27172 2092 27228
rect 2092 27172 2096 27228
rect 2032 27168 2096 27172
rect 2112 27228 2176 27232
rect 2112 27172 2116 27228
rect 2116 27172 2172 27228
rect 2172 27172 2176 27228
rect 2112 27168 2176 27172
rect 2192 27228 2256 27232
rect 2192 27172 2196 27228
rect 2196 27172 2252 27228
rect 2252 27172 2256 27228
rect 2192 27168 2256 27172
rect 85952 27228 86016 27232
rect 85952 27172 85956 27228
rect 85956 27172 86012 27228
rect 86012 27172 86016 27228
rect 85952 27168 86016 27172
rect 86032 27228 86096 27232
rect 86032 27172 86036 27228
rect 86036 27172 86092 27228
rect 86092 27172 86096 27228
rect 86032 27168 86096 27172
rect 86112 27228 86176 27232
rect 86112 27172 86116 27228
rect 86116 27172 86172 27228
rect 86172 27172 86176 27228
rect 86112 27168 86176 27172
rect 86192 27228 86256 27232
rect 86192 27172 86196 27228
rect 86196 27172 86252 27228
rect 86252 27172 86256 27228
rect 86192 27168 86256 27172
rect 89952 27228 90016 27232
rect 89952 27172 89956 27228
rect 89956 27172 90012 27228
rect 90012 27172 90016 27228
rect 89952 27168 90016 27172
rect 90032 27228 90096 27232
rect 90032 27172 90036 27228
rect 90036 27172 90092 27228
rect 90092 27172 90096 27228
rect 90032 27168 90096 27172
rect 90112 27228 90176 27232
rect 90112 27172 90116 27228
rect 90116 27172 90172 27228
rect 90172 27172 90176 27228
rect 90112 27168 90176 27172
rect 90192 27228 90256 27232
rect 90192 27172 90196 27228
rect 90196 27172 90252 27228
rect 90252 27172 90256 27228
rect 90192 27168 90256 27172
rect 3952 26684 4016 26688
rect 3952 26628 3956 26684
rect 3956 26628 4012 26684
rect 4012 26628 4016 26684
rect 3952 26624 4016 26628
rect 4032 26684 4096 26688
rect 4032 26628 4036 26684
rect 4036 26628 4092 26684
rect 4092 26628 4096 26684
rect 4032 26624 4096 26628
rect 4112 26684 4176 26688
rect 4112 26628 4116 26684
rect 4116 26628 4172 26684
rect 4172 26628 4176 26684
rect 4112 26624 4176 26628
rect 4192 26684 4256 26688
rect 4192 26628 4196 26684
rect 4196 26628 4252 26684
rect 4252 26628 4256 26684
rect 4192 26624 4256 26628
rect 87952 26684 88016 26688
rect 87952 26628 87956 26684
rect 87956 26628 88012 26684
rect 88012 26628 88016 26684
rect 87952 26624 88016 26628
rect 88032 26684 88096 26688
rect 88032 26628 88036 26684
rect 88036 26628 88092 26684
rect 88092 26628 88096 26684
rect 88032 26624 88096 26628
rect 88112 26684 88176 26688
rect 88112 26628 88116 26684
rect 88116 26628 88172 26684
rect 88172 26628 88176 26684
rect 88112 26624 88176 26628
rect 88192 26684 88256 26688
rect 88192 26628 88196 26684
rect 88196 26628 88252 26684
rect 88252 26628 88256 26684
rect 88192 26624 88256 26628
rect 1952 26140 2016 26144
rect 1952 26084 1956 26140
rect 1956 26084 2012 26140
rect 2012 26084 2016 26140
rect 1952 26080 2016 26084
rect 2032 26140 2096 26144
rect 2032 26084 2036 26140
rect 2036 26084 2092 26140
rect 2092 26084 2096 26140
rect 2032 26080 2096 26084
rect 2112 26140 2176 26144
rect 2112 26084 2116 26140
rect 2116 26084 2172 26140
rect 2172 26084 2176 26140
rect 2112 26080 2176 26084
rect 2192 26140 2256 26144
rect 2192 26084 2196 26140
rect 2196 26084 2252 26140
rect 2252 26084 2256 26140
rect 2192 26080 2256 26084
rect 85952 26140 86016 26144
rect 85952 26084 85956 26140
rect 85956 26084 86012 26140
rect 86012 26084 86016 26140
rect 85952 26080 86016 26084
rect 86032 26140 86096 26144
rect 86032 26084 86036 26140
rect 86036 26084 86092 26140
rect 86092 26084 86096 26140
rect 86032 26080 86096 26084
rect 86112 26140 86176 26144
rect 86112 26084 86116 26140
rect 86116 26084 86172 26140
rect 86172 26084 86176 26140
rect 86112 26080 86176 26084
rect 86192 26140 86256 26144
rect 86192 26084 86196 26140
rect 86196 26084 86252 26140
rect 86252 26084 86256 26140
rect 86192 26080 86256 26084
rect 89952 26140 90016 26144
rect 89952 26084 89956 26140
rect 89956 26084 90012 26140
rect 90012 26084 90016 26140
rect 89952 26080 90016 26084
rect 90032 26140 90096 26144
rect 90032 26084 90036 26140
rect 90036 26084 90092 26140
rect 90092 26084 90096 26140
rect 90032 26080 90096 26084
rect 90112 26140 90176 26144
rect 90112 26084 90116 26140
rect 90116 26084 90172 26140
rect 90172 26084 90176 26140
rect 90112 26080 90176 26084
rect 90192 26140 90256 26144
rect 90192 26084 90196 26140
rect 90196 26084 90252 26140
rect 90252 26084 90256 26140
rect 90192 26080 90256 26084
rect 3952 25596 4016 25600
rect 3952 25540 3956 25596
rect 3956 25540 4012 25596
rect 4012 25540 4016 25596
rect 3952 25536 4016 25540
rect 4032 25596 4096 25600
rect 4032 25540 4036 25596
rect 4036 25540 4092 25596
rect 4092 25540 4096 25596
rect 4032 25536 4096 25540
rect 4112 25596 4176 25600
rect 4112 25540 4116 25596
rect 4116 25540 4172 25596
rect 4172 25540 4176 25596
rect 4112 25536 4176 25540
rect 4192 25596 4256 25600
rect 4192 25540 4196 25596
rect 4196 25540 4252 25596
rect 4252 25540 4256 25596
rect 4192 25536 4256 25540
rect 87952 25596 88016 25600
rect 87952 25540 87956 25596
rect 87956 25540 88012 25596
rect 88012 25540 88016 25596
rect 87952 25536 88016 25540
rect 88032 25596 88096 25600
rect 88032 25540 88036 25596
rect 88036 25540 88092 25596
rect 88092 25540 88096 25596
rect 88032 25536 88096 25540
rect 88112 25596 88176 25600
rect 88112 25540 88116 25596
rect 88116 25540 88172 25596
rect 88172 25540 88176 25596
rect 88112 25536 88176 25540
rect 88192 25596 88256 25600
rect 88192 25540 88196 25596
rect 88196 25540 88252 25596
rect 88252 25540 88256 25596
rect 88192 25536 88256 25540
rect 1952 25052 2016 25056
rect 1952 24996 1956 25052
rect 1956 24996 2012 25052
rect 2012 24996 2016 25052
rect 1952 24992 2016 24996
rect 2032 25052 2096 25056
rect 2032 24996 2036 25052
rect 2036 24996 2092 25052
rect 2092 24996 2096 25052
rect 2032 24992 2096 24996
rect 2112 25052 2176 25056
rect 2112 24996 2116 25052
rect 2116 24996 2172 25052
rect 2172 24996 2176 25052
rect 2112 24992 2176 24996
rect 2192 25052 2256 25056
rect 2192 24996 2196 25052
rect 2196 24996 2252 25052
rect 2252 24996 2256 25052
rect 2192 24992 2256 24996
rect 85952 25052 86016 25056
rect 85952 24996 85956 25052
rect 85956 24996 86012 25052
rect 86012 24996 86016 25052
rect 85952 24992 86016 24996
rect 86032 25052 86096 25056
rect 86032 24996 86036 25052
rect 86036 24996 86092 25052
rect 86092 24996 86096 25052
rect 86032 24992 86096 24996
rect 86112 25052 86176 25056
rect 86112 24996 86116 25052
rect 86116 24996 86172 25052
rect 86172 24996 86176 25052
rect 86112 24992 86176 24996
rect 86192 25052 86256 25056
rect 86192 24996 86196 25052
rect 86196 24996 86252 25052
rect 86252 24996 86256 25052
rect 86192 24992 86256 24996
rect 89952 25052 90016 25056
rect 89952 24996 89956 25052
rect 89956 24996 90012 25052
rect 90012 24996 90016 25052
rect 89952 24992 90016 24996
rect 90032 25052 90096 25056
rect 90032 24996 90036 25052
rect 90036 24996 90092 25052
rect 90092 24996 90096 25052
rect 90032 24992 90096 24996
rect 90112 25052 90176 25056
rect 90112 24996 90116 25052
rect 90116 24996 90172 25052
rect 90172 24996 90176 25052
rect 90112 24992 90176 24996
rect 90192 25052 90256 25056
rect 90192 24996 90196 25052
rect 90196 24996 90252 25052
rect 90252 24996 90256 25052
rect 90192 24992 90256 24996
rect 3952 24508 4016 24512
rect 3952 24452 3956 24508
rect 3956 24452 4012 24508
rect 4012 24452 4016 24508
rect 3952 24448 4016 24452
rect 4032 24508 4096 24512
rect 4032 24452 4036 24508
rect 4036 24452 4092 24508
rect 4092 24452 4096 24508
rect 4032 24448 4096 24452
rect 4112 24508 4176 24512
rect 4112 24452 4116 24508
rect 4116 24452 4172 24508
rect 4172 24452 4176 24508
rect 4112 24448 4176 24452
rect 4192 24508 4256 24512
rect 4192 24452 4196 24508
rect 4196 24452 4252 24508
rect 4252 24452 4256 24508
rect 4192 24448 4256 24452
rect 87952 24508 88016 24512
rect 87952 24452 87956 24508
rect 87956 24452 88012 24508
rect 88012 24452 88016 24508
rect 87952 24448 88016 24452
rect 88032 24508 88096 24512
rect 88032 24452 88036 24508
rect 88036 24452 88092 24508
rect 88092 24452 88096 24508
rect 88032 24448 88096 24452
rect 88112 24508 88176 24512
rect 88112 24452 88116 24508
rect 88116 24452 88172 24508
rect 88172 24452 88176 24508
rect 88112 24448 88176 24452
rect 88192 24508 88256 24512
rect 88192 24452 88196 24508
rect 88196 24452 88252 24508
rect 88252 24452 88256 24508
rect 88192 24448 88256 24452
rect 1952 23964 2016 23968
rect 1952 23908 1956 23964
rect 1956 23908 2012 23964
rect 2012 23908 2016 23964
rect 1952 23904 2016 23908
rect 2032 23964 2096 23968
rect 2032 23908 2036 23964
rect 2036 23908 2092 23964
rect 2092 23908 2096 23964
rect 2032 23904 2096 23908
rect 2112 23964 2176 23968
rect 2112 23908 2116 23964
rect 2116 23908 2172 23964
rect 2172 23908 2176 23964
rect 2112 23904 2176 23908
rect 2192 23964 2256 23968
rect 2192 23908 2196 23964
rect 2196 23908 2252 23964
rect 2252 23908 2256 23964
rect 2192 23904 2256 23908
rect 85952 23964 86016 23968
rect 85952 23908 85956 23964
rect 85956 23908 86012 23964
rect 86012 23908 86016 23964
rect 85952 23904 86016 23908
rect 86032 23964 86096 23968
rect 86032 23908 86036 23964
rect 86036 23908 86092 23964
rect 86092 23908 86096 23964
rect 86032 23904 86096 23908
rect 86112 23964 86176 23968
rect 86112 23908 86116 23964
rect 86116 23908 86172 23964
rect 86172 23908 86176 23964
rect 86112 23904 86176 23908
rect 86192 23964 86256 23968
rect 86192 23908 86196 23964
rect 86196 23908 86252 23964
rect 86252 23908 86256 23964
rect 86192 23904 86256 23908
rect 89952 23964 90016 23968
rect 89952 23908 89956 23964
rect 89956 23908 90012 23964
rect 90012 23908 90016 23964
rect 89952 23904 90016 23908
rect 90032 23964 90096 23968
rect 90032 23908 90036 23964
rect 90036 23908 90092 23964
rect 90092 23908 90096 23964
rect 90032 23904 90096 23908
rect 90112 23964 90176 23968
rect 90112 23908 90116 23964
rect 90116 23908 90172 23964
rect 90172 23908 90176 23964
rect 90112 23904 90176 23908
rect 90192 23964 90256 23968
rect 90192 23908 90196 23964
rect 90196 23908 90252 23964
rect 90252 23908 90256 23964
rect 90192 23904 90256 23908
rect 3952 23420 4016 23424
rect 3952 23364 3956 23420
rect 3956 23364 4012 23420
rect 4012 23364 4016 23420
rect 3952 23360 4016 23364
rect 4032 23420 4096 23424
rect 4032 23364 4036 23420
rect 4036 23364 4092 23420
rect 4092 23364 4096 23420
rect 4032 23360 4096 23364
rect 4112 23420 4176 23424
rect 4112 23364 4116 23420
rect 4116 23364 4172 23420
rect 4172 23364 4176 23420
rect 4112 23360 4176 23364
rect 4192 23420 4256 23424
rect 4192 23364 4196 23420
rect 4196 23364 4252 23420
rect 4252 23364 4256 23420
rect 4192 23360 4256 23364
rect 87952 23420 88016 23424
rect 87952 23364 87956 23420
rect 87956 23364 88012 23420
rect 88012 23364 88016 23420
rect 87952 23360 88016 23364
rect 88032 23420 88096 23424
rect 88032 23364 88036 23420
rect 88036 23364 88092 23420
rect 88092 23364 88096 23420
rect 88032 23360 88096 23364
rect 88112 23420 88176 23424
rect 88112 23364 88116 23420
rect 88116 23364 88172 23420
rect 88172 23364 88176 23420
rect 88112 23360 88176 23364
rect 88192 23420 88256 23424
rect 88192 23364 88196 23420
rect 88196 23364 88252 23420
rect 88252 23364 88256 23420
rect 88192 23360 88256 23364
rect 1952 22876 2016 22880
rect 1952 22820 1956 22876
rect 1956 22820 2012 22876
rect 2012 22820 2016 22876
rect 1952 22816 2016 22820
rect 2032 22876 2096 22880
rect 2032 22820 2036 22876
rect 2036 22820 2092 22876
rect 2092 22820 2096 22876
rect 2032 22816 2096 22820
rect 2112 22876 2176 22880
rect 2112 22820 2116 22876
rect 2116 22820 2172 22876
rect 2172 22820 2176 22876
rect 2112 22816 2176 22820
rect 2192 22876 2256 22880
rect 2192 22820 2196 22876
rect 2196 22820 2252 22876
rect 2252 22820 2256 22876
rect 2192 22816 2256 22820
rect 85952 22876 86016 22880
rect 85952 22820 85956 22876
rect 85956 22820 86012 22876
rect 86012 22820 86016 22876
rect 85952 22816 86016 22820
rect 86032 22876 86096 22880
rect 86032 22820 86036 22876
rect 86036 22820 86092 22876
rect 86092 22820 86096 22876
rect 86032 22816 86096 22820
rect 86112 22876 86176 22880
rect 86112 22820 86116 22876
rect 86116 22820 86172 22876
rect 86172 22820 86176 22876
rect 86112 22816 86176 22820
rect 86192 22876 86256 22880
rect 86192 22820 86196 22876
rect 86196 22820 86252 22876
rect 86252 22820 86256 22876
rect 86192 22816 86256 22820
rect 89952 22876 90016 22880
rect 89952 22820 89956 22876
rect 89956 22820 90012 22876
rect 90012 22820 90016 22876
rect 89952 22816 90016 22820
rect 90032 22876 90096 22880
rect 90032 22820 90036 22876
rect 90036 22820 90092 22876
rect 90092 22820 90096 22876
rect 90032 22816 90096 22820
rect 90112 22876 90176 22880
rect 90112 22820 90116 22876
rect 90116 22820 90172 22876
rect 90172 22820 90176 22876
rect 90112 22816 90176 22820
rect 90192 22876 90256 22880
rect 90192 22820 90196 22876
rect 90196 22820 90252 22876
rect 90252 22820 90256 22876
rect 90192 22816 90256 22820
rect 3952 22332 4016 22336
rect 3952 22276 3956 22332
rect 3956 22276 4012 22332
rect 4012 22276 4016 22332
rect 3952 22272 4016 22276
rect 4032 22332 4096 22336
rect 4032 22276 4036 22332
rect 4036 22276 4092 22332
rect 4092 22276 4096 22332
rect 4032 22272 4096 22276
rect 4112 22332 4176 22336
rect 4112 22276 4116 22332
rect 4116 22276 4172 22332
rect 4172 22276 4176 22332
rect 4112 22272 4176 22276
rect 4192 22332 4256 22336
rect 4192 22276 4196 22332
rect 4196 22276 4252 22332
rect 4252 22276 4256 22332
rect 4192 22272 4256 22276
rect 87952 22332 88016 22336
rect 87952 22276 87956 22332
rect 87956 22276 88012 22332
rect 88012 22276 88016 22332
rect 87952 22272 88016 22276
rect 88032 22332 88096 22336
rect 88032 22276 88036 22332
rect 88036 22276 88092 22332
rect 88092 22276 88096 22332
rect 88032 22272 88096 22276
rect 88112 22332 88176 22336
rect 88112 22276 88116 22332
rect 88116 22276 88172 22332
rect 88172 22276 88176 22332
rect 88112 22272 88176 22276
rect 88192 22332 88256 22336
rect 88192 22276 88196 22332
rect 88196 22276 88252 22332
rect 88252 22276 88256 22332
rect 88192 22272 88256 22276
rect 1952 21788 2016 21792
rect 1952 21732 1956 21788
rect 1956 21732 2012 21788
rect 2012 21732 2016 21788
rect 1952 21728 2016 21732
rect 2032 21788 2096 21792
rect 2032 21732 2036 21788
rect 2036 21732 2092 21788
rect 2092 21732 2096 21788
rect 2032 21728 2096 21732
rect 2112 21788 2176 21792
rect 2112 21732 2116 21788
rect 2116 21732 2172 21788
rect 2172 21732 2176 21788
rect 2112 21728 2176 21732
rect 2192 21788 2256 21792
rect 2192 21732 2196 21788
rect 2196 21732 2252 21788
rect 2252 21732 2256 21788
rect 2192 21728 2256 21732
rect 85952 21788 86016 21792
rect 85952 21732 85956 21788
rect 85956 21732 86012 21788
rect 86012 21732 86016 21788
rect 85952 21728 86016 21732
rect 86032 21788 86096 21792
rect 86032 21732 86036 21788
rect 86036 21732 86092 21788
rect 86092 21732 86096 21788
rect 86032 21728 86096 21732
rect 86112 21788 86176 21792
rect 86112 21732 86116 21788
rect 86116 21732 86172 21788
rect 86172 21732 86176 21788
rect 86112 21728 86176 21732
rect 86192 21788 86256 21792
rect 86192 21732 86196 21788
rect 86196 21732 86252 21788
rect 86252 21732 86256 21788
rect 86192 21728 86256 21732
rect 89952 21788 90016 21792
rect 89952 21732 89956 21788
rect 89956 21732 90012 21788
rect 90012 21732 90016 21788
rect 89952 21728 90016 21732
rect 90032 21788 90096 21792
rect 90032 21732 90036 21788
rect 90036 21732 90092 21788
rect 90092 21732 90096 21788
rect 90032 21728 90096 21732
rect 90112 21788 90176 21792
rect 90112 21732 90116 21788
rect 90116 21732 90172 21788
rect 90172 21732 90176 21788
rect 90112 21728 90176 21732
rect 90192 21788 90256 21792
rect 90192 21732 90196 21788
rect 90196 21732 90252 21788
rect 90252 21732 90256 21788
rect 90192 21728 90256 21732
rect 3952 21244 4016 21248
rect 3952 21188 3956 21244
rect 3956 21188 4012 21244
rect 4012 21188 4016 21244
rect 3952 21184 4016 21188
rect 4032 21244 4096 21248
rect 4032 21188 4036 21244
rect 4036 21188 4092 21244
rect 4092 21188 4096 21244
rect 4032 21184 4096 21188
rect 4112 21244 4176 21248
rect 4112 21188 4116 21244
rect 4116 21188 4172 21244
rect 4172 21188 4176 21244
rect 4112 21184 4176 21188
rect 4192 21244 4256 21248
rect 4192 21188 4196 21244
rect 4196 21188 4252 21244
rect 4252 21188 4256 21244
rect 4192 21184 4256 21188
rect 87952 21244 88016 21248
rect 87952 21188 87956 21244
rect 87956 21188 88012 21244
rect 88012 21188 88016 21244
rect 87952 21184 88016 21188
rect 88032 21244 88096 21248
rect 88032 21188 88036 21244
rect 88036 21188 88092 21244
rect 88092 21188 88096 21244
rect 88032 21184 88096 21188
rect 88112 21244 88176 21248
rect 88112 21188 88116 21244
rect 88116 21188 88172 21244
rect 88172 21188 88176 21244
rect 88112 21184 88176 21188
rect 88192 21244 88256 21248
rect 88192 21188 88196 21244
rect 88196 21188 88252 21244
rect 88252 21188 88256 21244
rect 88192 21184 88256 21188
rect 1952 20700 2016 20704
rect 1952 20644 1956 20700
rect 1956 20644 2012 20700
rect 2012 20644 2016 20700
rect 1952 20640 2016 20644
rect 2032 20700 2096 20704
rect 2032 20644 2036 20700
rect 2036 20644 2092 20700
rect 2092 20644 2096 20700
rect 2032 20640 2096 20644
rect 2112 20700 2176 20704
rect 2112 20644 2116 20700
rect 2116 20644 2172 20700
rect 2172 20644 2176 20700
rect 2112 20640 2176 20644
rect 2192 20700 2256 20704
rect 2192 20644 2196 20700
rect 2196 20644 2252 20700
rect 2252 20644 2256 20700
rect 2192 20640 2256 20644
rect 85952 20700 86016 20704
rect 85952 20644 85956 20700
rect 85956 20644 86012 20700
rect 86012 20644 86016 20700
rect 85952 20640 86016 20644
rect 86032 20700 86096 20704
rect 86032 20644 86036 20700
rect 86036 20644 86092 20700
rect 86092 20644 86096 20700
rect 86032 20640 86096 20644
rect 86112 20700 86176 20704
rect 86112 20644 86116 20700
rect 86116 20644 86172 20700
rect 86172 20644 86176 20700
rect 86112 20640 86176 20644
rect 86192 20700 86256 20704
rect 86192 20644 86196 20700
rect 86196 20644 86252 20700
rect 86252 20644 86256 20700
rect 86192 20640 86256 20644
rect 89952 20700 90016 20704
rect 89952 20644 89956 20700
rect 89956 20644 90012 20700
rect 90012 20644 90016 20700
rect 89952 20640 90016 20644
rect 90032 20700 90096 20704
rect 90032 20644 90036 20700
rect 90036 20644 90092 20700
rect 90092 20644 90096 20700
rect 90032 20640 90096 20644
rect 90112 20700 90176 20704
rect 90112 20644 90116 20700
rect 90116 20644 90172 20700
rect 90172 20644 90176 20700
rect 90112 20640 90176 20644
rect 90192 20700 90256 20704
rect 90192 20644 90196 20700
rect 90196 20644 90252 20700
rect 90252 20644 90256 20700
rect 90192 20640 90256 20644
rect 3952 20156 4016 20160
rect 3952 20100 3956 20156
rect 3956 20100 4012 20156
rect 4012 20100 4016 20156
rect 3952 20096 4016 20100
rect 4032 20156 4096 20160
rect 4032 20100 4036 20156
rect 4036 20100 4092 20156
rect 4092 20100 4096 20156
rect 4032 20096 4096 20100
rect 4112 20156 4176 20160
rect 4112 20100 4116 20156
rect 4116 20100 4172 20156
rect 4172 20100 4176 20156
rect 4112 20096 4176 20100
rect 4192 20156 4256 20160
rect 4192 20100 4196 20156
rect 4196 20100 4252 20156
rect 4252 20100 4256 20156
rect 4192 20096 4256 20100
rect 87952 20156 88016 20160
rect 87952 20100 87956 20156
rect 87956 20100 88012 20156
rect 88012 20100 88016 20156
rect 87952 20096 88016 20100
rect 88032 20156 88096 20160
rect 88032 20100 88036 20156
rect 88036 20100 88092 20156
rect 88092 20100 88096 20156
rect 88032 20096 88096 20100
rect 88112 20156 88176 20160
rect 88112 20100 88116 20156
rect 88116 20100 88172 20156
rect 88172 20100 88176 20156
rect 88112 20096 88176 20100
rect 88192 20156 88256 20160
rect 88192 20100 88196 20156
rect 88196 20100 88252 20156
rect 88252 20100 88256 20156
rect 88192 20096 88256 20100
rect 1952 19612 2016 19616
rect 1952 19556 1956 19612
rect 1956 19556 2012 19612
rect 2012 19556 2016 19612
rect 1952 19552 2016 19556
rect 2032 19612 2096 19616
rect 2032 19556 2036 19612
rect 2036 19556 2092 19612
rect 2092 19556 2096 19612
rect 2032 19552 2096 19556
rect 2112 19612 2176 19616
rect 2112 19556 2116 19612
rect 2116 19556 2172 19612
rect 2172 19556 2176 19612
rect 2112 19552 2176 19556
rect 2192 19612 2256 19616
rect 2192 19556 2196 19612
rect 2196 19556 2252 19612
rect 2252 19556 2256 19612
rect 2192 19552 2256 19556
rect 85952 19612 86016 19616
rect 85952 19556 85956 19612
rect 85956 19556 86012 19612
rect 86012 19556 86016 19612
rect 85952 19552 86016 19556
rect 86032 19612 86096 19616
rect 86032 19556 86036 19612
rect 86036 19556 86092 19612
rect 86092 19556 86096 19612
rect 86032 19552 86096 19556
rect 86112 19612 86176 19616
rect 86112 19556 86116 19612
rect 86116 19556 86172 19612
rect 86172 19556 86176 19612
rect 86112 19552 86176 19556
rect 86192 19612 86256 19616
rect 86192 19556 86196 19612
rect 86196 19556 86252 19612
rect 86252 19556 86256 19612
rect 86192 19552 86256 19556
rect 89952 19612 90016 19616
rect 89952 19556 89956 19612
rect 89956 19556 90012 19612
rect 90012 19556 90016 19612
rect 89952 19552 90016 19556
rect 90032 19612 90096 19616
rect 90032 19556 90036 19612
rect 90036 19556 90092 19612
rect 90092 19556 90096 19612
rect 90032 19552 90096 19556
rect 90112 19612 90176 19616
rect 90112 19556 90116 19612
rect 90116 19556 90172 19612
rect 90172 19556 90176 19612
rect 90112 19552 90176 19556
rect 90192 19612 90256 19616
rect 90192 19556 90196 19612
rect 90196 19556 90252 19612
rect 90252 19556 90256 19612
rect 90192 19552 90256 19556
rect 3952 19068 4016 19072
rect 3952 19012 3956 19068
rect 3956 19012 4012 19068
rect 4012 19012 4016 19068
rect 3952 19008 4016 19012
rect 4032 19068 4096 19072
rect 4032 19012 4036 19068
rect 4036 19012 4092 19068
rect 4092 19012 4096 19068
rect 4032 19008 4096 19012
rect 4112 19068 4176 19072
rect 4112 19012 4116 19068
rect 4116 19012 4172 19068
rect 4172 19012 4176 19068
rect 4112 19008 4176 19012
rect 4192 19068 4256 19072
rect 4192 19012 4196 19068
rect 4196 19012 4252 19068
rect 4252 19012 4256 19068
rect 4192 19008 4256 19012
rect 87952 19068 88016 19072
rect 87952 19012 87956 19068
rect 87956 19012 88012 19068
rect 88012 19012 88016 19068
rect 87952 19008 88016 19012
rect 88032 19068 88096 19072
rect 88032 19012 88036 19068
rect 88036 19012 88092 19068
rect 88092 19012 88096 19068
rect 88032 19008 88096 19012
rect 88112 19068 88176 19072
rect 88112 19012 88116 19068
rect 88116 19012 88172 19068
rect 88172 19012 88176 19068
rect 88112 19008 88176 19012
rect 88192 19068 88256 19072
rect 88192 19012 88196 19068
rect 88196 19012 88252 19068
rect 88252 19012 88256 19068
rect 88192 19008 88256 19012
rect 1952 18524 2016 18528
rect 1952 18468 1956 18524
rect 1956 18468 2012 18524
rect 2012 18468 2016 18524
rect 1952 18464 2016 18468
rect 2032 18524 2096 18528
rect 2032 18468 2036 18524
rect 2036 18468 2092 18524
rect 2092 18468 2096 18524
rect 2032 18464 2096 18468
rect 2112 18524 2176 18528
rect 2112 18468 2116 18524
rect 2116 18468 2172 18524
rect 2172 18468 2176 18524
rect 2112 18464 2176 18468
rect 2192 18524 2256 18528
rect 2192 18468 2196 18524
rect 2196 18468 2252 18524
rect 2252 18468 2256 18524
rect 2192 18464 2256 18468
rect 85952 18524 86016 18528
rect 85952 18468 85956 18524
rect 85956 18468 86012 18524
rect 86012 18468 86016 18524
rect 85952 18464 86016 18468
rect 86032 18524 86096 18528
rect 86032 18468 86036 18524
rect 86036 18468 86092 18524
rect 86092 18468 86096 18524
rect 86032 18464 86096 18468
rect 86112 18524 86176 18528
rect 86112 18468 86116 18524
rect 86116 18468 86172 18524
rect 86172 18468 86176 18524
rect 86112 18464 86176 18468
rect 86192 18524 86256 18528
rect 86192 18468 86196 18524
rect 86196 18468 86252 18524
rect 86252 18468 86256 18524
rect 86192 18464 86256 18468
rect 89952 18524 90016 18528
rect 89952 18468 89956 18524
rect 89956 18468 90012 18524
rect 90012 18468 90016 18524
rect 89952 18464 90016 18468
rect 90032 18524 90096 18528
rect 90032 18468 90036 18524
rect 90036 18468 90092 18524
rect 90092 18468 90096 18524
rect 90032 18464 90096 18468
rect 90112 18524 90176 18528
rect 90112 18468 90116 18524
rect 90116 18468 90172 18524
rect 90172 18468 90176 18524
rect 90112 18464 90176 18468
rect 90192 18524 90256 18528
rect 90192 18468 90196 18524
rect 90196 18468 90252 18524
rect 90252 18468 90256 18524
rect 90192 18464 90256 18468
rect 3952 17980 4016 17984
rect 3952 17924 3956 17980
rect 3956 17924 4012 17980
rect 4012 17924 4016 17980
rect 3952 17920 4016 17924
rect 4032 17980 4096 17984
rect 4032 17924 4036 17980
rect 4036 17924 4092 17980
rect 4092 17924 4096 17980
rect 4032 17920 4096 17924
rect 4112 17980 4176 17984
rect 4112 17924 4116 17980
rect 4116 17924 4172 17980
rect 4172 17924 4176 17980
rect 4112 17920 4176 17924
rect 4192 17980 4256 17984
rect 4192 17924 4196 17980
rect 4196 17924 4252 17980
rect 4252 17924 4256 17980
rect 4192 17920 4256 17924
rect 87952 17980 88016 17984
rect 87952 17924 87956 17980
rect 87956 17924 88012 17980
rect 88012 17924 88016 17980
rect 87952 17920 88016 17924
rect 88032 17980 88096 17984
rect 88032 17924 88036 17980
rect 88036 17924 88092 17980
rect 88092 17924 88096 17980
rect 88032 17920 88096 17924
rect 88112 17980 88176 17984
rect 88112 17924 88116 17980
rect 88116 17924 88172 17980
rect 88172 17924 88176 17980
rect 88112 17920 88176 17924
rect 88192 17980 88256 17984
rect 88192 17924 88196 17980
rect 88196 17924 88252 17980
rect 88252 17924 88256 17980
rect 88192 17920 88256 17924
rect 1952 17436 2016 17440
rect 1952 17380 1956 17436
rect 1956 17380 2012 17436
rect 2012 17380 2016 17436
rect 1952 17376 2016 17380
rect 2032 17436 2096 17440
rect 2032 17380 2036 17436
rect 2036 17380 2092 17436
rect 2092 17380 2096 17436
rect 2032 17376 2096 17380
rect 2112 17436 2176 17440
rect 2112 17380 2116 17436
rect 2116 17380 2172 17436
rect 2172 17380 2176 17436
rect 2112 17376 2176 17380
rect 2192 17436 2256 17440
rect 2192 17380 2196 17436
rect 2196 17380 2252 17436
rect 2252 17380 2256 17436
rect 2192 17376 2256 17380
rect 85952 17436 86016 17440
rect 85952 17380 85956 17436
rect 85956 17380 86012 17436
rect 86012 17380 86016 17436
rect 85952 17376 86016 17380
rect 86032 17436 86096 17440
rect 86032 17380 86036 17436
rect 86036 17380 86092 17436
rect 86092 17380 86096 17436
rect 86032 17376 86096 17380
rect 86112 17436 86176 17440
rect 86112 17380 86116 17436
rect 86116 17380 86172 17436
rect 86172 17380 86176 17436
rect 86112 17376 86176 17380
rect 86192 17436 86256 17440
rect 86192 17380 86196 17436
rect 86196 17380 86252 17436
rect 86252 17380 86256 17436
rect 86192 17376 86256 17380
rect 89952 17436 90016 17440
rect 89952 17380 89956 17436
rect 89956 17380 90012 17436
rect 90012 17380 90016 17436
rect 89952 17376 90016 17380
rect 90032 17436 90096 17440
rect 90032 17380 90036 17436
rect 90036 17380 90092 17436
rect 90092 17380 90096 17436
rect 90032 17376 90096 17380
rect 90112 17436 90176 17440
rect 90112 17380 90116 17436
rect 90116 17380 90172 17436
rect 90172 17380 90176 17436
rect 90112 17376 90176 17380
rect 90192 17436 90256 17440
rect 90192 17380 90196 17436
rect 90196 17380 90252 17436
rect 90252 17380 90256 17436
rect 90192 17376 90256 17380
rect 3952 16892 4016 16896
rect 3952 16836 3956 16892
rect 3956 16836 4012 16892
rect 4012 16836 4016 16892
rect 3952 16832 4016 16836
rect 4032 16892 4096 16896
rect 4032 16836 4036 16892
rect 4036 16836 4092 16892
rect 4092 16836 4096 16892
rect 4032 16832 4096 16836
rect 4112 16892 4176 16896
rect 4112 16836 4116 16892
rect 4116 16836 4172 16892
rect 4172 16836 4176 16892
rect 4112 16832 4176 16836
rect 4192 16892 4256 16896
rect 4192 16836 4196 16892
rect 4196 16836 4252 16892
rect 4252 16836 4256 16892
rect 4192 16832 4256 16836
rect 87952 16892 88016 16896
rect 87952 16836 87956 16892
rect 87956 16836 88012 16892
rect 88012 16836 88016 16892
rect 87952 16832 88016 16836
rect 88032 16892 88096 16896
rect 88032 16836 88036 16892
rect 88036 16836 88092 16892
rect 88092 16836 88096 16892
rect 88032 16832 88096 16836
rect 88112 16892 88176 16896
rect 88112 16836 88116 16892
rect 88116 16836 88172 16892
rect 88172 16836 88176 16892
rect 88112 16832 88176 16836
rect 88192 16892 88256 16896
rect 88192 16836 88196 16892
rect 88196 16836 88252 16892
rect 88252 16836 88256 16892
rect 88192 16832 88256 16836
rect 84148 16628 84212 16692
rect 1952 16348 2016 16352
rect 1952 16292 1956 16348
rect 1956 16292 2012 16348
rect 2012 16292 2016 16348
rect 1952 16288 2016 16292
rect 2032 16348 2096 16352
rect 2032 16292 2036 16348
rect 2036 16292 2092 16348
rect 2092 16292 2096 16348
rect 2032 16288 2096 16292
rect 2112 16348 2176 16352
rect 2112 16292 2116 16348
rect 2116 16292 2172 16348
rect 2172 16292 2176 16348
rect 2112 16288 2176 16292
rect 2192 16348 2256 16352
rect 2192 16292 2196 16348
rect 2196 16292 2252 16348
rect 2252 16292 2256 16348
rect 2192 16288 2256 16292
rect 85952 16348 86016 16352
rect 85952 16292 85956 16348
rect 85956 16292 86012 16348
rect 86012 16292 86016 16348
rect 85952 16288 86016 16292
rect 86032 16348 86096 16352
rect 86032 16292 86036 16348
rect 86036 16292 86092 16348
rect 86092 16292 86096 16348
rect 86032 16288 86096 16292
rect 86112 16348 86176 16352
rect 86112 16292 86116 16348
rect 86116 16292 86172 16348
rect 86172 16292 86176 16348
rect 86112 16288 86176 16292
rect 86192 16348 86256 16352
rect 86192 16292 86196 16348
rect 86196 16292 86252 16348
rect 86252 16292 86256 16348
rect 86192 16288 86256 16292
rect 89952 16348 90016 16352
rect 89952 16292 89956 16348
rect 89956 16292 90012 16348
rect 90012 16292 90016 16348
rect 89952 16288 90016 16292
rect 90032 16348 90096 16352
rect 90032 16292 90036 16348
rect 90036 16292 90092 16348
rect 90092 16292 90096 16348
rect 90032 16288 90096 16292
rect 90112 16348 90176 16352
rect 90112 16292 90116 16348
rect 90116 16292 90172 16348
rect 90172 16292 90176 16348
rect 90112 16288 90176 16292
rect 90192 16348 90256 16352
rect 90192 16292 90196 16348
rect 90196 16292 90252 16348
rect 90252 16292 90256 16348
rect 90192 16288 90256 16292
rect 3952 15804 4016 15808
rect 3952 15748 3956 15804
rect 3956 15748 4012 15804
rect 4012 15748 4016 15804
rect 3952 15744 4016 15748
rect 4032 15804 4096 15808
rect 4032 15748 4036 15804
rect 4036 15748 4092 15804
rect 4092 15748 4096 15804
rect 4032 15744 4096 15748
rect 4112 15804 4176 15808
rect 4112 15748 4116 15804
rect 4116 15748 4172 15804
rect 4172 15748 4176 15804
rect 4112 15744 4176 15748
rect 4192 15804 4256 15808
rect 4192 15748 4196 15804
rect 4196 15748 4252 15804
rect 4252 15748 4256 15804
rect 4192 15744 4256 15748
rect 87952 15804 88016 15808
rect 87952 15748 87956 15804
rect 87956 15748 88012 15804
rect 88012 15748 88016 15804
rect 87952 15744 88016 15748
rect 88032 15804 88096 15808
rect 88032 15748 88036 15804
rect 88036 15748 88092 15804
rect 88092 15748 88096 15804
rect 88032 15744 88096 15748
rect 88112 15804 88176 15808
rect 88112 15748 88116 15804
rect 88116 15748 88172 15804
rect 88172 15748 88176 15804
rect 88112 15744 88176 15748
rect 88192 15804 88256 15808
rect 88192 15748 88196 15804
rect 88196 15748 88252 15804
rect 88252 15748 88256 15804
rect 88192 15744 88256 15748
rect 1952 15260 2016 15264
rect 1952 15204 1956 15260
rect 1956 15204 2012 15260
rect 2012 15204 2016 15260
rect 1952 15200 2016 15204
rect 2032 15260 2096 15264
rect 2032 15204 2036 15260
rect 2036 15204 2092 15260
rect 2092 15204 2096 15260
rect 2032 15200 2096 15204
rect 2112 15260 2176 15264
rect 2112 15204 2116 15260
rect 2116 15204 2172 15260
rect 2172 15204 2176 15260
rect 2112 15200 2176 15204
rect 2192 15260 2256 15264
rect 2192 15204 2196 15260
rect 2196 15204 2252 15260
rect 2252 15204 2256 15260
rect 2192 15200 2256 15204
rect 85952 15260 86016 15264
rect 85952 15204 85956 15260
rect 85956 15204 86012 15260
rect 86012 15204 86016 15260
rect 85952 15200 86016 15204
rect 86032 15260 86096 15264
rect 86032 15204 86036 15260
rect 86036 15204 86092 15260
rect 86092 15204 86096 15260
rect 86032 15200 86096 15204
rect 86112 15260 86176 15264
rect 86112 15204 86116 15260
rect 86116 15204 86172 15260
rect 86172 15204 86176 15260
rect 86112 15200 86176 15204
rect 86192 15260 86256 15264
rect 86192 15204 86196 15260
rect 86196 15204 86252 15260
rect 86252 15204 86256 15260
rect 86192 15200 86256 15204
rect 89952 15260 90016 15264
rect 89952 15204 89956 15260
rect 89956 15204 90012 15260
rect 90012 15204 90016 15260
rect 89952 15200 90016 15204
rect 90032 15260 90096 15264
rect 90032 15204 90036 15260
rect 90036 15204 90092 15260
rect 90092 15204 90096 15260
rect 90032 15200 90096 15204
rect 90112 15260 90176 15264
rect 90112 15204 90116 15260
rect 90116 15204 90172 15260
rect 90172 15204 90176 15260
rect 90112 15200 90176 15204
rect 90192 15260 90256 15264
rect 90192 15204 90196 15260
rect 90196 15204 90252 15260
rect 90252 15204 90256 15260
rect 90192 15200 90256 15204
rect 3952 14716 4016 14720
rect 3952 14660 3956 14716
rect 3956 14660 4012 14716
rect 4012 14660 4016 14716
rect 3952 14656 4016 14660
rect 4032 14716 4096 14720
rect 4032 14660 4036 14716
rect 4036 14660 4092 14716
rect 4092 14660 4096 14716
rect 4032 14656 4096 14660
rect 4112 14716 4176 14720
rect 4112 14660 4116 14716
rect 4116 14660 4172 14716
rect 4172 14660 4176 14716
rect 4112 14656 4176 14660
rect 4192 14716 4256 14720
rect 4192 14660 4196 14716
rect 4196 14660 4252 14716
rect 4252 14660 4256 14716
rect 4192 14656 4256 14660
rect 87952 14716 88016 14720
rect 87952 14660 87956 14716
rect 87956 14660 88012 14716
rect 88012 14660 88016 14716
rect 87952 14656 88016 14660
rect 88032 14716 88096 14720
rect 88032 14660 88036 14716
rect 88036 14660 88092 14716
rect 88092 14660 88096 14716
rect 88032 14656 88096 14660
rect 88112 14716 88176 14720
rect 88112 14660 88116 14716
rect 88116 14660 88172 14716
rect 88172 14660 88176 14716
rect 88112 14656 88176 14660
rect 88192 14716 88256 14720
rect 88192 14660 88196 14716
rect 88196 14660 88252 14716
rect 88252 14660 88256 14716
rect 88192 14656 88256 14660
rect 1952 14172 2016 14176
rect 1952 14116 1956 14172
rect 1956 14116 2012 14172
rect 2012 14116 2016 14172
rect 1952 14112 2016 14116
rect 2032 14172 2096 14176
rect 2032 14116 2036 14172
rect 2036 14116 2092 14172
rect 2092 14116 2096 14172
rect 2032 14112 2096 14116
rect 2112 14172 2176 14176
rect 2112 14116 2116 14172
rect 2116 14116 2172 14172
rect 2172 14116 2176 14172
rect 2112 14112 2176 14116
rect 2192 14172 2256 14176
rect 2192 14116 2196 14172
rect 2196 14116 2252 14172
rect 2252 14116 2256 14172
rect 2192 14112 2256 14116
rect 85952 14172 86016 14176
rect 85952 14116 85956 14172
rect 85956 14116 86012 14172
rect 86012 14116 86016 14172
rect 85952 14112 86016 14116
rect 86032 14172 86096 14176
rect 86032 14116 86036 14172
rect 86036 14116 86092 14172
rect 86092 14116 86096 14172
rect 86032 14112 86096 14116
rect 86112 14172 86176 14176
rect 86112 14116 86116 14172
rect 86116 14116 86172 14172
rect 86172 14116 86176 14172
rect 86112 14112 86176 14116
rect 86192 14172 86256 14176
rect 86192 14116 86196 14172
rect 86196 14116 86252 14172
rect 86252 14116 86256 14172
rect 86192 14112 86256 14116
rect 89952 14172 90016 14176
rect 89952 14116 89956 14172
rect 89956 14116 90012 14172
rect 90012 14116 90016 14172
rect 89952 14112 90016 14116
rect 90032 14172 90096 14176
rect 90032 14116 90036 14172
rect 90036 14116 90092 14172
rect 90092 14116 90096 14172
rect 90032 14112 90096 14116
rect 90112 14172 90176 14176
rect 90112 14116 90116 14172
rect 90116 14116 90172 14172
rect 90172 14116 90176 14172
rect 90112 14112 90176 14116
rect 90192 14172 90256 14176
rect 90192 14116 90196 14172
rect 90196 14116 90252 14172
rect 90252 14116 90256 14172
rect 90192 14112 90256 14116
rect 3952 13628 4016 13632
rect 3952 13572 3956 13628
rect 3956 13572 4012 13628
rect 4012 13572 4016 13628
rect 3952 13568 4016 13572
rect 4032 13628 4096 13632
rect 4032 13572 4036 13628
rect 4036 13572 4092 13628
rect 4092 13572 4096 13628
rect 4032 13568 4096 13572
rect 4112 13628 4176 13632
rect 4112 13572 4116 13628
rect 4116 13572 4172 13628
rect 4172 13572 4176 13628
rect 4112 13568 4176 13572
rect 4192 13628 4256 13632
rect 4192 13572 4196 13628
rect 4196 13572 4252 13628
rect 4252 13572 4256 13628
rect 4192 13568 4256 13572
rect 87952 13628 88016 13632
rect 87952 13572 87956 13628
rect 87956 13572 88012 13628
rect 88012 13572 88016 13628
rect 87952 13568 88016 13572
rect 88032 13628 88096 13632
rect 88032 13572 88036 13628
rect 88036 13572 88092 13628
rect 88092 13572 88096 13628
rect 88032 13568 88096 13572
rect 88112 13628 88176 13632
rect 88112 13572 88116 13628
rect 88116 13572 88172 13628
rect 88172 13572 88176 13628
rect 88112 13568 88176 13572
rect 88192 13628 88256 13632
rect 88192 13572 88196 13628
rect 88196 13572 88252 13628
rect 88252 13572 88256 13628
rect 88192 13568 88256 13572
rect 1952 13084 2016 13088
rect 1952 13028 1956 13084
rect 1956 13028 2012 13084
rect 2012 13028 2016 13084
rect 1952 13024 2016 13028
rect 2032 13084 2096 13088
rect 2032 13028 2036 13084
rect 2036 13028 2092 13084
rect 2092 13028 2096 13084
rect 2032 13024 2096 13028
rect 2112 13084 2176 13088
rect 2112 13028 2116 13084
rect 2116 13028 2172 13084
rect 2172 13028 2176 13084
rect 2112 13024 2176 13028
rect 2192 13084 2256 13088
rect 2192 13028 2196 13084
rect 2196 13028 2252 13084
rect 2252 13028 2256 13084
rect 2192 13024 2256 13028
rect 85952 13084 86016 13088
rect 85952 13028 85956 13084
rect 85956 13028 86012 13084
rect 86012 13028 86016 13084
rect 85952 13024 86016 13028
rect 86032 13084 86096 13088
rect 86032 13028 86036 13084
rect 86036 13028 86092 13084
rect 86092 13028 86096 13084
rect 86032 13024 86096 13028
rect 86112 13084 86176 13088
rect 86112 13028 86116 13084
rect 86116 13028 86172 13084
rect 86172 13028 86176 13084
rect 86112 13024 86176 13028
rect 86192 13084 86256 13088
rect 86192 13028 86196 13084
rect 86196 13028 86252 13084
rect 86252 13028 86256 13084
rect 86192 13024 86256 13028
rect 89952 13084 90016 13088
rect 89952 13028 89956 13084
rect 89956 13028 90012 13084
rect 90012 13028 90016 13084
rect 89952 13024 90016 13028
rect 90032 13084 90096 13088
rect 90032 13028 90036 13084
rect 90036 13028 90092 13084
rect 90092 13028 90096 13084
rect 90032 13024 90096 13028
rect 90112 13084 90176 13088
rect 90112 13028 90116 13084
rect 90116 13028 90172 13084
rect 90172 13028 90176 13084
rect 90112 13024 90176 13028
rect 90192 13084 90256 13088
rect 90192 13028 90196 13084
rect 90196 13028 90252 13084
rect 90252 13028 90256 13084
rect 90192 13024 90256 13028
rect 3952 12540 4016 12544
rect 3952 12484 3956 12540
rect 3956 12484 4012 12540
rect 4012 12484 4016 12540
rect 3952 12480 4016 12484
rect 4032 12540 4096 12544
rect 4032 12484 4036 12540
rect 4036 12484 4092 12540
rect 4092 12484 4096 12540
rect 4032 12480 4096 12484
rect 4112 12540 4176 12544
rect 4112 12484 4116 12540
rect 4116 12484 4172 12540
rect 4172 12484 4176 12540
rect 4112 12480 4176 12484
rect 4192 12540 4256 12544
rect 4192 12484 4196 12540
rect 4196 12484 4252 12540
rect 4252 12484 4256 12540
rect 4192 12480 4256 12484
rect 87952 12540 88016 12544
rect 87952 12484 87956 12540
rect 87956 12484 88012 12540
rect 88012 12484 88016 12540
rect 87952 12480 88016 12484
rect 88032 12540 88096 12544
rect 88032 12484 88036 12540
rect 88036 12484 88092 12540
rect 88092 12484 88096 12540
rect 88032 12480 88096 12484
rect 88112 12540 88176 12544
rect 88112 12484 88116 12540
rect 88116 12484 88172 12540
rect 88172 12484 88176 12540
rect 88112 12480 88176 12484
rect 88192 12540 88256 12544
rect 88192 12484 88196 12540
rect 88196 12484 88252 12540
rect 88252 12484 88256 12540
rect 88192 12480 88256 12484
rect 1952 11996 2016 12000
rect 1952 11940 1956 11996
rect 1956 11940 2012 11996
rect 2012 11940 2016 11996
rect 1952 11936 2016 11940
rect 2032 11996 2096 12000
rect 2032 11940 2036 11996
rect 2036 11940 2092 11996
rect 2092 11940 2096 11996
rect 2032 11936 2096 11940
rect 2112 11996 2176 12000
rect 2112 11940 2116 11996
rect 2116 11940 2172 11996
rect 2172 11940 2176 11996
rect 2112 11936 2176 11940
rect 2192 11996 2256 12000
rect 2192 11940 2196 11996
rect 2196 11940 2252 11996
rect 2252 11940 2256 11996
rect 2192 11936 2256 11940
rect 85952 11996 86016 12000
rect 85952 11940 85956 11996
rect 85956 11940 86012 11996
rect 86012 11940 86016 11996
rect 85952 11936 86016 11940
rect 86032 11996 86096 12000
rect 86032 11940 86036 11996
rect 86036 11940 86092 11996
rect 86092 11940 86096 11996
rect 86032 11936 86096 11940
rect 86112 11996 86176 12000
rect 86112 11940 86116 11996
rect 86116 11940 86172 11996
rect 86172 11940 86176 11996
rect 86112 11936 86176 11940
rect 86192 11996 86256 12000
rect 86192 11940 86196 11996
rect 86196 11940 86252 11996
rect 86252 11940 86256 11996
rect 86192 11936 86256 11940
rect 89952 11996 90016 12000
rect 89952 11940 89956 11996
rect 89956 11940 90012 11996
rect 90012 11940 90016 11996
rect 89952 11936 90016 11940
rect 90032 11996 90096 12000
rect 90032 11940 90036 11996
rect 90036 11940 90092 11996
rect 90092 11940 90096 11996
rect 90032 11936 90096 11940
rect 90112 11996 90176 12000
rect 90112 11940 90116 11996
rect 90116 11940 90172 11996
rect 90172 11940 90176 11996
rect 90112 11936 90176 11940
rect 90192 11996 90256 12000
rect 90192 11940 90196 11996
rect 90196 11940 90252 11996
rect 90252 11940 90256 11996
rect 90192 11936 90256 11940
rect 3952 11452 4016 11456
rect 3952 11396 3956 11452
rect 3956 11396 4012 11452
rect 4012 11396 4016 11452
rect 3952 11392 4016 11396
rect 4032 11452 4096 11456
rect 4032 11396 4036 11452
rect 4036 11396 4092 11452
rect 4092 11396 4096 11452
rect 4032 11392 4096 11396
rect 4112 11452 4176 11456
rect 4112 11396 4116 11452
rect 4116 11396 4172 11452
rect 4172 11396 4176 11452
rect 4112 11392 4176 11396
rect 4192 11452 4256 11456
rect 4192 11396 4196 11452
rect 4196 11396 4252 11452
rect 4252 11396 4256 11452
rect 4192 11392 4256 11396
rect 87952 11452 88016 11456
rect 87952 11396 87956 11452
rect 87956 11396 88012 11452
rect 88012 11396 88016 11452
rect 87952 11392 88016 11396
rect 88032 11452 88096 11456
rect 88032 11396 88036 11452
rect 88036 11396 88092 11452
rect 88092 11396 88096 11452
rect 88032 11392 88096 11396
rect 88112 11452 88176 11456
rect 88112 11396 88116 11452
rect 88116 11396 88172 11452
rect 88172 11396 88176 11452
rect 88112 11392 88176 11396
rect 88192 11452 88256 11456
rect 88192 11396 88196 11452
rect 88196 11396 88252 11452
rect 88252 11396 88256 11452
rect 88192 11392 88256 11396
rect 1952 10908 2016 10912
rect 1952 10852 1956 10908
rect 1956 10852 2012 10908
rect 2012 10852 2016 10908
rect 1952 10848 2016 10852
rect 2032 10908 2096 10912
rect 2032 10852 2036 10908
rect 2036 10852 2092 10908
rect 2092 10852 2096 10908
rect 2032 10848 2096 10852
rect 2112 10908 2176 10912
rect 2112 10852 2116 10908
rect 2116 10852 2172 10908
rect 2172 10852 2176 10908
rect 2112 10848 2176 10852
rect 2192 10908 2256 10912
rect 2192 10852 2196 10908
rect 2196 10852 2252 10908
rect 2252 10852 2256 10908
rect 2192 10848 2256 10852
rect 85952 10908 86016 10912
rect 85952 10852 85956 10908
rect 85956 10852 86012 10908
rect 86012 10852 86016 10908
rect 85952 10848 86016 10852
rect 86032 10908 86096 10912
rect 86032 10852 86036 10908
rect 86036 10852 86092 10908
rect 86092 10852 86096 10908
rect 86032 10848 86096 10852
rect 86112 10908 86176 10912
rect 86112 10852 86116 10908
rect 86116 10852 86172 10908
rect 86172 10852 86176 10908
rect 86112 10848 86176 10852
rect 86192 10908 86256 10912
rect 86192 10852 86196 10908
rect 86196 10852 86252 10908
rect 86252 10852 86256 10908
rect 86192 10848 86256 10852
rect 89952 10908 90016 10912
rect 89952 10852 89956 10908
rect 89956 10852 90012 10908
rect 90012 10852 90016 10908
rect 89952 10848 90016 10852
rect 90032 10908 90096 10912
rect 90032 10852 90036 10908
rect 90036 10852 90092 10908
rect 90092 10852 90096 10908
rect 90032 10848 90096 10852
rect 90112 10908 90176 10912
rect 90112 10852 90116 10908
rect 90116 10852 90172 10908
rect 90172 10852 90176 10908
rect 90112 10848 90176 10852
rect 90192 10908 90256 10912
rect 90192 10852 90196 10908
rect 90196 10852 90252 10908
rect 90252 10852 90256 10908
rect 90192 10848 90256 10852
rect 3952 10364 4016 10368
rect 3952 10308 3956 10364
rect 3956 10308 4012 10364
rect 4012 10308 4016 10364
rect 3952 10304 4016 10308
rect 4032 10364 4096 10368
rect 4032 10308 4036 10364
rect 4036 10308 4092 10364
rect 4092 10308 4096 10364
rect 4032 10304 4096 10308
rect 4112 10364 4176 10368
rect 4112 10308 4116 10364
rect 4116 10308 4172 10364
rect 4172 10308 4176 10364
rect 4112 10304 4176 10308
rect 4192 10364 4256 10368
rect 4192 10308 4196 10364
rect 4196 10308 4252 10364
rect 4252 10308 4256 10364
rect 4192 10304 4256 10308
rect 87952 10364 88016 10368
rect 87952 10308 87956 10364
rect 87956 10308 88012 10364
rect 88012 10308 88016 10364
rect 87952 10304 88016 10308
rect 88032 10364 88096 10368
rect 88032 10308 88036 10364
rect 88036 10308 88092 10364
rect 88092 10308 88096 10364
rect 88032 10304 88096 10308
rect 88112 10364 88176 10368
rect 88112 10308 88116 10364
rect 88116 10308 88172 10364
rect 88172 10308 88176 10364
rect 88112 10304 88176 10308
rect 88192 10364 88256 10368
rect 88192 10308 88196 10364
rect 88196 10308 88252 10364
rect 88252 10308 88256 10364
rect 88192 10304 88256 10308
rect 4476 10160 4540 10164
rect 4476 10104 4490 10160
rect 4490 10104 4540 10160
rect 4476 10100 4540 10104
rect 1952 9820 2016 9824
rect 1952 9764 1956 9820
rect 1956 9764 2012 9820
rect 2012 9764 2016 9820
rect 1952 9760 2016 9764
rect 2032 9820 2096 9824
rect 2032 9764 2036 9820
rect 2036 9764 2092 9820
rect 2092 9764 2096 9820
rect 2032 9760 2096 9764
rect 2112 9820 2176 9824
rect 2112 9764 2116 9820
rect 2116 9764 2172 9820
rect 2172 9764 2176 9820
rect 2112 9760 2176 9764
rect 2192 9820 2256 9824
rect 2192 9764 2196 9820
rect 2196 9764 2252 9820
rect 2252 9764 2256 9820
rect 2192 9760 2256 9764
rect 85952 9820 86016 9824
rect 85952 9764 85956 9820
rect 85956 9764 86012 9820
rect 86012 9764 86016 9820
rect 85952 9760 86016 9764
rect 86032 9820 86096 9824
rect 86032 9764 86036 9820
rect 86036 9764 86092 9820
rect 86092 9764 86096 9820
rect 86032 9760 86096 9764
rect 86112 9820 86176 9824
rect 86112 9764 86116 9820
rect 86116 9764 86172 9820
rect 86172 9764 86176 9820
rect 86112 9760 86176 9764
rect 86192 9820 86256 9824
rect 86192 9764 86196 9820
rect 86196 9764 86252 9820
rect 86252 9764 86256 9820
rect 86192 9760 86256 9764
rect 89952 9820 90016 9824
rect 89952 9764 89956 9820
rect 89956 9764 90012 9820
rect 90012 9764 90016 9820
rect 89952 9760 90016 9764
rect 90032 9820 90096 9824
rect 90032 9764 90036 9820
rect 90036 9764 90092 9820
rect 90092 9764 90096 9820
rect 90032 9760 90096 9764
rect 90112 9820 90176 9824
rect 90112 9764 90116 9820
rect 90116 9764 90172 9820
rect 90172 9764 90176 9820
rect 90112 9760 90176 9764
rect 90192 9820 90256 9824
rect 90192 9764 90196 9820
rect 90196 9764 90252 9820
rect 90252 9764 90256 9820
rect 90192 9760 90256 9764
rect 3952 9276 4016 9280
rect 3952 9220 3956 9276
rect 3956 9220 4012 9276
rect 4012 9220 4016 9276
rect 3952 9216 4016 9220
rect 4032 9276 4096 9280
rect 4032 9220 4036 9276
rect 4036 9220 4092 9276
rect 4092 9220 4096 9276
rect 4032 9216 4096 9220
rect 4112 9276 4176 9280
rect 4112 9220 4116 9276
rect 4116 9220 4172 9276
rect 4172 9220 4176 9276
rect 4112 9216 4176 9220
rect 4192 9276 4256 9280
rect 4192 9220 4196 9276
rect 4196 9220 4252 9276
rect 4252 9220 4256 9276
rect 4192 9216 4256 9220
rect 87952 9276 88016 9280
rect 87952 9220 87956 9276
rect 87956 9220 88012 9276
rect 88012 9220 88016 9276
rect 87952 9216 88016 9220
rect 88032 9276 88096 9280
rect 88032 9220 88036 9276
rect 88036 9220 88092 9276
rect 88092 9220 88096 9276
rect 88032 9216 88096 9220
rect 88112 9276 88176 9280
rect 88112 9220 88116 9276
rect 88116 9220 88172 9276
rect 88172 9220 88176 9276
rect 88112 9216 88176 9220
rect 88192 9276 88256 9280
rect 88192 9220 88196 9276
rect 88196 9220 88252 9276
rect 88252 9220 88256 9276
rect 88192 9216 88256 9220
rect 1952 8732 2016 8736
rect 1952 8676 1956 8732
rect 1956 8676 2012 8732
rect 2012 8676 2016 8732
rect 1952 8672 2016 8676
rect 2032 8732 2096 8736
rect 2032 8676 2036 8732
rect 2036 8676 2092 8732
rect 2092 8676 2096 8732
rect 2032 8672 2096 8676
rect 2112 8732 2176 8736
rect 2112 8676 2116 8732
rect 2116 8676 2172 8732
rect 2172 8676 2176 8732
rect 2112 8672 2176 8676
rect 2192 8732 2256 8736
rect 2192 8676 2196 8732
rect 2196 8676 2252 8732
rect 2252 8676 2256 8732
rect 2192 8672 2256 8676
rect 85952 8732 86016 8736
rect 85952 8676 85956 8732
rect 85956 8676 86012 8732
rect 86012 8676 86016 8732
rect 85952 8672 86016 8676
rect 86032 8732 86096 8736
rect 86032 8676 86036 8732
rect 86036 8676 86092 8732
rect 86092 8676 86096 8732
rect 86032 8672 86096 8676
rect 86112 8732 86176 8736
rect 86112 8676 86116 8732
rect 86116 8676 86172 8732
rect 86172 8676 86176 8732
rect 86112 8672 86176 8676
rect 86192 8732 86256 8736
rect 86192 8676 86196 8732
rect 86196 8676 86252 8732
rect 86252 8676 86256 8732
rect 86192 8672 86256 8676
rect 89952 8732 90016 8736
rect 89952 8676 89956 8732
rect 89956 8676 90012 8732
rect 90012 8676 90016 8732
rect 89952 8672 90016 8676
rect 90032 8732 90096 8736
rect 90032 8676 90036 8732
rect 90036 8676 90092 8732
rect 90092 8676 90096 8732
rect 90032 8672 90096 8676
rect 90112 8732 90176 8736
rect 90112 8676 90116 8732
rect 90116 8676 90172 8732
rect 90172 8676 90176 8732
rect 90112 8672 90176 8676
rect 90192 8732 90256 8736
rect 90192 8676 90196 8732
rect 90196 8676 90252 8732
rect 90252 8676 90256 8732
rect 90192 8672 90256 8676
rect 3952 8188 4016 8192
rect 3952 8132 3956 8188
rect 3956 8132 4012 8188
rect 4012 8132 4016 8188
rect 3952 8128 4016 8132
rect 4032 8188 4096 8192
rect 4032 8132 4036 8188
rect 4036 8132 4092 8188
rect 4092 8132 4096 8188
rect 4032 8128 4096 8132
rect 4112 8188 4176 8192
rect 4112 8132 4116 8188
rect 4116 8132 4172 8188
rect 4172 8132 4176 8188
rect 4112 8128 4176 8132
rect 4192 8188 4256 8192
rect 4192 8132 4196 8188
rect 4196 8132 4252 8188
rect 4252 8132 4256 8188
rect 4192 8128 4256 8132
rect 87952 8188 88016 8192
rect 87952 8132 87956 8188
rect 87956 8132 88012 8188
rect 88012 8132 88016 8188
rect 87952 8128 88016 8132
rect 88032 8188 88096 8192
rect 88032 8132 88036 8188
rect 88036 8132 88092 8188
rect 88092 8132 88096 8188
rect 88032 8128 88096 8132
rect 88112 8188 88176 8192
rect 88112 8132 88116 8188
rect 88116 8132 88172 8188
rect 88172 8132 88176 8188
rect 88112 8128 88176 8132
rect 88192 8188 88256 8192
rect 88192 8132 88196 8188
rect 88196 8132 88252 8188
rect 88252 8132 88256 8188
rect 88192 8128 88256 8132
rect 1952 7644 2016 7648
rect 1952 7588 1956 7644
rect 1956 7588 2012 7644
rect 2012 7588 2016 7644
rect 1952 7584 2016 7588
rect 2032 7644 2096 7648
rect 2032 7588 2036 7644
rect 2036 7588 2092 7644
rect 2092 7588 2096 7644
rect 2032 7584 2096 7588
rect 2112 7644 2176 7648
rect 2112 7588 2116 7644
rect 2116 7588 2172 7644
rect 2172 7588 2176 7644
rect 2112 7584 2176 7588
rect 2192 7644 2256 7648
rect 2192 7588 2196 7644
rect 2196 7588 2252 7644
rect 2252 7588 2256 7644
rect 2192 7584 2256 7588
rect 85952 7644 86016 7648
rect 85952 7588 85956 7644
rect 85956 7588 86012 7644
rect 86012 7588 86016 7644
rect 85952 7584 86016 7588
rect 86032 7644 86096 7648
rect 86032 7588 86036 7644
rect 86036 7588 86092 7644
rect 86092 7588 86096 7644
rect 86032 7584 86096 7588
rect 86112 7644 86176 7648
rect 86112 7588 86116 7644
rect 86116 7588 86172 7644
rect 86172 7588 86176 7644
rect 86112 7584 86176 7588
rect 86192 7644 86256 7648
rect 86192 7588 86196 7644
rect 86196 7588 86252 7644
rect 86252 7588 86256 7644
rect 86192 7584 86256 7588
rect 89952 7644 90016 7648
rect 89952 7588 89956 7644
rect 89956 7588 90012 7644
rect 90012 7588 90016 7644
rect 89952 7584 90016 7588
rect 90032 7644 90096 7648
rect 90032 7588 90036 7644
rect 90036 7588 90092 7644
rect 90092 7588 90096 7644
rect 90032 7584 90096 7588
rect 90112 7644 90176 7648
rect 90112 7588 90116 7644
rect 90116 7588 90172 7644
rect 90172 7588 90176 7644
rect 90112 7584 90176 7588
rect 90192 7644 90256 7648
rect 90192 7588 90196 7644
rect 90196 7588 90252 7644
rect 90252 7588 90256 7644
rect 90192 7584 90256 7588
rect 3952 7100 4016 7104
rect 3952 7044 3956 7100
rect 3956 7044 4012 7100
rect 4012 7044 4016 7100
rect 3952 7040 4016 7044
rect 4032 7100 4096 7104
rect 4032 7044 4036 7100
rect 4036 7044 4092 7100
rect 4092 7044 4096 7100
rect 4032 7040 4096 7044
rect 4112 7100 4176 7104
rect 4112 7044 4116 7100
rect 4116 7044 4172 7100
rect 4172 7044 4176 7100
rect 4112 7040 4176 7044
rect 4192 7100 4256 7104
rect 4192 7044 4196 7100
rect 4196 7044 4252 7100
rect 4252 7044 4256 7100
rect 4192 7040 4256 7044
rect 87952 7100 88016 7104
rect 87952 7044 87956 7100
rect 87956 7044 88012 7100
rect 88012 7044 88016 7100
rect 87952 7040 88016 7044
rect 88032 7100 88096 7104
rect 88032 7044 88036 7100
rect 88036 7044 88092 7100
rect 88092 7044 88096 7100
rect 88032 7040 88096 7044
rect 88112 7100 88176 7104
rect 88112 7044 88116 7100
rect 88116 7044 88172 7100
rect 88172 7044 88176 7100
rect 88112 7040 88176 7044
rect 88192 7100 88256 7104
rect 88192 7044 88196 7100
rect 88196 7044 88252 7100
rect 88252 7044 88256 7100
rect 88192 7040 88256 7044
rect 1952 6556 2016 6560
rect 1952 6500 1956 6556
rect 1956 6500 2012 6556
rect 2012 6500 2016 6556
rect 1952 6496 2016 6500
rect 2032 6556 2096 6560
rect 2032 6500 2036 6556
rect 2036 6500 2092 6556
rect 2092 6500 2096 6556
rect 2032 6496 2096 6500
rect 2112 6556 2176 6560
rect 2112 6500 2116 6556
rect 2116 6500 2172 6556
rect 2172 6500 2176 6556
rect 2112 6496 2176 6500
rect 2192 6556 2256 6560
rect 2192 6500 2196 6556
rect 2196 6500 2252 6556
rect 2252 6500 2256 6556
rect 2192 6496 2256 6500
rect 85952 6556 86016 6560
rect 85952 6500 85956 6556
rect 85956 6500 86012 6556
rect 86012 6500 86016 6556
rect 85952 6496 86016 6500
rect 86032 6556 86096 6560
rect 86032 6500 86036 6556
rect 86036 6500 86092 6556
rect 86092 6500 86096 6556
rect 86032 6496 86096 6500
rect 86112 6556 86176 6560
rect 86112 6500 86116 6556
rect 86116 6500 86172 6556
rect 86172 6500 86176 6556
rect 86112 6496 86176 6500
rect 86192 6556 86256 6560
rect 86192 6500 86196 6556
rect 86196 6500 86252 6556
rect 86252 6500 86256 6556
rect 86192 6496 86256 6500
rect 89952 6556 90016 6560
rect 89952 6500 89956 6556
rect 89956 6500 90012 6556
rect 90012 6500 90016 6556
rect 89952 6496 90016 6500
rect 90032 6556 90096 6560
rect 90032 6500 90036 6556
rect 90036 6500 90092 6556
rect 90092 6500 90096 6556
rect 90032 6496 90096 6500
rect 90112 6556 90176 6560
rect 90112 6500 90116 6556
rect 90116 6500 90172 6556
rect 90172 6500 90176 6556
rect 90112 6496 90176 6500
rect 90192 6556 90256 6560
rect 90192 6500 90196 6556
rect 90196 6500 90252 6556
rect 90252 6500 90256 6556
rect 90192 6496 90256 6500
rect 3952 6012 4016 6016
rect 3952 5956 3956 6012
rect 3956 5956 4012 6012
rect 4012 5956 4016 6012
rect 3952 5952 4016 5956
rect 4032 6012 4096 6016
rect 4032 5956 4036 6012
rect 4036 5956 4092 6012
rect 4092 5956 4096 6012
rect 4032 5952 4096 5956
rect 4112 6012 4176 6016
rect 4112 5956 4116 6012
rect 4116 5956 4172 6012
rect 4172 5956 4176 6012
rect 4112 5952 4176 5956
rect 4192 6012 4256 6016
rect 4192 5956 4196 6012
rect 4196 5956 4252 6012
rect 4252 5956 4256 6012
rect 4192 5952 4256 5956
rect 87952 6012 88016 6016
rect 87952 5956 87956 6012
rect 87956 5956 88012 6012
rect 88012 5956 88016 6012
rect 87952 5952 88016 5956
rect 88032 6012 88096 6016
rect 88032 5956 88036 6012
rect 88036 5956 88092 6012
rect 88092 5956 88096 6012
rect 88032 5952 88096 5956
rect 88112 6012 88176 6016
rect 88112 5956 88116 6012
rect 88116 5956 88172 6012
rect 88172 5956 88176 6012
rect 88112 5952 88176 5956
rect 88192 6012 88256 6016
rect 88192 5956 88196 6012
rect 88196 5956 88252 6012
rect 88252 5956 88256 6012
rect 88192 5952 88256 5956
rect 1952 5468 2016 5472
rect 1952 5412 1956 5468
rect 1956 5412 2012 5468
rect 2012 5412 2016 5468
rect 1952 5408 2016 5412
rect 2032 5468 2096 5472
rect 2032 5412 2036 5468
rect 2036 5412 2092 5468
rect 2092 5412 2096 5468
rect 2032 5408 2096 5412
rect 2112 5468 2176 5472
rect 2112 5412 2116 5468
rect 2116 5412 2172 5468
rect 2172 5412 2176 5468
rect 2112 5408 2176 5412
rect 2192 5468 2256 5472
rect 2192 5412 2196 5468
rect 2196 5412 2252 5468
rect 2252 5412 2256 5468
rect 2192 5408 2256 5412
rect 85952 5468 86016 5472
rect 85952 5412 85956 5468
rect 85956 5412 86012 5468
rect 86012 5412 86016 5468
rect 85952 5408 86016 5412
rect 86032 5468 86096 5472
rect 86032 5412 86036 5468
rect 86036 5412 86092 5468
rect 86092 5412 86096 5468
rect 86032 5408 86096 5412
rect 86112 5468 86176 5472
rect 86112 5412 86116 5468
rect 86116 5412 86172 5468
rect 86172 5412 86176 5468
rect 86112 5408 86176 5412
rect 86192 5468 86256 5472
rect 86192 5412 86196 5468
rect 86196 5412 86252 5468
rect 86252 5412 86256 5468
rect 86192 5408 86256 5412
rect 89952 5468 90016 5472
rect 89952 5412 89956 5468
rect 89956 5412 90012 5468
rect 90012 5412 90016 5468
rect 89952 5408 90016 5412
rect 90032 5468 90096 5472
rect 90032 5412 90036 5468
rect 90036 5412 90092 5468
rect 90092 5412 90096 5468
rect 90032 5408 90096 5412
rect 90112 5468 90176 5472
rect 90112 5412 90116 5468
rect 90116 5412 90172 5468
rect 90172 5412 90176 5468
rect 90112 5408 90176 5412
rect 90192 5468 90256 5472
rect 90192 5412 90196 5468
rect 90196 5412 90252 5468
rect 90252 5412 90256 5468
rect 90192 5408 90256 5412
rect 3952 4924 4016 4928
rect 3952 4868 3956 4924
rect 3956 4868 4012 4924
rect 4012 4868 4016 4924
rect 3952 4864 4016 4868
rect 4032 4924 4096 4928
rect 4032 4868 4036 4924
rect 4036 4868 4092 4924
rect 4092 4868 4096 4924
rect 4032 4864 4096 4868
rect 4112 4924 4176 4928
rect 4112 4868 4116 4924
rect 4116 4868 4172 4924
rect 4172 4868 4176 4924
rect 4112 4864 4176 4868
rect 4192 4924 4256 4928
rect 4192 4868 4196 4924
rect 4196 4868 4252 4924
rect 4252 4868 4256 4924
rect 4192 4864 4256 4868
rect 87952 4924 88016 4928
rect 87952 4868 87956 4924
rect 87956 4868 88012 4924
rect 88012 4868 88016 4924
rect 87952 4864 88016 4868
rect 88032 4924 88096 4928
rect 88032 4868 88036 4924
rect 88036 4868 88092 4924
rect 88092 4868 88096 4924
rect 88032 4864 88096 4868
rect 88112 4924 88176 4928
rect 88112 4868 88116 4924
rect 88116 4868 88172 4924
rect 88172 4868 88176 4924
rect 88112 4864 88176 4868
rect 88192 4924 88256 4928
rect 88192 4868 88196 4924
rect 88196 4868 88252 4924
rect 88252 4868 88256 4924
rect 88192 4864 88256 4868
rect 1952 4380 2016 4384
rect 1952 4324 1956 4380
rect 1956 4324 2012 4380
rect 2012 4324 2016 4380
rect 1952 4320 2016 4324
rect 2032 4380 2096 4384
rect 2032 4324 2036 4380
rect 2036 4324 2092 4380
rect 2092 4324 2096 4380
rect 2032 4320 2096 4324
rect 2112 4380 2176 4384
rect 2112 4324 2116 4380
rect 2116 4324 2172 4380
rect 2172 4324 2176 4380
rect 2112 4320 2176 4324
rect 2192 4380 2256 4384
rect 2192 4324 2196 4380
rect 2196 4324 2252 4380
rect 2252 4324 2256 4380
rect 2192 4320 2256 4324
rect 85952 4380 86016 4384
rect 85952 4324 85956 4380
rect 85956 4324 86012 4380
rect 86012 4324 86016 4380
rect 85952 4320 86016 4324
rect 86032 4380 86096 4384
rect 86032 4324 86036 4380
rect 86036 4324 86092 4380
rect 86092 4324 86096 4380
rect 86032 4320 86096 4324
rect 86112 4380 86176 4384
rect 86112 4324 86116 4380
rect 86116 4324 86172 4380
rect 86172 4324 86176 4380
rect 86112 4320 86176 4324
rect 86192 4380 86256 4384
rect 86192 4324 86196 4380
rect 86196 4324 86252 4380
rect 86252 4324 86256 4380
rect 86192 4320 86256 4324
rect 89952 4380 90016 4384
rect 89952 4324 89956 4380
rect 89956 4324 90012 4380
rect 90012 4324 90016 4380
rect 89952 4320 90016 4324
rect 90032 4380 90096 4384
rect 90032 4324 90036 4380
rect 90036 4324 90092 4380
rect 90092 4324 90096 4380
rect 90032 4320 90096 4324
rect 90112 4380 90176 4384
rect 90112 4324 90116 4380
rect 90116 4324 90172 4380
rect 90172 4324 90176 4380
rect 90112 4320 90176 4324
rect 90192 4380 90256 4384
rect 90192 4324 90196 4380
rect 90196 4324 90252 4380
rect 90252 4324 90256 4380
rect 90192 4320 90256 4324
rect 4844 3904 4908 3908
rect 4844 3848 4858 3904
rect 4858 3848 4908 3904
rect 4844 3844 4908 3848
rect 3952 3836 4016 3840
rect 3952 3780 3956 3836
rect 3956 3780 4012 3836
rect 4012 3780 4016 3836
rect 3952 3776 4016 3780
rect 4032 3836 4096 3840
rect 4032 3780 4036 3836
rect 4036 3780 4092 3836
rect 4092 3780 4096 3836
rect 4032 3776 4096 3780
rect 4112 3836 4176 3840
rect 4112 3780 4116 3836
rect 4116 3780 4172 3836
rect 4172 3780 4176 3836
rect 4112 3776 4176 3780
rect 4192 3836 4256 3840
rect 4192 3780 4196 3836
rect 4196 3780 4252 3836
rect 4252 3780 4256 3836
rect 4192 3776 4256 3780
rect 87952 3836 88016 3840
rect 87952 3780 87956 3836
rect 87956 3780 88012 3836
rect 88012 3780 88016 3836
rect 87952 3776 88016 3780
rect 88032 3836 88096 3840
rect 88032 3780 88036 3836
rect 88036 3780 88092 3836
rect 88092 3780 88096 3836
rect 88032 3776 88096 3780
rect 88112 3836 88176 3840
rect 88112 3780 88116 3836
rect 88116 3780 88172 3836
rect 88172 3780 88176 3836
rect 88112 3776 88176 3780
rect 88192 3836 88256 3840
rect 88192 3780 88196 3836
rect 88196 3780 88252 3836
rect 88252 3780 88256 3836
rect 88192 3776 88256 3780
rect 1952 3292 2016 3296
rect 1952 3236 1956 3292
rect 1956 3236 2012 3292
rect 2012 3236 2016 3292
rect 1952 3232 2016 3236
rect 2032 3292 2096 3296
rect 2032 3236 2036 3292
rect 2036 3236 2092 3292
rect 2092 3236 2096 3292
rect 2032 3232 2096 3236
rect 2112 3292 2176 3296
rect 2112 3236 2116 3292
rect 2116 3236 2172 3292
rect 2172 3236 2176 3292
rect 2112 3232 2176 3236
rect 2192 3292 2256 3296
rect 2192 3236 2196 3292
rect 2196 3236 2252 3292
rect 2252 3236 2256 3292
rect 2192 3232 2256 3236
rect 85952 3292 86016 3296
rect 85952 3236 85956 3292
rect 85956 3236 86012 3292
rect 86012 3236 86016 3292
rect 85952 3232 86016 3236
rect 86032 3292 86096 3296
rect 86032 3236 86036 3292
rect 86036 3236 86092 3292
rect 86092 3236 86096 3292
rect 86032 3232 86096 3236
rect 86112 3292 86176 3296
rect 86112 3236 86116 3292
rect 86116 3236 86172 3292
rect 86172 3236 86176 3292
rect 86112 3232 86176 3236
rect 86192 3292 86256 3296
rect 86192 3236 86196 3292
rect 86196 3236 86252 3292
rect 86252 3236 86256 3292
rect 86192 3232 86256 3236
rect 89952 3292 90016 3296
rect 89952 3236 89956 3292
rect 89956 3236 90012 3292
rect 90012 3236 90016 3292
rect 89952 3232 90016 3236
rect 90032 3292 90096 3296
rect 90032 3236 90036 3292
rect 90036 3236 90092 3292
rect 90092 3236 90096 3292
rect 90032 3232 90096 3236
rect 90112 3292 90176 3296
rect 90112 3236 90116 3292
rect 90116 3236 90172 3292
rect 90172 3236 90176 3292
rect 90112 3232 90176 3236
rect 90192 3292 90256 3296
rect 90192 3236 90196 3292
rect 90196 3236 90252 3292
rect 90252 3236 90256 3292
rect 90192 3232 90256 3236
rect 39068 3164 39132 3228
rect 45324 3164 45388 3228
rect 40172 3028 40236 3092
rect 47716 3224 47780 3228
rect 47716 3168 47766 3224
rect 47766 3168 47780 3224
rect 47716 3164 47780 3168
rect 37964 2892 38028 2956
rect 44036 2892 44100 2956
rect 49924 2952 49988 2956
rect 49924 2896 49974 2952
rect 49974 2896 49988 2952
rect 49924 2892 49988 2896
rect 53420 2952 53484 2956
rect 53420 2896 53470 2952
rect 53470 2896 53484 2952
rect 53420 2892 53484 2896
rect 26004 2756 26068 2820
rect 46244 2756 46308 2820
rect 3952 2748 4016 2752
rect 3952 2692 3956 2748
rect 3956 2692 4012 2748
rect 4012 2692 4016 2748
rect 3952 2688 4016 2692
rect 4032 2748 4096 2752
rect 4032 2692 4036 2748
rect 4036 2692 4092 2748
rect 4092 2692 4096 2748
rect 4032 2688 4096 2692
rect 4112 2748 4176 2752
rect 4112 2692 4116 2748
rect 4116 2692 4172 2748
rect 4172 2692 4176 2748
rect 4112 2688 4176 2692
rect 4192 2748 4256 2752
rect 4192 2692 4196 2748
rect 4196 2692 4252 2748
rect 4252 2692 4256 2748
rect 4192 2688 4256 2692
rect 87952 2748 88016 2752
rect 87952 2692 87956 2748
rect 87956 2692 88012 2748
rect 88012 2692 88016 2748
rect 87952 2688 88016 2692
rect 88032 2748 88096 2752
rect 88032 2692 88036 2748
rect 88036 2692 88092 2748
rect 88092 2692 88096 2748
rect 88032 2688 88096 2692
rect 88112 2748 88176 2752
rect 88112 2692 88116 2748
rect 88116 2692 88172 2748
rect 88172 2692 88176 2748
rect 88112 2688 88176 2692
rect 88192 2748 88256 2752
rect 88192 2692 88196 2748
rect 88196 2692 88252 2748
rect 88252 2692 88256 2748
rect 88192 2688 88256 2692
rect 8156 2680 8220 2684
rect 8156 2624 8170 2680
rect 8170 2624 8220 2680
rect 8156 2620 8220 2624
rect 15332 2680 15396 2684
rect 15332 2624 15346 2680
rect 15346 2624 15396 2680
rect 15332 2620 15396 2624
rect 20668 2680 20732 2684
rect 20668 2624 20718 2680
rect 20718 2624 20732 2680
rect 20668 2620 20732 2624
rect 25084 2680 25148 2684
rect 25084 2624 25098 2680
rect 25098 2624 25148 2680
rect 25084 2620 25148 2624
rect 22692 2544 22756 2548
rect 22692 2488 22706 2544
rect 22706 2488 22756 2544
rect 22692 2484 22756 2488
rect 9801 2272 9865 2276
rect 9801 2216 9826 2272
rect 9826 2216 9865 2272
rect 9801 2212 9865 2216
rect 13968 2212 14032 2276
rect 16304 2272 16368 2276
rect 16304 2216 16358 2272
rect 16358 2216 16368 2272
rect 16304 2212 16368 2216
rect 22144 2272 22208 2276
rect 22144 2216 22154 2272
rect 22154 2216 22208 2272
rect 22144 2212 22208 2216
rect 24480 2212 24544 2276
rect 32656 2272 32720 2276
rect 32656 2216 32678 2272
rect 32678 2216 32720 2272
rect 32656 2212 32720 2216
rect 36160 2272 36224 2276
rect 36160 2216 36174 2272
rect 36174 2216 36224 2272
rect 36160 2212 36224 2216
rect 37452 2272 37516 2276
rect 37452 2216 37462 2272
rect 37462 2216 37516 2272
rect 37452 2212 37516 2216
rect 51344 2272 51408 2276
rect 51344 2216 51354 2272
rect 51354 2216 51408 2272
rect 51344 2212 51408 2216
rect 52512 2272 52576 2276
rect 52512 2216 52550 2272
rect 52550 2216 52576 2272
rect 52512 2212 52576 2216
rect 1952 2204 2016 2208
rect 1952 2148 1956 2204
rect 1956 2148 2012 2204
rect 2012 2148 2016 2204
rect 1952 2144 2016 2148
rect 2032 2204 2096 2208
rect 2032 2148 2036 2204
rect 2036 2148 2092 2204
rect 2092 2148 2096 2204
rect 2032 2144 2096 2148
rect 2112 2204 2176 2208
rect 2112 2148 2116 2204
rect 2116 2148 2172 2204
rect 2172 2148 2176 2204
rect 2112 2144 2176 2148
rect 2192 2204 2256 2208
rect 2192 2148 2196 2204
rect 2196 2148 2252 2204
rect 2252 2148 2256 2204
rect 2192 2144 2256 2148
rect 85952 2204 86016 2208
rect 85952 2148 85956 2204
rect 85956 2148 86012 2204
rect 86012 2148 86016 2204
rect 85952 2144 86016 2148
rect 86032 2204 86096 2208
rect 86032 2148 86036 2204
rect 86036 2148 86092 2204
rect 86092 2148 86096 2204
rect 86032 2144 86096 2148
rect 86112 2204 86176 2208
rect 86112 2148 86116 2204
rect 86116 2148 86172 2204
rect 86172 2148 86176 2204
rect 86112 2144 86176 2148
rect 86192 2204 86256 2208
rect 86192 2148 86196 2204
rect 86196 2148 86252 2204
rect 86252 2148 86256 2204
rect 86192 2144 86256 2148
rect 89952 2204 90016 2208
rect 89952 2148 89956 2204
rect 89956 2148 90012 2204
rect 90012 2148 90016 2204
rect 89952 2144 90016 2148
rect 90032 2204 90096 2208
rect 90032 2148 90036 2204
rect 90036 2148 90092 2204
rect 90092 2148 90096 2204
rect 90032 2144 90096 2148
rect 90112 2204 90176 2208
rect 90112 2148 90116 2204
rect 90116 2148 90172 2204
rect 90172 2148 90176 2204
rect 90112 2144 90176 2148
rect 90192 2204 90256 2208
rect 90192 2148 90196 2204
rect 90196 2148 90252 2204
rect 90252 2148 90256 2204
rect 90192 2144 90256 2148
rect 32780 2136 32844 2140
rect 32780 2080 32826 2136
rect 32826 2080 32844 2136
rect 32780 2076 32844 2080
rect 33948 2136 34012 2140
rect 33948 2080 33966 2136
rect 33966 2080 34012 2136
rect 33948 2076 34012 2080
rect 36284 2136 36348 2140
rect 36284 2080 36322 2136
rect 36322 2080 36348 2136
rect 36284 2076 36348 2080
rect 29152 1940 29216 2004
rect 30444 2000 30508 2004
rect 30444 1944 30470 2000
rect 30470 1944 30508 2000
rect 30444 1940 30508 1944
rect 31612 2000 31676 2004
rect 31612 1944 31666 2000
rect 31666 1944 31676 2000
rect 31612 1940 31676 1944
rect 17472 1864 17536 1868
rect 17472 1808 17498 1864
rect 17498 1808 17536 1864
rect 17472 1804 17536 1808
rect 21100 1864 21164 1868
rect 21100 1808 21142 1864
rect 21142 1808 21164 1864
rect 21100 1804 21164 1808
rect 22268 1864 22332 1868
rect 22268 1808 22282 1864
rect 22282 1808 22332 1864
rect 22268 1804 22332 1808
rect 25772 1864 25836 1868
rect 25772 1808 25778 1864
rect 25778 1808 25834 1864
rect 25834 1808 25836 1864
rect 25772 1804 25836 1808
rect 26940 1864 27004 1868
rect 26940 1808 26974 1864
rect 26974 1808 27004 1864
rect 26940 1804 27004 1808
rect 28108 1864 28172 1868
rect 28108 1808 28170 1864
rect 28170 1808 28172 1864
rect 28108 1804 28172 1808
rect 49004 1532 49068 1596
rect 83412 1396 83476 1460
rect 12756 1260 12820 1324
rect 18828 1260 18892 1324
rect 29316 1260 29380 1324
rect 35204 1260 35268 1324
rect 39252 1260 39316 1324
rect 44772 1260 44836 1324
rect 48084 1260 48148 1324
rect 18644 1124 18708 1188
rect 19748 1124 19812 1188
rect 29684 1124 29748 1188
rect 34836 1124 34900 1188
rect 39804 1124 39868 1188
rect 52132 1124 52196 1188
rect 24716 1048 24780 1052
rect 24716 992 24766 1048
rect 24766 992 24780 1048
rect 24716 988 24780 992
rect 30972 988 31036 1052
rect 41276 1048 41340 1052
rect 41276 992 41326 1048
rect 41326 992 41340 1048
rect 41276 988 41340 992
rect 42564 988 42628 1052
rect 45692 988 45756 1052
rect 49188 988 49252 1052
rect 53788 988 53852 1052
rect 27660 912 27724 916
rect 27660 856 27674 912
rect 27674 856 27724 912
rect 27660 852 27724 856
rect 43116 852 43180 916
rect 43300 852 43364 916
rect 46796 912 46860 916
rect 46796 856 46846 912
rect 46846 856 46860 912
rect 46796 852 46860 856
rect 23428 716 23492 780
rect 33732 716 33796 780
rect 50292 716 50356 780
rect 54708 716 54772 780
rect 52684 444 52748 508
rect 55076 504 55140 508
rect 55076 448 55126 504
rect 55126 448 55140 504
rect 55076 444 55140 448
rect 19932 172 19996 236
<< metal4 >>
rect 89299 191452 89365 191453
rect 89299 191388 89300 191452
rect 89364 191388 89365 191452
rect 89299 191387 89365 191388
rect 88931 190228 88997 190229
rect 88931 190164 88932 190228
rect 88996 190164 88997 190228
rect 88931 190163 88997 190164
rect 1944 189344 2264 189360
rect 1944 189280 1952 189344
rect 2016 189280 2032 189344
rect 2096 189280 2112 189344
rect 2176 189280 2192 189344
rect 2256 189280 2264 189344
rect 1944 188256 2264 189280
rect 1944 188192 1952 188256
rect 2016 188192 2032 188256
rect 2096 188192 2112 188256
rect 2176 188192 2192 188256
rect 2256 188192 2264 188256
rect 1944 187168 2264 188192
rect 1944 187104 1952 187168
rect 2016 187104 2032 187168
rect 2096 187104 2112 187168
rect 2176 187104 2192 187168
rect 2256 187104 2264 187168
rect 1944 186080 2264 187104
rect 1944 186016 1952 186080
rect 2016 186016 2032 186080
rect 2096 186016 2112 186080
rect 2176 186016 2192 186080
rect 2256 186016 2264 186080
rect 1944 185576 2264 186016
rect 1944 185340 1986 185576
rect 2222 185340 2264 185576
rect 1944 184992 2264 185340
rect 1944 184928 1952 184992
rect 2016 184928 2032 184992
rect 2096 184928 2112 184992
rect 2176 184928 2192 184992
rect 2256 184928 2264 184992
rect 1944 183904 2264 184928
rect 1944 183840 1952 183904
rect 2016 183840 2032 183904
rect 2096 183840 2112 183904
rect 2176 183840 2192 183904
rect 2256 183840 2264 183904
rect 1944 182816 2264 183840
rect 1944 182752 1952 182816
rect 2016 182752 2032 182816
rect 2096 182752 2112 182816
rect 2176 182752 2192 182816
rect 2256 182752 2264 182816
rect 1944 181728 2264 182752
rect 1944 181664 1952 181728
rect 2016 181664 2032 181728
rect 2096 181664 2112 181728
rect 2176 181664 2192 181728
rect 2256 181664 2264 181728
rect 1944 180640 2264 181664
rect 1944 180576 1952 180640
rect 2016 180576 2032 180640
rect 2096 180576 2112 180640
rect 2176 180576 2192 180640
rect 2256 180576 2264 180640
rect 1944 179552 2264 180576
rect 1944 179488 1952 179552
rect 2016 179488 2032 179552
rect 2096 179488 2112 179552
rect 2176 179488 2192 179552
rect 2256 179488 2264 179552
rect 1944 178464 2264 179488
rect 1944 178400 1952 178464
rect 2016 178400 2032 178464
rect 2096 178400 2112 178464
rect 2176 178400 2192 178464
rect 2256 178400 2264 178464
rect 1944 177376 2264 178400
rect 1944 177312 1952 177376
rect 2016 177312 2032 177376
rect 2096 177312 2112 177376
rect 2176 177312 2192 177376
rect 2256 177312 2264 177376
rect 1944 176288 2264 177312
rect 1944 176224 1952 176288
rect 2016 176224 2032 176288
rect 2096 176224 2112 176288
rect 2176 176224 2192 176288
rect 2256 176224 2264 176288
rect 1944 175576 2264 176224
rect 1944 175340 1986 175576
rect 2222 175340 2264 175576
rect 1944 175200 2264 175340
rect 1944 175136 1952 175200
rect 2016 175136 2032 175200
rect 2096 175136 2112 175200
rect 2176 175136 2192 175200
rect 2256 175136 2264 175200
rect 1944 174112 2264 175136
rect 1944 174048 1952 174112
rect 2016 174048 2032 174112
rect 2096 174048 2112 174112
rect 2176 174048 2192 174112
rect 2256 174048 2264 174112
rect 1944 173024 2264 174048
rect 1944 172960 1952 173024
rect 2016 172960 2032 173024
rect 2096 172960 2112 173024
rect 2176 172960 2192 173024
rect 2256 172960 2264 173024
rect 1944 171936 2264 172960
rect 1944 171872 1952 171936
rect 2016 171872 2032 171936
rect 2096 171872 2112 171936
rect 2176 171872 2192 171936
rect 2256 171872 2264 171936
rect 1944 170848 2264 171872
rect 1944 170784 1952 170848
rect 2016 170784 2032 170848
rect 2096 170784 2112 170848
rect 2176 170784 2192 170848
rect 2256 170784 2264 170848
rect 1944 169760 2264 170784
rect 1944 169696 1952 169760
rect 2016 169696 2032 169760
rect 2096 169696 2112 169760
rect 2176 169696 2192 169760
rect 2256 169696 2264 169760
rect 1944 168672 2264 169696
rect 1944 168608 1952 168672
rect 2016 168608 2032 168672
rect 2096 168608 2112 168672
rect 2176 168608 2192 168672
rect 2256 168608 2264 168672
rect 1944 167584 2264 168608
rect 1944 167520 1952 167584
rect 2016 167520 2032 167584
rect 2096 167520 2112 167584
rect 2176 167520 2192 167584
rect 2256 167520 2264 167584
rect 1944 166496 2264 167520
rect 1944 166432 1952 166496
rect 2016 166432 2032 166496
rect 2096 166432 2112 166496
rect 2176 166432 2192 166496
rect 2256 166432 2264 166496
rect 1944 165576 2264 166432
rect 1944 165408 1986 165576
rect 2222 165408 2264 165576
rect 1944 165344 1952 165408
rect 2256 165344 2264 165408
rect 1944 165340 1986 165344
rect 2222 165340 2264 165344
rect 1944 164320 2264 165340
rect 1944 164256 1952 164320
rect 2016 164256 2032 164320
rect 2096 164256 2112 164320
rect 2176 164256 2192 164320
rect 2256 164256 2264 164320
rect 1944 163232 2264 164256
rect 1944 163168 1952 163232
rect 2016 163168 2032 163232
rect 2096 163168 2112 163232
rect 2176 163168 2192 163232
rect 2256 163168 2264 163232
rect 1944 162144 2264 163168
rect 1944 162080 1952 162144
rect 2016 162080 2032 162144
rect 2096 162080 2112 162144
rect 2176 162080 2192 162144
rect 2256 162080 2264 162144
rect 1944 161056 2264 162080
rect 1944 160992 1952 161056
rect 2016 160992 2032 161056
rect 2096 160992 2112 161056
rect 2176 160992 2192 161056
rect 2256 160992 2264 161056
rect 1944 159968 2264 160992
rect 1944 159904 1952 159968
rect 2016 159904 2032 159968
rect 2096 159904 2112 159968
rect 2176 159904 2192 159968
rect 2256 159904 2264 159968
rect 1944 158880 2264 159904
rect 1944 158816 1952 158880
rect 2016 158816 2032 158880
rect 2096 158816 2112 158880
rect 2176 158816 2192 158880
rect 2256 158816 2264 158880
rect 1944 157792 2264 158816
rect 1944 157728 1952 157792
rect 2016 157728 2032 157792
rect 2096 157728 2112 157792
rect 2176 157728 2192 157792
rect 2256 157728 2264 157792
rect 1944 156704 2264 157728
rect 1944 156640 1952 156704
rect 2016 156640 2032 156704
rect 2096 156640 2112 156704
rect 2176 156640 2192 156704
rect 2256 156640 2264 156704
rect 1944 155616 2264 156640
rect 1944 155552 1952 155616
rect 2016 155576 2032 155616
rect 2096 155576 2112 155616
rect 2176 155576 2192 155616
rect 2256 155552 2264 155616
rect 1944 155340 1986 155552
rect 2222 155340 2264 155552
rect 1944 154528 2264 155340
rect 1944 154464 1952 154528
rect 2016 154464 2032 154528
rect 2096 154464 2112 154528
rect 2176 154464 2192 154528
rect 2256 154464 2264 154528
rect 1944 153440 2264 154464
rect 1944 153376 1952 153440
rect 2016 153376 2032 153440
rect 2096 153376 2112 153440
rect 2176 153376 2192 153440
rect 2256 153376 2264 153440
rect 1944 152352 2264 153376
rect 1944 152288 1952 152352
rect 2016 152288 2032 152352
rect 2096 152288 2112 152352
rect 2176 152288 2192 152352
rect 2256 152288 2264 152352
rect 1944 151264 2264 152288
rect 1944 151200 1952 151264
rect 2016 151200 2032 151264
rect 2096 151200 2112 151264
rect 2176 151200 2192 151264
rect 2256 151200 2264 151264
rect 1944 150176 2264 151200
rect 1944 150112 1952 150176
rect 2016 150112 2032 150176
rect 2096 150112 2112 150176
rect 2176 150112 2192 150176
rect 2256 150112 2264 150176
rect 1944 149088 2264 150112
rect 1944 149024 1952 149088
rect 2016 149024 2032 149088
rect 2096 149024 2112 149088
rect 2176 149024 2192 149088
rect 2256 149024 2264 149088
rect 1944 148000 2264 149024
rect 1944 147936 1952 148000
rect 2016 147936 2032 148000
rect 2096 147936 2112 148000
rect 2176 147936 2192 148000
rect 2256 147936 2264 148000
rect 1944 146912 2264 147936
rect 1944 146848 1952 146912
rect 2016 146848 2032 146912
rect 2096 146848 2112 146912
rect 2176 146848 2192 146912
rect 2256 146848 2264 146912
rect 1944 145824 2264 146848
rect 1944 145760 1952 145824
rect 2016 145760 2032 145824
rect 2096 145760 2112 145824
rect 2176 145760 2192 145824
rect 2256 145760 2264 145824
rect 1944 145576 2264 145760
rect 1944 145340 1986 145576
rect 2222 145340 2264 145576
rect 1944 144736 2264 145340
rect 1944 144672 1952 144736
rect 2016 144672 2032 144736
rect 2096 144672 2112 144736
rect 2176 144672 2192 144736
rect 2256 144672 2264 144736
rect 1944 143648 2264 144672
rect 1944 143584 1952 143648
rect 2016 143584 2032 143648
rect 2096 143584 2112 143648
rect 2176 143584 2192 143648
rect 2256 143584 2264 143648
rect 1944 142560 2264 143584
rect 1944 142496 1952 142560
rect 2016 142496 2032 142560
rect 2096 142496 2112 142560
rect 2176 142496 2192 142560
rect 2256 142496 2264 142560
rect 1944 141472 2264 142496
rect 1944 141408 1952 141472
rect 2016 141408 2032 141472
rect 2096 141408 2112 141472
rect 2176 141408 2192 141472
rect 2256 141408 2264 141472
rect 1944 140384 2264 141408
rect 1944 140320 1952 140384
rect 2016 140320 2032 140384
rect 2096 140320 2112 140384
rect 2176 140320 2192 140384
rect 2256 140320 2264 140384
rect 1944 139296 2264 140320
rect 1944 139232 1952 139296
rect 2016 139232 2032 139296
rect 2096 139232 2112 139296
rect 2176 139232 2192 139296
rect 2256 139232 2264 139296
rect 1944 138208 2264 139232
rect 1944 138144 1952 138208
rect 2016 138144 2032 138208
rect 2096 138144 2112 138208
rect 2176 138144 2192 138208
rect 2256 138144 2264 138208
rect 1944 137120 2264 138144
rect 1944 137056 1952 137120
rect 2016 137056 2032 137120
rect 2096 137056 2112 137120
rect 2176 137056 2192 137120
rect 2256 137056 2264 137120
rect 1944 136032 2264 137056
rect 1944 135968 1952 136032
rect 2016 135968 2032 136032
rect 2096 135968 2112 136032
rect 2176 135968 2192 136032
rect 2256 135968 2264 136032
rect 1944 135576 2264 135968
rect 1944 135340 1986 135576
rect 2222 135340 2264 135576
rect 1944 134944 2264 135340
rect 1944 134880 1952 134944
rect 2016 134880 2032 134944
rect 2096 134880 2112 134944
rect 2176 134880 2192 134944
rect 2256 134880 2264 134944
rect 1944 133856 2264 134880
rect 1944 133792 1952 133856
rect 2016 133792 2032 133856
rect 2096 133792 2112 133856
rect 2176 133792 2192 133856
rect 2256 133792 2264 133856
rect 1944 132768 2264 133792
rect 1944 132704 1952 132768
rect 2016 132704 2032 132768
rect 2096 132704 2112 132768
rect 2176 132704 2192 132768
rect 2256 132704 2264 132768
rect 1944 131680 2264 132704
rect 1944 131616 1952 131680
rect 2016 131616 2032 131680
rect 2096 131616 2112 131680
rect 2176 131616 2192 131680
rect 2256 131616 2264 131680
rect 1944 130592 2264 131616
rect 1944 130528 1952 130592
rect 2016 130528 2032 130592
rect 2096 130528 2112 130592
rect 2176 130528 2192 130592
rect 2256 130528 2264 130592
rect 1944 129504 2264 130528
rect 1944 129440 1952 129504
rect 2016 129440 2032 129504
rect 2096 129440 2112 129504
rect 2176 129440 2192 129504
rect 2256 129440 2264 129504
rect 1944 128416 2264 129440
rect 1944 128352 1952 128416
rect 2016 128352 2032 128416
rect 2096 128352 2112 128416
rect 2176 128352 2192 128416
rect 2256 128352 2264 128416
rect 1944 127328 2264 128352
rect 1944 127264 1952 127328
rect 2016 127264 2032 127328
rect 2096 127264 2112 127328
rect 2176 127264 2192 127328
rect 2256 127264 2264 127328
rect 1944 126240 2264 127264
rect 1944 126176 1952 126240
rect 2016 126176 2032 126240
rect 2096 126176 2112 126240
rect 2176 126176 2192 126240
rect 2256 126176 2264 126240
rect 1944 125576 2264 126176
rect 1944 125340 1986 125576
rect 2222 125340 2264 125576
rect 1944 125152 2264 125340
rect 1944 125088 1952 125152
rect 2016 125088 2032 125152
rect 2096 125088 2112 125152
rect 2176 125088 2192 125152
rect 2256 125088 2264 125152
rect 1944 124064 2264 125088
rect 1944 124000 1952 124064
rect 2016 124000 2032 124064
rect 2096 124000 2112 124064
rect 2176 124000 2192 124064
rect 2256 124000 2264 124064
rect 1944 122976 2264 124000
rect 1944 122912 1952 122976
rect 2016 122912 2032 122976
rect 2096 122912 2112 122976
rect 2176 122912 2192 122976
rect 2256 122912 2264 122976
rect 1944 121888 2264 122912
rect 1944 121824 1952 121888
rect 2016 121824 2032 121888
rect 2096 121824 2112 121888
rect 2176 121824 2192 121888
rect 2256 121824 2264 121888
rect 1944 120800 2264 121824
rect 1944 120736 1952 120800
rect 2016 120736 2032 120800
rect 2096 120736 2112 120800
rect 2176 120736 2192 120800
rect 2256 120736 2264 120800
rect 1944 119712 2264 120736
rect 1944 119648 1952 119712
rect 2016 119648 2032 119712
rect 2096 119648 2112 119712
rect 2176 119648 2192 119712
rect 2256 119648 2264 119712
rect 1944 118624 2264 119648
rect 1944 118560 1952 118624
rect 2016 118560 2032 118624
rect 2096 118560 2112 118624
rect 2176 118560 2192 118624
rect 2256 118560 2264 118624
rect 1944 117536 2264 118560
rect 1944 117472 1952 117536
rect 2016 117472 2032 117536
rect 2096 117472 2112 117536
rect 2176 117472 2192 117536
rect 2256 117472 2264 117536
rect 1944 116448 2264 117472
rect 1944 116384 1952 116448
rect 2016 116384 2032 116448
rect 2096 116384 2112 116448
rect 2176 116384 2192 116448
rect 2256 116384 2264 116448
rect 1944 115576 2264 116384
rect 1944 115360 1986 115576
rect 2222 115360 2264 115576
rect 1944 115296 1952 115360
rect 2016 115296 2032 115340
rect 2096 115296 2112 115340
rect 2176 115296 2192 115340
rect 2256 115296 2264 115360
rect 1944 114272 2264 115296
rect 1944 114208 1952 114272
rect 2016 114208 2032 114272
rect 2096 114208 2112 114272
rect 2176 114208 2192 114272
rect 2256 114208 2264 114272
rect 1944 113184 2264 114208
rect 1944 113120 1952 113184
rect 2016 113120 2032 113184
rect 2096 113120 2112 113184
rect 2176 113120 2192 113184
rect 2256 113120 2264 113184
rect 1944 112096 2264 113120
rect 1944 112032 1952 112096
rect 2016 112032 2032 112096
rect 2096 112032 2112 112096
rect 2176 112032 2192 112096
rect 2256 112032 2264 112096
rect 1944 111008 2264 112032
rect 1944 110944 1952 111008
rect 2016 110944 2032 111008
rect 2096 110944 2112 111008
rect 2176 110944 2192 111008
rect 2256 110944 2264 111008
rect 1944 109920 2264 110944
rect 1944 109856 1952 109920
rect 2016 109856 2032 109920
rect 2096 109856 2112 109920
rect 2176 109856 2192 109920
rect 2256 109856 2264 109920
rect 1944 108832 2264 109856
rect 1944 108768 1952 108832
rect 2016 108768 2032 108832
rect 2096 108768 2112 108832
rect 2176 108768 2192 108832
rect 2256 108768 2264 108832
rect 1944 107744 2264 108768
rect 1944 107680 1952 107744
rect 2016 107680 2032 107744
rect 2096 107680 2112 107744
rect 2176 107680 2192 107744
rect 2256 107680 2264 107744
rect 1944 106656 2264 107680
rect 1944 106592 1952 106656
rect 2016 106592 2032 106656
rect 2096 106592 2112 106656
rect 2176 106592 2192 106656
rect 2256 106592 2264 106656
rect 1944 105576 2264 106592
rect 1944 105568 1986 105576
rect 2222 105568 2264 105576
rect 1944 105504 1952 105568
rect 2256 105504 2264 105568
rect 1944 105340 1986 105504
rect 2222 105340 2264 105504
rect 1944 104480 2264 105340
rect 1944 104416 1952 104480
rect 2016 104416 2032 104480
rect 2096 104416 2112 104480
rect 2176 104416 2192 104480
rect 2256 104416 2264 104480
rect 1944 103392 2264 104416
rect 1944 103328 1952 103392
rect 2016 103328 2032 103392
rect 2096 103328 2112 103392
rect 2176 103328 2192 103392
rect 2256 103328 2264 103392
rect 1944 102304 2264 103328
rect 1944 102240 1952 102304
rect 2016 102240 2032 102304
rect 2096 102240 2112 102304
rect 2176 102240 2192 102304
rect 2256 102240 2264 102304
rect 1944 101216 2264 102240
rect 1944 101152 1952 101216
rect 2016 101152 2032 101216
rect 2096 101152 2112 101216
rect 2176 101152 2192 101216
rect 2256 101152 2264 101216
rect 1944 100128 2264 101152
rect 1944 100064 1952 100128
rect 2016 100064 2032 100128
rect 2096 100064 2112 100128
rect 2176 100064 2192 100128
rect 2256 100064 2264 100128
rect 1944 99040 2264 100064
rect 1944 98976 1952 99040
rect 2016 98976 2032 99040
rect 2096 98976 2112 99040
rect 2176 98976 2192 99040
rect 2256 98976 2264 99040
rect 1944 97952 2264 98976
rect 1944 97888 1952 97952
rect 2016 97888 2032 97952
rect 2096 97888 2112 97952
rect 2176 97888 2192 97952
rect 2256 97888 2264 97952
rect 1944 96864 2264 97888
rect 1944 96800 1952 96864
rect 2016 96800 2032 96864
rect 2096 96800 2112 96864
rect 2176 96800 2192 96864
rect 2256 96800 2264 96864
rect 1944 95776 2264 96800
rect 1944 95712 1952 95776
rect 2016 95712 2032 95776
rect 2096 95712 2112 95776
rect 2176 95712 2192 95776
rect 2256 95712 2264 95776
rect 1944 95576 2264 95712
rect 1944 95340 1986 95576
rect 2222 95340 2264 95576
rect 1944 94688 2264 95340
rect 1944 94624 1952 94688
rect 2016 94624 2032 94688
rect 2096 94624 2112 94688
rect 2176 94624 2192 94688
rect 2256 94624 2264 94688
rect 1944 93600 2264 94624
rect 1944 93536 1952 93600
rect 2016 93536 2032 93600
rect 2096 93536 2112 93600
rect 2176 93536 2192 93600
rect 2256 93536 2264 93600
rect 1944 92512 2264 93536
rect 1944 92448 1952 92512
rect 2016 92448 2032 92512
rect 2096 92448 2112 92512
rect 2176 92448 2192 92512
rect 2256 92448 2264 92512
rect 1944 91424 2264 92448
rect 1944 91360 1952 91424
rect 2016 91360 2032 91424
rect 2096 91360 2112 91424
rect 2176 91360 2192 91424
rect 2256 91360 2264 91424
rect 1944 90336 2264 91360
rect 1944 90272 1952 90336
rect 2016 90272 2032 90336
rect 2096 90272 2112 90336
rect 2176 90272 2192 90336
rect 2256 90272 2264 90336
rect 1944 89248 2264 90272
rect 1944 89184 1952 89248
rect 2016 89184 2032 89248
rect 2096 89184 2112 89248
rect 2176 89184 2192 89248
rect 2256 89184 2264 89248
rect 1944 88160 2264 89184
rect 1944 88096 1952 88160
rect 2016 88096 2032 88160
rect 2096 88096 2112 88160
rect 2176 88096 2192 88160
rect 2256 88096 2264 88160
rect 1944 87072 2264 88096
rect 1944 87008 1952 87072
rect 2016 87008 2032 87072
rect 2096 87008 2112 87072
rect 2176 87008 2192 87072
rect 2256 87008 2264 87072
rect 1944 85984 2264 87008
rect 1944 85920 1952 85984
rect 2016 85920 2032 85984
rect 2096 85920 2112 85984
rect 2176 85920 2192 85984
rect 2256 85920 2264 85984
rect 1944 85576 2264 85920
rect 1944 85340 1986 85576
rect 2222 85340 2264 85576
rect 1944 84896 2264 85340
rect 1944 84832 1952 84896
rect 2016 84832 2032 84896
rect 2096 84832 2112 84896
rect 2176 84832 2192 84896
rect 2256 84832 2264 84896
rect 1944 83808 2264 84832
rect 1944 83744 1952 83808
rect 2016 83744 2032 83808
rect 2096 83744 2112 83808
rect 2176 83744 2192 83808
rect 2256 83744 2264 83808
rect 1944 82720 2264 83744
rect 1944 82656 1952 82720
rect 2016 82656 2032 82720
rect 2096 82656 2112 82720
rect 2176 82656 2192 82720
rect 2256 82656 2264 82720
rect 1944 81632 2264 82656
rect 1944 81568 1952 81632
rect 2016 81568 2032 81632
rect 2096 81568 2112 81632
rect 2176 81568 2192 81632
rect 2256 81568 2264 81632
rect 1944 80544 2264 81568
rect 1944 80480 1952 80544
rect 2016 80480 2032 80544
rect 2096 80480 2112 80544
rect 2176 80480 2192 80544
rect 2256 80480 2264 80544
rect 1944 79456 2264 80480
rect 1944 79392 1952 79456
rect 2016 79392 2032 79456
rect 2096 79392 2112 79456
rect 2176 79392 2192 79456
rect 2256 79392 2264 79456
rect 1944 78368 2264 79392
rect 1944 78304 1952 78368
rect 2016 78304 2032 78368
rect 2096 78304 2112 78368
rect 2176 78304 2192 78368
rect 2256 78304 2264 78368
rect 1944 77280 2264 78304
rect 1944 77216 1952 77280
rect 2016 77216 2032 77280
rect 2096 77216 2112 77280
rect 2176 77216 2192 77280
rect 2256 77216 2264 77280
rect 1944 76192 2264 77216
rect 1944 76128 1952 76192
rect 2016 76128 2032 76192
rect 2096 76128 2112 76192
rect 2176 76128 2192 76192
rect 2256 76128 2264 76192
rect 1944 75576 2264 76128
rect 1944 75340 1986 75576
rect 2222 75340 2264 75576
rect 1944 75104 2264 75340
rect 1944 75040 1952 75104
rect 2016 75040 2032 75104
rect 2096 75040 2112 75104
rect 2176 75040 2192 75104
rect 2256 75040 2264 75104
rect 1944 74016 2264 75040
rect 1944 73952 1952 74016
rect 2016 73952 2032 74016
rect 2096 73952 2112 74016
rect 2176 73952 2192 74016
rect 2256 73952 2264 74016
rect 1944 72928 2264 73952
rect 1944 72864 1952 72928
rect 2016 72864 2032 72928
rect 2096 72864 2112 72928
rect 2176 72864 2192 72928
rect 2256 72864 2264 72928
rect 1944 71840 2264 72864
rect 1944 71776 1952 71840
rect 2016 71776 2032 71840
rect 2096 71776 2112 71840
rect 2176 71776 2192 71840
rect 2256 71776 2264 71840
rect 1944 70752 2264 71776
rect 1944 70688 1952 70752
rect 2016 70688 2032 70752
rect 2096 70688 2112 70752
rect 2176 70688 2192 70752
rect 2256 70688 2264 70752
rect 1944 69664 2264 70688
rect 1944 69600 1952 69664
rect 2016 69600 2032 69664
rect 2096 69600 2112 69664
rect 2176 69600 2192 69664
rect 2256 69600 2264 69664
rect 1944 68576 2264 69600
rect 1944 68512 1952 68576
rect 2016 68512 2032 68576
rect 2096 68512 2112 68576
rect 2176 68512 2192 68576
rect 2256 68512 2264 68576
rect 1944 67488 2264 68512
rect 1944 67424 1952 67488
rect 2016 67424 2032 67488
rect 2096 67424 2112 67488
rect 2176 67424 2192 67488
rect 2256 67424 2264 67488
rect 1944 66400 2264 67424
rect 1944 66336 1952 66400
rect 2016 66336 2032 66400
rect 2096 66336 2112 66400
rect 2176 66336 2192 66400
rect 2256 66336 2264 66400
rect 1944 65576 2264 66336
rect 1944 65340 1986 65576
rect 2222 65340 2264 65576
rect 1944 65312 2264 65340
rect 1944 65248 1952 65312
rect 2016 65248 2032 65312
rect 2096 65248 2112 65312
rect 2176 65248 2192 65312
rect 2256 65248 2264 65312
rect 1944 64224 2264 65248
rect 1944 64160 1952 64224
rect 2016 64160 2032 64224
rect 2096 64160 2112 64224
rect 2176 64160 2192 64224
rect 2256 64160 2264 64224
rect 1944 63136 2264 64160
rect 1944 63072 1952 63136
rect 2016 63072 2032 63136
rect 2096 63072 2112 63136
rect 2176 63072 2192 63136
rect 2256 63072 2264 63136
rect 1944 62048 2264 63072
rect 1944 61984 1952 62048
rect 2016 61984 2032 62048
rect 2096 61984 2112 62048
rect 2176 61984 2192 62048
rect 2256 61984 2264 62048
rect 1944 60960 2264 61984
rect 1944 60896 1952 60960
rect 2016 60896 2032 60960
rect 2096 60896 2112 60960
rect 2176 60896 2192 60960
rect 2256 60896 2264 60960
rect 1944 59872 2264 60896
rect 1944 59808 1952 59872
rect 2016 59808 2032 59872
rect 2096 59808 2112 59872
rect 2176 59808 2192 59872
rect 2256 59808 2264 59872
rect 1944 58784 2264 59808
rect 1944 58720 1952 58784
rect 2016 58720 2032 58784
rect 2096 58720 2112 58784
rect 2176 58720 2192 58784
rect 2256 58720 2264 58784
rect 1944 57696 2264 58720
rect 1944 57632 1952 57696
rect 2016 57632 2032 57696
rect 2096 57632 2112 57696
rect 2176 57632 2192 57696
rect 2256 57632 2264 57696
rect 1944 56608 2264 57632
rect 1944 56544 1952 56608
rect 2016 56544 2032 56608
rect 2096 56544 2112 56608
rect 2176 56544 2192 56608
rect 2256 56544 2264 56608
rect 1944 55576 2264 56544
rect 1944 55520 1986 55576
rect 2222 55520 2264 55576
rect 1944 55456 1952 55520
rect 2256 55456 2264 55520
rect 1944 55340 1986 55456
rect 2222 55340 2264 55456
rect 1944 54432 2264 55340
rect 1944 54368 1952 54432
rect 2016 54368 2032 54432
rect 2096 54368 2112 54432
rect 2176 54368 2192 54432
rect 2256 54368 2264 54432
rect 1944 53344 2264 54368
rect 1944 53280 1952 53344
rect 2016 53280 2032 53344
rect 2096 53280 2112 53344
rect 2176 53280 2192 53344
rect 2256 53280 2264 53344
rect 1944 52256 2264 53280
rect 1944 52192 1952 52256
rect 2016 52192 2032 52256
rect 2096 52192 2112 52256
rect 2176 52192 2192 52256
rect 2256 52192 2264 52256
rect 1944 51168 2264 52192
rect 1944 51104 1952 51168
rect 2016 51104 2032 51168
rect 2096 51104 2112 51168
rect 2176 51104 2192 51168
rect 2256 51104 2264 51168
rect 1944 50080 2264 51104
rect 1944 50016 1952 50080
rect 2016 50016 2032 50080
rect 2096 50016 2112 50080
rect 2176 50016 2192 50080
rect 2256 50016 2264 50080
rect 1944 48992 2264 50016
rect 1944 48928 1952 48992
rect 2016 48928 2032 48992
rect 2096 48928 2112 48992
rect 2176 48928 2192 48992
rect 2256 48928 2264 48992
rect 1944 47904 2264 48928
rect 1944 47840 1952 47904
rect 2016 47840 2032 47904
rect 2096 47840 2112 47904
rect 2176 47840 2192 47904
rect 2256 47840 2264 47904
rect 1944 46816 2264 47840
rect 1944 46752 1952 46816
rect 2016 46752 2032 46816
rect 2096 46752 2112 46816
rect 2176 46752 2192 46816
rect 2256 46752 2264 46816
rect 1944 45728 2264 46752
rect 1944 45664 1952 45728
rect 2016 45664 2032 45728
rect 2096 45664 2112 45728
rect 2176 45664 2192 45728
rect 2256 45664 2264 45728
rect 1944 45576 2264 45664
rect 1944 45340 1986 45576
rect 2222 45340 2264 45576
rect 1944 44640 2264 45340
rect 1944 44576 1952 44640
rect 2016 44576 2032 44640
rect 2096 44576 2112 44640
rect 2176 44576 2192 44640
rect 2256 44576 2264 44640
rect 1944 43552 2264 44576
rect 1944 43488 1952 43552
rect 2016 43488 2032 43552
rect 2096 43488 2112 43552
rect 2176 43488 2192 43552
rect 2256 43488 2264 43552
rect 1944 42464 2264 43488
rect 1944 42400 1952 42464
rect 2016 42400 2032 42464
rect 2096 42400 2112 42464
rect 2176 42400 2192 42464
rect 2256 42400 2264 42464
rect 1944 41376 2264 42400
rect 1944 41312 1952 41376
rect 2016 41312 2032 41376
rect 2096 41312 2112 41376
rect 2176 41312 2192 41376
rect 2256 41312 2264 41376
rect 1944 40288 2264 41312
rect 1944 40224 1952 40288
rect 2016 40224 2032 40288
rect 2096 40224 2112 40288
rect 2176 40224 2192 40288
rect 2256 40224 2264 40288
rect 1944 39200 2264 40224
rect 1944 39136 1952 39200
rect 2016 39136 2032 39200
rect 2096 39136 2112 39200
rect 2176 39136 2192 39200
rect 2256 39136 2264 39200
rect 1944 38112 2264 39136
rect 1944 38048 1952 38112
rect 2016 38048 2032 38112
rect 2096 38048 2112 38112
rect 2176 38048 2192 38112
rect 2256 38048 2264 38112
rect 1944 37024 2264 38048
rect 1944 36960 1952 37024
rect 2016 36960 2032 37024
rect 2096 36960 2112 37024
rect 2176 36960 2192 37024
rect 2256 36960 2264 37024
rect 1944 35936 2264 36960
rect 1944 35872 1952 35936
rect 2016 35872 2032 35936
rect 2096 35872 2112 35936
rect 2176 35872 2192 35936
rect 2256 35872 2264 35936
rect 1944 35576 2264 35872
rect 1944 35340 1986 35576
rect 2222 35340 2264 35576
rect 1944 34848 2264 35340
rect 1944 34784 1952 34848
rect 2016 34784 2032 34848
rect 2096 34784 2112 34848
rect 2176 34784 2192 34848
rect 2256 34784 2264 34848
rect 1944 33760 2264 34784
rect 1944 33696 1952 33760
rect 2016 33696 2032 33760
rect 2096 33696 2112 33760
rect 2176 33696 2192 33760
rect 2256 33696 2264 33760
rect 1944 32672 2264 33696
rect 1944 32608 1952 32672
rect 2016 32608 2032 32672
rect 2096 32608 2112 32672
rect 2176 32608 2192 32672
rect 2256 32608 2264 32672
rect 1944 31584 2264 32608
rect 1944 31520 1952 31584
rect 2016 31520 2032 31584
rect 2096 31520 2112 31584
rect 2176 31520 2192 31584
rect 2256 31520 2264 31584
rect 1944 30496 2264 31520
rect 1944 30432 1952 30496
rect 2016 30432 2032 30496
rect 2096 30432 2112 30496
rect 2176 30432 2192 30496
rect 2256 30432 2264 30496
rect 1944 29408 2264 30432
rect 1944 29344 1952 29408
rect 2016 29344 2032 29408
rect 2096 29344 2112 29408
rect 2176 29344 2192 29408
rect 2256 29344 2264 29408
rect 1944 28320 2264 29344
rect 1944 28256 1952 28320
rect 2016 28256 2032 28320
rect 2096 28256 2112 28320
rect 2176 28256 2192 28320
rect 2256 28256 2264 28320
rect 1944 27232 2264 28256
rect 1944 27168 1952 27232
rect 2016 27168 2032 27232
rect 2096 27168 2112 27232
rect 2176 27168 2192 27232
rect 2256 27168 2264 27232
rect 1944 26144 2264 27168
rect 1944 26080 1952 26144
rect 2016 26080 2032 26144
rect 2096 26080 2112 26144
rect 2176 26080 2192 26144
rect 2256 26080 2264 26144
rect 1944 25576 2264 26080
rect 1944 25340 1986 25576
rect 2222 25340 2264 25576
rect 1944 25056 2264 25340
rect 1944 24992 1952 25056
rect 2016 24992 2032 25056
rect 2096 24992 2112 25056
rect 2176 24992 2192 25056
rect 2256 24992 2264 25056
rect 1944 23968 2264 24992
rect 1944 23904 1952 23968
rect 2016 23904 2032 23968
rect 2096 23904 2112 23968
rect 2176 23904 2192 23968
rect 2256 23904 2264 23968
rect 1944 22880 2264 23904
rect 1944 22816 1952 22880
rect 2016 22816 2032 22880
rect 2096 22816 2112 22880
rect 2176 22816 2192 22880
rect 2256 22816 2264 22880
rect 1944 21792 2264 22816
rect 1944 21728 1952 21792
rect 2016 21728 2032 21792
rect 2096 21728 2112 21792
rect 2176 21728 2192 21792
rect 2256 21728 2264 21792
rect 1944 20704 2264 21728
rect 1944 20640 1952 20704
rect 2016 20640 2032 20704
rect 2096 20640 2112 20704
rect 2176 20640 2192 20704
rect 2256 20640 2264 20704
rect 1944 19616 2264 20640
rect 1944 19552 1952 19616
rect 2016 19552 2032 19616
rect 2096 19552 2112 19616
rect 2176 19552 2192 19616
rect 2256 19552 2264 19616
rect 1944 18528 2264 19552
rect 1944 18464 1952 18528
rect 2016 18464 2032 18528
rect 2096 18464 2112 18528
rect 2176 18464 2192 18528
rect 2256 18464 2264 18528
rect 1944 17440 2264 18464
rect 1944 17376 1952 17440
rect 2016 17376 2032 17440
rect 2096 17376 2112 17440
rect 2176 17376 2192 17440
rect 2256 17376 2264 17440
rect 1944 16352 2264 17376
rect 1944 16288 1952 16352
rect 2016 16288 2032 16352
rect 2096 16288 2112 16352
rect 2176 16288 2192 16352
rect 2256 16288 2264 16352
rect 1944 15576 2264 16288
rect 1944 15340 1986 15576
rect 2222 15340 2264 15576
rect 1944 15264 2264 15340
rect 1944 15200 1952 15264
rect 2016 15200 2032 15264
rect 2096 15200 2112 15264
rect 2176 15200 2192 15264
rect 2256 15200 2264 15264
rect 1944 14176 2264 15200
rect 1944 14112 1952 14176
rect 2016 14112 2032 14176
rect 2096 14112 2112 14176
rect 2176 14112 2192 14176
rect 2256 14112 2264 14176
rect 1944 13088 2264 14112
rect 1944 13024 1952 13088
rect 2016 13024 2032 13088
rect 2096 13024 2112 13088
rect 2176 13024 2192 13088
rect 2256 13024 2264 13088
rect 1944 12000 2264 13024
rect 1944 11936 1952 12000
rect 2016 11936 2032 12000
rect 2096 11936 2112 12000
rect 2176 11936 2192 12000
rect 2256 11936 2264 12000
rect 1944 10912 2264 11936
rect 1944 10848 1952 10912
rect 2016 10848 2032 10912
rect 2096 10848 2112 10912
rect 2176 10848 2192 10912
rect 2256 10848 2264 10912
rect 1944 9824 2264 10848
rect 1944 9760 1952 9824
rect 2016 9760 2032 9824
rect 2096 9760 2112 9824
rect 2176 9760 2192 9824
rect 2256 9760 2264 9824
rect 1944 8736 2264 9760
rect 1944 8672 1952 8736
rect 2016 8672 2032 8736
rect 2096 8672 2112 8736
rect 2176 8672 2192 8736
rect 2256 8672 2264 8736
rect 1944 7648 2264 8672
rect 1944 7584 1952 7648
rect 2016 7584 2032 7648
rect 2096 7584 2112 7648
rect 2176 7584 2192 7648
rect 2256 7584 2264 7648
rect 1944 6560 2264 7584
rect 1944 6496 1952 6560
rect 2016 6496 2032 6560
rect 2096 6496 2112 6560
rect 2176 6496 2192 6560
rect 2256 6496 2264 6560
rect 1944 5576 2264 6496
rect 1944 5472 1986 5576
rect 2222 5472 2264 5576
rect 1944 5408 1952 5472
rect 2256 5408 2264 5472
rect 1944 5340 1986 5408
rect 2222 5340 2264 5408
rect 1944 4384 2264 5340
rect 1944 4320 1952 4384
rect 2016 4320 2032 4384
rect 2096 4320 2112 4384
rect 2176 4320 2192 4384
rect 2256 4320 2264 4384
rect 1944 3296 2264 4320
rect 1944 3232 1952 3296
rect 2016 3232 2032 3296
rect 2096 3232 2112 3296
rect 2176 3232 2192 3296
rect 2256 3232 2264 3296
rect 1944 2208 2264 3232
rect 1944 2144 1952 2208
rect 2016 2144 2032 2208
rect 2096 2144 2112 2208
rect 2176 2144 2192 2208
rect 2256 2144 2264 2208
rect 1944 2128 2264 2144
rect 3944 188800 4264 189360
rect 85944 189344 86264 189360
rect 85944 189280 85952 189344
rect 86016 189280 86032 189344
rect 86096 189280 86112 189344
rect 86176 189280 86192 189344
rect 86256 189280 86264 189344
rect 75131 189140 75197 189141
rect 75131 189076 75132 189140
rect 75196 189076 75197 189140
rect 75131 189075 75197 189076
rect 3944 188736 3952 188800
rect 4016 188736 4032 188800
rect 4096 188736 4112 188800
rect 4176 188736 4192 188800
rect 4256 188736 4264 188800
rect 3944 187712 4264 188736
rect 3944 187648 3952 187712
rect 4016 187648 4032 187712
rect 4096 187648 4112 187712
rect 4176 187648 4192 187712
rect 4256 187648 4264 187712
rect 3944 186624 4264 187648
rect 75134 187370 75194 189075
rect 74608 187310 75194 187370
rect 85944 188256 86264 189280
rect 85944 188192 85952 188256
rect 86016 188192 86032 188256
rect 86096 188192 86112 188256
rect 86176 188192 86192 188256
rect 86256 188192 86264 188256
rect 79366 187205 79603 187265
rect 79366 187101 79426 187205
rect 85944 187168 86264 188192
rect 85944 187104 85952 187168
rect 86016 187104 86032 187168
rect 86096 187104 86112 187168
rect 86176 187104 86192 187168
rect 86256 187104 86264 187168
rect 79363 187100 79429 187101
rect 79363 187036 79364 187100
rect 79428 187036 79429 187100
rect 79363 187035 79429 187036
rect 3944 186560 3952 186624
rect 4016 186560 4032 186624
rect 4096 186560 4112 186624
rect 4176 186560 4192 186624
rect 4256 186560 4264 186624
rect 3944 185536 4264 186560
rect 3944 185472 3952 185536
rect 4016 185472 4032 185536
rect 4096 185472 4112 185536
rect 4176 185472 4192 185536
rect 4256 185472 4264 185536
rect 3944 184448 4264 185472
rect 3944 184384 3952 184448
rect 4016 184384 4032 184448
rect 4096 184384 4112 184448
rect 4176 184384 4192 184448
rect 4256 184384 4264 184448
rect 3944 183360 4264 184384
rect 3944 183296 3952 183360
rect 4016 183296 4032 183360
rect 4096 183296 4112 183360
rect 4176 183296 4192 183360
rect 4256 183296 4264 183360
rect 3944 182272 4264 183296
rect 3944 182208 3952 182272
rect 4016 182208 4032 182272
rect 4096 182208 4112 182272
rect 4176 182208 4192 182272
rect 4256 182208 4264 182272
rect 3944 181184 4264 182208
rect 3944 181120 3952 181184
rect 4016 181120 4032 181184
rect 4096 181120 4112 181184
rect 4176 181120 4192 181184
rect 4256 181120 4264 181184
rect 3944 180576 4264 181120
rect 85944 186080 86264 187104
rect 85944 186016 85952 186080
rect 86016 186016 86032 186080
rect 86096 186016 86112 186080
rect 86176 186016 86192 186080
rect 86256 186016 86264 186080
rect 85944 185576 86264 186016
rect 85944 185340 85986 185576
rect 86222 185340 86264 185576
rect 85944 184992 86264 185340
rect 85944 184928 85952 184992
rect 86016 184928 86032 184992
rect 86096 184928 86112 184992
rect 86176 184928 86192 184992
rect 86256 184928 86264 184992
rect 85944 183904 86264 184928
rect 87944 188800 88264 189360
rect 87944 188736 87952 188800
rect 88016 188736 88032 188800
rect 88096 188736 88112 188800
rect 88176 188736 88192 188800
rect 88256 188736 88264 188800
rect 87944 187712 88264 188736
rect 87944 187648 87952 187712
rect 88016 187648 88032 187712
rect 88096 187648 88112 187712
rect 88176 187648 88192 187712
rect 88256 187648 88264 187712
rect 87944 186624 88264 187648
rect 87944 186560 87952 186624
rect 88016 186560 88032 186624
rect 88096 186560 88112 186624
rect 88176 186560 88192 186624
rect 88256 186560 88264 186624
rect 87944 185536 88264 186560
rect 88747 186556 88813 186557
rect 88747 186492 88748 186556
rect 88812 186492 88813 186556
rect 88747 186491 88813 186492
rect 87944 185472 87952 185536
rect 88016 185472 88032 185536
rect 88096 185472 88112 185536
rect 88176 185472 88192 185536
rect 88256 185472 88264 185536
rect 87944 184448 88264 185472
rect 88379 185332 88445 185333
rect 88379 185268 88380 185332
rect 88444 185268 88445 185332
rect 88379 185267 88445 185268
rect 87944 184384 87952 184448
rect 88016 184384 88032 184448
rect 88096 184384 88112 184448
rect 88176 184384 88192 184448
rect 88256 184384 88264 184448
rect 87459 184108 87525 184109
rect 87459 184044 87460 184108
rect 87524 184044 87525 184108
rect 87459 184043 87525 184044
rect 85944 183840 85952 183904
rect 86016 183840 86032 183904
rect 86096 183840 86112 183904
rect 86176 183840 86192 183904
rect 86256 183840 86264 183904
rect 85944 182816 86264 183840
rect 85944 182752 85952 182816
rect 86016 182752 86032 182816
rect 86096 182752 86112 182816
rect 86176 182752 86192 182816
rect 86256 182752 86264 182816
rect 85944 181728 86264 182752
rect 87091 182612 87157 182613
rect 87091 182548 87092 182612
rect 87156 182548 87157 182612
rect 87091 182547 87157 182548
rect 85944 181664 85952 181728
rect 86016 181664 86032 181728
rect 86096 181664 86112 181728
rect 86176 181664 86192 181728
rect 86256 181664 86264 181728
rect 85944 180640 86264 181664
rect 3944 180340 3986 180576
rect 4222 180340 4264 180576
rect 3944 180096 4264 180340
rect 82938 180576 83262 180618
rect 82938 180340 82982 180576
rect 83218 180340 83262 180576
rect 82938 180298 83262 180340
rect 85944 180576 85952 180640
rect 86016 180576 86032 180640
rect 86096 180576 86112 180640
rect 86176 180576 86192 180640
rect 86256 180576 86264 180640
rect 3944 180032 3952 180096
rect 4016 180032 4032 180096
rect 4096 180032 4112 180096
rect 4176 180032 4192 180096
rect 4256 180032 4264 180096
rect 3944 179008 4264 180032
rect 3944 178944 3952 179008
rect 4016 178944 4032 179008
rect 4096 178944 4112 179008
rect 4176 178944 4192 179008
rect 4256 178944 4264 179008
rect 3944 177920 4264 178944
rect 3944 177856 3952 177920
rect 4016 177856 4032 177920
rect 4096 177856 4112 177920
rect 4176 177856 4192 177920
rect 4256 177856 4264 177920
rect 3944 176832 4264 177856
rect 85944 179552 86264 180576
rect 85944 179488 85952 179552
rect 86016 179488 86032 179552
rect 86096 179488 86112 179552
rect 86176 179488 86192 179552
rect 86256 179488 86264 179552
rect 85944 178464 86264 179488
rect 85944 178400 85952 178464
rect 86016 178400 86032 178464
rect 86096 178400 86112 178464
rect 86176 178400 86192 178464
rect 86256 178400 86264 178464
rect 85944 177376 86264 178400
rect 85944 177312 85952 177376
rect 86016 177312 86032 177376
rect 86096 177312 86112 177376
rect 86176 177312 86192 177376
rect 86256 177312 86264 177376
rect 83411 177036 83477 177037
rect 83411 176972 83412 177036
rect 83476 176972 83477 177036
rect 83411 176971 83477 176972
rect 3944 176768 3952 176832
rect 4016 176768 4032 176832
rect 4096 176768 4112 176832
rect 4176 176768 4192 176832
rect 4256 176768 4264 176832
rect 3944 175744 4264 176768
rect 3944 175680 3952 175744
rect 4016 175680 4032 175744
rect 4096 175680 4112 175744
rect 4176 175680 4192 175744
rect 4256 175680 4264 175744
rect 3944 174656 4264 175680
rect 82494 175576 82814 175618
rect 82494 175340 82536 175576
rect 82772 175340 82814 175576
rect 82494 175298 82814 175340
rect 3944 174592 3952 174656
rect 4016 174592 4032 174656
rect 4096 174592 4112 174656
rect 4176 174592 4192 174656
rect 4256 174592 4264 174656
rect 3944 173568 4264 174592
rect 3944 173504 3952 173568
rect 4016 173504 4032 173568
rect 4096 173504 4112 173568
rect 4176 173504 4192 173568
rect 4256 173504 4264 173568
rect 3944 172480 4264 173504
rect 3944 172416 3952 172480
rect 4016 172416 4032 172480
rect 4096 172416 4112 172480
rect 4176 172416 4192 172480
rect 4256 172416 4264 172480
rect 3944 171392 4264 172416
rect 3944 171328 3952 171392
rect 4016 171328 4032 171392
rect 4096 171328 4112 171392
rect 4176 171328 4192 171392
rect 4256 171328 4264 171392
rect 3944 170576 4264 171328
rect 3944 170340 3986 170576
rect 4222 170340 4264 170576
rect 3944 170304 4264 170340
rect 3944 170240 3952 170304
rect 4016 170240 4032 170304
rect 4096 170240 4112 170304
rect 4176 170240 4192 170304
rect 4256 170240 4264 170304
rect 82938 170576 83262 170618
rect 82938 170340 82982 170576
rect 83218 170340 83262 170576
rect 82938 170298 83262 170340
rect 3944 169216 4264 170240
rect 3944 169152 3952 169216
rect 4016 169152 4032 169216
rect 4096 169152 4112 169216
rect 4176 169152 4192 169216
rect 4256 169152 4264 169216
rect 3944 168128 4264 169152
rect 3944 168064 3952 168128
rect 4016 168064 4032 168128
rect 4096 168064 4112 168128
rect 4176 168064 4192 168128
rect 4256 168064 4264 168128
rect 3944 167040 4264 168064
rect 3944 166976 3952 167040
rect 4016 166976 4032 167040
rect 4096 166976 4112 167040
rect 4176 166976 4192 167040
rect 4256 166976 4264 167040
rect 3944 165952 4264 166976
rect 3944 165888 3952 165952
rect 4016 165888 4032 165952
rect 4096 165888 4112 165952
rect 4176 165888 4192 165952
rect 4256 165888 4264 165952
rect 3944 164864 4264 165888
rect 82494 165576 82814 165618
rect 82494 165340 82536 165576
rect 82772 165340 82814 165576
rect 82494 165298 82814 165340
rect 3944 164800 3952 164864
rect 4016 164800 4032 164864
rect 4096 164800 4112 164864
rect 4176 164800 4192 164864
rect 4256 164800 4264 164864
rect 3944 163776 4264 164800
rect 3944 163712 3952 163776
rect 4016 163712 4032 163776
rect 4096 163712 4112 163776
rect 4176 163712 4192 163776
rect 4256 163712 4264 163776
rect 3944 162688 4264 163712
rect 3944 162624 3952 162688
rect 4016 162624 4032 162688
rect 4096 162624 4112 162688
rect 4176 162624 4192 162688
rect 4256 162624 4264 162688
rect 3944 161600 4264 162624
rect 3944 161536 3952 161600
rect 4016 161536 4032 161600
rect 4096 161536 4112 161600
rect 4176 161536 4192 161600
rect 4256 161536 4264 161600
rect 3944 160576 4264 161536
rect 3944 160512 3986 160576
rect 4222 160512 4264 160576
rect 3944 160448 3952 160512
rect 4256 160448 4264 160512
rect 3944 160340 3986 160448
rect 4222 160340 4264 160448
rect 3944 159424 4264 160340
rect 82938 160576 83262 160618
rect 82938 160340 82982 160576
rect 83218 160340 83262 160576
rect 82938 160298 83262 160340
rect 3944 159360 3952 159424
rect 4016 159360 4032 159424
rect 4096 159360 4112 159424
rect 4176 159360 4192 159424
rect 4256 159360 4264 159424
rect 3944 158336 4264 159360
rect 3944 158272 3952 158336
rect 4016 158272 4032 158336
rect 4096 158272 4112 158336
rect 4176 158272 4192 158336
rect 4256 158272 4264 158336
rect 3944 157248 4264 158272
rect 3944 157184 3952 157248
rect 4016 157184 4032 157248
rect 4096 157184 4112 157248
rect 4176 157184 4192 157248
rect 4256 157184 4264 157248
rect 3944 156160 4264 157184
rect 3944 156096 3952 156160
rect 4016 156096 4032 156160
rect 4096 156096 4112 156160
rect 4176 156096 4192 156160
rect 4256 156096 4264 156160
rect 3944 155072 4264 156096
rect 82494 155576 82814 155618
rect 82494 155340 82536 155576
rect 82772 155340 82814 155576
rect 82494 155298 82814 155340
rect 3944 155008 3952 155072
rect 4016 155008 4032 155072
rect 4096 155008 4112 155072
rect 4176 155008 4192 155072
rect 4256 155008 4264 155072
rect 3944 153984 4264 155008
rect 3944 153920 3952 153984
rect 4016 153920 4032 153984
rect 4096 153920 4112 153984
rect 4176 153920 4192 153984
rect 4256 153920 4264 153984
rect 3944 152896 4264 153920
rect 3944 152832 3952 152896
rect 4016 152832 4032 152896
rect 4096 152832 4112 152896
rect 4176 152832 4192 152896
rect 4256 152832 4264 152896
rect 3944 151808 4264 152832
rect 3944 151744 3952 151808
rect 4016 151744 4032 151808
rect 4096 151744 4112 151808
rect 4176 151744 4192 151808
rect 4256 151744 4264 151808
rect 3944 150720 4264 151744
rect 3944 150656 3952 150720
rect 4016 150656 4032 150720
rect 4096 150656 4112 150720
rect 4176 150656 4192 150720
rect 4256 150656 4264 150720
rect 3944 150576 4264 150656
rect 3944 150340 3986 150576
rect 4222 150340 4264 150576
rect 3944 149632 4264 150340
rect 82938 150576 83262 150618
rect 82938 150340 82982 150576
rect 83218 150340 83262 150576
rect 82938 150298 83262 150340
rect 3944 149568 3952 149632
rect 4016 149568 4032 149632
rect 4096 149568 4112 149632
rect 4176 149568 4192 149632
rect 4256 149568 4264 149632
rect 3944 148544 4264 149568
rect 3944 148480 3952 148544
rect 4016 148480 4032 148544
rect 4096 148480 4112 148544
rect 4176 148480 4192 148544
rect 4256 148480 4264 148544
rect 3944 147456 4264 148480
rect 3944 147392 3952 147456
rect 4016 147392 4032 147456
rect 4096 147392 4112 147456
rect 4176 147392 4192 147456
rect 4256 147392 4264 147456
rect 3944 146368 4264 147392
rect 3944 146304 3952 146368
rect 4016 146304 4032 146368
rect 4096 146304 4112 146368
rect 4176 146304 4192 146368
rect 4256 146304 4264 146368
rect 3944 145280 4264 146304
rect 82494 145576 82814 145618
rect 82494 145340 82536 145576
rect 82772 145340 82814 145576
rect 82494 145298 82814 145340
rect 3944 145216 3952 145280
rect 4016 145216 4032 145280
rect 4096 145216 4112 145280
rect 4176 145216 4192 145280
rect 4256 145216 4264 145280
rect 3944 144192 4264 145216
rect 3944 144128 3952 144192
rect 4016 144128 4032 144192
rect 4096 144128 4112 144192
rect 4176 144128 4192 144192
rect 4256 144128 4264 144192
rect 3944 143104 4264 144128
rect 3944 143040 3952 143104
rect 4016 143040 4032 143104
rect 4096 143040 4112 143104
rect 4176 143040 4192 143104
rect 4256 143040 4264 143104
rect 3944 142016 4264 143040
rect 3944 141952 3952 142016
rect 4016 141952 4032 142016
rect 4096 141952 4112 142016
rect 4176 141952 4192 142016
rect 4256 141952 4264 142016
rect 3944 140928 4264 141952
rect 3944 140864 3952 140928
rect 4016 140864 4032 140928
rect 4096 140864 4112 140928
rect 4176 140864 4192 140928
rect 4256 140864 4264 140928
rect 3944 140576 4264 140864
rect 3944 140340 3986 140576
rect 4222 140340 4264 140576
rect 3944 139840 4264 140340
rect 82938 140576 83262 140618
rect 82938 140340 82982 140576
rect 83218 140340 83262 140576
rect 82938 140298 83262 140340
rect 3944 139776 3952 139840
rect 4016 139776 4032 139840
rect 4096 139776 4112 139840
rect 4176 139776 4192 139840
rect 4256 139776 4264 139840
rect 3944 138752 4264 139776
rect 3944 138688 3952 138752
rect 4016 138688 4032 138752
rect 4096 138688 4112 138752
rect 4176 138688 4192 138752
rect 4256 138688 4264 138752
rect 3944 137664 4264 138688
rect 3944 137600 3952 137664
rect 4016 137600 4032 137664
rect 4096 137600 4112 137664
rect 4176 137600 4192 137664
rect 4256 137600 4264 137664
rect 3944 136576 4264 137600
rect 3944 136512 3952 136576
rect 4016 136512 4032 136576
rect 4096 136512 4112 136576
rect 4176 136512 4192 136576
rect 4256 136512 4264 136576
rect 3944 135488 4264 136512
rect 3944 135424 3952 135488
rect 4016 135424 4032 135488
rect 4096 135424 4112 135488
rect 4176 135424 4192 135488
rect 4256 135424 4264 135488
rect 3944 134400 4264 135424
rect 82494 135576 82814 135618
rect 82494 135340 82536 135576
rect 82772 135340 82814 135576
rect 82494 135298 82814 135340
rect 3944 134336 3952 134400
rect 4016 134336 4032 134400
rect 4096 134336 4112 134400
rect 4176 134336 4192 134400
rect 4256 134336 4264 134400
rect 3944 133312 4264 134336
rect 3944 133248 3952 133312
rect 4016 133248 4032 133312
rect 4096 133248 4112 133312
rect 4176 133248 4192 133312
rect 4256 133248 4264 133312
rect 3944 132224 4264 133248
rect 83414 132429 83474 176971
rect 85944 176288 86264 177312
rect 85944 176224 85952 176288
rect 86016 176224 86032 176288
rect 86096 176224 86112 176288
rect 86176 176224 86192 176288
rect 86256 176224 86264 176288
rect 85944 175576 86264 176224
rect 83595 175404 83661 175405
rect 83595 175340 83596 175404
rect 83660 175340 83661 175404
rect 83595 175339 83661 175340
rect 85944 175340 85986 175576
rect 86222 175340 86264 175576
rect 83411 132428 83477 132429
rect 83411 132364 83412 132428
rect 83476 132364 83477 132428
rect 83411 132363 83477 132364
rect 83411 132292 83477 132293
rect 83411 132228 83412 132292
rect 83476 132228 83477 132292
rect 83411 132227 83477 132228
rect 3944 132160 3952 132224
rect 4016 132160 4032 132224
rect 4096 132160 4112 132224
rect 4176 132160 4192 132224
rect 4256 132160 4264 132224
rect 3944 131136 4264 132160
rect 3944 131072 3952 131136
rect 4016 131072 4032 131136
rect 4096 131072 4112 131136
rect 4176 131072 4192 131136
rect 4256 131072 4264 131136
rect 3944 130576 4264 131072
rect 3944 130340 3986 130576
rect 4222 130340 4264 130576
rect 3944 130048 4264 130340
rect 82938 130576 83262 130618
rect 82938 130340 82982 130576
rect 83218 130340 83262 130576
rect 82938 130298 83262 130340
rect 3944 129984 3952 130048
rect 4016 129984 4032 130048
rect 4096 129984 4112 130048
rect 4176 129984 4192 130048
rect 4256 129984 4264 130048
rect 3944 128960 4264 129984
rect 3944 128896 3952 128960
rect 4016 128896 4032 128960
rect 4096 128896 4112 128960
rect 4176 128896 4192 128960
rect 4256 128896 4264 128960
rect 3944 127872 4264 128896
rect 3944 127808 3952 127872
rect 4016 127808 4032 127872
rect 4096 127808 4112 127872
rect 4176 127808 4192 127872
rect 4256 127808 4264 127872
rect 3944 126784 4264 127808
rect 3944 126720 3952 126784
rect 4016 126720 4032 126784
rect 4096 126720 4112 126784
rect 4176 126720 4192 126784
rect 4256 126720 4264 126784
rect 3944 125696 4264 126720
rect 3944 125632 3952 125696
rect 4016 125632 4032 125696
rect 4096 125632 4112 125696
rect 4176 125632 4192 125696
rect 4256 125632 4264 125696
rect 3944 124608 4264 125632
rect 3944 124544 3952 124608
rect 4016 124544 4032 124608
rect 4096 124544 4112 124608
rect 4176 124544 4192 124608
rect 4256 124544 4264 124608
rect 3944 123520 4264 124544
rect 3944 123456 3952 123520
rect 4016 123456 4032 123520
rect 4096 123456 4112 123520
rect 4176 123456 4192 123520
rect 4256 123456 4264 123520
rect 3944 122432 4264 123456
rect 3944 122368 3952 122432
rect 4016 122368 4032 122432
rect 4096 122368 4112 122432
rect 4176 122368 4192 122432
rect 4256 122368 4264 122432
rect 3944 121344 4264 122368
rect 6134 121549 6194 126022
rect 82494 125576 82814 125618
rect 82494 125340 82536 125576
rect 82772 125340 82814 125576
rect 82494 125298 82814 125340
rect 6131 121548 6197 121549
rect 6131 121484 6132 121548
rect 6196 121484 6197 121548
rect 6131 121483 6197 121484
rect 3944 121280 3952 121344
rect 4016 121280 4032 121344
rect 4096 121280 4112 121344
rect 4176 121280 4192 121344
rect 4256 121280 4264 121344
rect 3944 120576 4264 121280
rect 3944 120340 3986 120576
rect 4222 120340 4264 120576
rect 3944 120256 4264 120340
rect 82938 120576 83262 120618
rect 82938 120340 82982 120576
rect 83218 120340 83262 120576
rect 82938 120298 83262 120340
rect 3944 120192 3952 120256
rect 4016 120192 4032 120256
rect 4096 120192 4112 120256
rect 4176 120192 4192 120256
rect 4256 120192 4264 120256
rect 3944 119168 4264 120192
rect 3944 119104 3952 119168
rect 4016 119104 4032 119168
rect 4096 119104 4112 119168
rect 4176 119104 4192 119168
rect 4256 119104 4264 119168
rect 3944 118080 4264 119104
rect 3944 118016 3952 118080
rect 4016 118016 4032 118080
rect 4096 118016 4112 118080
rect 4176 118016 4192 118080
rect 4256 118016 4264 118080
rect 3944 116992 4264 118016
rect 3944 116928 3952 116992
rect 4016 116928 4032 116992
rect 4096 116928 4112 116992
rect 4176 116928 4192 116992
rect 4256 116928 4264 116992
rect 3944 115904 4264 116928
rect 3944 115840 3952 115904
rect 4016 115840 4032 115904
rect 4096 115840 4112 115904
rect 4176 115840 4192 115904
rect 4256 115840 4264 115904
rect 3944 114816 4264 115840
rect 82494 115576 82814 115618
rect 82494 115340 82536 115576
rect 82772 115340 82814 115576
rect 82494 115298 82814 115340
rect 3944 114752 3952 114816
rect 4016 114752 4032 114816
rect 4096 114752 4112 114816
rect 4176 114752 4192 114816
rect 4256 114752 4264 114816
rect 3944 113728 4264 114752
rect 83414 114341 83474 132227
rect 83411 114340 83477 114341
rect 83411 114276 83412 114340
rect 83476 114276 83477 114340
rect 83411 114275 83477 114276
rect 83411 113932 83477 113933
rect 83411 113868 83412 113932
rect 83476 113868 83477 113932
rect 83411 113867 83477 113868
rect 3944 113664 3952 113728
rect 4016 113664 4032 113728
rect 4096 113664 4112 113728
rect 4176 113664 4192 113728
rect 4256 113664 4264 113728
rect 3944 112640 4264 113664
rect 3944 112576 3952 112640
rect 4016 112576 4032 112640
rect 4096 112576 4112 112640
rect 4176 112576 4192 112640
rect 4256 112576 4264 112640
rect 3944 111552 4264 112576
rect 3944 111488 3952 111552
rect 4016 111488 4032 111552
rect 4096 111488 4112 111552
rect 4176 111488 4192 111552
rect 4256 111488 4264 111552
rect 3944 110576 4264 111488
rect 3944 110464 3986 110576
rect 4222 110464 4264 110576
rect 3944 110400 3952 110464
rect 4256 110400 4264 110464
rect 3944 110340 3986 110400
rect 4222 110340 4264 110400
rect 3944 109376 4264 110340
rect 82938 110576 83262 110618
rect 82938 110340 82982 110576
rect 83218 110340 83262 110576
rect 82938 110298 83262 110340
rect 3944 109312 3952 109376
rect 4016 109312 4032 109376
rect 4096 109312 4112 109376
rect 4176 109312 4192 109376
rect 4256 109312 4264 109376
rect 3944 108288 4264 109312
rect 3944 108224 3952 108288
rect 4016 108224 4032 108288
rect 4096 108224 4112 108288
rect 4176 108224 4192 108288
rect 4256 108224 4264 108288
rect 3944 107200 4264 108224
rect 3944 107136 3952 107200
rect 4016 107136 4032 107200
rect 4096 107136 4112 107200
rect 4176 107136 4192 107200
rect 4256 107136 4264 107200
rect 3944 106112 4264 107136
rect 3944 106048 3952 106112
rect 4016 106048 4032 106112
rect 4096 106048 4112 106112
rect 4176 106048 4192 106112
rect 4256 106048 4264 106112
rect 3944 105024 4264 106048
rect 82494 105576 82814 105618
rect 82494 105340 82536 105576
rect 82772 105340 82814 105576
rect 82494 105298 82814 105340
rect 3944 104960 3952 105024
rect 4016 104960 4032 105024
rect 4096 104960 4112 105024
rect 4176 104960 4192 105024
rect 4256 104960 4264 105024
rect 3944 103936 4264 104960
rect 3944 103872 3952 103936
rect 4016 103872 4032 103936
rect 4096 103872 4112 103936
rect 4176 103872 4192 103936
rect 4256 103872 4264 103936
rect 3944 102848 4264 103872
rect 3944 102784 3952 102848
rect 4016 102784 4032 102848
rect 4096 102784 4112 102848
rect 4176 102784 4192 102848
rect 4256 102784 4264 102848
rect 3944 101760 4264 102784
rect 3944 101696 3952 101760
rect 4016 101696 4032 101760
rect 4096 101696 4112 101760
rect 4176 101696 4192 101760
rect 4256 101696 4264 101760
rect 3944 100672 4264 101696
rect 3944 100608 3952 100672
rect 4016 100608 4032 100672
rect 4096 100608 4112 100672
rect 4176 100608 4192 100672
rect 4256 100608 4264 100672
rect 3944 100576 4264 100608
rect 3944 100340 3986 100576
rect 4222 100340 4264 100576
rect 3944 99584 4264 100340
rect 82938 100576 83262 100618
rect 82938 100340 82982 100576
rect 83218 100340 83262 100576
rect 82938 100298 83262 100340
rect 3944 99520 3952 99584
rect 4016 99520 4032 99584
rect 4096 99520 4112 99584
rect 4176 99520 4192 99584
rect 4256 99520 4264 99584
rect 3944 98496 4264 99520
rect 3944 98432 3952 98496
rect 4016 98432 4032 98496
rect 4096 98432 4112 98496
rect 4176 98432 4192 98496
rect 4256 98432 4264 98496
rect 3944 97408 4264 98432
rect 3944 97344 3952 97408
rect 4016 97344 4032 97408
rect 4096 97344 4112 97408
rect 4176 97344 4192 97408
rect 4256 97344 4264 97408
rect 3944 96320 4264 97344
rect 22691 97204 22757 97205
rect 22691 97140 22692 97204
rect 22756 97140 22757 97204
rect 22691 97139 22757 97140
rect 40355 97204 40421 97205
rect 40355 97140 40356 97204
rect 40420 97140 40421 97204
rect 40355 97139 40421 97140
rect 79915 97204 79981 97205
rect 79915 97140 79916 97204
rect 79980 97140 79981 97204
rect 79915 97139 79981 97140
rect 14595 97068 14661 97069
rect 14595 97004 14596 97068
rect 14660 97004 14661 97068
rect 14595 97003 14661 97004
rect 17171 97068 17237 97069
rect 17171 97004 17172 97068
rect 17236 97004 17237 97068
rect 17171 97003 17237 97004
rect 18091 97068 18157 97069
rect 18091 97004 18092 97068
rect 18156 97004 18157 97068
rect 18091 97003 18157 97004
rect 14598 96930 14658 97003
rect 17174 96930 17234 97003
rect 18094 96930 18154 97003
rect 22694 96930 22754 97139
rect 24347 97068 24413 97069
rect 24347 97004 24348 97068
rect 24412 97004 24413 97068
rect 24347 97003 24413 97004
rect 25451 97068 25517 97069
rect 25451 97004 25452 97068
rect 25516 97004 25517 97068
rect 25451 97003 25517 97004
rect 30051 97068 30117 97069
rect 30051 97004 30052 97068
rect 30116 97004 30117 97068
rect 30051 97003 30117 97004
rect 32075 97068 32141 97069
rect 32075 97004 32076 97068
rect 32140 97004 32141 97068
rect 32075 97003 32141 97004
rect 33179 97068 33245 97069
rect 33179 97004 33180 97068
rect 33244 97004 33245 97068
rect 33179 97003 33245 97004
rect 24350 96930 24410 97003
rect 25454 96930 25514 97003
rect 30054 96930 30114 97003
rect 32078 96930 32138 97003
rect 33182 96930 33242 97003
rect 35939 96932 36005 96933
rect 14000 96870 14658 96930
rect 16336 96870 16498 96930
rect 17174 96870 17504 96930
rect 18094 96870 18672 96930
rect 22694 96870 23344 96930
rect 24350 96870 24512 96930
rect 25454 96870 25680 96930
rect 30054 96870 30352 96930
rect 32078 96870 32688 96930
rect 33182 96870 33856 96930
rect 3944 96256 3952 96320
rect 4016 96256 4032 96320
rect 4096 96256 4112 96320
rect 4176 96256 4192 96320
rect 4256 96256 4264 96320
rect 3944 95232 4264 96256
rect 9630 96530 9833 96590
rect 12758 96530 12832 96590
rect 15168 96530 15762 96590
rect 9630 96253 9690 96530
rect 9627 96252 9693 96253
rect 9627 96188 9628 96252
rect 9692 96188 9693 96252
rect 9627 96187 9693 96188
rect 3944 95168 3952 95232
rect 4016 95168 4032 95232
rect 4096 95168 4112 95232
rect 4176 95168 4192 95232
rect 4256 95168 4264 95232
rect 3944 94144 4264 95168
rect 12758 95165 12818 96530
rect 15702 96389 15762 96530
rect 16438 96525 16498 96870
rect 35939 96868 35940 96932
rect 36004 96930 36005 96932
rect 40358 96930 40418 97139
rect 42931 97068 42997 97069
rect 42931 97004 42932 97068
rect 42996 97004 42997 97068
rect 42931 97003 42997 97004
rect 42934 96930 42994 97003
rect 36004 96870 36192 96930
rect 40358 96870 40864 96930
rect 42750 96870 43200 96930
rect 46828 96870 47226 96930
rect 51500 96870 52194 96930
rect 52668 96870 53150 96930
rect 36004 96868 36005 96870
rect 35939 96867 36005 96868
rect 40542 96797 40602 96870
rect 40539 96796 40605 96797
rect 40539 96732 40540 96796
rect 40604 96732 40605 96796
rect 40539 96731 40605 96732
rect 42750 96661 42810 96870
rect 47166 96797 47226 96870
rect 52134 96797 52194 96870
rect 47163 96796 47229 96797
rect 47163 96732 47164 96796
rect 47228 96732 47229 96796
rect 47163 96731 47229 96732
rect 52131 96796 52197 96797
rect 52131 96732 52132 96796
rect 52196 96732 52197 96796
rect 56550 96870 58082 96930
rect 52131 96731 52197 96732
rect 42747 96660 42813 96661
rect 42747 96596 42748 96660
rect 42812 96596 42813 96660
rect 42747 96595 42813 96596
rect 18796 96530 19258 96590
rect 16435 96524 16501 96525
rect 16435 96460 16436 96524
rect 16500 96460 16501 96524
rect 16435 96459 16501 96460
rect 15699 96388 15765 96389
rect 15699 96324 15700 96388
rect 15764 96324 15765 96388
rect 15699 96323 15765 96324
rect 12755 95164 12821 95165
rect 12755 95100 12756 95164
rect 12820 95100 12821 95164
rect 12755 95099 12821 95100
rect 3944 94080 3952 94144
rect 4016 94080 4032 94144
rect 4096 94080 4112 94144
rect 4176 94080 4192 94144
rect 4256 94080 4264 94144
rect 3944 93056 4264 94080
rect 3944 92992 3952 93056
rect 4016 92992 4032 93056
rect 4096 92992 4112 93056
rect 4176 92992 4192 93056
rect 4256 92992 4264 93056
rect 3944 91968 4264 92992
rect 3944 91904 3952 91968
rect 4016 91904 4032 91968
rect 4096 91904 4112 91968
rect 4176 91904 4192 91968
rect 4256 91904 4264 91968
rect 3944 90880 4264 91904
rect 3944 90816 3952 90880
rect 4016 90816 4032 90880
rect 4096 90816 4112 90880
rect 4176 90816 4192 90880
rect 4256 90816 4264 90880
rect 3944 90576 4264 90816
rect 3944 90340 3986 90576
rect 4222 90340 4264 90576
rect 3944 89792 4264 90340
rect 3944 89728 3952 89792
rect 4016 89728 4032 89792
rect 4096 89728 4112 89792
rect 4176 89728 4192 89792
rect 4256 89728 4264 89792
rect 3944 88704 4264 89728
rect 3944 88640 3952 88704
rect 4016 88640 4032 88704
rect 4096 88640 4112 88704
rect 4176 88640 4192 88704
rect 4256 88640 4264 88704
rect 3944 87616 4264 88640
rect 3944 87552 3952 87616
rect 4016 87552 4032 87616
rect 4096 87552 4112 87616
rect 4176 87552 4192 87616
rect 4256 87552 4264 87616
rect 3944 86528 4264 87552
rect 3944 86464 3952 86528
rect 4016 86464 4032 86528
rect 4096 86464 4112 86528
rect 4176 86464 4192 86528
rect 4256 86464 4264 86528
rect 3944 85440 4264 86464
rect 3944 85376 3952 85440
rect 4016 85376 4032 85440
rect 4096 85376 4112 85440
rect 4176 85376 4192 85440
rect 4256 85376 4264 85440
rect 3944 84352 4264 85376
rect 3944 84288 3952 84352
rect 4016 84288 4032 84352
rect 4096 84288 4112 84352
rect 4176 84288 4192 84352
rect 4256 84288 4264 84352
rect 3944 83264 4264 84288
rect 3944 83200 3952 83264
rect 4016 83200 4032 83264
rect 4096 83200 4112 83264
rect 4176 83200 4192 83264
rect 4256 83200 4264 83264
rect 3944 82176 4264 83200
rect 3944 82112 3952 82176
rect 4016 82112 4032 82176
rect 4096 82112 4112 82176
rect 4176 82112 4192 82176
rect 4256 82112 4264 82176
rect 3944 81088 4264 82112
rect 3944 81024 3952 81088
rect 4016 81024 4032 81088
rect 4096 81024 4112 81088
rect 4176 81024 4192 81088
rect 4256 81024 4264 81088
rect 3944 80576 4264 81024
rect 3944 80340 3986 80576
rect 4222 80340 4264 80576
rect 3944 80000 4264 80340
rect 3944 79936 3952 80000
rect 4016 79936 4032 80000
rect 4096 79936 4112 80000
rect 4176 79936 4192 80000
rect 4256 79936 4264 80000
rect 3944 78912 4264 79936
rect 3944 78848 3952 78912
rect 4016 78848 4032 78912
rect 4096 78848 4112 78912
rect 4176 78848 4192 78912
rect 4256 78848 4264 78912
rect 3944 77824 4264 78848
rect 3944 77760 3952 77824
rect 4016 77760 4032 77824
rect 4096 77760 4112 77824
rect 4176 77760 4192 77824
rect 4256 77760 4264 77824
rect 3944 76736 4264 77760
rect 3944 76672 3952 76736
rect 4016 76672 4032 76736
rect 4096 76672 4112 76736
rect 4176 76672 4192 76736
rect 4256 76672 4264 76736
rect 3944 75648 4264 76672
rect 3944 75584 3952 75648
rect 4016 75584 4032 75648
rect 4096 75584 4112 75648
rect 4176 75584 4192 75648
rect 4256 75584 4264 75648
rect 3944 74560 4264 75584
rect 3944 74496 3952 74560
rect 4016 74496 4032 74560
rect 4096 74496 4112 74560
rect 4176 74496 4192 74560
rect 4256 74496 4264 74560
rect 3944 73472 4264 74496
rect 3944 73408 3952 73472
rect 4016 73408 4032 73472
rect 4096 73408 4112 73472
rect 4176 73408 4192 73472
rect 4256 73408 4264 73472
rect 3944 72384 4264 73408
rect 3944 72320 3952 72384
rect 4016 72320 4032 72384
rect 4096 72320 4112 72384
rect 4176 72320 4192 72384
rect 4256 72320 4264 72384
rect 3944 71296 4264 72320
rect 3944 71232 3952 71296
rect 4016 71232 4032 71296
rect 4096 71232 4112 71296
rect 4176 71232 4192 71296
rect 4256 71232 4264 71296
rect 3944 70576 4264 71232
rect 3944 70340 3986 70576
rect 4222 70340 4264 70576
rect 3944 70208 4264 70340
rect 3944 70144 3952 70208
rect 4016 70144 4032 70208
rect 4096 70144 4112 70208
rect 4176 70144 4192 70208
rect 4256 70144 4264 70208
rect 3944 69120 4264 70144
rect 3944 69056 3952 69120
rect 4016 69056 4032 69120
rect 4096 69056 4112 69120
rect 4176 69056 4192 69120
rect 4256 69056 4264 69120
rect 3944 68032 4264 69056
rect 3944 67968 3952 68032
rect 4016 67968 4032 68032
rect 4096 67968 4112 68032
rect 4176 67968 4192 68032
rect 4256 67968 4264 68032
rect 3944 66944 4264 67968
rect 3944 66880 3952 66944
rect 4016 66880 4032 66944
rect 4096 66880 4112 66944
rect 4176 66880 4192 66944
rect 4256 66880 4264 66944
rect 3944 65856 4264 66880
rect 3944 65792 3952 65856
rect 4016 65792 4032 65856
rect 4096 65792 4112 65856
rect 4176 65792 4192 65856
rect 4256 65792 4264 65856
rect 3944 64768 4264 65792
rect 3944 64704 3952 64768
rect 4016 64704 4032 64768
rect 4096 64704 4112 64768
rect 4176 64704 4192 64768
rect 4256 64704 4264 64768
rect 3944 63680 4264 64704
rect 3944 63616 3952 63680
rect 4016 63616 4032 63680
rect 4096 63616 4112 63680
rect 4176 63616 4192 63680
rect 4256 63616 4264 63680
rect 3944 62592 4264 63616
rect 3944 62528 3952 62592
rect 4016 62528 4032 62592
rect 4096 62528 4112 62592
rect 4176 62528 4192 62592
rect 4256 62528 4264 62592
rect 3944 61504 4264 62528
rect 3944 61440 3952 61504
rect 4016 61440 4032 61504
rect 4096 61440 4112 61504
rect 4176 61440 4192 61504
rect 4256 61440 4264 61504
rect 3944 60576 4264 61440
rect 3944 60416 3986 60576
rect 4222 60416 4264 60576
rect 3944 60352 3952 60416
rect 4256 60352 4264 60416
rect 3944 60340 3986 60352
rect 4222 60340 4264 60352
rect 3944 59328 4264 60340
rect 3944 59264 3952 59328
rect 4016 59264 4032 59328
rect 4096 59264 4112 59328
rect 4176 59264 4192 59328
rect 4256 59264 4264 59328
rect 3944 58240 4264 59264
rect 3944 58176 3952 58240
rect 4016 58176 4032 58240
rect 4096 58176 4112 58240
rect 4176 58176 4192 58240
rect 4256 58176 4264 58240
rect 3944 57152 4264 58176
rect 3944 57088 3952 57152
rect 4016 57088 4032 57152
rect 4096 57088 4112 57152
rect 4176 57088 4192 57152
rect 4256 57088 4264 57152
rect 3944 56064 4264 57088
rect 3944 56000 3952 56064
rect 4016 56000 4032 56064
rect 4096 56000 4112 56064
rect 4176 56000 4192 56064
rect 4256 56000 4264 56064
rect 3944 54976 4264 56000
rect 3944 54912 3952 54976
rect 4016 54912 4032 54976
rect 4096 54912 4112 54976
rect 4176 54912 4192 54976
rect 4256 54912 4264 54976
rect 3944 53888 4264 54912
rect 3944 53824 3952 53888
rect 4016 53824 4032 53888
rect 4096 53824 4112 53888
rect 4176 53824 4192 53888
rect 4256 53824 4264 53888
rect 3944 52800 4264 53824
rect 3944 52736 3952 52800
rect 4016 52736 4032 52800
rect 4096 52736 4112 52800
rect 4176 52736 4192 52800
rect 4256 52736 4264 52800
rect 3944 51712 4264 52736
rect 3944 51648 3952 51712
rect 4016 51648 4032 51712
rect 4096 51648 4112 51712
rect 4176 51648 4192 51712
rect 4256 51648 4264 51712
rect 3944 50624 4264 51648
rect 3944 50560 3952 50624
rect 4016 50576 4032 50624
rect 4096 50576 4112 50624
rect 4176 50576 4192 50624
rect 4256 50560 4264 50624
rect 3944 50340 3986 50560
rect 4222 50340 4264 50560
rect 3944 49536 4264 50340
rect 3944 49472 3952 49536
rect 4016 49472 4032 49536
rect 4096 49472 4112 49536
rect 4176 49472 4192 49536
rect 4256 49472 4264 49536
rect 3944 48448 4264 49472
rect 3944 48384 3952 48448
rect 4016 48384 4032 48448
rect 4096 48384 4112 48448
rect 4176 48384 4192 48448
rect 4256 48384 4264 48448
rect 3944 47360 4264 48384
rect 3944 47296 3952 47360
rect 4016 47296 4032 47360
rect 4096 47296 4112 47360
rect 4176 47296 4192 47360
rect 4256 47296 4264 47360
rect 3944 46272 4264 47296
rect 3944 46208 3952 46272
rect 4016 46208 4032 46272
rect 4096 46208 4112 46272
rect 4176 46208 4192 46272
rect 4256 46208 4264 46272
rect 3944 45184 4264 46208
rect 3944 45120 3952 45184
rect 4016 45120 4032 45184
rect 4096 45120 4112 45184
rect 4176 45120 4192 45184
rect 4256 45120 4264 45184
rect 3944 44096 4264 45120
rect 3944 44032 3952 44096
rect 4016 44032 4032 44096
rect 4096 44032 4112 44096
rect 4176 44032 4192 44096
rect 4256 44032 4264 44096
rect 3944 43008 4264 44032
rect 3944 42944 3952 43008
rect 4016 42944 4032 43008
rect 4096 42944 4112 43008
rect 4176 42944 4192 43008
rect 4256 42944 4264 43008
rect 3944 41920 4264 42944
rect 3944 41856 3952 41920
rect 4016 41856 4032 41920
rect 4096 41856 4112 41920
rect 4176 41856 4192 41920
rect 4256 41856 4264 41920
rect 3944 40832 4264 41856
rect 3944 40768 3952 40832
rect 4016 40768 4032 40832
rect 4096 40768 4112 40832
rect 4176 40768 4192 40832
rect 4256 40768 4264 40832
rect 3944 40576 4264 40768
rect 3944 40340 3986 40576
rect 4222 40340 4264 40576
rect 3944 39744 4264 40340
rect 3944 39680 3952 39744
rect 4016 39680 4032 39744
rect 4096 39680 4112 39744
rect 4176 39680 4192 39744
rect 4256 39680 4264 39744
rect 3944 38656 4264 39680
rect 3944 38592 3952 38656
rect 4016 38592 4032 38656
rect 4096 38592 4112 38656
rect 4176 38592 4192 38656
rect 4256 38592 4264 38656
rect 3944 37568 4264 38592
rect 3944 37504 3952 37568
rect 4016 37504 4032 37568
rect 4096 37504 4112 37568
rect 4176 37504 4192 37568
rect 4256 37504 4264 37568
rect 3944 36480 4264 37504
rect 3944 36416 3952 36480
rect 4016 36416 4032 36480
rect 4096 36416 4112 36480
rect 4176 36416 4192 36480
rect 4256 36416 4264 36480
rect 3944 35392 4264 36416
rect 3944 35328 3952 35392
rect 4016 35328 4032 35392
rect 4096 35328 4112 35392
rect 4176 35328 4192 35392
rect 4256 35328 4264 35392
rect 3944 34304 4264 35328
rect 3944 34240 3952 34304
rect 4016 34240 4032 34304
rect 4096 34240 4112 34304
rect 4176 34240 4192 34304
rect 4256 34240 4264 34304
rect 3944 33216 4264 34240
rect 3944 33152 3952 33216
rect 4016 33152 4032 33216
rect 4096 33152 4112 33216
rect 4176 33152 4192 33216
rect 4256 33152 4264 33216
rect 3944 32128 4264 33152
rect 3944 32064 3952 32128
rect 4016 32064 4032 32128
rect 4096 32064 4112 32128
rect 4176 32064 4192 32128
rect 4256 32064 4264 32128
rect 3944 31040 4264 32064
rect 3944 30976 3952 31040
rect 4016 30976 4032 31040
rect 4096 30976 4112 31040
rect 4176 30976 4192 31040
rect 4256 30976 4264 31040
rect 3944 30576 4264 30976
rect 3944 30340 3986 30576
rect 4222 30340 4264 30576
rect 3944 29952 4264 30340
rect 3944 29888 3952 29952
rect 4016 29888 4032 29952
rect 4096 29888 4112 29952
rect 4176 29888 4192 29952
rect 4256 29888 4264 29952
rect 3944 28864 4264 29888
rect 3944 28800 3952 28864
rect 4016 28800 4032 28864
rect 4096 28800 4112 28864
rect 4176 28800 4192 28864
rect 4256 28800 4264 28864
rect 3944 27776 4264 28800
rect 3944 27712 3952 27776
rect 4016 27712 4032 27776
rect 4096 27712 4112 27776
rect 4176 27712 4192 27776
rect 4256 27712 4264 27776
rect 3944 26688 4264 27712
rect 3944 26624 3952 26688
rect 4016 26624 4032 26688
rect 4096 26624 4112 26688
rect 4176 26624 4192 26688
rect 4256 26624 4264 26688
rect 3944 25600 4264 26624
rect 3944 25536 3952 25600
rect 4016 25536 4032 25600
rect 4096 25536 4112 25600
rect 4176 25536 4192 25600
rect 4256 25536 4264 25600
rect 3944 24512 4264 25536
rect 3944 24448 3952 24512
rect 4016 24448 4032 24512
rect 4096 24448 4112 24512
rect 4176 24448 4192 24512
rect 4256 24448 4264 24512
rect 3944 23424 4264 24448
rect 3944 23360 3952 23424
rect 4016 23360 4032 23424
rect 4096 23360 4112 23424
rect 4176 23360 4192 23424
rect 4256 23360 4264 23424
rect 3944 22336 4264 23360
rect 3944 22272 3952 22336
rect 4016 22272 4032 22336
rect 4096 22272 4112 22336
rect 4176 22272 4192 22336
rect 4256 22272 4264 22336
rect 3944 21248 4264 22272
rect 3944 21184 3952 21248
rect 4016 21184 4032 21248
rect 4096 21184 4112 21248
rect 4176 21184 4192 21248
rect 4256 21184 4264 21248
rect 3944 20576 4264 21184
rect 3944 20340 3986 20576
rect 4222 20340 4264 20576
rect 3944 20160 4264 20340
rect 3944 20096 3952 20160
rect 4016 20096 4032 20160
rect 4096 20096 4112 20160
rect 4176 20096 4192 20160
rect 4256 20096 4264 20160
rect 3944 19072 4264 20096
rect 3944 19008 3952 19072
rect 4016 19008 4032 19072
rect 4096 19008 4112 19072
rect 4176 19008 4192 19072
rect 4256 19008 4264 19072
rect 3944 17984 4264 19008
rect 3944 17920 3952 17984
rect 4016 17920 4032 17984
rect 4096 17920 4112 17984
rect 4176 17920 4192 17984
rect 4256 17920 4264 17984
rect 3944 16896 4264 17920
rect 3944 16832 3952 16896
rect 4016 16832 4032 16896
rect 4096 16832 4112 16896
rect 4176 16832 4192 16896
rect 4256 16832 4264 16896
rect 3944 15808 4264 16832
rect 3944 15744 3952 15808
rect 4016 15744 4032 15808
rect 4096 15744 4112 15808
rect 4176 15744 4192 15808
rect 4256 15744 4264 15808
rect 3944 14720 4264 15744
rect 3944 14656 3952 14720
rect 4016 14656 4032 14720
rect 4096 14656 4112 14720
rect 4176 14656 4192 14720
rect 4256 14656 4264 14720
rect 3944 13632 4264 14656
rect 3944 13568 3952 13632
rect 4016 13568 4032 13632
rect 4096 13568 4112 13632
rect 4176 13568 4192 13632
rect 4256 13568 4264 13632
rect 3944 12544 4264 13568
rect 3944 12480 3952 12544
rect 4016 12480 4032 12544
rect 4096 12480 4112 12544
rect 4176 12480 4192 12544
rect 4256 12480 4264 12544
rect 3944 11456 4264 12480
rect 3944 11392 3952 11456
rect 4016 11392 4032 11456
rect 4096 11392 4112 11456
rect 4176 11392 4192 11456
rect 4256 11392 4264 11456
rect 3944 10576 4264 11392
rect 3944 10368 3986 10576
rect 4222 10368 4264 10576
rect 3944 10304 3952 10368
rect 4016 10304 4032 10340
rect 4096 10304 4112 10340
rect 4176 10304 4192 10340
rect 4256 10304 4264 10368
rect 3944 9280 4264 10304
rect 4478 10165 4538 94062
rect 19198 93941 19258 96530
rect 19382 96530 19840 96590
rect 19382 95165 19442 96530
rect 19379 95164 19445 95165
rect 19379 95100 19380 95164
rect 19444 95100 19445 95164
rect 19379 95099 19445 95100
rect 19934 94893 19994 96560
rect 20978 96117 21038 96560
rect 21132 96530 21282 96590
rect 21222 96389 21282 96530
rect 21219 96388 21285 96389
rect 21219 96324 21220 96388
rect 21284 96324 21285 96388
rect 21219 96323 21285 96324
rect 22142 96253 22202 96590
rect 22300 96530 22938 96590
rect 23468 96530 24042 96590
rect 22139 96252 22205 96253
rect 22139 96188 22140 96252
rect 22204 96188 22205 96252
rect 22139 96187 22205 96188
rect 20975 96116 21041 96117
rect 20975 96052 20976 96116
rect 21040 96052 21041 96116
rect 20975 96051 21041 96052
rect 22878 95029 22938 96530
rect 23982 95437 24042 96530
rect 24606 96250 24666 96560
rect 25804 96530 25882 96590
rect 24606 96190 24778 96250
rect 23979 95436 24045 95437
rect 23979 95372 23980 95436
rect 24044 95372 24045 95436
rect 23979 95371 24045 95372
rect 24531 95300 24597 95301
rect 24531 95236 24532 95300
rect 24596 95236 24597 95300
rect 24531 95235 24597 95236
rect 22875 95028 22941 95029
rect 22875 94964 22876 95028
rect 22940 94964 22941 95028
rect 22875 94963 22941 94964
rect 19931 94892 19997 94893
rect 19931 94828 19932 94892
rect 19996 94828 19997 94892
rect 19931 94827 19997 94828
rect 19195 93940 19261 93941
rect 19195 93876 19196 93940
rect 19260 93876 19261 93940
rect 19195 93875 19261 93876
rect 24534 93530 24594 95235
rect 24718 95165 24778 96190
rect 25822 95165 25882 96530
rect 26818 96117 26878 96560
rect 26972 96530 27538 96590
rect 26815 96116 26881 96117
rect 26815 96052 26816 96116
rect 26880 96052 26881 96116
rect 26815 96051 26881 96052
rect 27478 95165 27538 96530
rect 27986 96253 28046 96560
rect 28140 96530 28826 96590
rect 27983 96252 28049 96253
rect 27983 96188 27984 96252
rect 28048 96188 28049 96252
rect 27983 96187 28049 96188
rect 28766 95573 28826 96530
rect 29154 96253 29214 96560
rect 29308 96530 29930 96590
rect 30476 96530 31034 96590
rect 29151 96252 29217 96253
rect 29151 96188 29152 96252
rect 29216 96188 29217 96252
rect 29151 96187 29217 96188
rect 28763 95572 28829 95573
rect 28763 95508 28764 95572
rect 28828 95508 28829 95572
rect 28763 95507 28829 95508
rect 24715 95164 24781 95165
rect 24715 95100 24716 95164
rect 24780 95100 24781 95164
rect 24715 95099 24781 95100
rect 25819 95164 25885 95165
rect 25819 95100 25820 95164
rect 25884 95100 25885 95164
rect 25819 95099 25885 95100
rect 27475 95164 27541 95165
rect 27475 95100 27476 95164
rect 27540 95100 27541 95164
rect 27475 95099 27541 95100
rect 29870 95029 29930 96530
rect 30974 95029 31034 96530
rect 31490 96117 31550 96560
rect 31614 96250 31674 96560
rect 32812 96530 33058 96590
rect 33980 96530 34530 96590
rect 31614 96190 31770 96250
rect 31487 96116 31553 96117
rect 31487 96052 31488 96116
rect 31552 96052 31553 96116
rect 31487 96051 31553 96052
rect 29867 95028 29933 95029
rect 29867 94964 29868 95028
rect 29932 94964 29933 95028
rect 29867 94963 29933 94964
rect 30971 95028 31037 95029
rect 30971 94964 30972 95028
rect 31036 94964 31037 95028
rect 30971 94963 31037 94964
rect 31710 94893 31770 96190
rect 32998 95709 33058 96530
rect 32995 95708 33061 95709
rect 32995 95644 32996 95708
rect 33060 95644 33061 95708
rect 32995 95643 33061 95644
rect 31707 94892 31773 94893
rect 31707 94828 31708 94892
rect 31772 94828 31773 94892
rect 31707 94827 31773 94828
rect 34470 94757 34530 96530
rect 34994 96117 35054 96560
rect 35148 96530 35818 96590
rect 36316 96530 36922 96590
rect 34991 96116 35057 96117
rect 34991 96052 34992 96116
rect 35056 96052 35057 96116
rect 34991 96051 35057 96052
rect 34467 94756 34533 94757
rect 34467 94692 34468 94756
rect 34532 94692 34533 94756
rect 34467 94691 34533 94692
rect 35758 93805 35818 96530
rect 36862 94485 36922 96530
rect 37330 96250 37390 96560
rect 37484 96530 38026 96590
rect 37230 96190 37390 96250
rect 37230 94621 37290 96190
rect 37779 95300 37845 95301
rect 37779 95236 37780 95300
rect 37844 95236 37845 95300
rect 37779 95235 37845 95236
rect 37227 94620 37293 94621
rect 37227 94556 37228 94620
rect 37292 94556 37293 94620
rect 37227 94555 37293 94556
rect 36859 94484 36925 94485
rect 36859 94420 36860 94484
rect 36924 94420 36925 94484
rect 36859 94419 36925 94420
rect 35755 93804 35821 93805
rect 35755 93740 35756 93804
rect 35820 93740 35821 93804
rect 35755 93739 35821 93740
rect 31707 93668 31773 93669
rect 31707 93604 31708 93668
rect 31772 93604 31773 93668
rect 31707 93603 31773 93604
rect 31710 93530 31770 93603
rect 37782 93530 37842 95235
rect 37966 95165 38026 96530
rect 38498 96250 38558 96560
rect 38652 96530 39314 96590
rect 38498 96190 38578 96250
rect 38518 95845 38578 96190
rect 38515 95844 38581 95845
rect 38515 95780 38516 95844
rect 38580 95780 38581 95844
rect 38515 95779 38581 95780
rect 37963 95164 38029 95165
rect 37963 95100 37964 95164
rect 38028 95100 38029 95164
rect 37963 95099 38029 95100
rect 39254 94213 39314 96530
rect 39622 96530 39696 96590
rect 39820 96530 40050 96590
rect 40988 96530 41338 96590
rect 39622 95981 39682 96530
rect 39619 95980 39685 95981
rect 39619 95916 39620 95980
rect 39684 95916 39685 95980
rect 39619 95915 39685 95916
rect 39990 94349 40050 96530
rect 41091 95300 41157 95301
rect 41091 95236 41092 95300
rect 41156 95236 41157 95300
rect 41091 95235 41157 95236
rect 39987 94348 40053 94349
rect 39987 94284 39988 94348
rect 40052 94284 40053 94348
rect 39987 94283 40053 94284
rect 39251 94212 39317 94213
rect 39251 94148 39252 94212
rect 39316 94148 39317 94212
rect 39251 94147 39317 94148
rect 41094 93870 41154 95235
rect 41278 94077 41338 96530
rect 42002 96253 42062 96560
rect 42156 96530 42626 96590
rect 43324 96530 43914 96590
rect 41999 96252 42065 96253
rect 41999 96188 42000 96252
rect 42064 96188 42065 96252
rect 41999 96187 42065 96188
rect 42566 94485 42626 96530
rect 43854 95165 43914 96530
rect 44338 96250 44398 96560
rect 44492 96530 45018 96590
rect 44338 96190 44466 96250
rect 44406 95165 44466 96190
rect 43851 95164 43917 95165
rect 43851 95100 43852 95164
rect 43916 95100 43917 95164
rect 43851 95099 43917 95100
rect 44403 95164 44469 95165
rect 44403 95100 44404 95164
rect 44468 95100 44469 95164
rect 44403 95099 44469 95100
rect 44958 94485 45018 96530
rect 45506 96250 45566 96560
rect 45660 96530 46306 96590
rect 45506 96190 45570 96250
rect 45323 95300 45389 95301
rect 45323 95236 45324 95300
rect 45388 95236 45389 95300
rect 45323 95235 45389 95236
rect 42563 94484 42629 94485
rect 42563 94420 42564 94484
rect 42628 94420 42629 94484
rect 42563 94419 42629 94420
rect 44955 94484 45021 94485
rect 44955 94420 44956 94484
rect 45020 94420 45021 94484
rect 44955 94419 45021 94420
rect 41275 94076 41341 94077
rect 41275 94012 41276 94076
rect 41340 94012 41341 94076
rect 41275 94011 41341 94012
rect 24534 93470 24835 93530
rect 27331 93470 27538 93530
rect 29827 93470 30298 93530
rect 31075 93470 31770 93530
rect 37315 93470 37842 93530
rect 41029 93810 41154 93870
rect 41029 93500 41089 93810
rect 42563 93668 42629 93669
rect 42563 93604 42564 93668
rect 42628 93604 42629 93668
rect 42563 93603 42629 93604
rect 44035 93668 44101 93669
rect 44035 93604 44036 93668
rect 44100 93604 44101 93668
rect 44035 93603 44101 93604
rect 42566 93530 42626 93603
rect 44038 93530 44098 93603
rect 45326 93530 45386 95235
rect 45510 95165 45570 96190
rect 45507 95164 45573 95165
rect 45507 95100 45508 95164
rect 45572 95100 45573 95164
rect 45507 95099 45573 95100
rect 46246 94485 46306 96530
rect 46614 96530 46704 96590
rect 46614 95165 46674 96530
rect 47842 96250 47902 96560
rect 47996 96530 48146 96590
rect 47842 96190 47962 96250
rect 47902 95301 47962 96190
rect 47899 95300 47965 95301
rect 47899 95236 47900 95300
rect 47964 95236 47965 95300
rect 47899 95235 47965 95236
rect 48086 95165 48146 96530
rect 46611 95164 46677 95165
rect 46611 95100 46612 95164
rect 46676 95100 46677 95164
rect 46611 95099 46677 95100
rect 48083 95164 48149 95165
rect 48083 95100 48084 95164
rect 48148 95100 48149 95164
rect 48083 95099 48149 95100
rect 46243 94484 46309 94485
rect 46243 94420 46244 94484
rect 46308 94420 46309 94484
rect 46243 94419 46309 94420
rect 49006 93669 49066 96590
rect 49164 96530 49250 96590
rect 49190 93870 49250 96530
rect 49926 96530 50208 96590
rect 50332 96530 50538 96590
rect 49190 93810 49434 93870
rect 46611 93668 46677 93669
rect 46611 93604 46612 93668
rect 46676 93604 46677 93668
rect 46611 93603 46677 93604
rect 47899 93668 47965 93669
rect 47899 93604 47900 93668
rect 47964 93604 47965 93668
rect 48267 93668 48333 93669
rect 48267 93618 48268 93668
rect 48332 93618 48333 93668
rect 49003 93668 49069 93669
rect 47899 93603 47965 93604
rect 46614 93530 46674 93603
rect 47902 93530 47962 93603
rect 42307 93470 42626 93530
rect 43555 93470 44098 93530
rect 44803 93470 45386 93530
rect 46051 93470 46674 93530
rect 47299 93470 47962 93530
rect 27478 93261 27538 93470
rect 30238 93397 30298 93470
rect 30235 93396 30301 93397
rect 30235 93332 30236 93396
rect 30300 93332 30301 93396
rect 49003 93604 49004 93668
rect 49068 93604 49069 93668
rect 49003 93603 49069 93604
rect 49187 93668 49253 93669
rect 49187 93604 49188 93668
rect 49252 93604 49253 93668
rect 49187 93603 49253 93604
rect 49190 93530 49250 93603
rect 48547 93470 49250 93530
rect 30235 93331 30301 93332
rect 49374 93278 49434 93810
rect 49926 93669 49986 96530
rect 50478 96389 50538 96530
rect 50475 96388 50541 96389
rect 50475 96324 50476 96388
rect 50540 96324 50541 96388
rect 51027 96388 51093 96389
rect 51027 96338 51028 96388
rect 51092 96338 51093 96388
rect 50475 96323 50541 96324
rect 51346 96250 51406 96560
rect 51346 96190 51458 96250
rect 51398 93669 51458 96190
rect 52502 93669 52562 96590
rect 53682 96250 53742 96560
rect 53836 96530 54402 96590
rect 54974 96570 55322 96630
rect 54974 96560 55034 96570
rect 53682 96190 53850 96250
rect 53790 94210 53850 96190
rect 53790 94150 54034 94210
rect 53974 93669 54034 94150
rect 54342 93669 54402 96530
rect 54850 96250 54910 96560
rect 54850 96190 54954 96250
rect 54894 93669 54954 96190
rect 55262 93669 55322 96570
rect 49923 93668 49989 93669
rect 49923 93604 49924 93668
rect 49988 93604 49989 93668
rect 49923 93603 49989 93604
rect 50291 93668 50357 93669
rect 50291 93604 50292 93668
rect 50356 93604 50357 93668
rect 50291 93603 50357 93604
rect 51211 93668 51277 93669
rect 51211 93604 51212 93668
rect 51276 93604 51277 93668
rect 51211 93603 51277 93604
rect 51395 93668 51461 93669
rect 51395 93604 51396 93668
rect 51460 93604 51461 93668
rect 51395 93603 51461 93604
rect 52131 93668 52197 93669
rect 52131 93604 52132 93668
rect 52196 93604 52197 93668
rect 52131 93603 52197 93604
rect 52499 93668 52565 93669
rect 52499 93604 52500 93668
rect 52564 93604 52565 93668
rect 53235 93668 53301 93669
rect 53235 93618 53236 93668
rect 53300 93618 53301 93668
rect 53787 93668 53853 93669
rect 52499 93603 52565 93604
rect 50294 93530 50354 93603
rect 51214 93530 51274 93603
rect 49795 93470 50354 93530
rect 51030 93470 51274 93530
rect 52134 93530 52194 93603
rect 52134 93470 52291 93530
rect 53787 93604 53788 93668
rect 53852 93604 53853 93668
rect 53787 93603 53853 93604
rect 53971 93668 54037 93669
rect 53971 93604 53972 93668
rect 54036 93604 54037 93668
rect 53971 93603 54037 93604
rect 54339 93668 54405 93669
rect 54339 93604 54340 93668
rect 54404 93604 54405 93668
rect 54339 93603 54405 93604
rect 54523 93668 54589 93669
rect 54523 93604 54524 93668
rect 54588 93604 54589 93668
rect 54523 93603 54589 93604
rect 54891 93668 54957 93669
rect 54891 93604 54892 93668
rect 54956 93604 54957 93668
rect 54891 93603 54957 93604
rect 55259 93668 55325 93669
rect 55259 93604 55260 93668
rect 55324 93604 55325 93668
rect 55259 93603 55325 93604
rect 53790 93530 53850 93603
rect 53539 93470 53850 93530
rect 54526 93530 54586 93603
rect 56550 93530 56610 96870
rect 58022 96661 58082 96870
rect 60595 96796 60661 96797
rect 58206 96734 58634 96794
rect 57835 96660 57901 96661
rect 57835 96596 57836 96660
rect 57900 96596 57901 96660
rect 57835 96595 57901 96596
rect 58019 96660 58085 96661
rect 58019 96596 58020 96660
rect 58084 96596 58085 96660
rect 58019 96595 58085 96596
rect 57838 93530 57898 96595
rect 58206 93618 58266 96734
rect 58387 96660 58453 96661
rect 58387 96596 58388 96660
rect 58452 96596 58453 96660
rect 58574 96658 58634 96734
rect 60595 96732 60596 96796
rect 60660 96732 60661 96796
rect 60595 96731 60661 96732
rect 61515 96796 61581 96797
rect 61515 96732 61516 96796
rect 61580 96732 61581 96796
rect 61515 96731 61581 96732
rect 61699 96796 61765 96797
rect 61699 96732 61700 96796
rect 61764 96794 61765 96796
rect 61764 96734 62130 96794
rect 61764 96732 61765 96734
rect 61699 96731 61765 96732
rect 59675 96660 59741 96661
rect 59675 96658 59676 96660
rect 58574 96598 59002 96658
rect 58387 96595 58453 96596
rect 54526 93470 54787 93530
rect 56035 93470 56610 93530
rect 57283 93470 57898 93530
rect 58216 93470 58266 93618
rect 58390 93666 58450 96595
rect 58390 93606 58561 93666
rect 58501 93500 58561 93606
rect 58942 93530 59002 96598
rect 59494 96598 59676 96658
rect 59494 94890 59554 96598
rect 59675 96596 59676 96598
rect 59740 96596 59741 96660
rect 59675 96595 59741 96596
rect 60227 96660 60293 96661
rect 60227 96596 60228 96660
rect 60292 96658 60293 96660
rect 60292 96598 60474 96658
rect 60292 96596 60293 96598
rect 60227 96595 60293 96596
rect 60414 96250 60474 96598
rect 60598 96630 60658 96731
rect 60598 96570 61026 96630
rect 60414 96190 60658 96250
rect 59494 94830 60290 94890
rect 58942 93470 59406 93530
rect 60230 93530 60290 94830
rect 60598 93618 60658 96190
rect 60966 94298 61026 96570
rect 59779 93470 60290 93530
rect 61518 93530 61578 96731
rect 61027 93470 61578 93530
rect 62070 93530 62130 96734
rect 79918 96630 79978 97139
rect 82491 96796 82557 96797
rect 82491 96732 82492 96796
rect 82556 96732 82557 96796
rect 82491 96731 82557 96732
rect 79918 96570 80162 96630
rect 80102 96250 80162 96570
rect 80102 96190 80530 96250
rect 75131 95572 75197 95573
rect 75131 95508 75132 95572
rect 75196 95508 75197 95572
rect 75131 95507 75197 95508
rect 79179 95572 79245 95573
rect 79179 95508 79180 95572
rect 79244 95570 79245 95572
rect 79244 95510 79794 95570
rect 79244 95508 79245 95510
rect 79179 95507 79245 95508
rect 64091 95300 64157 95301
rect 64091 95236 64092 95300
rect 64156 95236 64157 95300
rect 64091 95235 64157 95236
rect 64094 93530 64154 95235
rect 75134 93530 75194 95507
rect 79734 95029 79794 95510
rect 80470 95029 80530 96190
rect 79731 95028 79797 95029
rect 79731 94964 79732 95028
rect 79796 94964 79797 95028
rect 79731 94963 79797 94964
rect 80467 95028 80533 95029
rect 80467 94964 80468 95028
rect 80532 94964 80533 95028
rect 80467 94963 80533 94964
rect 77250 94150 77438 94210
rect 76790 93666 76850 94062
rect 77250 93666 77310 94150
rect 82494 93805 82554 96731
rect 83414 94213 83474 113867
rect 83598 94349 83658 175339
rect 85944 175200 86264 175340
rect 85944 175136 85952 175200
rect 86016 175136 86032 175200
rect 86096 175136 86112 175200
rect 86176 175136 86192 175200
rect 86256 175136 86264 175200
rect 85944 174112 86264 175136
rect 85944 174048 85952 174112
rect 86016 174048 86032 174112
rect 86096 174048 86112 174112
rect 86176 174048 86192 174112
rect 86256 174048 86264 174112
rect 85944 173024 86264 174048
rect 85944 172960 85952 173024
rect 86016 172960 86032 173024
rect 86096 172960 86112 173024
rect 86176 172960 86192 173024
rect 86256 172960 86264 173024
rect 85944 171936 86264 172960
rect 85944 171872 85952 171936
rect 86016 171872 86032 171936
rect 86096 171872 86112 171936
rect 86176 171872 86192 171936
rect 86256 171872 86264 171936
rect 85944 170848 86264 171872
rect 85944 170784 85952 170848
rect 86016 170784 86032 170848
rect 86096 170784 86112 170848
rect 86176 170784 86192 170848
rect 86256 170784 86264 170848
rect 85944 169760 86264 170784
rect 85944 169696 85952 169760
rect 86016 169696 86032 169760
rect 86096 169696 86112 169760
rect 86176 169696 86192 169760
rect 86256 169696 86264 169760
rect 85944 168672 86264 169696
rect 85944 168608 85952 168672
rect 86016 168608 86032 168672
rect 86096 168608 86112 168672
rect 86176 168608 86192 168672
rect 86256 168608 86264 168672
rect 85944 167584 86264 168608
rect 85944 167520 85952 167584
rect 86016 167520 86032 167584
rect 86096 167520 86112 167584
rect 86176 167520 86192 167584
rect 86256 167520 86264 167584
rect 83779 167380 83845 167381
rect 83779 167316 83780 167380
rect 83844 167316 83845 167380
rect 83779 167315 83845 167316
rect 83782 94893 83842 167315
rect 85944 166496 86264 167520
rect 85944 166432 85952 166496
rect 86016 166432 86032 166496
rect 86096 166432 86112 166496
rect 86176 166432 86192 166496
rect 86256 166432 86264 166496
rect 85944 165576 86264 166432
rect 85944 165408 85986 165576
rect 86222 165408 86264 165576
rect 85944 165344 85952 165408
rect 86256 165344 86264 165408
rect 85944 165340 85986 165344
rect 86222 165340 86264 165344
rect 85944 164320 86264 165340
rect 85944 164256 85952 164320
rect 86016 164256 86032 164320
rect 86096 164256 86112 164320
rect 86176 164256 86192 164320
rect 86256 164256 86264 164320
rect 84331 164116 84397 164117
rect 84331 164052 84332 164116
rect 84396 164052 84397 164116
rect 84331 164051 84397 164052
rect 84334 154053 84394 164051
rect 85944 163232 86264 164256
rect 85944 163168 85952 163232
rect 86016 163168 86032 163232
rect 86096 163168 86112 163232
rect 86176 163168 86192 163232
rect 86256 163168 86264 163232
rect 85944 162144 86264 163168
rect 85944 162080 85952 162144
rect 86016 162080 86032 162144
rect 86096 162080 86112 162144
rect 86176 162080 86192 162144
rect 86256 162080 86264 162144
rect 85067 161804 85133 161805
rect 85067 161740 85068 161804
rect 85132 161740 85133 161804
rect 85067 161739 85133 161740
rect 84331 154052 84397 154053
rect 84331 153988 84332 154052
rect 84396 153988 84397 154052
rect 84331 153987 84397 153988
rect 84883 133108 84949 133109
rect 84883 133044 84884 133108
rect 84948 133044 84949 133108
rect 84883 133043 84949 133044
rect 83963 132428 84029 132429
rect 83963 132364 83964 132428
rect 84028 132364 84029 132428
rect 83963 132363 84029 132364
rect 83966 113933 84026 132363
rect 84515 126988 84581 126989
rect 84515 126924 84516 126988
rect 84580 126924 84581 126988
rect 84515 126923 84581 126924
rect 84518 126258 84578 126923
rect 84699 125764 84765 125765
rect 84699 125700 84700 125764
rect 84764 125700 84765 125764
rect 84699 125699 84765 125700
rect 84331 120188 84397 120189
rect 84331 120124 84332 120188
rect 84396 120124 84397 120188
rect 84331 120123 84397 120124
rect 83963 113932 84029 113933
rect 83963 113868 83964 113932
rect 84028 113868 84029 113932
rect 83963 113867 84029 113868
rect 83779 94892 83845 94893
rect 83779 94828 83780 94892
rect 83844 94828 83845 94892
rect 83779 94827 83845 94828
rect 84147 94484 84213 94485
rect 84147 94420 84148 94484
rect 84212 94420 84213 94484
rect 84147 94419 84213 94420
rect 83595 94348 83661 94349
rect 83595 94284 83596 94348
rect 83660 94284 83661 94348
rect 83595 94283 83661 94284
rect 83411 94212 83477 94213
rect 83411 94148 83412 94212
rect 83476 94148 83477 94212
rect 83411 94147 83477 94148
rect 82491 93804 82557 93805
rect 82491 93740 82492 93804
rect 82556 93740 82557 93804
rect 82491 93739 82557 93740
rect 83411 93804 83477 93805
rect 83411 93740 83412 93804
rect 83476 93740 83477 93804
rect 83411 93739 83477 93740
rect 76790 93606 77310 93666
rect 62070 93470 62275 93530
rect 63523 93470 64154 93530
rect 74608 93470 75194 93530
rect 27475 93260 27541 93261
rect 27475 93196 27476 93260
rect 27540 93196 27541 93260
rect 27475 93195 27541 93196
rect 28947 93124 29013 93125
rect 28947 93060 28948 93124
rect 29012 93060 29013 93124
rect 28947 93059 29013 93060
rect 26187 92988 26253 92989
rect 26187 92924 26188 92988
rect 26252 92924 26253 92988
rect 26187 92923 26253 92924
rect 26190 92850 26250 92923
rect 28950 92850 29010 93059
rect 32811 92852 32877 92853
rect 32811 92850 32812 92852
rect 26083 92790 26250 92850
rect 28579 92790 29010 92850
rect 32323 92790 32812 92850
rect 32811 92788 32812 92790
rect 32876 92788 32877 92852
rect 34099 92852 34165 92853
rect 34099 92850 34100 92852
rect 33571 92790 34100 92850
rect 32811 92787 32877 92788
rect 34099 92788 34100 92790
rect 34164 92788 34165 92852
rect 35203 92852 35269 92853
rect 35203 92850 35204 92852
rect 34819 92790 35204 92850
rect 34099 92787 34165 92788
rect 35203 92788 35204 92790
rect 35268 92788 35269 92852
rect 36675 92852 36741 92853
rect 36675 92850 36676 92852
rect 36067 92790 36676 92850
rect 35203 92787 35269 92788
rect 36675 92788 36676 92790
rect 36740 92788 36741 92852
rect 36675 92787 36741 92788
rect 38331 92852 38397 92853
rect 38331 92788 38332 92852
rect 38396 92850 38397 92852
rect 39987 92852 40053 92853
rect 39987 92850 39988 92852
rect 38396 92790 38563 92850
rect 39811 92790 39988 92850
rect 38396 92788 38397 92790
rect 38331 92787 38397 92788
rect 39987 92788 39988 92790
rect 40052 92788 40053 92852
rect 80099 92852 80165 92853
rect 80099 92850 80100 92852
rect 79603 92790 80100 92850
rect 39987 92787 40053 92788
rect 80099 92788 80100 92790
rect 80164 92788 80165 92852
rect 80099 92787 80165 92788
rect 4843 92444 4909 92445
rect 4843 92380 4844 92444
rect 4908 92380 4909 92444
rect 4843 92379 4909 92380
rect 4846 91578 4906 92379
rect 4846 88909 4906 91342
rect 82938 90576 83262 90618
rect 82938 90340 82982 90576
rect 83218 90340 83262 90576
rect 82938 90298 83262 90340
rect 5211 89452 5277 89453
rect 5211 89388 5212 89452
rect 5276 89388 5277 89452
rect 5211 89387 5277 89388
rect 4843 88908 4909 88909
rect 4843 88844 4844 88908
rect 4908 88844 4909 88908
rect 5214 88858 5274 89387
rect 5582 89181 5642 89302
rect 5579 89180 5645 89181
rect 5579 89116 5580 89180
rect 5644 89116 5645 89180
rect 5579 89115 5645 89116
rect 4843 88843 4909 88844
rect 82494 85576 82814 85618
rect 82494 85340 82536 85576
rect 82772 85340 82814 85576
rect 82494 85298 82814 85340
rect 82938 80576 83262 80618
rect 82938 80340 82982 80576
rect 83218 80340 83262 80576
rect 82938 80298 83262 80340
rect 82494 75576 82814 75618
rect 82494 75340 82536 75576
rect 82772 75340 82814 75576
rect 82494 75298 82814 75340
rect 82938 70576 83262 70618
rect 82938 70340 82982 70576
rect 83218 70340 83262 70576
rect 82938 70298 83262 70340
rect 82494 65576 82814 65618
rect 82494 65340 82536 65576
rect 82772 65340 82814 65576
rect 82494 65298 82814 65340
rect 82938 60576 83262 60618
rect 82938 60340 82982 60576
rect 83218 60340 83262 60576
rect 82938 60298 83262 60340
rect 82494 55576 82814 55618
rect 82494 55340 82536 55576
rect 82772 55340 82814 55576
rect 82494 55298 82814 55340
rect 82938 50576 83262 50618
rect 82938 50340 82982 50576
rect 83218 50340 83262 50576
rect 82938 50298 83262 50340
rect 83414 49330 83474 93739
rect 83779 93396 83845 93397
rect 83779 93332 83780 93396
rect 83844 93332 83845 93396
rect 83779 93331 83845 93332
rect 83595 93124 83661 93125
rect 83595 93060 83596 93124
rect 83660 93060 83661 93124
rect 83595 93059 83661 93060
rect 83598 49741 83658 93059
rect 83782 51373 83842 93331
rect 84150 55317 84210 94419
rect 84334 93669 84394 120123
rect 84515 99516 84581 99517
rect 84515 99452 84516 99516
rect 84580 99452 84581 99516
rect 84515 99451 84581 99452
rect 84518 99381 84578 99451
rect 84515 99380 84581 99381
rect 84515 99316 84516 99380
rect 84580 99316 84581 99380
rect 84515 99315 84581 99316
rect 84331 93668 84397 93669
rect 84331 93604 84332 93668
rect 84396 93604 84397 93668
rect 84331 93603 84397 93604
rect 84702 92258 84762 125699
rect 84886 96933 84946 133043
rect 84883 96932 84949 96933
rect 84883 96868 84884 96932
rect 84948 96868 84949 96932
rect 84883 96867 84949 96868
rect 85070 93669 85130 161739
rect 85944 161056 86264 162080
rect 86355 161940 86421 161941
rect 86355 161876 86356 161940
rect 86420 161876 86421 161940
rect 86355 161875 86421 161876
rect 85944 160992 85952 161056
rect 86016 160992 86032 161056
rect 86096 160992 86112 161056
rect 86176 160992 86192 161056
rect 86256 160992 86264 161056
rect 85944 159968 86264 160992
rect 85944 159904 85952 159968
rect 86016 159904 86032 159968
rect 86096 159904 86112 159968
rect 86176 159904 86192 159968
rect 86256 159904 86264 159968
rect 85944 158880 86264 159904
rect 85944 158816 85952 158880
rect 86016 158816 86032 158880
rect 86096 158816 86112 158880
rect 86176 158816 86192 158880
rect 86256 158816 86264 158880
rect 85944 157792 86264 158816
rect 85944 157728 85952 157792
rect 86016 157728 86032 157792
rect 86096 157728 86112 157792
rect 86176 157728 86192 157792
rect 86256 157728 86264 157792
rect 85944 156704 86264 157728
rect 85944 156640 85952 156704
rect 86016 156640 86032 156704
rect 86096 156640 86112 156704
rect 86176 156640 86192 156704
rect 86256 156640 86264 156704
rect 85803 156364 85869 156365
rect 85803 156300 85804 156364
rect 85868 156300 85869 156364
rect 85803 156299 85869 156300
rect 85251 130388 85317 130389
rect 85251 130324 85252 130388
rect 85316 130324 85317 130388
rect 85251 130323 85317 130324
rect 85254 97341 85314 130323
rect 85619 108628 85685 108629
rect 85619 108564 85620 108628
rect 85684 108564 85685 108628
rect 85619 108563 85685 108564
rect 85435 99516 85501 99517
rect 85435 99452 85436 99516
rect 85500 99452 85501 99516
rect 85435 99451 85501 99452
rect 85438 99109 85498 99451
rect 85435 99108 85501 99109
rect 85435 99044 85436 99108
rect 85500 99044 85501 99108
rect 85435 99043 85501 99044
rect 85251 97340 85317 97341
rect 85251 97276 85252 97340
rect 85316 97276 85317 97340
rect 85251 97275 85317 97276
rect 85622 95301 85682 108563
rect 85806 96525 85866 156299
rect 85944 155616 86264 156640
rect 85944 155552 85952 155616
rect 86016 155576 86032 155616
rect 86096 155576 86112 155616
rect 86176 155576 86192 155616
rect 86256 155552 86264 155616
rect 85944 155340 85986 155552
rect 86222 155340 86264 155552
rect 85944 154528 86264 155340
rect 85944 154464 85952 154528
rect 86016 154464 86032 154528
rect 86096 154464 86112 154528
rect 86176 154464 86192 154528
rect 86256 154464 86264 154528
rect 85944 153440 86264 154464
rect 85944 153376 85952 153440
rect 86016 153376 86032 153440
rect 86096 153376 86112 153440
rect 86176 153376 86192 153440
rect 86256 153376 86264 153440
rect 85944 152352 86264 153376
rect 85944 152288 85952 152352
rect 86016 152288 86032 152352
rect 86096 152288 86112 152352
rect 86176 152288 86192 152352
rect 86256 152288 86264 152352
rect 85944 151264 86264 152288
rect 85944 151200 85952 151264
rect 86016 151200 86032 151264
rect 86096 151200 86112 151264
rect 86176 151200 86192 151264
rect 86256 151200 86264 151264
rect 85944 150176 86264 151200
rect 85944 150112 85952 150176
rect 86016 150112 86032 150176
rect 86096 150112 86112 150176
rect 86176 150112 86192 150176
rect 86256 150112 86264 150176
rect 85944 149088 86264 150112
rect 85944 149024 85952 149088
rect 86016 149024 86032 149088
rect 86096 149024 86112 149088
rect 86176 149024 86192 149088
rect 86256 149024 86264 149088
rect 85944 148000 86264 149024
rect 85944 147936 85952 148000
rect 86016 147936 86032 148000
rect 86096 147936 86112 148000
rect 86176 147936 86192 148000
rect 86256 147936 86264 148000
rect 85944 146912 86264 147936
rect 85944 146848 85952 146912
rect 86016 146848 86032 146912
rect 86096 146848 86112 146912
rect 86176 146848 86192 146912
rect 86256 146848 86264 146912
rect 85944 145824 86264 146848
rect 85944 145760 85952 145824
rect 86016 145760 86032 145824
rect 86096 145760 86112 145824
rect 86176 145760 86192 145824
rect 86256 145760 86264 145824
rect 85944 145576 86264 145760
rect 85944 145340 85986 145576
rect 86222 145340 86264 145576
rect 85944 144736 86264 145340
rect 85944 144672 85952 144736
rect 86016 144672 86032 144736
rect 86096 144672 86112 144736
rect 86176 144672 86192 144736
rect 86256 144672 86264 144736
rect 85944 143648 86264 144672
rect 85944 143584 85952 143648
rect 86016 143584 86032 143648
rect 86096 143584 86112 143648
rect 86176 143584 86192 143648
rect 86256 143584 86264 143648
rect 85944 142560 86264 143584
rect 85944 142496 85952 142560
rect 86016 142496 86032 142560
rect 86096 142496 86112 142560
rect 86176 142496 86192 142560
rect 86256 142496 86264 142560
rect 85944 141472 86264 142496
rect 85944 141408 85952 141472
rect 86016 141408 86032 141472
rect 86096 141408 86112 141472
rect 86176 141408 86192 141472
rect 86256 141408 86264 141472
rect 85944 140384 86264 141408
rect 85944 140320 85952 140384
rect 86016 140320 86032 140384
rect 86096 140320 86112 140384
rect 86176 140320 86192 140384
rect 86256 140320 86264 140384
rect 85944 139296 86264 140320
rect 85944 139232 85952 139296
rect 86016 139232 86032 139296
rect 86096 139232 86112 139296
rect 86176 139232 86192 139296
rect 86256 139232 86264 139296
rect 85944 138208 86264 139232
rect 85944 138144 85952 138208
rect 86016 138144 86032 138208
rect 86096 138144 86112 138208
rect 86176 138144 86192 138208
rect 86256 138144 86264 138208
rect 85944 137120 86264 138144
rect 85944 137056 85952 137120
rect 86016 137056 86032 137120
rect 86096 137056 86112 137120
rect 86176 137056 86192 137120
rect 86256 137056 86264 137120
rect 85944 136032 86264 137056
rect 85944 135968 85952 136032
rect 86016 135968 86032 136032
rect 86096 135968 86112 136032
rect 86176 135968 86192 136032
rect 86256 135968 86264 136032
rect 85944 135576 86264 135968
rect 85944 135340 85986 135576
rect 86222 135340 86264 135576
rect 85944 134944 86264 135340
rect 85944 134880 85952 134944
rect 86016 134880 86032 134944
rect 86096 134880 86112 134944
rect 86176 134880 86192 134944
rect 86256 134880 86264 134944
rect 85944 133856 86264 134880
rect 85944 133792 85952 133856
rect 86016 133792 86032 133856
rect 86096 133792 86112 133856
rect 86176 133792 86192 133856
rect 86256 133792 86264 133856
rect 85944 132768 86264 133792
rect 85944 132704 85952 132768
rect 86016 132704 86032 132768
rect 86096 132704 86112 132768
rect 86176 132704 86192 132768
rect 86256 132704 86264 132768
rect 85944 131680 86264 132704
rect 85944 131616 85952 131680
rect 86016 131616 86032 131680
rect 86096 131616 86112 131680
rect 86176 131616 86192 131680
rect 86256 131616 86264 131680
rect 85944 130592 86264 131616
rect 85944 130528 85952 130592
rect 86016 130528 86032 130592
rect 86096 130528 86112 130592
rect 86176 130528 86192 130592
rect 86256 130528 86264 130592
rect 85944 129504 86264 130528
rect 85944 129440 85952 129504
rect 86016 129440 86032 129504
rect 86096 129440 86112 129504
rect 86176 129440 86192 129504
rect 86256 129440 86264 129504
rect 85944 128416 86264 129440
rect 85944 128352 85952 128416
rect 86016 128352 86032 128416
rect 86096 128352 86112 128416
rect 86176 128352 86192 128416
rect 86256 128352 86264 128416
rect 85944 127328 86264 128352
rect 85944 127264 85952 127328
rect 86016 127264 86032 127328
rect 86096 127264 86112 127328
rect 86176 127264 86192 127328
rect 86256 127264 86264 127328
rect 85944 126240 86264 127264
rect 85944 126176 85952 126240
rect 86016 126176 86032 126240
rect 86096 126176 86112 126240
rect 86176 126176 86192 126240
rect 86256 126176 86264 126240
rect 85944 125576 86264 126176
rect 85944 125340 85986 125576
rect 86222 125340 86264 125576
rect 85944 125152 86264 125340
rect 85944 125088 85952 125152
rect 86016 125088 86032 125152
rect 86096 125088 86112 125152
rect 86176 125088 86192 125152
rect 86256 125088 86264 125152
rect 85944 124064 86264 125088
rect 85944 124000 85952 124064
rect 86016 124000 86032 124064
rect 86096 124000 86112 124064
rect 86176 124000 86192 124064
rect 86256 124000 86264 124064
rect 85944 122976 86264 124000
rect 85944 122912 85952 122976
rect 86016 122912 86032 122976
rect 86096 122912 86112 122976
rect 86176 122912 86192 122976
rect 86256 122912 86264 122976
rect 85944 121888 86264 122912
rect 85944 121824 85952 121888
rect 86016 121824 86032 121888
rect 86096 121824 86112 121888
rect 86176 121824 86192 121888
rect 86256 121824 86264 121888
rect 85944 120800 86264 121824
rect 85944 120736 85952 120800
rect 86016 120736 86032 120800
rect 86096 120736 86112 120800
rect 86176 120736 86192 120800
rect 86256 120736 86264 120800
rect 85944 119712 86264 120736
rect 85944 119648 85952 119712
rect 86016 119648 86032 119712
rect 86096 119648 86112 119712
rect 86176 119648 86192 119712
rect 86256 119648 86264 119712
rect 85944 118624 86264 119648
rect 85944 118560 85952 118624
rect 86016 118560 86032 118624
rect 86096 118560 86112 118624
rect 86176 118560 86192 118624
rect 86256 118560 86264 118624
rect 85944 117536 86264 118560
rect 85944 117472 85952 117536
rect 86016 117472 86032 117536
rect 86096 117472 86112 117536
rect 86176 117472 86192 117536
rect 86256 117472 86264 117536
rect 85944 116448 86264 117472
rect 85944 116384 85952 116448
rect 86016 116384 86032 116448
rect 86096 116384 86112 116448
rect 86176 116384 86192 116448
rect 86256 116384 86264 116448
rect 85944 115576 86264 116384
rect 85944 115360 85986 115576
rect 86222 115360 86264 115576
rect 85944 115296 85952 115360
rect 86016 115296 86032 115340
rect 86096 115296 86112 115340
rect 86176 115296 86192 115340
rect 86256 115296 86264 115360
rect 85944 114272 86264 115296
rect 85944 114208 85952 114272
rect 86016 114208 86032 114272
rect 86096 114208 86112 114272
rect 86176 114208 86192 114272
rect 86256 114208 86264 114272
rect 85944 113184 86264 114208
rect 85944 113120 85952 113184
rect 86016 113120 86032 113184
rect 86096 113120 86112 113184
rect 86176 113120 86192 113184
rect 86256 113120 86264 113184
rect 85944 112096 86264 113120
rect 85944 112032 85952 112096
rect 86016 112032 86032 112096
rect 86096 112032 86112 112096
rect 86176 112032 86192 112096
rect 86256 112032 86264 112096
rect 85944 111008 86264 112032
rect 85944 110944 85952 111008
rect 86016 110944 86032 111008
rect 86096 110944 86112 111008
rect 86176 110944 86192 111008
rect 86256 110944 86264 111008
rect 85944 109920 86264 110944
rect 85944 109856 85952 109920
rect 86016 109856 86032 109920
rect 86096 109856 86112 109920
rect 86176 109856 86192 109920
rect 86256 109856 86264 109920
rect 85944 108832 86264 109856
rect 85944 108768 85952 108832
rect 86016 108768 86032 108832
rect 86096 108768 86112 108832
rect 86176 108768 86192 108832
rect 86256 108768 86264 108832
rect 85944 107744 86264 108768
rect 85944 107680 85952 107744
rect 86016 107680 86032 107744
rect 86096 107680 86112 107744
rect 86176 107680 86192 107744
rect 86256 107680 86264 107744
rect 85944 106656 86264 107680
rect 85944 106592 85952 106656
rect 86016 106592 86032 106656
rect 86096 106592 86112 106656
rect 86176 106592 86192 106656
rect 86256 106592 86264 106656
rect 85944 105576 86264 106592
rect 85944 105568 85986 105576
rect 86222 105568 86264 105576
rect 85944 105504 85952 105568
rect 86256 105504 86264 105568
rect 85944 105340 85986 105504
rect 86222 105340 86264 105504
rect 85944 104480 86264 105340
rect 85944 104416 85952 104480
rect 86016 104416 86032 104480
rect 86096 104416 86112 104480
rect 86176 104416 86192 104480
rect 86256 104416 86264 104480
rect 85944 103392 86264 104416
rect 85944 103328 85952 103392
rect 86016 103328 86032 103392
rect 86096 103328 86112 103392
rect 86176 103328 86192 103392
rect 86256 103328 86264 103392
rect 85944 102304 86264 103328
rect 85944 102240 85952 102304
rect 86016 102240 86032 102304
rect 86096 102240 86112 102304
rect 86176 102240 86192 102304
rect 86256 102240 86264 102304
rect 85944 101216 86264 102240
rect 85944 101152 85952 101216
rect 86016 101152 86032 101216
rect 86096 101152 86112 101216
rect 86176 101152 86192 101216
rect 86256 101152 86264 101216
rect 85944 100128 86264 101152
rect 85944 100064 85952 100128
rect 86016 100064 86032 100128
rect 86096 100064 86112 100128
rect 86176 100064 86192 100128
rect 86256 100064 86264 100128
rect 85944 99040 86264 100064
rect 85944 98976 85952 99040
rect 86016 98976 86032 99040
rect 86096 98976 86112 99040
rect 86176 98976 86192 99040
rect 86256 98976 86264 99040
rect 85944 97952 86264 98976
rect 85944 97888 85952 97952
rect 86016 97888 86032 97952
rect 86096 97888 86112 97952
rect 86176 97888 86192 97952
rect 86256 97888 86264 97952
rect 85944 96864 86264 97888
rect 85944 96800 85952 96864
rect 86016 96800 86032 96864
rect 86096 96800 86112 96864
rect 86176 96800 86192 96864
rect 86256 96800 86264 96864
rect 85803 96524 85869 96525
rect 85803 96460 85804 96524
rect 85868 96460 85869 96524
rect 85803 96459 85869 96460
rect 85944 95776 86264 96800
rect 85944 95712 85952 95776
rect 86016 95712 86032 95776
rect 86096 95712 86112 95776
rect 86176 95712 86192 95776
rect 86256 95712 86264 95776
rect 85944 95576 86264 95712
rect 85944 95340 85986 95576
rect 86222 95340 86264 95576
rect 85619 95300 85685 95301
rect 85619 95236 85620 95300
rect 85684 95236 85685 95300
rect 85619 95235 85685 95236
rect 85944 94688 86264 95340
rect 85944 94624 85952 94688
rect 86016 94624 86032 94688
rect 86096 94624 86112 94688
rect 86176 94624 86192 94688
rect 86256 94624 86264 94688
rect 85067 93668 85133 93669
rect 85067 93604 85068 93668
rect 85132 93604 85133 93668
rect 85067 93603 85133 93604
rect 85944 93600 86264 94624
rect 86358 93941 86418 161875
rect 86539 153780 86605 153781
rect 86539 153716 86540 153780
rect 86604 153716 86605 153780
rect 86539 153715 86605 153716
rect 86542 94077 86602 153715
rect 86907 147660 86973 147661
rect 86907 147596 86908 147660
rect 86972 147596 86973 147660
rect 86907 147595 86973 147596
rect 86910 122637 86970 147595
rect 86907 122636 86973 122637
rect 86907 122572 86908 122636
rect 86972 122572 86973 122636
rect 86907 122571 86973 122572
rect 86907 122364 86973 122365
rect 86907 122300 86908 122364
rect 86972 122300 86973 122364
rect 86907 122299 86973 122300
rect 86910 118557 86970 122299
rect 86907 118556 86973 118557
rect 86907 118492 86908 118556
rect 86972 118492 86973 118556
rect 86907 118491 86973 118492
rect 86907 109172 86973 109173
rect 86907 109108 86908 109172
rect 86972 109108 86973 109172
rect 86907 109107 86973 109108
rect 86910 108765 86970 109107
rect 86907 108764 86973 108765
rect 86907 108700 86908 108764
rect 86972 108700 86973 108764
rect 86907 108699 86973 108700
rect 86723 103732 86789 103733
rect 86723 103668 86724 103732
rect 86788 103668 86789 103732
rect 86723 103667 86789 103668
rect 86726 99381 86786 103667
rect 86907 102644 86973 102645
rect 86907 102580 86908 102644
rect 86972 102580 86973 102644
rect 86907 102579 86973 102580
rect 86910 99517 86970 102579
rect 86907 99516 86973 99517
rect 86907 99452 86908 99516
rect 86972 99452 86973 99516
rect 86907 99451 86973 99452
rect 86723 99380 86789 99381
rect 86723 99316 86724 99380
rect 86788 99316 86789 99380
rect 86723 99315 86789 99316
rect 87094 97018 87154 182547
rect 87275 179212 87341 179213
rect 87275 179148 87276 179212
rect 87340 179148 87341 179212
rect 87275 179147 87341 179148
rect 87278 97205 87338 179147
rect 87275 97204 87341 97205
rect 87275 97140 87276 97204
rect 87340 97140 87341 97204
rect 87275 97139 87341 97140
rect 87462 97069 87522 184043
rect 87944 183360 88264 184384
rect 87944 183296 87952 183360
rect 88016 183296 88032 183360
rect 88096 183296 88112 183360
rect 88176 183296 88192 183360
rect 88256 183296 88264 183360
rect 87944 182272 88264 183296
rect 87944 182208 87952 182272
rect 88016 182208 88032 182272
rect 88096 182208 88112 182272
rect 88176 182208 88192 182272
rect 88256 182208 88264 182272
rect 87944 181184 88264 182208
rect 87944 181120 87952 181184
rect 88016 181120 88032 181184
rect 88096 181120 88112 181184
rect 88176 181120 88192 181184
rect 88256 181120 88264 181184
rect 87944 180576 88264 181120
rect 87643 180436 87709 180437
rect 87643 180372 87644 180436
rect 87708 180372 87709 180436
rect 87643 180371 87709 180372
rect 87459 97068 87525 97069
rect 87459 97004 87460 97068
rect 87524 97004 87525 97068
rect 87459 97003 87525 97004
rect 87646 96797 87706 180371
rect 87944 180340 87986 180576
rect 88222 180340 88264 180576
rect 87944 180096 88264 180340
rect 87944 180032 87952 180096
rect 88016 180032 88032 180096
rect 88096 180032 88112 180096
rect 88176 180032 88192 180096
rect 88256 180032 88264 180096
rect 87944 179008 88264 180032
rect 87944 178944 87952 179008
rect 88016 178944 88032 179008
rect 88096 178944 88112 179008
rect 88176 178944 88192 179008
rect 88256 178944 88264 179008
rect 87944 177920 88264 178944
rect 87944 177856 87952 177920
rect 88016 177856 88032 177920
rect 88096 177856 88112 177920
rect 88176 177856 88192 177920
rect 88256 177856 88264 177920
rect 87944 176832 88264 177856
rect 87944 176768 87952 176832
rect 88016 176768 88032 176832
rect 88096 176768 88112 176832
rect 88176 176768 88192 176832
rect 88256 176768 88264 176832
rect 87944 175744 88264 176768
rect 87944 175680 87952 175744
rect 88016 175680 88032 175744
rect 88096 175680 88112 175744
rect 88176 175680 88192 175744
rect 88256 175680 88264 175744
rect 87944 174656 88264 175680
rect 87944 174592 87952 174656
rect 88016 174592 88032 174656
rect 88096 174592 88112 174656
rect 88176 174592 88192 174656
rect 88256 174592 88264 174656
rect 87944 173568 88264 174592
rect 87944 173504 87952 173568
rect 88016 173504 88032 173568
rect 88096 173504 88112 173568
rect 88176 173504 88192 173568
rect 88256 173504 88264 173568
rect 87944 172480 88264 173504
rect 87944 172416 87952 172480
rect 88016 172416 88032 172480
rect 88096 172416 88112 172480
rect 88176 172416 88192 172480
rect 88256 172416 88264 172480
rect 87944 171392 88264 172416
rect 87944 171328 87952 171392
rect 88016 171328 88032 171392
rect 88096 171328 88112 171392
rect 88176 171328 88192 171392
rect 88256 171328 88264 171392
rect 87944 170576 88264 171328
rect 87944 170340 87986 170576
rect 88222 170340 88264 170576
rect 87944 170304 88264 170340
rect 87944 170240 87952 170304
rect 88016 170240 88032 170304
rect 88096 170240 88112 170304
rect 88176 170240 88192 170304
rect 88256 170240 88264 170304
rect 87944 169216 88264 170240
rect 87944 169152 87952 169216
rect 88016 169152 88032 169216
rect 88096 169152 88112 169216
rect 88176 169152 88192 169216
rect 88256 169152 88264 169216
rect 87944 168128 88264 169152
rect 87944 168064 87952 168128
rect 88016 168064 88032 168128
rect 88096 168064 88112 168128
rect 88176 168064 88192 168128
rect 88256 168064 88264 168128
rect 87944 167040 88264 168064
rect 87944 166976 87952 167040
rect 88016 166976 88032 167040
rect 88096 166976 88112 167040
rect 88176 166976 88192 167040
rect 88256 166976 88264 167040
rect 87944 165952 88264 166976
rect 87944 165888 87952 165952
rect 88016 165888 88032 165952
rect 88096 165888 88112 165952
rect 88176 165888 88192 165952
rect 88256 165888 88264 165952
rect 87944 164864 88264 165888
rect 87944 164800 87952 164864
rect 88016 164800 88032 164864
rect 88096 164800 88112 164864
rect 88176 164800 88192 164864
rect 88256 164800 88264 164864
rect 87944 163776 88264 164800
rect 87944 163712 87952 163776
rect 88016 163712 88032 163776
rect 88096 163712 88112 163776
rect 88176 163712 88192 163776
rect 88256 163712 88264 163776
rect 87944 162688 88264 163712
rect 87944 162624 87952 162688
rect 88016 162624 88032 162688
rect 88096 162624 88112 162688
rect 88176 162624 88192 162688
rect 88256 162624 88264 162688
rect 87944 161600 88264 162624
rect 87944 161536 87952 161600
rect 88016 161536 88032 161600
rect 88096 161536 88112 161600
rect 88176 161536 88192 161600
rect 88256 161536 88264 161600
rect 87944 160576 88264 161536
rect 87944 160512 87986 160576
rect 88222 160512 88264 160576
rect 87944 160448 87952 160512
rect 88256 160448 88264 160512
rect 87944 160340 87986 160448
rect 88222 160340 88264 160448
rect 87944 159424 88264 160340
rect 87944 159360 87952 159424
rect 88016 159360 88032 159424
rect 88096 159360 88112 159424
rect 88176 159360 88192 159424
rect 88256 159360 88264 159424
rect 87944 158336 88264 159360
rect 87944 158272 87952 158336
rect 88016 158272 88032 158336
rect 88096 158272 88112 158336
rect 88176 158272 88192 158336
rect 88256 158272 88264 158336
rect 87944 157248 88264 158272
rect 87944 157184 87952 157248
rect 88016 157184 88032 157248
rect 88096 157184 88112 157248
rect 88176 157184 88192 157248
rect 88256 157184 88264 157248
rect 87944 156160 88264 157184
rect 87944 156096 87952 156160
rect 88016 156096 88032 156160
rect 88096 156096 88112 156160
rect 88176 156096 88192 156160
rect 88256 156096 88264 156160
rect 87944 155072 88264 156096
rect 87944 155008 87952 155072
rect 88016 155008 88032 155072
rect 88096 155008 88112 155072
rect 88176 155008 88192 155072
rect 88256 155008 88264 155072
rect 87944 153984 88264 155008
rect 87944 153920 87952 153984
rect 88016 153920 88032 153984
rect 88096 153920 88112 153984
rect 88176 153920 88192 153984
rect 88256 153920 88264 153984
rect 87944 152896 88264 153920
rect 87944 152832 87952 152896
rect 88016 152832 88032 152896
rect 88096 152832 88112 152896
rect 88176 152832 88192 152896
rect 88256 152832 88264 152896
rect 87944 151808 88264 152832
rect 87944 151744 87952 151808
rect 88016 151744 88032 151808
rect 88096 151744 88112 151808
rect 88176 151744 88192 151808
rect 88256 151744 88264 151808
rect 87944 150720 88264 151744
rect 87944 150656 87952 150720
rect 88016 150656 88032 150720
rect 88096 150656 88112 150720
rect 88176 150656 88192 150720
rect 88256 150656 88264 150720
rect 87944 150576 88264 150656
rect 87944 150340 87986 150576
rect 88222 150340 88264 150576
rect 87944 149632 88264 150340
rect 87944 149568 87952 149632
rect 88016 149568 88032 149632
rect 88096 149568 88112 149632
rect 88176 149568 88192 149632
rect 88256 149568 88264 149632
rect 87944 148544 88264 149568
rect 87944 148480 87952 148544
rect 88016 148480 88032 148544
rect 88096 148480 88112 148544
rect 88176 148480 88192 148544
rect 88256 148480 88264 148544
rect 87944 147456 88264 148480
rect 87944 147392 87952 147456
rect 88016 147392 88032 147456
rect 88096 147392 88112 147456
rect 88176 147392 88192 147456
rect 88256 147392 88264 147456
rect 87944 146368 88264 147392
rect 87944 146304 87952 146368
rect 88016 146304 88032 146368
rect 88096 146304 88112 146368
rect 88176 146304 88192 146368
rect 88256 146304 88264 146368
rect 87944 145280 88264 146304
rect 87944 145216 87952 145280
rect 88016 145216 88032 145280
rect 88096 145216 88112 145280
rect 88176 145216 88192 145280
rect 88256 145216 88264 145280
rect 87944 144192 88264 145216
rect 87944 144128 87952 144192
rect 88016 144128 88032 144192
rect 88096 144128 88112 144192
rect 88176 144128 88192 144192
rect 88256 144128 88264 144192
rect 87944 143104 88264 144128
rect 87944 143040 87952 143104
rect 88016 143040 88032 143104
rect 88096 143040 88112 143104
rect 88176 143040 88192 143104
rect 88256 143040 88264 143104
rect 87944 142016 88264 143040
rect 87944 141952 87952 142016
rect 88016 141952 88032 142016
rect 88096 141952 88112 142016
rect 88176 141952 88192 142016
rect 88256 141952 88264 142016
rect 87944 140928 88264 141952
rect 87944 140864 87952 140928
rect 88016 140864 88032 140928
rect 88096 140864 88112 140928
rect 88176 140864 88192 140928
rect 88256 140864 88264 140928
rect 87944 140576 88264 140864
rect 87944 140340 87986 140576
rect 88222 140340 88264 140576
rect 87944 139840 88264 140340
rect 87944 139776 87952 139840
rect 88016 139776 88032 139840
rect 88096 139776 88112 139840
rect 88176 139776 88192 139840
rect 88256 139776 88264 139840
rect 87944 138752 88264 139776
rect 87944 138688 87952 138752
rect 88016 138688 88032 138752
rect 88096 138688 88112 138752
rect 88176 138688 88192 138752
rect 88256 138688 88264 138752
rect 87944 137664 88264 138688
rect 87944 137600 87952 137664
rect 88016 137600 88032 137664
rect 88096 137600 88112 137664
rect 88176 137600 88192 137664
rect 88256 137600 88264 137664
rect 87944 136576 88264 137600
rect 87944 136512 87952 136576
rect 88016 136512 88032 136576
rect 88096 136512 88112 136576
rect 88176 136512 88192 136576
rect 88256 136512 88264 136576
rect 87944 135488 88264 136512
rect 87944 135424 87952 135488
rect 88016 135424 88032 135488
rect 88096 135424 88112 135488
rect 88176 135424 88192 135488
rect 88256 135424 88264 135488
rect 87944 134400 88264 135424
rect 87944 134336 87952 134400
rect 88016 134336 88032 134400
rect 88096 134336 88112 134400
rect 88176 134336 88192 134400
rect 88256 134336 88264 134400
rect 87944 133312 88264 134336
rect 87944 133248 87952 133312
rect 88016 133248 88032 133312
rect 88096 133248 88112 133312
rect 88176 133248 88192 133312
rect 88256 133248 88264 133312
rect 87944 132224 88264 133248
rect 87944 132160 87952 132224
rect 88016 132160 88032 132224
rect 88096 132160 88112 132224
rect 88176 132160 88192 132224
rect 88256 132160 88264 132224
rect 87944 131136 88264 132160
rect 87944 131072 87952 131136
rect 88016 131072 88032 131136
rect 88096 131072 88112 131136
rect 88176 131072 88192 131136
rect 88256 131072 88264 131136
rect 87944 130576 88264 131072
rect 87944 130340 87986 130576
rect 88222 130340 88264 130576
rect 87944 130048 88264 130340
rect 87944 129984 87952 130048
rect 88016 129984 88032 130048
rect 88096 129984 88112 130048
rect 88176 129984 88192 130048
rect 88256 129984 88264 130048
rect 87944 128960 88264 129984
rect 87944 128896 87952 128960
rect 88016 128896 88032 128960
rect 88096 128896 88112 128960
rect 88176 128896 88192 128960
rect 88256 128896 88264 128960
rect 87944 127872 88264 128896
rect 87944 127808 87952 127872
rect 88016 127808 88032 127872
rect 88096 127808 88112 127872
rect 88176 127808 88192 127872
rect 88256 127808 88264 127872
rect 87944 126784 88264 127808
rect 87944 126720 87952 126784
rect 88016 126720 88032 126784
rect 88096 126720 88112 126784
rect 88176 126720 88192 126784
rect 88256 126720 88264 126784
rect 87944 125696 88264 126720
rect 87944 125632 87952 125696
rect 88016 125632 88032 125696
rect 88096 125632 88112 125696
rect 88176 125632 88192 125696
rect 88256 125632 88264 125696
rect 87944 124608 88264 125632
rect 87944 124544 87952 124608
rect 88016 124544 88032 124608
rect 88096 124544 88112 124608
rect 88176 124544 88192 124608
rect 88256 124544 88264 124608
rect 87944 123520 88264 124544
rect 87944 123456 87952 123520
rect 88016 123456 88032 123520
rect 88096 123456 88112 123520
rect 88176 123456 88192 123520
rect 88256 123456 88264 123520
rect 87944 122432 88264 123456
rect 87944 122368 87952 122432
rect 88016 122368 88032 122432
rect 88096 122368 88112 122432
rect 88176 122368 88192 122432
rect 88256 122368 88264 122432
rect 87944 121344 88264 122368
rect 87944 121280 87952 121344
rect 88016 121280 88032 121344
rect 88096 121280 88112 121344
rect 88176 121280 88192 121344
rect 88256 121280 88264 121344
rect 87944 120576 88264 121280
rect 87944 120340 87986 120576
rect 88222 120340 88264 120576
rect 87944 120256 88264 120340
rect 87944 120192 87952 120256
rect 88016 120192 88032 120256
rect 88096 120192 88112 120256
rect 88176 120192 88192 120256
rect 88256 120192 88264 120256
rect 87944 119168 88264 120192
rect 87944 119104 87952 119168
rect 88016 119104 88032 119168
rect 88096 119104 88112 119168
rect 88176 119104 88192 119168
rect 88256 119104 88264 119168
rect 87944 118080 88264 119104
rect 87944 118016 87952 118080
rect 88016 118016 88032 118080
rect 88096 118016 88112 118080
rect 88176 118016 88192 118080
rect 88256 118016 88264 118080
rect 87944 116992 88264 118016
rect 87944 116928 87952 116992
rect 88016 116928 88032 116992
rect 88096 116928 88112 116992
rect 88176 116928 88192 116992
rect 88256 116928 88264 116992
rect 87944 115904 88264 116928
rect 87944 115840 87952 115904
rect 88016 115840 88032 115904
rect 88096 115840 88112 115904
rect 88176 115840 88192 115904
rect 88256 115840 88264 115904
rect 87944 114816 88264 115840
rect 87944 114752 87952 114816
rect 88016 114752 88032 114816
rect 88096 114752 88112 114816
rect 88176 114752 88192 114816
rect 88256 114752 88264 114816
rect 87944 113728 88264 114752
rect 87944 113664 87952 113728
rect 88016 113664 88032 113728
rect 88096 113664 88112 113728
rect 88176 113664 88192 113728
rect 88256 113664 88264 113728
rect 87944 112640 88264 113664
rect 87944 112576 87952 112640
rect 88016 112576 88032 112640
rect 88096 112576 88112 112640
rect 88176 112576 88192 112640
rect 88256 112576 88264 112640
rect 87944 111552 88264 112576
rect 87944 111488 87952 111552
rect 88016 111488 88032 111552
rect 88096 111488 88112 111552
rect 88176 111488 88192 111552
rect 88256 111488 88264 111552
rect 87944 110576 88264 111488
rect 87944 110464 87986 110576
rect 88222 110464 88264 110576
rect 87944 110400 87952 110464
rect 88256 110400 88264 110464
rect 87944 110340 87986 110400
rect 88222 110340 88264 110400
rect 87944 109376 88264 110340
rect 87944 109312 87952 109376
rect 88016 109312 88032 109376
rect 88096 109312 88112 109376
rect 88176 109312 88192 109376
rect 88256 109312 88264 109376
rect 87944 108288 88264 109312
rect 87944 108224 87952 108288
rect 88016 108224 88032 108288
rect 88096 108224 88112 108288
rect 88176 108224 88192 108288
rect 88256 108224 88264 108288
rect 87944 107200 88264 108224
rect 87944 107136 87952 107200
rect 88016 107136 88032 107200
rect 88096 107136 88112 107200
rect 88176 107136 88192 107200
rect 88256 107136 88264 107200
rect 87944 106112 88264 107136
rect 87944 106048 87952 106112
rect 88016 106048 88032 106112
rect 88096 106048 88112 106112
rect 88176 106048 88192 106112
rect 88256 106048 88264 106112
rect 87944 105024 88264 106048
rect 87944 104960 87952 105024
rect 88016 104960 88032 105024
rect 88096 104960 88112 105024
rect 88176 104960 88192 105024
rect 88256 104960 88264 105024
rect 87944 103936 88264 104960
rect 87944 103872 87952 103936
rect 88016 103872 88032 103936
rect 88096 103872 88112 103936
rect 88176 103872 88192 103936
rect 88256 103872 88264 103936
rect 87944 102848 88264 103872
rect 87944 102784 87952 102848
rect 88016 102784 88032 102848
rect 88096 102784 88112 102848
rect 88176 102784 88192 102848
rect 88256 102784 88264 102848
rect 87944 101760 88264 102784
rect 87944 101696 87952 101760
rect 88016 101696 88032 101760
rect 88096 101696 88112 101760
rect 88176 101696 88192 101760
rect 88256 101696 88264 101760
rect 87944 100672 88264 101696
rect 87944 100608 87952 100672
rect 88016 100608 88032 100672
rect 88096 100608 88112 100672
rect 88176 100608 88192 100672
rect 88256 100608 88264 100672
rect 87944 100576 88264 100608
rect 87944 100340 87986 100576
rect 88222 100340 88264 100576
rect 87944 99584 88264 100340
rect 87944 99520 87952 99584
rect 88016 99520 88032 99584
rect 88096 99520 88112 99584
rect 88176 99520 88192 99584
rect 88256 99520 88264 99584
rect 87944 98496 88264 99520
rect 87944 98432 87952 98496
rect 88016 98432 88032 98496
rect 88096 98432 88112 98496
rect 88176 98432 88192 98496
rect 88256 98432 88264 98496
rect 87944 97408 88264 98432
rect 87944 97344 87952 97408
rect 88016 97344 88032 97408
rect 88096 97344 88112 97408
rect 88176 97344 88192 97408
rect 88256 97344 88264 97408
rect 87643 96796 87709 96797
rect 87643 96732 87644 96796
rect 87708 96732 87709 96796
rect 87643 96731 87709 96732
rect 87944 96320 88264 97344
rect 87944 96256 87952 96320
rect 88016 96256 88032 96320
rect 88096 96256 88112 96320
rect 88176 96256 88192 96320
rect 88256 96256 88264 96320
rect 87944 95232 88264 96256
rect 87944 95168 87952 95232
rect 88016 95168 88032 95232
rect 88096 95168 88112 95232
rect 88176 95168 88192 95232
rect 88256 95168 88264 95232
rect 87944 94144 88264 95168
rect 88382 94890 88442 185267
rect 88750 96338 88810 186491
rect 88934 96930 88994 190163
rect 89115 189004 89181 189005
rect 89115 188940 89116 189004
rect 89180 188940 89181 189004
rect 89115 188939 89181 188940
rect 89118 98157 89178 188939
rect 89115 98156 89181 98157
rect 89115 98092 89116 98156
rect 89180 98092 89181 98156
rect 89115 98091 89181 98092
rect 89302 97885 89362 191387
rect 89944 189344 90264 189360
rect 89944 189280 89952 189344
rect 90016 189280 90032 189344
rect 90096 189280 90112 189344
rect 90176 189280 90192 189344
rect 90256 189280 90264 189344
rect 89944 188256 90264 189280
rect 89944 188192 89952 188256
rect 90016 188192 90032 188256
rect 90096 188192 90112 188256
rect 90176 188192 90192 188256
rect 90256 188192 90264 188256
rect 89483 187780 89549 187781
rect 89483 187716 89484 187780
rect 89548 187716 89549 187780
rect 89483 187715 89549 187716
rect 89486 109050 89546 187715
rect 89944 187168 90264 188192
rect 89944 187104 89952 187168
rect 90016 187104 90032 187168
rect 90096 187104 90112 187168
rect 90176 187104 90192 187168
rect 90256 187104 90264 187168
rect 89944 186080 90264 187104
rect 89944 186016 89952 186080
rect 90016 186016 90032 186080
rect 90096 186016 90112 186080
rect 90176 186016 90192 186080
rect 90256 186016 90264 186080
rect 89944 185576 90264 186016
rect 89944 185340 89986 185576
rect 90222 185340 90264 185576
rect 89944 184992 90264 185340
rect 89944 184928 89952 184992
rect 90016 184928 90032 184992
rect 90096 184928 90112 184992
rect 90176 184928 90192 184992
rect 90256 184928 90264 184992
rect 89944 183904 90264 184928
rect 89944 183840 89952 183904
rect 90016 183840 90032 183904
rect 90096 183840 90112 183904
rect 90176 183840 90192 183904
rect 90256 183840 90264 183904
rect 89944 182816 90264 183840
rect 89944 182752 89952 182816
rect 90016 182752 90032 182816
rect 90096 182752 90112 182816
rect 90176 182752 90192 182816
rect 90256 182752 90264 182816
rect 89944 181728 90264 182752
rect 89944 181664 89952 181728
rect 90016 181664 90032 181728
rect 90096 181664 90112 181728
rect 90176 181664 90192 181728
rect 90256 181664 90264 181728
rect 89944 180640 90264 181664
rect 89944 180576 89952 180640
rect 90016 180576 90032 180640
rect 90096 180576 90112 180640
rect 90176 180576 90192 180640
rect 90256 180576 90264 180640
rect 89944 179552 90264 180576
rect 89944 179488 89952 179552
rect 90016 179488 90032 179552
rect 90096 179488 90112 179552
rect 90176 179488 90192 179552
rect 90256 179488 90264 179552
rect 89944 178464 90264 179488
rect 89944 178400 89952 178464
rect 90016 178400 90032 178464
rect 90096 178400 90112 178464
rect 90176 178400 90192 178464
rect 90256 178400 90264 178464
rect 89944 177376 90264 178400
rect 89944 177312 89952 177376
rect 90016 177312 90032 177376
rect 90096 177312 90112 177376
rect 90176 177312 90192 177376
rect 90256 177312 90264 177376
rect 89944 176288 90264 177312
rect 89944 176224 89952 176288
rect 90016 176224 90032 176288
rect 90096 176224 90112 176288
rect 90176 176224 90192 176288
rect 90256 176224 90264 176288
rect 89944 175576 90264 176224
rect 89944 175340 89986 175576
rect 90222 175340 90264 175576
rect 89944 175200 90264 175340
rect 89944 175136 89952 175200
rect 90016 175136 90032 175200
rect 90096 175136 90112 175200
rect 90176 175136 90192 175200
rect 90256 175136 90264 175200
rect 89944 174112 90264 175136
rect 89944 174048 89952 174112
rect 90016 174048 90032 174112
rect 90096 174048 90112 174112
rect 90176 174048 90192 174112
rect 90256 174048 90264 174112
rect 89944 173024 90264 174048
rect 89944 172960 89952 173024
rect 90016 172960 90032 173024
rect 90096 172960 90112 173024
rect 90176 172960 90192 173024
rect 90256 172960 90264 173024
rect 89944 171936 90264 172960
rect 89944 171872 89952 171936
rect 90016 171872 90032 171936
rect 90096 171872 90112 171936
rect 90176 171872 90192 171936
rect 90256 171872 90264 171936
rect 89944 170848 90264 171872
rect 89944 170784 89952 170848
rect 90016 170784 90032 170848
rect 90096 170784 90112 170848
rect 90176 170784 90192 170848
rect 90256 170784 90264 170848
rect 89944 169760 90264 170784
rect 89944 169696 89952 169760
rect 90016 169696 90032 169760
rect 90096 169696 90112 169760
rect 90176 169696 90192 169760
rect 90256 169696 90264 169760
rect 89944 168672 90264 169696
rect 89944 168608 89952 168672
rect 90016 168608 90032 168672
rect 90096 168608 90112 168672
rect 90176 168608 90192 168672
rect 90256 168608 90264 168672
rect 89944 167584 90264 168608
rect 89944 167520 89952 167584
rect 90016 167520 90032 167584
rect 90096 167520 90112 167584
rect 90176 167520 90192 167584
rect 90256 167520 90264 167584
rect 89944 166496 90264 167520
rect 89944 166432 89952 166496
rect 90016 166432 90032 166496
rect 90096 166432 90112 166496
rect 90176 166432 90192 166496
rect 90256 166432 90264 166496
rect 89944 165576 90264 166432
rect 89944 165408 89986 165576
rect 90222 165408 90264 165576
rect 89944 165344 89952 165408
rect 90256 165344 90264 165408
rect 89944 165340 89986 165344
rect 90222 165340 90264 165344
rect 89944 164320 90264 165340
rect 89944 164256 89952 164320
rect 90016 164256 90032 164320
rect 90096 164256 90112 164320
rect 90176 164256 90192 164320
rect 90256 164256 90264 164320
rect 89944 163232 90264 164256
rect 89944 163168 89952 163232
rect 90016 163168 90032 163232
rect 90096 163168 90112 163232
rect 90176 163168 90192 163232
rect 90256 163168 90264 163232
rect 89944 162144 90264 163168
rect 89944 162080 89952 162144
rect 90016 162080 90032 162144
rect 90096 162080 90112 162144
rect 90176 162080 90192 162144
rect 90256 162080 90264 162144
rect 89944 161056 90264 162080
rect 89944 160992 89952 161056
rect 90016 160992 90032 161056
rect 90096 160992 90112 161056
rect 90176 160992 90192 161056
rect 90256 160992 90264 161056
rect 89944 159968 90264 160992
rect 89944 159904 89952 159968
rect 90016 159904 90032 159968
rect 90096 159904 90112 159968
rect 90176 159904 90192 159968
rect 90256 159904 90264 159968
rect 89944 158880 90264 159904
rect 89944 158816 89952 158880
rect 90016 158816 90032 158880
rect 90096 158816 90112 158880
rect 90176 158816 90192 158880
rect 90256 158816 90264 158880
rect 89944 157792 90264 158816
rect 89944 157728 89952 157792
rect 90016 157728 90032 157792
rect 90096 157728 90112 157792
rect 90176 157728 90192 157792
rect 90256 157728 90264 157792
rect 89944 156704 90264 157728
rect 89944 156640 89952 156704
rect 90016 156640 90032 156704
rect 90096 156640 90112 156704
rect 90176 156640 90192 156704
rect 90256 156640 90264 156704
rect 89944 155616 90264 156640
rect 89944 155552 89952 155616
rect 90016 155576 90032 155616
rect 90096 155576 90112 155616
rect 90176 155576 90192 155616
rect 90256 155552 90264 155616
rect 89944 155340 89986 155552
rect 90222 155340 90264 155552
rect 89944 154528 90264 155340
rect 89944 154464 89952 154528
rect 90016 154464 90032 154528
rect 90096 154464 90112 154528
rect 90176 154464 90192 154528
rect 90256 154464 90264 154528
rect 89944 153440 90264 154464
rect 89944 153376 89952 153440
rect 90016 153376 90032 153440
rect 90096 153376 90112 153440
rect 90176 153376 90192 153440
rect 90256 153376 90264 153440
rect 89944 152352 90264 153376
rect 89944 152288 89952 152352
rect 90016 152288 90032 152352
rect 90096 152288 90112 152352
rect 90176 152288 90192 152352
rect 90256 152288 90264 152352
rect 89944 151264 90264 152288
rect 89944 151200 89952 151264
rect 90016 151200 90032 151264
rect 90096 151200 90112 151264
rect 90176 151200 90192 151264
rect 90256 151200 90264 151264
rect 89944 150176 90264 151200
rect 89944 150112 89952 150176
rect 90016 150112 90032 150176
rect 90096 150112 90112 150176
rect 90176 150112 90192 150176
rect 90256 150112 90264 150176
rect 89944 149088 90264 150112
rect 89944 149024 89952 149088
rect 90016 149024 90032 149088
rect 90096 149024 90112 149088
rect 90176 149024 90192 149088
rect 90256 149024 90264 149088
rect 89944 148000 90264 149024
rect 89944 147936 89952 148000
rect 90016 147936 90032 148000
rect 90096 147936 90112 148000
rect 90176 147936 90192 148000
rect 90256 147936 90264 148000
rect 89944 146912 90264 147936
rect 89944 146848 89952 146912
rect 90016 146848 90032 146912
rect 90096 146848 90112 146912
rect 90176 146848 90192 146912
rect 90256 146848 90264 146912
rect 89944 145824 90264 146848
rect 89944 145760 89952 145824
rect 90016 145760 90032 145824
rect 90096 145760 90112 145824
rect 90176 145760 90192 145824
rect 90256 145760 90264 145824
rect 89944 145576 90264 145760
rect 89944 145340 89986 145576
rect 90222 145340 90264 145576
rect 89944 144736 90264 145340
rect 89944 144672 89952 144736
rect 90016 144672 90032 144736
rect 90096 144672 90112 144736
rect 90176 144672 90192 144736
rect 90256 144672 90264 144736
rect 89944 143648 90264 144672
rect 89944 143584 89952 143648
rect 90016 143584 90032 143648
rect 90096 143584 90112 143648
rect 90176 143584 90192 143648
rect 90256 143584 90264 143648
rect 89944 142560 90264 143584
rect 89944 142496 89952 142560
rect 90016 142496 90032 142560
rect 90096 142496 90112 142560
rect 90176 142496 90192 142560
rect 90256 142496 90264 142560
rect 89944 141472 90264 142496
rect 89944 141408 89952 141472
rect 90016 141408 90032 141472
rect 90096 141408 90112 141472
rect 90176 141408 90192 141472
rect 90256 141408 90264 141472
rect 89944 140384 90264 141408
rect 89944 140320 89952 140384
rect 90016 140320 90032 140384
rect 90096 140320 90112 140384
rect 90176 140320 90192 140384
rect 90256 140320 90264 140384
rect 89944 139296 90264 140320
rect 89944 139232 89952 139296
rect 90016 139232 90032 139296
rect 90096 139232 90112 139296
rect 90176 139232 90192 139296
rect 90256 139232 90264 139296
rect 89944 138208 90264 139232
rect 89944 138144 89952 138208
rect 90016 138144 90032 138208
rect 90096 138144 90112 138208
rect 90176 138144 90192 138208
rect 90256 138144 90264 138208
rect 89944 137120 90264 138144
rect 89944 137056 89952 137120
rect 90016 137056 90032 137120
rect 90096 137056 90112 137120
rect 90176 137056 90192 137120
rect 90256 137056 90264 137120
rect 89944 136032 90264 137056
rect 89944 135968 89952 136032
rect 90016 135968 90032 136032
rect 90096 135968 90112 136032
rect 90176 135968 90192 136032
rect 90256 135968 90264 136032
rect 89944 135576 90264 135968
rect 89944 135340 89986 135576
rect 90222 135340 90264 135576
rect 89944 134944 90264 135340
rect 89944 134880 89952 134944
rect 90016 134880 90032 134944
rect 90096 134880 90112 134944
rect 90176 134880 90192 134944
rect 90256 134880 90264 134944
rect 89944 133856 90264 134880
rect 89944 133792 89952 133856
rect 90016 133792 90032 133856
rect 90096 133792 90112 133856
rect 90176 133792 90192 133856
rect 90256 133792 90264 133856
rect 89944 132768 90264 133792
rect 89944 132704 89952 132768
rect 90016 132704 90032 132768
rect 90096 132704 90112 132768
rect 90176 132704 90192 132768
rect 90256 132704 90264 132768
rect 89944 131680 90264 132704
rect 89944 131616 89952 131680
rect 90016 131616 90032 131680
rect 90096 131616 90112 131680
rect 90176 131616 90192 131680
rect 90256 131616 90264 131680
rect 89944 130592 90264 131616
rect 89944 130528 89952 130592
rect 90016 130528 90032 130592
rect 90096 130528 90112 130592
rect 90176 130528 90192 130592
rect 90256 130528 90264 130592
rect 89944 129504 90264 130528
rect 89944 129440 89952 129504
rect 90016 129440 90032 129504
rect 90096 129440 90112 129504
rect 90176 129440 90192 129504
rect 90256 129440 90264 129504
rect 89944 128416 90264 129440
rect 89944 128352 89952 128416
rect 90016 128352 90032 128416
rect 90096 128352 90112 128416
rect 90176 128352 90192 128416
rect 90256 128352 90264 128416
rect 89944 127328 90264 128352
rect 89944 127264 89952 127328
rect 90016 127264 90032 127328
rect 90096 127264 90112 127328
rect 90176 127264 90192 127328
rect 90256 127264 90264 127328
rect 89944 126240 90264 127264
rect 89944 126176 89952 126240
rect 90016 126176 90032 126240
rect 90096 126176 90112 126240
rect 90176 126176 90192 126240
rect 90256 126176 90264 126240
rect 89944 125576 90264 126176
rect 89944 125340 89986 125576
rect 90222 125340 90264 125576
rect 89944 125152 90264 125340
rect 89944 125088 89952 125152
rect 90016 125088 90032 125152
rect 90096 125088 90112 125152
rect 90176 125088 90192 125152
rect 90256 125088 90264 125152
rect 89944 124064 90264 125088
rect 89944 124000 89952 124064
rect 90016 124000 90032 124064
rect 90096 124000 90112 124064
rect 90176 124000 90192 124064
rect 90256 124000 90264 124064
rect 89944 122976 90264 124000
rect 89944 122912 89952 122976
rect 90016 122912 90032 122976
rect 90096 122912 90112 122976
rect 90176 122912 90192 122976
rect 90256 122912 90264 122976
rect 89944 121888 90264 122912
rect 90587 122636 90653 122637
rect 90587 122572 90588 122636
rect 90652 122572 90653 122636
rect 90587 122571 90653 122572
rect 89944 121824 89952 121888
rect 90016 121824 90032 121888
rect 90096 121824 90112 121888
rect 90176 121824 90192 121888
rect 90256 121824 90264 121888
rect 89944 120800 90264 121824
rect 89944 120736 89952 120800
rect 90016 120736 90032 120800
rect 90096 120736 90112 120800
rect 90176 120736 90192 120800
rect 90256 120736 90264 120800
rect 89944 119712 90264 120736
rect 89944 119648 89952 119712
rect 90016 119648 90032 119712
rect 90096 119648 90112 119712
rect 90176 119648 90192 119712
rect 90256 119648 90264 119712
rect 89944 118624 90264 119648
rect 89944 118560 89952 118624
rect 90016 118560 90032 118624
rect 90096 118560 90112 118624
rect 90176 118560 90192 118624
rect 90256 118560 90264 118624
rect 89944 117536 90264 118560
rect 89944 117472 89952 117536
rect 90016 117472 90032 117536
rect 90096 117472 90112 117536
rect 90176 117472 90192 117536
rect 90256 117472 90264 117536
rect 89944 116448 90264 117472
rect 90590 116738 90650 122571
rect 89944 116384 89952 116448
rect 90016 116384 90032 116448
rect 90096 116384 90112 116448
rect 90176 116384 90192 116448
rect 90256 116384 90264 116448
rect 89944 115576 90264 116384
rect 89944 115360 89986 115576
rect 90222 115360 90264 115576
rect 89944 115296 89952 115360
rect 90016 115296 90032 115340
rect 90096 115296 90112 115340
rect 90176 115296 90192 115340
rect 90256 115296 90264 115360
rect 89944 114272 90264 115296
rect 89944 114208 89952 114272
rect 90016 114208 90032 114272
rect 90096 114208 90112 114272
rect 90176 114208 90192 114272
rect 90256 114208 90264 114272
rect 89944 113184 90264 114208
rect 89944 113120 89952 113184
rect 90016 113120 90032 113184
rect 90096 113120 90112 113184
rect 90176 113120 90192 113184
rect 90256 113120 90264 113184
rect 89944 112096 90264 113120
rect 89944 112032 89952 112096
rect 90016 112032 90032 112096
rect 90096 112032 90112 112096
rect 90176 112032 90192 112096
rect 90256 112032 90264 112096
rect 89944 111008 90264 112032
rect 89944 110944 89952 111008
rect 90016 110944 90032 111008
rect 90096 110944 90112 111008
rect 90176 110944 90192 111008
rect 90256 110944 90264 111008
rect 89944 109920 90264 110944
rect 89944 109856 89952 109920
rect 90016 109856 90032 109920
rect 90096 109856 90112 109920
rect 90176 109856 90192 109920
rect 90256 109856 90264 109920
rect 89486 108990 89730 109050
rect 89299 97884 89365 97885
rect 89299 97820 89300 97884
rect 89364 97820 89365 97884
rect 89299 97819 89365 97820
rect 88934 96870 89178 96930
rect 88382 94830 88810 94890
rect 87944 94080 87952 94144
rect 88016 94080 88032 94144
rect 88096 94080 88112 94144
rect 88176 94080 88192 94144
rect 88256 94080 88264 94144
rect 86539 94076 86605 94077
rect 86539 94012 86540 94076
rect 86604 94012 86605 94076
rect 86539 94011 86605 94012
rect 86355 93940 86421 93941
rect 86355 93876 86356 93940
rect 86420 93876 86421 93940
rect 86355 93875 86421 93876
rect 85944 93536 85952 93600
rect 86016 93536 86032 93600
rect 86096 93536 86112 93600
rect 86176 93536 86192 93600
rect 86256 93536 86264 93600
rect 85944 92512 86264 93536
rect 87944 93056 88264 94080
rect 88750 93618 88810 94830
rect 87944 92992 87952 93056
rect 88016 92992 88032 93056
rect 88096 92992 88112 93056
rect 88176 92992 88192 93056
rect 88256 92992 88264 93056
rect 87275 92852 87341 92853
rect 87275 92788 87276 92852
rect 87340 92788 87341 92852
rect 87275 92787 87341 92788
rect 85944 92448 85952 92512
rect 86016 92448 86032 92512
rect 86096 92448 86112 92512
rect 86176 92448 86192 92512
rect 86256 92448 86264 92512
rect 85944 91424 86264 92448
rect 86907 91764 86973 91765
rect 86907 91700 86908 91764
rect 86972 91700 86973 91764
rect 86907 91699 86973 91700
rect 86910 91578 86970 91699
rect 85944 91360 85952 91424
rect 86016 91360 86032 91424
rect 86096 91360 86112 91424
rect 86176 91360 86192 91424
rect 86256 91360 86264 91424
rect 85944 90336 86264 91360
rect 86907 90540 86973 90541
rect 86907 90476 86908 90540
rect 86972 90476 86973 90540
rect 86907 90475 86973 90476
rect 85944 90272 85952 90336
rect 86016 90272 86032 90336
rect 86096 90272 86112 90336
rect 86176 90272 86192 90336
rect 86256 90272 86264 90336
rect 85944 89248 86264 90272
rect 86910 89538 86970 90475
rect 85944 89184 85952 89248
rect 86016 89184 86032 89248
rect 86096 89184 86112 89248
rect 86176 89184 86192 89248
rect 86256 89184 86264 89248
rect 85944 88160 86264 89184
rect 86907 89044 86973 89045
rect 86907 88980 86908 89044
rect 86972 88980 86973 89044
rect 86907 88979 86973 88980
rect 86910 88858 86970 88979
rect 85944 88096 85952 88160
rect 86016 88096 86032 88160
rect 86096 88096 86112 88160
rect 86176 88096 86192 88160
rect 86256 88096 86264 88160
rect 85944 87072 86264 88096
rect 85944 87008 85952 87072
rect 86016 87008 86032 87072
rect 86096 87008 86112 87072
rect 86176 87008 86192 87072
rect 86256 87008 86264 87072
rect 85944 85984 86264 87008
rect 87278 86818 87338 92787
rect 87944 91968 88264 92992
rect 89118 92938 89178 96870
rect 89670 94298 89730 108990
rect 89944 108832 90264 109856
rect 89944 108768 89952 108832
rect 90016 108768 90032 108832
rect 90096 108768 90112 108832
rect 90176 108768 90192 108832
rect 90256 108768 90264 108832
rect 89944 107744 90264 108768
rect 89944 107680 89952 107744
rect 90016 107680 90032 107744
rect 90096 107680 90112 107744
rect 90176 107680 90192 107744
rect 90256 107680 90264 107744
rect 89944 106656 90264 107680
rect 89944 106592 89952 106656
rect 90016 106592 90032 106656
rect 90096 106592 90112 106656
rect 90176 106592 90192 106656
rect 90256 106592 90264 106656
rect 89944 105576 90264 106592
rect 89944 105568 89986 105576
rect 90222 105568 90264 105576
rect 89944 105504 89952 105568
rect 90256 105504 90264 105568
rect 89944 105340 89986 105504
rect 90222 105340 90264 105504
rect 89944 104480 90264 105340
rect 89944 104416 89952 104480
rect 90016 104416 90032 104480
rect 90096 104416 90112 104480
rect 90176 104416 90192 104480
rect 90256 104416 90264 104480
rect 89944 103392 90264 104416
rect 89944 103328 89952 103392
rect 90016 103328 90032 103392
rect 90096 103328 90112 103392
rect 90176 103328 90192 103392
rect 90256 103328 90264 103392
rect 89944 102304 90264 103328
rect 89944 102240 89952 102304
rect 90016 102240 90032 102304
rect 90096 102240 90112 102304
rect 90176 102240 90192 102304
rect 90256 102240 90264 102304
rect 89944 101216 90264 102240
rect 89944 101152 89952 101216
rect 90016 101152 90032 101216
rect 90096 101152 90112 101216
rect 90176 101152 90192 101216
rect 90256 101152 90264 101216
rect 89944 100128 90264 101152
rect 89944 100064 89952 100128
rect 90016 100064 90032 100128
rect 90096 100064 90112 100128
rect 90176 100064 90192 100128
rect 90256 100064 90264 100128
rect 89944 99040 90264 100064
rect 89944 98976 89952 99040
rect 90016 98976 90032 99040
rect 90096 98976 90112 99040
rect 90176 98976 90192 99040
rect 90256 98976 90264 99040
rect 89944 97952 90264 98976
rect 90587 98156 90653 98157
rect 90587 98092 90588 98156
rect 90652 98092 90653 98156
rect 90587 98091 90653 98092
rect 89944 97888 89952 97952
rect 90016 97888 90032 97952
rect 90096 97888 90112 97952
rect 90176 97888 90192 97952
rect 90256 97888 90264 97952
rect 89944 96864 90264 97888
rect 90590 97698 90650 98091
rect 89944 96800 89952 96864
rect 90016 96800 90032 96864
rect 90096 96800 90112 96864
rect 90176 96800 90192 96864
rect 90256 96800 90264 96864
rect 89944 95776 90264 96800
rect 89944 95712 89952 95776
rect 90016 95712 90032 95776
rect 90096 95712 90112 95776
rect 90176 95712 90192 95776
rect 90256 95712 90264 95776
rect 89944 95576 90264 95712
rect 89944 95340 89986 95576
rect 90222 95340 90264 95576
rect 89944 94688 90264 95340
rect 89944 94624 89952 94688
rect 90016 94624 90032 94688
rect 90096 94624 90112 94688
rect 90176 94624 90192 94688
rect 90256 94624 90264 94688
rect 89944 93600 90264 94624
rect 89944 93536 89952 93600
rect 90016 93536 90032 93600
rect 90096 93536 90112 93600
rect 90176 93536 90192 93600
rect 90256 93536 90264 93600
rect 87944 91904 87952 91968
rect 88016 91904 88032 91968
rect 88096 91904 88112 91968
rect 88176 91904 88192 91968
rect 88256 91904 88264 91968
rect 87944 90880 88264 91904
rect 87944 90816 87952 90880
rect 88016 90816 88032 90880
rect 88096 90816 88112 90880
rect 88176 90816 88192 90880
rect 88256 90816 88264 90880
rect 87944 90576 88264 90816
rect 87944 90340 87986 90576
rect 88222 90340 88264 90576
rect 87944 89792 88264 90340
rect 87944 89728 87952 89792
rect 88016 89728 88032 89792
rect 88096 89728 88112 89792
rect 88176 89728 88192 89792
rect 88256 89728 88264 89792
rect 87944 88704 88264 89728
rect 87944 88640 87952 88704
rect 88016 88640 88032 88704
rect 88096 88640 88112 88704
rect 88176 88640 88192 88704
rect 88256 88640 88264 88704
rect 87944 87616 88264 88640
rect 87944 87552 87952 87616
rect 88016 87552 88032 87616
rect 88096 87552 88112 87616
rect 88176 87552 88192 87616
rect 88256 87552 88264 87616
rect 85944 85920 85952 85984
rect 86016 85920 86032 85984
rect 86096 85920 86112 85984
rect 86176 85920 86192 85984
rect 86256 85920 86264 85984
rect 85944 85576 86264 85920
rect 85944 85340 85986 85576
rect 86222 85340 86264 85576
rect 85944 84896 86264 85340
rect 85944 84832 85952 84896
rect 86016 84832 86032 84896
rect 86096 84832 86112 84896
rect 86176 84832 86192 84896
rect 86256 84832 86264 84896
rect 85944 83808 86264 84832
rect 85944 83744 85952 83808
rect 86016 83744 86032 83808
rect 86096 83744 86112 83808
rect 86176 83744 86192 83808
rect 86256 83744 86264 83808
rect 85944 82720 86264 83744
rect 85944 82656 85952 82720
rect 86016 82656 86032 82720
rect 86096 82656 86112 82720
rect 86176 82656 86192 82720
rect 86256 82656 86264 82720
rect 85944 81632 86264 82656
rect 85944 81568 85952 81632
rect 86016 81568 86032 81632
rect 86096 81568 86112 81632
rect 86176 81568 86192 81632
rect 86256 81568 86264 81632
rect 85944 80544 86264 81568
rect 85944 80480 85952 80544
rect 86016 80480 86032 80544
rect 86096 80480 86112 80544
rect 86176 80480 86192 80544
rect 86256 80480 86264 80544
rect 85944 79456 86264 80480
rect 85944 79392 85952 79456
rect 86016 79392 86032 79456
rect 86096 79392 86112 79456
rect 86176 79392 86192 79456
rect 86256 79392 86264 79456
rect 85944 78368 86264 79392
rect 85944 78304 85952 78368
rect 86016 78304 86032 78368
rect 86096 78304 86112 78368
rect 86176 78304 86192 78368
rect 86256 78304 86264 78368
rect 85944 77280 86264 78304
rect 85944 77216 85952 77280
rect 86016 77216 86032 77280
rect 86096 77216 86112 77280
rect 86176 77216 86192 77280
rect 86256 77216 86264 77280
rect 85944 76192 86264 77216
rect 85944 76128 85952 76192
rect 86016 76128 86032 76192
rect 86096 76128 86112 76192
rect 86176 76128 86192 76192
rect 86256 76128 86264 76192
rect 85944 75576 86264 76128
rect 85944 75340 85986 75576
rect 86222 75340 86264 75576
rect 85944 75104 86264 75340
rect 85944 75040 85952 75104
rect 86016 75040 86032 75104
rect 86096 75040 86112 75104
rect 86176 75040 86192 75104
rect 86256 75040 86264 75104
rect 85944 74016 86264 75040
rect 85944 73952 85952 74016
rect 86016 73952 86032 74016
rect 86096 73952 86112 74016
rect 86176 73952 86192 74016
rect 86256 73952 86264 74016
rect 85944 72928 86264 73952
rect 85944 72864 85952 72928
rect 86016 72864 86032 72928
rect 86096 72864 86112 72928
rect 86176 72864 86192 72928
rect 86256 72864 86264 72928
rect 85944 71840 86264 72864
rect 85944 71776 85952 71840
rect 86016 71776 86032 71840
rect 86096 71776 86112 71840
rect 86176 71776 86192 71840
rect 86256 71776 86264 71840
rect 85944 70752 86264 71776
rect 85944 70688 85952 70752
rect 86016 70688 86032 70752
rect 86096 70688 86112 70752
rect 86176 70688 86192 70752
rect 86256 70688 86264 70752
rect 85944 69664 86264 70688
rect 85944 69600 85952 69664
rect 86016 69600 86032 69664
rect 86096 69600 86112 69664
rect 86176 69600 86192 69664
rect 86256 69600 86264 69664
rect 85944 68576 86264 69600
rect 85944 68512 85952 68576
rect 86016 68512 86032 68576
rect 86096 68512 86112 68576
rect 86176 68512 86192 68576
rect 86256 68512 86264 68576
rect 85944 67488 86264 68512
rect 85944 67424 85952 67488
rect 86016 67424 86032 67488
rect 86096 67424 86112 67488
rect 86176 67424 86192 67488
rect 86256 67424 86264 67488
rect 85944 66400 86264 67424
rect 85944 66336 85952 66400
rect 86016 66336 86032 66400
rect 86096 66336 86112 66400
rect 86176 66336 86192 66400
rect 86256 66336 86264 66400
rect 85944 65576 86264 66336
rect 85944 65340 85986 65576
rect 86222 65340 86264 65576
rect 85944 65312 86264 65340
rect 85944 65248 85952 65312
rect 86016 65248 86032 65312
rect 86096 65248 86112 65312
rect 86176 65248 86192 65312
rect 86256 65248 86264 65312
rect 85944 64224 86264 65248
rect 85944 64160 85952 64224
rect 86016 64160 86032 64224
rect 86096 64160 86112 64224
rect 86176 64160 86192 64224
rect 86256 64160 86264 64224
rect 85944 63136 86264 64160
rect 85944 63072 85952 63136
rect 86016 63072 86032 63136
rect 86096 63072 86112 63136
rect 86176 63072 86192 63136
rect 86256 63072 86264 63136
rect 85944 62048 86264 63072
rect 85944 61984 85952 62048
rect 86016 61984 86032 62048
rect 86096 61984 86112 62048
rect 86176 61984 86192 62048
rect 86256 61984 86264 62048
rect 85944 60960 86264 61984
rect 85944 60896 85952 60960
rect 86016 60896 86032 60960
rect 86096 60896 86112 60960
rect 86176 60896 86192 60960
rect 86256 60896 86264 60960
rect 85944 59872 86264 60896
rect 85944 59808 85952 59872
rect 86016 59808 86032 59872
rect 86096 59808 86112 59872
rect 86176 59808 86192 59872
rect 86256 59808 86264 59872
rect 85944 58784 86264 59808
rect 85944 58720 85952 58784
rect 86016 58720 86032 58784
rect 86096 58720 86112 58784
rect 86176 58720 86192 58784
rect 86256 58720 86264 58784
rect 85944 57696 86264 58720
rect 85944 57632 85952 57696
rect 86016 57632 86032 57696
rect 86096 57632 86112 57696
rect 86176 57632 86192 57696
rect 86256 57632 86264 57696
rect 85944 56608 86264 57632
rect 85944 56544 85952 56608
rect 86016 56544 86032 56608
rect 86096 56544 86112 56608
rect 86176 56544 86192 56608
rect 86256 56544 86264 56608
rect 85944 55576 86264 56544
rect 85944 55520 85986 55576
rect 86222 55520 86264 55576
rect 85944 55456 85952 55520
rect 86256 55456 86264 55520
rect 85944 55340 85986 55456
rect 86222 55340 86264 55456
rect 84147 55316 84213 55317
rect 84147 55252 84148 55316
rect 84212 55252 84213 55316
rect 84147 55251 84213 55252
rect 85944 54432 86264 55340
rect 85944 54368 85952 54432
rect 86016 54368 86032 54432
rect 86096 54368 86112 54432
rect 86176 54368 86192 54432
rect 86256 54368 86264 54432
rect 85944 53344 86264 54368
rect 85944 53280 85952 53344
rect 86016 53280 86032 53344
rect 86096 53280 86112 53344
rect 86176 53280 86192 53344
rect 86256 53280 86264 53344
rect 85944 52256 86264 53280
rect 85944 52192 85952 52256
rect 86016 52192 86032 52256
rect 86096 52192 86112 52256
rect 86176 52192 86192 52256
rect 86256 52192 86264 52256
rect 83779 51372 83845 51373
rect 83779 51308 83780 51372
rect 83844 51308 83845 51372
rect 83779 51307 83845 51308
rect 85944 51168 86264 52192
rect 85944 51104 85952 51168
rect 86016 51104 86032 51168
rect 86096 51104 86112 51168
rect 86176 51104 86192 51168
rect 86256 51104 86264 51168
rect 85944 50080 86264 51104
rect 85944 50016 85952 50080
rect 86016 50016 86032 50080
rect 86096 50016 86112 50080
rect 86176 50016 86192 50080
rect 86256 50016 86264 50080
rect 83595 49740 83661 49741
rect 83595 49676 83596 49740
rect 83660 49676 83661 49740
rect 83595 49675 83661 49676
rect 83414 49270 83658 49330
rect 82494 45576 82814 45618
rect 82494 45340 82536 45576
rect 82772 45340 82814 45576
rect 83598 45570 83658 49270
rect 85944 48992 86264 50016
rect 85944 48928 85952 48992
rect 86016 48928 86032 48992
rect 86096 48928 86112 48992
rect 86176 48928 86192 48992
rect 86256 48928 86264 48992
rect 85944 47904 86264 48928
rect 85944 47840 85952 47904
rect 86016 47840 86032 47904
rect 86096 47840 86112 47904
rect 86176 47840 86192 47904
rect 86256 47840 86264 47904
rect 85944 46816 86264 47840
rect 85944 46752 85952 46816
rect 86016 46752 86032 46816
rect 86096 46752 86112 46816
rect 86176 46752 86192 46816
rect 86256 46752 86264 46816
rect 85944 45728 86264 46752
rect 85944 45664 85952 45728
rect 86016 45664 86032 45728
rect 86096 45664 86112 45728
rect 86176 45664 86192 45728
rect 86256 45664 86264 45728
rect 85944 45576 86264 45664
rect 83411 45524 83477 45525
rect 83411 45460 83412 45524
rect 83476 45460 83477 45524
rect 83598 45510 83842 45570
rect 83411 45459 83477 45460
rect 82494 45298 82814 45340
rect 82938 40576 83262 40618
rect 82938 40340 82982 40576
rect 83218 40340 83262 40576
rect 82938 40298 83262 40340
rect 82494 35576 82814 35618
rect 82494 35340 82536 35576
rect 82772 35340 82814 35576
rect 82494 35298 82814 35340
rect 83414 33829 83474 45459
rect 83782 38670 83842 45510
rect 83598 38610 83842 38670
rect 85944 45340 85986 45576
rect 86222 45340 86264 45576
rect 85944 44640 86264 45340
rect 85944 44576 85952 44640
rect 86016 44576 86032 44640
rect 86096 44576 86112 44640
rect 86176 44576 86192 44640
rect 86256 44576 86264 44640
rect 85944 43552 86264 44576
rect 85944 43488 85952 43552
rect 86016 43488 86032 43552
rect 86096 43488 86112 43552
rect 86176 43488 86192 43552
rect 86256 43488 86264 43552
rect 85944 42464 86264 43488
rect 85944 42400 85952 42464
rect 86016 42400 86032 42464
rect 86096 42400 86112 42464
rect 86176 42400 86192 42464
rect 86256 42400 86264 42464
rect 85944 41376 86264 42400
rect 85944 41312 85952 41376
rect 86016 41312 86032 41376
rect 86096 41312 86112 41376
rect 86176 41312 86192 41376
rect 86256 41312 86264 41376
rect 85944 40288 86264 41312
rect 85944 40224 85952 40288
rect 86016 40224 86032 40288
rect 86096 40224 86112 40288
rect 86176 40224 86192 40288
rect 86256 40224 86264 40288
rect 85944 39200 86264 40224
rect 85944 39136 85952 39200
rect 86016 39136 86032 39200
rect 86096 39136 86112 39200
rect 86176 39136 86192 39200
rect 86256 39136 86264 39200
rect 83411 33828 83477 33829
rect 83411 33764 83412 33828
rect 83476 33764 83477 33828
rect 83411 33763 83477 33764
rect 82938 30576 83262 30618
rect 82938 30340 82982 30576
rect 83218 30340 83262 30576
rect 82938 30298 83262 30340
rect 83598 29010 83658 38610
rect 85944 38112 86264 39136
rect 85944 38048 85952 38112
rect 86016 38048 86032 38112
rect 86096 38048 86112 38112
rect 86176 38048 86192 38112
rect 86256 38048 86264 38112
rect 85944 37024 86264 38048
rect 85944 36960 85952 37024
rect 86016 36960 86032 37024
rect 86096 36960 86112 37024
rect 86176 36960 86192 37024
rect 86256 36960 86264 37024
rect 85944 35936 86264 36960
rect 85944 35872 85952 35936
rect 86016 35872 86032 35936
rect 86096 35872 86112 35936
rect 86176 35872 86192 35936
rect 86256 35872 86264 35936
rect 85944 35576 86264 35872
rect 85944 35340 85986 35576
rect 86222 35340 86264 35576
rect 85944 34848 86264 35340
rect 85944 34784 85952 34848
rect 86016 34784 86032 34848
rect 86096 34784 86112 34848
rect 86176 34784 86192 34848
rect 86256 34784 86264 34848
rect 83963 33828 84029 33829
rect 83963 33764 83964 33828
rect 84028 33764 84029 33828
rect 83963 33763 84029 33764
rect 83598 28950 83842 29010
rect 82494 25576 82814 25618
rect 82494 25340 82536 25576
rect 82772 25340 82814 25576
rect 82494 25298 82814 25340
rect 82938 20576 83262 20618
rect 82938 20340 82982 20576
rect 83218 20340 83262 20576
rect 82938 20298 83262 20340
rect 82494 15576 82814 15618
rect 82494 15340 82536 15576
rect 82772 15340 82814 15576
rect 82494 15298 82814 15340
rect 82938 10576 83262 10618
rect 82938 10340 82982 10576
rect 83218 10340 83262 10576
rect 82938 10298 83262 10340
rect 4475 10164 4541 10165
rect 4475 10100 4476 10164
rect 4540 10100 4541 10164
rect 4475 10099 4541 10100
rect 3944 9216 3952 9280
rect 4016 9216 4032 9280
rect 4096 9216 4112 9280
rect 4176 9216 4192 9280
rect 4256 9216 4264 9280
rect 3944 8192 4264 9216
rect 3944 8128 3952 8192
rect 4016 8128 4032 8192
rect 4096 8128 4112 8192
rect 4176 8128 4192 8192
rect 4256 8128 4264 8192
rect 3944 7104 4264 8128
rect 3944 7040 3952 7104
rect 4016 7040 4032 7104
rect 4096 7040 4112 7104
rect 4176 7040 4192 7104
rect 4256 7040 4264 7104
rect 3944 6016 4264 7040
rect 3944 5952 3952 6016
rect 4016 5952 4032 6016
rect 4096 5952 4112 6016
rect 4176 5952 4192 6016
rect 4256 5952 4264 6016
rect 3944 4928 4264 5952
rect 82494 5576 82814 5618
rect 82494 5340 82536 5576
rect 82772 5340 82814 5576
rect 82494 5298 82814 5340
rect 3944 4864 3952 4928
rect 4016 4864 4032 4928
rect 4096 4864 4112 4928
rect 4176 4864 4192 4928
rect 4256 4864 4264 4928
rect 3944 3840 4264 4864
rect 4843 3908 4909 3909
rect 4843 3858 4844 3908
rect 4908 3858 4909 3908
rect 3944 3776 3952 3840
rect 4016 3776 4032 3840
rect 4096 3776 4112 3840
rect 4176 3776 4192 3840
rect 4256 3776 4264 3840
rect 3944 2752 4264 3776
rect 39067 3228 39133 3229
rect 15168 3030 15394 3090
rect 3944 2688 3952 2752
rect 4016 2688 4032 2752
rect 4096 2688 4112 2752
rect 4176 2688 4192 2752
rect 4256 2688 4264 2752
rect 3944 2128 4264 2688
rect 8158 2685 8218 2942
rect 15334 2685 15394 3030
rect 20670 3030 21008 3090
rect 25086 3030 25680 3090
rect 20670 2685 20730 3030
rect 22694 2690 23344 2750
rect 8155 2684 8221 2685
rect 8155 2620 8156 2684
rect 8220 2620 8221 2684
rect 8155 2619 8221 2620
rect 15331 2684 15397 2685
rect 15331 2620 15332 2684
rect 15396 2620 15397 2684
rect 15331 2619 15397 2620
rect 20667 2684 20733 2685
rect 20667 2620 20668 2684
rect 20732 2620 20733 2684
rect 20667 2619 20733 2620
rect 22694 2549 22754 2690
rect 25086 2685 25146 3030
rect 39067 3164 39068 3228
rect 39132 3164 39133 3228
rect 45323 3228 45389 3229
rect 39067 3163 39133 3164
rect 39070 3090 39130 3163
rect 40171 3092 40237 3093
rect 37194 3030 37360 3090
rect 37966 3030 38528 3090
rect 39070 3030 39696 3090
rect 37966 2957 38026 3030
rect 40171 3028 40172 3092
rect 40236 3090 40237 3092
rect 40236 3030 40864 3090
rect 40236 3028 40237 3030
rect 40171 3027 40237 3028
rect 37963 2956 38029 2957
rect 37963 2892 37964 2956
rect 38028 2892 38029 2956
rect 45323 3164 45324 3228
rect 45388 3164 45389 3228
rect 45323 3163 45389 3164
rect 47715 3228 47781 3229
rect 47715 3164 47716 3228
rect 47780 3164 47781 3228
rect 47715 3163 47781 3164
rect 45326 3090 45386 3163
rect 47718 3090 47778 3163
rect 41610 3030 42032 3090
rect 44038 3030 44368 3090
rect 45326 3030 45536 3090
rect 46246 3030 46704 3090
rect 47718 3030 47872 3090
rect 49926 3030 50208 3090
rect 53422 3030 53712 3090
rect 44038 2957 44098 3030
rect 44035 2956 44101 2957
rect 37963 2891 38029 2892
rect 44035 2892 44036 2956
rect 44100 2892 44101 2956
rect 44035 2891 44101 2892
rect 46246 2821 46306 3030
rect 49926 2957 49986 3030
rect 53422 2957 53482 3030
rect 49923 2956 49989 2957
rect 49923 2892 49924 2956
rect 49988 2892 49989 2956
rect 49923 2891 49989 2892
rect 53419 2956 53485 2957
rect 53419 2892 53420 2956
rect 53484 2892 53485 2956
rect 53419 2891 53485 2892
rect 26003 2820 26069 2821
rect 26003 2756 26004 2820
rect 26068 2790 26069 2820
rect 46243 2820 46309 2821
rect 26068 2756 26250 2790
rect 26003 2755 26250 2756
rect 46243 2756 46244 2820
rect 46308 2756 46309 2820
rect 83782 2790 83842 28950
rect 83966 22110 84026 33763
rect 85944 33760 86264 34784
rect 85944 33696 85952 33760
rect 86016 33696 86032 33760
rect 86096 33696 86112 33760
rect 86176 33696 86192 33760
rect 86256 33696 86264 33760
rect 85944 32672 86264 33696
rect 85944 32608 85952 32672
rect 86016 32608 86032 32672
rect 86096 32608 86112 32672
rect 86176 32608 86192 32672
rect 86256 32608 86264 32672
rect 85944 31584 86264 32608
rect 85944 31520 85952 31584
rect 86016 31520 86032 31584
rect 86096 31520 86112 31584
rect 86176 31520 86192 31584
rect 86256 31520 86264 31584
rect 85944 30496 86264 31520
rect 85944 30432 85952 30496
rect 86016 30432 86032 30496
rect 86096 30432 86112 30496
rect 86176 30432 86192 30496
rect 86256 30432 86264 30496
rect 85944 29408 86264 30432
rect 85944 29344 85952 29408
rect 86016 29344 86032 29408
rect 86096 29344 86112 29408
rect 86176 29344 86192 29408
rect 86256 29344 86264 29408
rect 85944 28320 86264 29344
rect 85944 28256 85952 28320
rect 86016 28256 86032 28320
rect 86096 28256 86112 28320
rect 86176 28256 86192 28320
rect 86256 28256 86264 28320
rect 85944 27232 86264 28256
rect 85944 27168 85952 27232
rect 86016 27168 86032 27232
rect 86096 27168 86112 27232
rect 86176 27168 86192 27232
rect 86256 27168 86264 27232
rect 85944 26144 86264 27168
rect 85944 26080 85952 26144
rect 86016 26080 86032 26144
rect 86096 26080 86112 26144
rect 86176 26080 86192 26144
rect 86256 26080 86264 26144
rect 85944 25576 86264 26080
rect 85944 25340 85986 25576
rect 86222 25340 86264 25576
rect 85944 25056 86264 25340
rect 85944 24992 85952 25056
rect 86016 24992 86032 25056
rect 86096 24992 86112 25056
rect 86176 24992 86192 25056
rect 86256 24992 86264 25056
rect 85944 23968 86264 24992
rect 85944 23904 85952 23968
rect 86016 23904 86032 23968
rect 86096 23904 86112 23968
rect 86176 23904 86192 23968
rect 86256 23904 86264 23968
rect 85944 22880 86264 23904
rect 85944 22816 85952 22880
rect 86016 22816 86032 22880
rect 86096 22816 86112 22880
rect 86176 22816 86192 22880
rect 86256 22816 86264 22880
rect 83966 22050 84210 22110
rect 84150 16693 84210 22050
rect 85944 21792 86264 22816
rect 85944 21728 85952 21792
rect 86016 21728 86032 21792
rect 86096 21728 86112 21792
rect 86176 21728 86192 21792
rect 86256 21728 86264 21792
rect 85944 20704 86264 21728
rect 85944 20640 85952 20704
rect 86016 20640 86032 20704
rect 86096 20640 86112 20704
rect 86176 20640 86192 20704
rect 86256 20640 86264 20704
rect 85944 19616 86264 20640
rect 85944 19552 85952 19616
rect 86016 19552 86032 19616
rect 86096 19552 86112 19616
rect 86176 19552 86192 19616
rect 86256 19552 86264 19616
rect 85944 18528 86264 19552
rect 85944 18464 85952 18528
rect 86016 18464 86032 18528
rect 86096 18464 86112 18528
rect 86176 18464 86192 18528
rect 86256 18464 86264 18528
rect 85944 17440 86264 18464
rect 85944 17376 85952 17440
rect 86016 17376 86032 17440
rect 86096 17376 86112 17440
rect 86176 17376 86192 17440
rect 86256 17376 86264 17440
rect 84147 16692 84213 16693
rect 84147 16628 84148 16692
rect 84212 16628 84213 16692
rect 84147 16627 84213 16628
rect 46243 2755 46309 2756
rect 26006 2750 26250 2755
rect 26006 2730 26848 2750
rect 26190 2690 26848 2730
rect 27662 2690 28016 2750
rect 29686 2690 30352 2750
rect 30974 2690 31520 2750
rect 38652 2690 39314 2750
rect 40988 2690 41338 2750
rect 42156 2690 42626 2750
rect 44492 2690 44834 2750
rect 47996 2690 48146 2750
rect 51500 2690 52194 2750
rect 25083 2684 25149 2685
rect 25083 2620 25084 2684
rect 25148 2620 25149 2684
rect 25083 2619 25149 2620
rect 22691 2548 22757 2549
rect 22691 2484 22692 2548
rect 22756 2484 22757 2548
rect 22691 2483 22757 2484
rect 9803 2277 9863 2380
rect 9800 2276 9866 2277
rect 9800 2212 9801 2276
rect 9865 2212 9866 2276
rect 9800 2211 9866 2212
rect 12802 1730 12862 2380
rect 13970 2277 14030 2380
rect 16306 2277 16366 2380
rect 13967 2276 14033 2277
rect 13967 2212 13968 2276
rect 14032 2212 14033 2276
rect 13967 2211 14033 2212
rect 16303 2276 16369 2277
rect 16303 2212 16304 2276
rect 16368 2212 16369 2276
rect 16303 2211 16369 2212
rect 17474 1869 17534 2380
rect 17471 1868 17537 1869
rect 17471 1804 17472 1868
rect 17536 1804 17537 1868
rect 17471 1803 17537 1804
rect 12758 1670 12862 1730
rect 18642 1730 18702 2380
rect 18766 1730 18826 2380
rect 19810 1730 19870 2380
rect 18642 1670 18706 1730
rect 18766 1670 18890 1730
rect 12758 1325 12818 1670
rect 12755 1324 12821 1325
rect 12755 1260 12756 1324
rect 12820 1260 12821 1324
rect 12755 1259 12821 1260
rect 18646 1189 18706 1670
rect 18830 1325 18890 1670
rect 19750 1670 19870 1730
rect 18827 1324 18893 1325
rect 18827 1260 18828 1324
rect 18892 1260 18893 1324
rect 18827 1259 18893 1260
rect 19750 1189 19810 1670
rect 18643 1188 18709 1189
rect 18643 1124 18644 1188
rect 18708 1124 18709 1188
rect 18643 1123 18709 1124
rect 19747 1188 19813 1189
rect 19747 1124 19748 1188
rect 19812 1124 19813 1188
rect 19747 1123 19813 1124
rect 19934 237 19994 2380
rect 21102 1869 21162 2380
rect 22146 2277 22206 2380
rect 22143 2276 22209 2277
rect 22143 2212 22144 2276
rect 22208 2212 22209 2276
rect 22143 2211 22209 2212
rect 22270 1869 22330 2380
rect 21099 1868 21165 1869
rect 21099 1804 21100 1868
rect 21164 1804 21165 1868
rect 21099 1803 21165 1804
rect 22267 1868 22333 1869
rect 22267 1804 22268 1868
rect 22332 1804 22333 1868
rect 22267 1803 22333 1804
rect 23438 1730 23498 2380
rect 24482 2277 24542 2380
rect 24479 2276 24545 2277
rect 24479 2212 24480 2276
rect 24544 2212 24545 2276
rect 24479 2211 24545 2212
rect 23430 1670 23498 1730
rect 24606 1730 24666 2380
rect 25774 1869 25834 2380
rect 26942 1869 27002 2380
rect 25771 1868 25837 1869
rect 25771 1804 25772 1868
rect 25836 1804 25837 1868
rect 25771 1803 25837 1804
rect 26939 1868 27005 1869
rect 26939 1804 26940 1868
rect 27004 1804 27005 1868
rect 26939 1803 27005 1804
rect 24606 1670 24778 1730
rect 23430 781 23490 1670
rect 24718 1053 24778 1670
rect 24715 1052 24781 1053
rect 24715 988 24716 1052
rect 24780 988 24781 1052
rect 24715 987 24781 988
rect 27662 917 27722 2690
rect 28110 1869 28170 2380
rect 29154 2005 29214 2380
rect 29151 2004 29217 2005
rect 29151 1940 29152 2004
rect 29216 1940 29217 2004
rect 29151 1939 29217 1940
rect 28107 1868 28173 1869
rect 28107 1804 28108 1868
rect 28172 1804 28173 1868
rect 28107 1803 28173 1804
rect 29278 1730 29338 2380
rect 29278 1670 29378 1730
rect 29318 1325 29378 1670
rect 29315 1324 29381 1325
rect 29315 1260 29316 1324
rect 29380 1260 29381 1324
rect 29315 1259 29381 1260
rect 29686 1189 29746 2690
rect 30446 2005 30506 2380
rect 30443 2004 30509 2005
rect 30443 1940 30444 2004
rect 30508 1940 30509 2004
rect 30443 1939 30509 1940
rect 29683 1188 29749 1189
rect 29683 1124 29684 1188
rect 29748 1124 29749 1188
rect 29683 1123 29749 1124
rect 30974 1053 31034 2690
rect 31614 2005 31674 2380
rect 32658 2277 32718 2380
rect 32655 2276 32721 2277
rect 32655 2212 32656 2276
rect 32720 2212 32721 2276
rect 32655 2211 32721 2212
rect 32782 2141 32842 2380
rect 32779 2140 32845 2141
rect 32779 2076 32780 2140
rect 32844 2076 32845 2140
rect 32779 2075 32845 2076
rect 31611 2004 31677 2005
rect 31611 1940 31612 2004
rect 31676 1940 31677 2004
rect 31611 1939 31677 1940
rect 33826 1866 33886 2380
rect 33950 2141 34010 2380
rect 33947 2140 34013 2141
rect 33947 2076 33948 2140
rect 34012 2076 34013 2140
rect 33947 2075 34013 2076
rect 34994 1866 35054 2380
rect 33734 1806 33886 1866
rect 34838 1806 35054 1866
rect 35118 1866 35178 2380
rect 36162 2277 36222 2380
rect 36159 2276 36225 2277
rect 36159 2212 36160 2276
rect 36224 2212 36225 2276
rect 36159 2211 36225 2212
rect 36286 2141 36346 2380
rect 37454 2277 37514 2380
rect 37451 2276 37517 2277
rect 37451 2212 37452 2276
rect 37516 2212 37517 2276
rect 37451 2211 37517 2212
rect 36283 2140 36349 2141
rect 36283 2076 36284 2140
rect 36348 2076 36349 2140
rect 36283 2075 36349 2076
rect 35118 1806 35266 1866
rect 30971 1052 31037 1053
rect 30971 988 30972 1052
rect 31036 988 31037 1052
rect 30971 987 31037 988
rect 27659 916 27725 917
rect 27659 852 27660 916
rect 27724 852 27725 916
rect 27659 851 27725 852
rect 33734 781 33794 1806
rect 34838 1189 34898 1806
rect 35206 1325 35266 1806
rect 39254 1325 39314 2690
rect 39790 1730 39850 2380
rect 39790 1670 39866 1730
rect 35203 1324 35269 1325
rect 35203 1260 35204 1324
rect 35268 1260 35269 1324
rect 35203 1259 35269 1260
rect 39251 1324 39317 1325
rect 39251 1260 39252 1324
rect 39316 1260 39317 1324
rect 39251 1259 39317 1260
rect 39806 1189 39866 1670
rect 34835 1188 34901 1189
rect 34835 1124 34836 1188
rect 34900 1124 34901 1188
rect 34835 1123 34901 1124
rect 39803 1188 39869 1189
rect 39803 1124 39804 1188
rect 39868 1124 39869 1188
rect 39803 1123 39869 1124
rect 41278 1053 41338 2690
rect 42566 1053 42626 2690
rect 43170 1730 43230 2380
rect 43118 1670 43230 1730
rect 43294 1730 43354 2380
rect 43294 1670 43362 1730
rect 41275 1052 41341 1053
rect 41275 988 41276 1052
rect 41340 988 41341 1052
rect 41275 987 41341 988
rect 42563 1052 42629 1053
rect 42563 988 42564 1052
rect 42628 988 42629 1052
rect 42563 987 42629 988
rect 43118 917 43178 1670
rect 43302 917 43362 1670
rect 44774 1325 44834 2690
rect 45630 1730 45690 2380
rect 45630 1670 45754 1730
rect 44771 1324 44837 1325
rect 44771 1260 44772 1324
rect 44836 1260 44837 1324
rect 44771 1259 44837 1260
rect 45694 1053 45754 1670
rect 45691 1052 45757 1053
rect 45691 988 45692 1052
rect 45756 988 45757 1052
rect 45691 987 45757 988
rect 46798 917 46858 2380
rect 48086 1325 48146 2690
rect 49010 1730 49070 2380
rect 49006 1670 49070 1730
rect 49134 1730 49194 2380
rect 50302 1730 50362 2380
rect 51346 2277 51406 2380
rect 51343 2276 51409 2277
rect 51343 2212 51344 2276
rect 51408 2212 51409 2276
rect 51343 2211 51409 2212
rect 49134 1670 49250 1730
rect 49006 1597 49066 1670
rect 49003 1596 49069 1597
rect 49003 1532 49004 1596
rect 49068 1532 49069 1596
rect 49003 1531 49069 1532
rect 48083 1324 48149 1325
rect 48083 1260 48084 1324
rect 48148 1260 48149 1324
rect 48083 1259 48149 1260
rect 49190 1053 49250 1670
rect 50294 1670 50362 1730
rect 49187 1052 49253 1053
rect 49187 988 49188 1052
rect 49252 988 49253 1052
rect 49187 987 49253 988
rect 43115 916 43181 917
rect 43115 852 43116 916
rect 43180 852 43181 916
rect 43115 851 43181 852
rect 43299 916 43365 917
rect 43299 852 43300 916
rect 43364 852 43365 916
rect 43299 851 43365 852
rect 46795 916 46861 917
rect 46795 852 46796 916
rect 46860 852 46861 916
rect 46795 851 46861 852
rect 50294 781 50354 1670
rect 52134 1189 52194 2690
rect 54710 2690 54880 2750
rect 83414 2730 83842 2790
rect 85944 16352 86264 17376
rect 85944 16288 85952 16352
rect 86016 16288 86032 16352
rect 86096 16288 86112 16352
rect 86176 16288 86192 16352
rect 86256 16288 86264 16352
rect 85944 15576 86264 16288
rect 85944 15340 85986 15576
rect 86222 15340 86264 15576
rect 85944 15264 86264 15340
rect 85944 15200 85952 15264
rect 86016 15200 86032 15264
rect 86096 15200 86112 15264
rect 86176 15200 86192 15264
rect 86256 15200 86264 15264
rect 85944 14176 86264 15200
rect 85944 14112 85952 14176
rect 86016 14112 86032 14176
rect 86096 14112 86112 14176
rect 86176 14112 86192 14176
rect 86256 14112 86264 14176
rect 85944 13088 86264 14112
rect 85944 13024 85952 13088
rect 86016 13024 86032 13088
rect 86096 13024 86112 13088
rect 86176 13024 86192 13088
rect 86256 13024 86264 13088
rect 85944 12000 86264 13024
rect 85944 11936 85952 12000
rect 86016 11936 86032 12000
rect 86096 11936 86112 12000
rect 86176 11936 86192 12000
rect 86256 11936 86264 12000
rect 85944 10912 86264 11936
rect 85944 10848 85952 10912
rect 86016 10848 86032 10912
rect 86096 10848 86112 10912
rect 86176 10848 86192 10912
rect 86256 10848 86264 10912
rect 85944 9824 86264 10848
rect 85944 9760 85952 9824
rect 86016 9760 86032 9824
rect 86096 9760 86112 9824
rect 86176 9760 86192 9824
rect 86256 9760 86264 9824
rect 85944 8736 86264 9760
rect 85944 8672 85952 8736
rect 86016 8672 86032 8736
rect 86096 8672 86112 8736
rect 86176 8672 86192 8736
rect 86256 8672 86264 8736
rect 85944 7648 86264 8672
rect 85944 7584 85952 7648
rect 86016 7584 86032 7648
rect 86096 7584 86112 7648
rect 86176 7584 86192 7648
rect 86256 7584 86264 7648
rect 85944 6560 86264 7584
rect 85944 6496 85952 6560
rect 86016 6496 86032 6560
rect 86096 6496 86112 6560
rect 86176 6496 86192 6560
rect 86256 6496 86264 6560
rect 85944 5576 86264 6496
rect 85944 5472 85986 5576
rect 86222 5472 86264 5576
rect 85944 5408 85952 5472
rect 86256 5408 86264 5472
rect 85944 5340 85986 5408
rect 86222 5340 86264 5408
rect 85944 4384 86264 5340
rect 85944 4320 85952 4384
rect 86016 4320 86032 4384
rect 86096 4320 86112 4384
rect 86176 4320 86192 4384
rect 86256 4320 86264 4384
rect 85944 3296 86264 4320
rect 85944 3232 85952 3296
rect 86016 3232 86032 3296
rect 86096 3232 86112 3296
rect 86176 3232 86192 3296
rect 86256 3232 86264 3296
rect 52514 2277 52574 2380
rect 52511 2276 52577 2277
rect 52511 2212 52512 2276
rect 52576 2212 52577 2276
rect 52511 2211 52577 2212
rect 52638 1730 52698 2380
rect 53806 1730 53866 2380
rect 52638 1670 52746 1730
rect 52131 1188 52197 1189
rect 52131 1124 52132 1188
rect 52196 1124 52197 1188
rect 52131 1123 52197 1124
rect 23427 780 23493 781
rect 23427 716 23428 780
rect 23492 716 23493 780
rect 23427 715 23493 716
rect 33731 780 33797 781
rect 33731 716 33732 780
rect 33796 716 33797 780
rect 33731 715 33797 716
rect 50291 780 50357 781
rect 50291 716 50292 780
rect 50356 716 50357 780
rect 50291 715 50357 716
rect 52686 509 52746 1670
rect 53790 1670 53866 1730
rect 53790 1053 53850 1670
rect 53787 1052 53853 1053
rect 53787 988 53788 1052
rect 53852 988 53853 1052
rect 53787 987 53853 988
rect 54710 781 54770 2690
rect 54974 1730 55034 2380
rect 54974 1670 55138 1730
rect 54707 780 54773 781
rect 54707 716 54708 780
rect 54772 716 54773 780
rect 54707 715 54773 716
rect 55078 509 55138 1670
rect 83414 1461 83474 2730
rect 85944 2208 86264 3232
rect 85944 2144 85952 2208
rect 86016 2144 86032 2208
rect 86096 2144 86112 2208
rect 86176 2144 86192 2208
rect 86256 2144 86264 2208
rect 85944 2128 86264 2144
rect 87944 86528 88264 87552
rect 87944 86464 87952 86528
rect 88016 86464 88032 86528
rect 88096 86464 88112 86528
rect 88176 86464 88192 86528
rect 88256 86464 88264 86528
rect 87944 85440 88264 86464
rect 87944 85376 87952 85440
rect 88016 85376 88032 85440
rect 88096 85376 88112 85440
rect 88176 85376 88192 85440
rect 88256 85376 88264 85440
rect 87944 84352 88264 85376
rect 87944 84288 87952 84352
rect 88016 84288 88032 84352
rect 88096 84288 88112 84352
rect 88176 84288 88192 84352
rect 88256 84288 88264 84352
rect 87944 83264 88264 84288
rect 87944 83200 87952 83264
rect 88016 83200 88032 83264
rect 88096 83200 88112 83264
rect 88176 83200 88192 83264
rect 88256 83200 88264 83264
rect 87944 82176 88264 83200
rect 87944 82112 87952 82176
rect 88016 82112 88032 82176
rect 88096 82112 88112 82176
rect 88176 82112 88192 82176
rect 88256 82112 88264 82176
rect 87944 81088 88264 82112
rect 87944 81024 87952 81088
rect 88016 81024 88032 81088
rect 88096 81024 88112 81088
rect 88176 81024 88192 81088
rect 88256 81024 88264 81088
rect 87944 80576 88264 81024
rect 87944 80340 87986 80576
rect 88222 80340 88264 80576
rect 87944 80000 88264 80340
rect 87944 79936 87952 80000
rect 88016 79936 88032 80000
rect 88096 79936 88112 80000
rect 88176 79936 88192 80000
rect 88256 79936 88264 80000
rect 87944 78912 88264 79936
rect 87944 78848 87952 78912
rect 88016 78848 88032 78912
rect 88096 78848 88112 78912
rect 88176 78848 88192 78912
rect 88256 78848 88264 78912
rect 87944 77824 88264 78848
rect 87944 77760 87952 77824
rect 88016 77760 88032 77824
rect 88096 77760 88112 77824
rect 88176 77760 88192 77824
rect 88256 77760 88264 77824
rect 87944 76736 88264 77760
rect 87944 76672 87952 76736
rect 88016 76672 88032 76736
rect 88096 76672 88112 76736
rect 88176 76672 88192 76736
rect 88256 76672 88264 76736
rect 87944 75648 88264 76672
rect 87944 75584 87952 75648
rect 88016 75584 88032 75648
rect 88096 75584 88112 75648
rect 88176 75584 88192 75648
rect 88256 75584 88264 75648
rect 87944 74560 88264 75584
rect 87944 74496 87952 74560
rect 88016 74496 88032 74560
rect 88096 74496 88112 74560
rect 88176 74496 88192 74560
rect 88256 74496 88264 74560
rect 87944 73472 88264 74496
rect 87944 73408 87952 73472
rect 88016 73408 88032 73472
rect 88096 73408 88112 73472
rect 88176 73408 88192 73472
rect 88256 73408 88264 73472
rect 87944 72384 88264 73408
rect 87944 72320 87952 72384
rect 88016 72320 88032 72384
rect 88096 72320 88112 72384
rect 88176 72320 88192 72384
rect 88256 72320 88264 72384
rect 87944 71296 88264 72320
rect 87944 71232 87952 71296
rect 88016 71232 88032 71296
rect 88096 71232 88112 71296
rect 88176 71232 88192 71296
rect 88256 71232 88264 71296
rect 87944 70576 88264 71232
rect 87944 70340 87986 70576
rect 88222 70340 88264 70576
rect 87944 70208 88264 70340
rect 87944 70144 87952 70208
rect 88016 70144 88032 70208
rect 88096 70144 88112 70208
rect 88176 70144 88192 70208
rect 88256 70144 88264 70208
rect 87944 69120 88264 70144
rect 87944 69056 87952 69120
rect 88016 69056 88032 69120
rect 88096 69056 88112 69120
rect 88176 69056 88192 69120
rect 88256 69056 88264 69120
rect 87944 68032 88264 69056
rect 87944 67968 87952 68032
rect 88016 67968 88032 68032
rect 88096 67968 88112 68032
rect 88176 67968 88192 68032
rect 88256 67968 88264 68032
rect 87944 66944 88264 67968
rect 87944 66880 87952 66944
rect 88016 66880 88032 66944
rect 88096 66880 88112 66944
rect 88176 66880 88192 66944
rect 88256 66880 88264 66944
rect 87944 65856 88264 66880
rect 87944 65792 87952 65856
rect 88016 65792 88032 65856
rect 88096 65792 88112 65856
rect 88176 65792 88192 65856
rect 88256 65792 88264 65856
rect 87944 64768 88264 65792
rect 87944 64704 87952 64768
rect 88016 64704 88032 64768
rect 88096 64704 88112 64768
rect 88176 64704 88192 64768
rect 88256 64704 88264 64768
rect 87944 63680 88264 64704
rect 87944 63616 87952 63680
rect 88016 63616 88032 63680
rect 88096 63616 88112 63680
rect 88176 63616 88192 63680
rect 88256 63616 88264 63680
rect 87944 62592 88264 63616
rect 87944 62528 87952 62592
rect 88016 62528 88032 62592
rect 88096 62528 88112 62592
rect 88176 62528 88192 62592
rect 88256 62528 88264 62592
rect 87944 61504 88264 62528
rect 87944 61440 87952 61504
rect 88016 61440 88032 61504
rect 88096 61440 88112 61504
rect 88176 61440 88192 61504
rect 88256 61440 88264 61504
rect 87944 60576 88264 61440
rect 87944 60416 87986 60576
rect 88222 60416 88264 60576
rect 87944 60352 87952 60416
rect 88256 60352 88264 60416
rect 87944 60340 87986 60352
rect 88222 60340 88264 60352
rect 87944 59328 88264 60340
rect 87944 59264 87952 59328
rect 88016 59264 88032 59328
rect 88096 59264 88112 59328
rect 88176 59264 88192 59328
rect 88256 59264 88264 59328
rect 87944 58240 88264 59264
rect 87944 58176 87952 58240
rect 88016 58176 88032 58240
rect 88096 58176 88112 58240
rect 88176 58176 88192 58240
rect 88256 58176 88264 58240
rect 87944 57152 88264 58176
rect 87944 57088 87952 57152
rect 88016 57088 88032 57152
rect 88096 57088 88112 57152
rect 88176 57088 88192 57152
rect 88256 57088 88264 57152
rect 87944 56064 88264 57088
rect 87944 56000 87952 56064
rect 88016 56000 88032 56064
rect 88096 56000 88112 56064
rect 88176 56000 88192 56064
rect 88256 56000 88264 56064
rect 87944 54976 88264 56000
rect 87944 54912 87952 54976
rect 88016 54912 88032 54976
rect 88096 54912 88112 54976
rect 88176 54912 88192 54976
rect 88256 54912 88264 54976
rect 87944 53888 88264 54912
rect 87944 53824 87952 53888
rect 88016 53824 88032 53888
rect 88096 53824 88112 53888
rect 88176 53824 88192 53888
rect 88256 53824 88264 53888
rect 87944 52800 88264 53824
rect 87944 52736 87952 52800
rect 88016 52736 88032 52800
rect 88096 52736 88112 52800
rect 88176 52736 88192 52800
rect 88256 52736 88264 52800
rect 87944 51712 88264 52736
rect 87944 51648 87952 51712
rect 88016 51648 88032 51712
rect 88096 51648 88112 51712
rect 88176 51648 88192 51712
rect 88256 51648 88264 51712
rect 87944 50624 88264 51648
rect 87944 50560 87952 50624
rect 88016 50576 88032 50624
rect 88096 50576 88112 50624
rect 88176 50576 88192 50624
rect 88256 50560 88264 50624
rect 87944 50340 87986 50560
rect 88222 50340 88264 50560
rect 87944 49536 88264 50340
rect 87944 49472 87952 49536
rect 88016 49472 88032 49536
rect 88096 49472 88112 49536
rect 88176 49472 88192 49536
rect 88256 49472 88264 49536
rect 87944 48448 88264 49472
rect 87944 48384 87952 48448
rect 88016 48384 88032 48448
rect 88096 48384 88112 48448
rect 88176 48384 88192 48448
rect 88256 48384 88264 48448
rect 87944 47360 88264 48384
rect 87944 47296 87952 47360
rect 88016 47296 88032 47360
rect 88096 47296 88112 47360
rect 88176 47296 88192 47360
rect 88256 47296 88264 47360
rect 87944 46272 88264 47296
rect 87944 46208 87952 46272
rect 88016 46208 88032 46272
rect 88096 46208 88112 46272
rect 88176 46208 88192 46272
rect 88256 46208 88264 46272
rect 87944 45184 88264 46208
rect 87944 45120 87952 45184
rect 88016 45120 88032 45184
rect 88096 45120 88112 45184
rect 88176 45120 88192 45184
rect 88256 45120 88264 45184
rect 87944 44096 88264 45120
rect 87944 44032 87952 44096
rect 88016 44032 88032 44096
rect 88096 44032 88112 44096
rect 88176 44032 88192 44096
rect 88256 44032 88264 44096
rect 87944 43008 88264 44032
rect 87944 42944 87952 43008
rect 88016 42944 88032 43008
rect 88096 42944 88112 43008
rect 88176 42944 88192 43008
rect 88256 42944 88264 43008
rect 87944 41920 88264 42944
rect 87944 41856 87952 41920
rect 88016 41856 88032 41920
rect 88096 41856 88112 41920
rect 88176 41856 88192 41920
rect 88256 41856 88264 41920
rect 87944 40832 88264 41856
rect 87944 40768 87952 40832
rect 88016 40768 88032 40832
rect 88096 40768 88112 40832
rect 88176 40768 88192 40832
rect 88256 40768 88264 40832
rect 87944 40576 88264 40768
rect 87944 40340 87986 40576
rect 88222 40340 88264 40576
rect 87944 39744 88264 40340
rect 87944 39680 87952 39744
rect 88016 39680 88032 39744
rect 88096 39680 88112 39744
rect 88176 39680 88192 39744
rect 88256 39680 88264 39744
rect 87944 38656 88264 39680
rect 87944 38592 87952 38656
rect 88016 38592 88032 38656
rect 88096 38592 88112 38656
rect 88176 38592 88192 38656
rect 88256 38592 88264 38656
rect 87944 37568 88264 38592
rect 87944 37504 87952 37568
rect 88016 37504 88032 37568
rect 88096 37504 88112 37568
rect 88176 37504 88192 37568
rect 88256 37504 88264 37568
rect 87944 36480 88264 37504
rect 87944 36416 87952 36480
rect 88016 36416 88032 36480
rect 88096 36416 88112 36480
rect 88176 36416 88192 36480
rect 88256 36416 88264 36480
rect 87944 35392 88264 36416
rect 87944 35328 87952 35392
rect 88016 35328 88032 35392
rect 88096 35328 88112 35392
rect 88176 35328 88192 35392
rect 88256 35328 88264 35392
rect 87944 34304 88264 35328
rect 87944 34240 87952 34304
rect 88016 34240 88032 34304
rect 88096 34240 88112 34304
rect 88176 34240 88192 34304
rect 88256 34240 88264 34304
rect 87944 33216 88264 34240
rect 87944 33152 87952 33216
rect 88016 33152 88032 33216
rect 88096 33152 88112 33216
rect 88176 33152 88192 33216
rect 88256 33152 88264 33216
rect 87944 32128 88264 33152
rect 87944 32064 87952 32128
rect 88016 32064 88032 32128
rect 88096 32064 88112 32128
rect 88176 32064 88192 32128
rect 88256 32064 88264 32128
rect 87944 31040 88264 32064
rect 87944 30976 87952 31040
rect 88016 30976 88032 31040
rect 88096 30976 88112 31040
rect 88176 30976 88192 31040
rect 88256 30976 88264 31040
rect 87944 30576 88264 30976
rect 87944 30340 87986 30576
rect 88222 30340 88264 30576
rect 87944 29952 88264 30340
rect 87944 29888 87952 29952
rect 88016 29888 88032 29952
rect 88096 29888 88112 29952
rect 88176 29888 88192 29952
rect 88256 29888 88264 29952
rect 87944 28864 88264 29888
rect 87944 28800 87952 28864
rect 88016 28800 88032 28864
rect 88096 28800 88112 28864
rect 88176 28800 88192 28864
rect 88256 28800 88264 28864
rect 87944 27776 88264 28800
rect 87944 27712 87952 27776
rect 88016 27712 88032 27776
rect 88096 27712 88112 27776
rect 88176 27712 88192 27776
rect 88256 27712 88264 27776
rect 87944 26688 88264 27712
rect 87944 26624 87952 26688
rect 88016 26624 88032 26688
rect 88096 26624 88112 26688
rect 88176 26624 88192 26688
rect 88256 26624 88264 26688
rect 87944 25600 88264 26624
rect 87944 25536 87952 25600
rect 88016 25536 88032 25600
rect 88096 25536 88112 25600
rect 88176 25536 88192 25600
rect 88256 25536 88264 25600
rect 87944 24512 88264 25536
rect 87944 24448 87952 24512
rect 88016 24448 88032 24512
rect 88096 24448 88112 24512
rect 88176 24448 88192 24512
rect 88256 24448 88264 24512
rect 87944 23424 88264 24448
rect 87944 23360 87952 23424
rect 88016 23360 88032 23424
rect 88096 23360 88112 23424
rect 88176 23360 88192 23424
rect 88256 23360 88264 23424
rect 87944 22336 88264 23360
rect 87944 22272 87952 22336
rect 88016 22272 88032 22336
rect 88096 22272 88112 22336
rect 88176 22272 88192 22336
rect 88256 22272 88264 22336
rect 87944 21248 88264 22272
rect 87944 21184 87952 21248
rect 88016 21184 88032 21248
rect 88096 21184 88112 21248
rect 88176 21184 88192 21248
rect 88256 21184 88264 21248
rect 87944 20576 88264 21184
rect 87944 20340 87986 20576
rect 88222 20340 88264 20576
rect 87944 20160 88264 20340
rect 87944 20096 87952 20160
rect 88016 20096 88032 20160
rect 88096 20096 88112 20160
rect 88176 20096 88192 20160
rect 88256 20096 88264 20160
rect 87944 19072 88264 20096
rect 87944 19008 87952 19072
rect 88016 19008 88032 19072
rect 88096 19008 88112 19072
rect 88176 19008 88192 19072
rect 88256 19008 88264 19072
rect 87944 17984 88264 19008
rect 87944 17920 87952 17984
rect 88016 17920 88032 17984
rect 88096 17920 88112 17984
rect 88176 17920 88192 17984
rect 88256 17920 88264 17984
rect 87944 16896 88264 17920
rect 87944 16832 87952 16896
rect 88016 16832 88032 16896
rect 88096 16832 88112 16896
rect 88176 16832 88192 16896
rect 88256 16832 88264 16896
rect 87944 15808 88264 16832
rect 87944 15744 87952 15808
rect 88016 15744 88032 15808
rect 88096 15744 88112 15808
rect 88176 15744 88192 15808
rect 88256 15744 88264 15808
rect 87944 14720 88264 15744
rect 87944 14656 87952 14720
rect 88016 14656 88032 14720
rect 88096 14656 88112 14720
rect 88176 14656 88192 14720
rect 88256 14656 88264 14720
rect 87944 13632 88264 14656
rect 87944 13568 87952 13632
rect 88016 13568 88032 13632
rect 88096 13568 88112 13632
rect 88176 13568 88192 13632
rect 88256 13568 88264 13632
rect 87944 12544 88264 13568
rect 87944 12480 87952 12544
rect 88016 12480 88032 12544
rect 88096 12480 88112 12544
rect 88176 12480 88192 12544
rect 88256 12480 88264 12544
rect 87944 11456 88264 12480
rect 87944 11392 87952 11456
rect 88016 11392 88032 11456
rect 88096 11392 88112 11456
rect 88176 11392 88192 11456
rect 88256 11392 88264 11456
rect 87944 10576 88264 11392
rect 87944 10368 87986 10576
rect 88222 10368 88264 10576
rect 87944 10304 87952 10368
rect 88016 10304 88032 10340
rect 88096 10304 88112 10340
rect 88176 10304 88192 10340
rect 88256 10304 88264 10368
rect 87944 9280 88264 10304
rect 87944 9216 87952 9280
rect 88016 9216 88032 9280
rect 88096 9216 88112 9280
rect 88176 9216 88192 9280
rect 88256 9216 88264 9280
rect 87944 8192 88264 9216
rect 87944 8128 87952 8192
rect 88016 8128 88032 8192
rect 88096 8128 88112 8192
rect 88176 8128 88192 8192
rect 88256 8128 88264 8192
rect 87944 7104 88264 8128
rect 87944 7040 87952 7104
rect 88016 7040 88032 7104
rect 88096 7040 88112 7104
rect 88176 7040 88192 7104
rect 88256 7040 88264 7104
rect 87944 6016 88264 7040
rect 87944 5952 87952 6016
rect 88016 5952 88032 6016
rect 88096 5952 88112 6016
rect 88176 5952 88192 6016
rect 88256 5952 88264 6016
rect 87944 4928 88264 5952
rect 87944 4864 87952 4928
rect 88016 4864 88032 4928
rect 88096 4864 88112 4928
rect 88176 4864 88192 4928
rect 88256 4864 88264 4928
rect 87944 3840 88264 4864
rect 87944 3776 87952 3840
rect 88016 3776 88032 3840
rect 88096 3776 88112 3840
rect 88176 3776 88192 3840
rect 88256 3776 88264 3840
rect 87944 2752 88264 3776
rect 87944 2688 87952 2752
rect 88016 2688 88032 2752
rect 88096 2688 88112 2752
rect 88176 2688 88192 2752
rect 88256 2688 88264 2752
rect 87944 2128 88264 2688
rect 89944 92512 90264 93536
rect 89944 92448 89952 92512
rect 90016 92448 90032 92512
rect 90096 92448 90112 92512
rect 90176 92448 90192 92512
rect 90256 92448 90264 92512
rect 89944 91424 90264 92448
rect 89944 91360 89952 91424
rect 90016 91360 90032 91424
rect 90096 91360 90112 91424
rect 90176 91360 90192 91424
rect 90256 91360 90264 91424
rect 89944 90336 90264 91360
rect 89944 90272 89952 90336
rect 90016 90272 90032 90336
rect 90096 90272 90112 90336
rect 90176 90272 90192 90336
rect 90256 90272 90264 90336
rect 89944 89248 90264 90272
rect 89944 89184 89952 89248
rect 90016 89184 90032 89248
rect 90096 89184 90112 89248
rect 90176 89184 90192 89248
rect 90256 89184 90264 89248
rect 89944 88160 90264 89184
rect 89944 88096 89952 88160
rect 90016 88096 90032 88160
rect 90096 88096 90112 88160
rect 90176 88096 90192 88160
rect 90256 88096 90264 88160
rect 89944 87072 90264 88096
rect 89944 87008 89952 87072
rect 90016 87008 90032 87072
rect 90096 87008 90112 87072
rect 90176 87008 90192 87072
rect 90256 87008 90264 87072
rect 89944 85984 90264 87008
rect 89944 85920 89952 85984
rect 90016 85920 90032 85984
rect 90096 85920 90112 85984
rect 90176 85920 90192 85984
rect 90256 85920 90264 85984
rect 89944 85576 90264 85920
rect 89944 85340 89986 85576
rect 90222 85340 90264 85576
rect 89944 84896 90264 85340
rect 89944 84832 89952 84896
rect 90016 84832 90032 84896
rect 90096 84832 90112 84896
rect 90176 84832 90192 84896
rect 90256 84832 90264 84896
rect 89944 83808 90264 84832
rect 89944 83744 89952 83808
rect 90016 83744 90032 83808
rect 90096 83744 90112 83808
rect 90176 83744 90192 83808
rect 90256 83744 90264 83808
rect 89944 82720 90264 83744
rect 89944 82656 89952 82720
rect 90016 82656 90032 82720
rect 90096 82656 90112 82720
rect 90176 82656 90192 82720
rect 90256 82656 90264 82720
rect 89944 81632 90264 82656
rect 89944 81568 89952 81632
rect 90016 81568 90032 81632
rect 90096 81568 90112 81632
rect 90176 81568 90192 81632
rect 90256 81568 90264 81632
rect 89944 80544 90264 81568
rect 89944 80480 89952 80544
rect 90016 80480 90032 80544
rect 90096 80480 90112 80544
rect 90176 80480 90192 80544
rect 90256 80480 90264 80544
rect 89944 79456 90264 80480
rect 89944 79392 89952 79456
rect 90016 79392 90032 79456
rect 90096 79392 90112 79456
rect 90176 79392 90192 79456
rect 90256 79392 90264 79456
rect 89944 78368 90264 79392
rect 89944 78304 89952 78368
rect 90016 78304 90032 78368
rect 90096 78304 90112 78368
rect 90176 78304 90192 78368
rect 90256 78304 90264 78368
rect 89944 77280 90264 78304
rect 89944 77216 89952 77280
rect 90016 77216 90032 77280
rect 90096 77216 90112 77280
rect 90176 77216 90192 77280
rect 90256 77216 90264 77280
rect 89944 76192 90264 77216
rect 89944 76128 89952 76192
rect 90016 76128 90032 76192
rect 90096 76128 90112 76192
rect 90176 76128 90192 76192
rect 90256 76128 90264 76192
rect 89944 75576 90264 76128
rect 89944 75340 89986 75576
rect 90222 75340 90264 75576
rect 89944 75104 90264 75340
rect 89944 75040 89952 75104
rect 90016 75040 90032 75104
rect 90096 75040 90112 75104
rect 90176 75040 90192 75104
rect 90256 75040 90264 75104
rect 89944 74016 90264 75040
rect 89944 73952 89952 74016
rect 90016 73952 90032 74016
rect 90096 73952 90112 74016
rect 90176 73952 90192 74016
rect 90256 73952 90264 74016
rect 89944 72928 90264 73952
rect 89944 72864 89952 72928
rect 90016 72864 90032 72928
rect 90096 72864 90112 72928
rect 90176 72864 90192 72928
rect 90256 72864 90264 72928
rect 89944 71840 90264 72864
rect 89944 71776 89952 71840
rect 90016 71776 90032 71840
rect 90096 71776 90112 71840
rect 90176 71776 90192 71840
rect 90256 71776 90264 71840
rect 89944 70752 90264 71776
rect 89944 70688 89952 70752
rect 90016 70688 90032 70752
rect 90096 70688 90112 70752
rect 90176 70688 90192 70752
rect 90256 70688 90264 70752
rect 89944 69664 90264 70688
rect 89944 69600 89952 69664
rect 90016 69600 90032 69664
rect 90096 69600 90112 69664
rect 90176 69600 90192 69664
rect 90256 69600 90264 69664
rect 89944 68576 90264 69600
rect 89944 68512 89952 68576
rect 90016 68512 90032 68576
rect 90096 68512 90112 68576
rect 90176 68512 90192 68576
rect 90256 68512 90264 68576
rect 89944 67488 90264 68512
rect 89944 67424 89952 67488
rect 90016 67424 90032 67488
rect 90096 67424 90112 67488
rect 90176 67424 90192 67488
rect 90256 67424 90264 67488
rect 89944 66400 90264 67424
rect 89944 66336 89952 66400
rect 90016 66336 90032 66400
rect 90096 66336 90112 66400
rect 90176 66336 90192 66400
rect 90256 66336 90264 66400
rect 89944 65576 90264 66336
rect 89944 65340 89986 65576
rect 90222 65340 90264 65576
rect 89944 65312 90264 65340
rect 89944 65248 89952 65312
rect 90016 65248 90032 65312
rect 90096 65248 90112 65312
rect 90176 65248 90192 65312
rect 90256 65248 90264 65312
rect 89944 64224 90264 65248
rect 89944 64160 89952 64224
rect 90016 64160 90032 64224
rect 90096 64160 90112 64224
rect 90176 64160 90192 64224
rect 90256 64160 90264 64224
rect 89944 63136 90264 64160
rect 89944 63072 89952 63136
rect 90016 63072 90032 63136
rect 90096 63072 90112 63136
rect 90176 63072 90192 63136
rect 90256 63072 90264 63136
rect 89944 62048 90264 63072
rect 89944 61984 89952 62048
rect 90016 61984 90032 62048
rect 90096 61984 90112 62048
rect 90176 61984 90192 62048
rect 90256 61984 90264 62048
rect 89944 60960 90264 61984
rect 89944 60896 89952 60960
rect 90016 60896 90032 60960
rect 90096 60896 90112 60960
rect 90176 60896 90192 60960
rect 90256 60896 90264 60960
rect 89944 59872 90264 60896
rect 89944 59808 89952 59872
rect 90016 59808 90032 59872
rect 90096 59808 90112 59872
rect 90176 59808 90192 59872
rect 90256 59808 90264 59872
rect 89944 58784 90264 59808
rect 89944 58720 89952 58784
rect 90016 58720 90032 58784
rect 90096 58720 90112 58784
rect 90176 58720 90192 58784
rect 90256 58720 90264 58784
rect 89944 57696 90264 58720
rect 89944 57632 89952 57696
rect 90016 57632 90032 57696
rect 90096 57632 90112 57696
rect 90176 57632 90192 57696
rect 90256 57632 90264 57696
rect 89944 56608 90264 57632
rect 89944 56544 89952 56608
rect 90016 56544 90032 56608
rect 90096 56544 90112 56608
rect 90176 56544 90192 56608
rect 90256 56544 90264 56608
rect 89944 55576 90264 56544
rect 89944 55520 89986 55576
rect 90222 55520 90264 55576
rect 89944 55456 89952 55520
rect 90256 55456 90264 55520
rect 89944 55340 89986 55456
rect 90222 55340 90264 55456
rect 89944 54432 90264 55340
rect 89944 54368 89952 54432
rect 90016 54368 90032 54432
rect 90096 54368 90112 54432
rect 90176 54368 90192 54432
rect 90256 54368 90264 54432
rect 89944 53344 90264 54368
rect 89944 53280 89952 53344
rect 90016 53280 90032 53344
rect 90096 53280 90112 53344
rect 90176 53280 90192 53344
rect 90256 53280 90264 53344
rect 89944 52256 90264 53280
rect 89944 52192 89952 52256
rect 90016 52192 90032 52256
rect 90096 52192 90112 52256
rect 90176 52192 90192 52256
rect 90256 52192 90264 52256
rect 89944 51168 90264 52192
rect 89944 51104 89952 51168
rect 90016 51104 90032 51168
rect 90096 51104 90112 51168
rect 90176 51104 90192 51168
rect 90256 51104 90264 51168
rect 89944 50080 90264 51104
rect 89944 50016 89952 50080
rect 90016 50016 90032 50080
rect 90096 50016 90112 50080
rect 90176 50016 90192 50080
rect 90256 50016 90264 50080
rect 89944 48992 90264 50016
rect 89944 48928 89952 48992
rect 90016 48928 90032 48992
rect 90096 48928 90112 48992
rect 90176 48928 90192 48992
rect 90256 48928 90264 48992
rect 89944 47904 90264 48928
rect 89944 47840 89952 47904
rect 90016 47840 90032 47904
rect 90096 47840 90112 47904
rect 90176 47840 90192 47904
rect 90256 47840 90264 47904
rect 89944 46816 90264 47840
rect 89944 46752 89952 46816
rect 90016 46752 90032 46816
rect 90096 46752 90112 46816
rect 90176 46752 90192 46816
rect 90256 46752 90264 46816
rect 89944 45728 90264 46752
rect 89944 45664 89952 45728
rect 90016 45664 90032 45728
rect 90096 45664 90112 45728
rect 90176 45664 90192 45728
rect 90256 45664 90264 45728
rect 89944 45576 90264 45664
rect 89944 45340 89986 45576
rect 90222 45340 90264 45576
rect 89944 44640 90264 45340
rect 89944 44576 89952 44640
rect 90016 44576 90032 44640
rect 90096 44576 90112 44640
rect 90176 44576 90192 44640
rect 90256 44576 90264 44640
rect 89944 43552 90264 44576
rect 89944 43488 89952 43552
rect 90016 43488 90032 43552
rect 90096 43488 90112 43552
rect 90176 43488 90192 43552
rect 90256 43488 90264 43552
rect 89944 42464 90264 43488
rect 89944 42400 89952 42464
rect 90016 42400 90032 42464
rect 90096 42400 90112 42464
rect 90176 42400 90192 42464
rect 90256 42400 90264 42464
rect 89944 41376 90264 42400
rect 89944 41312 89952 41376
rect 90016 41312 90032 41376
rect 90096 41312 90112 41376
rect 90176 41312 90192 41376
rect 90256 41312 90264 41376
rect 89944 40288 90264 41312
rect 89944 40224 89952 40288
rect 90016 40224 90032 40288
rect 90096 40224 90112 40288
rect 90176 40224 90192 40288
rect 90256 40224 90264 40288
rect 89944 39200 90264 40224
rect 89944 39136 89952 39200
rect 90016 39136 90032 39200
rect 90096 39136 90112 39200
rect 90176 39136 90192 39200
rect 90256 39136 90264 39200
rect 89944 38112 90264 39136
rect 89944 38048 89952 38112
rect 90016 38048 90032 38112
rect 90096 38048 90112 38112
rect 90176 38048 90192 38112
rect 90256 38048 90264 38112
rect 89944 37024 90264 38048
rect 89944 36960 89952 37024
rect 90016 36960 90032 37024
rect 90096 36960 90112 37024
rect 90176 36960 90192 37024
rect 90256 36960 90264 37024
rect 89944 35936 90264 36960
rect 89944 35872 89952 35936
rect 90016 35872 90032 35936
rect 90096 35872 90112 35936
rect 90176 35872 90192 35936
rect 90256 35872 90264 35936
rect 89944 35576 90264 35872
rect 89944 35340 89986 35576
rect 90222 35340 90264 35576
rect 89944 34848 90264 35340
rect 89944 34784 89952 34848
rect 90016 34784 90032 34848
rect 90096 34784 90112 34848
rect 90176 34784 90192 34848
rect 90256 34784 90264 34848
rect 89944 33760 90264 34784
rect 89944 33696 89952 33760
rect 90016 33696 90032 33760
rect 90096 33696 90112 33760
rect 90176 33696 90192 33760
rect 90256 33696 90264 33760
rect 89944 32672 90264 33696
rect 89944 32608 89952 32672
rect 90016 32608 90032 32672
rect 90096 32608 90112 32672
rect 90176 32608 90192 32672
rect 90256 32608 90264 32672
rect 89944 31584 90264 32608
rect 89944 31520 89952 31584
rect 90016 31520 90032 31584
rect 90096 31520 90112 31584
rect 90176 31520 90192 31584
rect 90256 31520 90264 31584
rect 89944 30496 90264 31520
rect 89944 30432 89952 30496
rect 90016 30432 90032 30496
rect 90096 30432 90112 30496
rect 90176 30432 90192 30496
rect 90256 30432 90264 30496
rect 89944 29408 90264 30432
rect 89944 29344 89952 29408
rect 90016 29344 90032 29408
rect 90096 29344 90112 29408
rect 90176 29344 90192 29408
rect 90256 29344 90264 29408
rect 89944 28320 90264 29344
rect 89944 28256 89952 28320
rect 90016 28256 90032 28320
rect 90096 28256 90112 28320
rect 90176 28256 90192 28320
rect 90256 28256 90264 28320
rect 89944 27232 90264 28256
rect 89944 27168 89952 27232
rect 90016 27168 90032 27232
rect 90096 27168 90112 27232
rect 90176 27168 90192 27232
rect 90256 27168 90264 27232
rect 89944 26144 90264 27168
rect 89944 26080 89952 26144
rect 90016 26080 90032 26144
rect 90096 26080 90112 26144
rect 90176 26080 90192 26144
rect 90256 26080 90264 26144
rect 89944 25576 90264 26080
rect 89944 25340 89986 25576
rect 90222 25340 90264 25576
rect 89944 25056 90264 25340
rect 89944 24992 89952 25056
rect 90016 24992 90032 25056
rect 90096 24992 90112 25056
rect 90176 24992 90192 25056
rect 90256 24992 90264 25056
rect 89944 23968 90264 24992
rect 89944 23904 89952 23968
rect 90016 23904 90032 23968
rect 90096 23904 90112 23968
rect 90176 23904 90192 23968
rect 90256 23904 90264 23968
rect 89944 22880 90264 23904
rect 89944 22816 89952 22880
rect 90016 22816 90032 22880
rect 90096 22816 90112 22880
rect 90176 22816 90192 22880
rect 90256 22816 90264 22880
rect 89944 21792 90264 22816
rect 89944 21728 89952 21792
rect 90016 21728 90032 21792
rect 90096 21728 90112 21792
rect 90176 21728 90192 21792
rect 90256 21728 90264 21792
rect 89944 20704 90264 21728
rect 89944 20640 89952 20704
rect 90016 20640 90032 20704
rect 90096 20640 90112 20704
rect 90176 20640 90192 20704
rect 90256 20640 90264 20704
rect 89944 19616 90264 20640
rect 89944 19552 89952 19616
rect 90016 19552 90032 19616
rect 90096 19552 90112 19616
rect 90176 19552 90192 19616
rect 90256 19552 90264 19616
rect 89944 18528 90264 19552
rect 89944 18464 89952 18528
rect 90016 18464 90032 18528
rect 90096 18464 90112 18528
rect 90176 18464 90192 18528
rect 90256 18464 90264 18528
rect 89944 17440 90264 18464
rect 89944 17376 89952 17440
rect 90016 17376 90032 17440
rect 90096 17376 90112 17440
rect 90176 17376 90192 17440
rect 90256 17376 90264 17440
rect 89944 16352 90264 17376
rect 89944 16288 89952 16352
rect 90016 16288 90032 16352
rect 90096 16288 90112 16352
rect 90176 16288 90192 16352
rect 90256 16288 90264 16352
rect 89944 15576 90264 16288
rect 89944 15340 89986 15576
rect 90222 15340 90264 15576
rect 89944 15264 90264 15340
rect 89944 15200 89952 15264
rect 90016 15200 90032 15264
rect 90096 15200 90112 15264
rect 90176 15200 90192 15264
rect 90256 15200 90264 15264
rect 89944 14176 90264 15200
rect 89944 14112 89952 14176
rect 90016 14112 90032 14176
rect 90096 14112 90112 14176
rect 90176 14112 90192 14176
rect 90256 14112 90264 14176
rect 89944 13088 90264 14112
rect 89944 13024 89952 13088
rect 90016 13024 90032 13088
rect 90096 13024 90112 13088
rect 90176 13024 90192 13088
rect 90256 13024 90264 13088
rect 89944 12000 90264 13024
rect 89944 11936 89952 12000
rect 90016 11936 90032 12000
rect 90096 11936 90112 12000
rect 90176 11936 90192 12000
rect 90256 11936 90264 12000
rect 89944 10912 90264 11936
rect 89944 10848 89952 10912
rect 90016 10848 90032 10912
rect 90096 10848 90112 10912
rect 90176 10848 90192 10912
rect 90256 10848 90264 10912
rect 89944 9824 90264 10848
rect 89944 9760 89952 9824
rect 90016 9760 90032 9824
rect 90096 9760 90112 9824
rect 90176 9760 90192 9824
rect 90256 9760 90264 9824
rect 89944 8736 90264 9760
rect 89944 8672 89952 8736
rect 90016 8672 90032 8736
rect 90096 8672 90112 8736
rect 90176 8672 90192 8736
rect 90256 8672 90264 8736
rect 89944 7648 90264 8672
rect 89944 7584 89952 7648
rect 90016 7584 90032 7648
rect 90096 7584 90112 7648
rect 90176 7584 90192 7648
rect 90256 7584 90264 7648
rect 89944 6560 90264 7584
rect 89944 6496 89952 6560
rect 90016 6496 90032 6560
rect 90096 6496 90112 6560
rect 90176 6496 90192 6560
rect 90256 6496 90264 6560
rect 89944 5576 90264 6496
rect 89944 5472 89986 5576
rect 90222 5472 90264 5576
rect 89944 5408 89952 5472
rect 90256 5408 90264 5472
rect 89944 5340 89986 5408
rect 90222 5340 90264 5408
rect 89944 4384 90264 5340
rect 89944 4320 89952 4384
rect 90016 4320 90032 4384
rect 90096 4320 90112 4384
rect 90176 4320 90192 4384
rect 90256 4320 90264 4384
rect 89944 3296 90264 4320
rect 89944 3232 89952 3296
rect 90016 3232 90032 3296
rect 90096 3232 90112 3296
rect 90176 3232 90192 3296
rect 90256 3232 90264 3296
rect 89944 2208 90264 3232
rect 89944 2144 89952 2208
rect 90016 2144 90032 2208
rect 90096 2144 90112 2208
rect 90176 2144 90192 2208
rect 90256 2144 90264 2208
rect 89944 2128 90264 2144
rect 83411 1460 83477 1461
rect 83411 1396 83412 1460
rect 83476 1396 83477 1460
rect 83411 1395 83477 1396
rect 52683 508 52749 509
rect 52683 444 52684 508
rect 52748 444 52749 508
rect 52683 443 52749 444
rect 55075 508 55141 509
rect 55075 444 55076 508
rect 55140 444 55141 508
rect 55075 443 55141 444
rect 19931 236 19997 237
rect 19931 172 19932 236
rect 19996 172 19997 236
rect 19931 171 19997 172
<< via4 >>
rect 1986 185340 2222 185576
rect 1986 175340 2222 175576
rect 1986 165408 2222 165576
rect 1986 165344 2016 165408
rect 2016 165344 2032 165408
rect 2032 165344 2096 165408
rect 2096 165344 2112 165408
rect 2112 165344 2176 165408
rect 2176 165344 2192 165408
rect 2192 165344 2222 165408
rect 1986 165340 2222 165344
rect 1986 155552 2016 155576
rect 2016 155552 2032 155576
rect 2032 155552 2096 155576
rect 2096 155552 2112 155576
rect 2112 155552 2176 155576
rect 2176 155552 2192 155576
rect 2192 155552 2222 155576
rect 1986 155340 2222 155552
rect 1986 145340 2222 145576
rect 1986 135340 2222 135576
rect 1986 125340 2222 125576
rect 1986 115360 2222 115576
rect 1986 115340 2016 115360
rect 2016 115340 2032 115360
rect 2032 115340 2096 115360
rect 2096 115340 2112 115360
rect 2112 115340 2176 115360
rect 2176 115340 2192 115360
rect 2192 115340 2222 115360
rect 1986 105568 2222 105576
rect 1986 105504 2016 105568
rect 2016 105504 2032 105568
rect 2032 105504 2096 105568
rect 2096 105504 2112 105568
rect 2112 105504 2176 105568
rect 2176 105504 2192 105568
rect 2192 105504 2222 105568
rect 1986 105340 2222 105504
rect 1986 95340 2222 95576
rect 1986 85340 2222 85576
rect 1986 75340 2222 75576
rect 1986 65340 2222 65576
rect 1986 55520 2222 55576
rect 1986 55456 2016 55520
rect 2016 55456 2032 55520
rect 2032 55456 2096 55520
rect 2096 55456 2112 55520
rect 2112 55456 2176 55520
rect 2176 55456 2192 55520
rect 2192 55456 2222 55520
rect 1986 55340 2222 55456
rect 1986 45340 2222 45576
rect 1986 35340 2222 35576
rect 1986 25340 2222 25576
rect 1986 15340 2222 15576
rect 1986 5472 2222 5576
rect 1986 5408 2016 5472
rect 2016 5408 2032 5472
rect 2032 5408 2096 5472
rect 2096 5408 2112 5472
rect 2112 5408 2176 5472
rect 2176 5408 2192 5472
rect 2192 5408 2222 5472
rect 1986 5340 2222 5408
rect 85986 185340 86222 185576
rect 3986 180340 4222 180576
rect 82982 180340 83218 180576
rect 82536 175340 82772 175576
rect 3986 170340 4222 170576
rect 82982 170340 83218 170576
rect 82536 165340 82772 165576
rect 3986 160512 4222 160576
rect 3986 160448 4016 160512
rect 4016 160448 4032 160512
rect 4032 160448 4096 160512
rect 4096 160448 4112 160512
rect 4112 160448 4176 160512
rect 4176 160448 4192 160512
rect 4192 160448 4222 160512
rect 3986 160340 4222 160448
rect 82982 160340 83218 160576
rect 82536 155340 82772 155576
rect 3986 150340 4222 150576
rect 82982 150340 83218 150576
rect 82536 145340 82772 145576
rect 3986 140340 4222 140576
rect 82982 140340 83218 140576
rect 82536 135340 82772 135576
rect 85986 175340 86222 175576
rect 3986 130340 4222 130576
rect 82982 130340 83218 130576
rect 6046 126022 6282 126258
rect 82536 125340 82772 125576
rect 3986 120340 4222 120576
rect 82982 120340 83218 120576
rect 5310 116652 5546 116738
rect 5310 116588 5396 116652
rect 5396 116588 5460 116652
rect 5460 116588 5546 116652
rect 5310 116502 5546 116588
rect 82536 115340 82772 115576
rect 3986 110464 4222 110576
rect 3986 110400 4016 110464
rect 4016 110400 4032 110464
rect 4032 110400 4096 110464
rect 4096 110400 4112 110464
rect 4112 110400 4176 110464
rect 4176 110400 4192 110464
rect 4192 110400 4222 110464
rect 3986 110340 4222 110400
rect 82982 110340 83218 110576
rect 82536 105340 82772 105576
rect 3986 100340 4222 100576
rect 82982 100340 83218 100576
rect 53150 96782 53386 97018
rect 54070 96932 54306 97018
rect 54070 96868 54156 96932
rect 54156 96868 54220 96932
rect 54220 96868 54306 96932
rect 54070 96782 54306 96868
rect 4390 94062 4626 94298
rect 3986 90340 4222 90576
rect 3986 80340 4222 80576
rect 3986 70340 4222 70576
rect 3986 60416 4222 60576
rect 3986 60352 4016 60416
rect 4016 60352 4032 60416
rect 4032 60352 4096 60416
rect 4096 60352 4112 60416
rect 4112 60352 4176 60416
rect 4176 60352 4192 60416
rect 4192 60352 4222 60416
rect 3986 60340 4222 60352
rect 3986 50560 4016 50576
rect 4016 50560 4032 50576
rect 4032 50560 4096 50576
rect 4096 50560 4112 50576
rect 4112 50560 4176 50576
rect 4176 50560 4192 50576
rect 4192 50560 4222 50576
rect 3986 50340 4222 50560
rect 3986 40340 4222 40576
rect 3986 30340 4222 30576
rect 3986 20340 4222 20576
rect 3986 10368 4222 10576
rect 3986 10340 4016 10368
rect 4016 10340 4032 10368
rect 4032 10340 4096 10368
rect 4096 10340 4112 10368
rect 4112 10340 4176 10368
rect 4176 10340 4192 10368
rect 4192 10340 4222 10368
rect 48182 93604 48268 93618
rect 48268 93604 48332 93618
rect 48332 93604 48418 93618
rect 48182 93382 48418 93604
rect 50942 96324 51028 96338
rect 51028 96324 51092 96338
rect 51092 96324 51178 96338
rect 50942 96102 51178 96324
rect 53150 93604 53236 93618
rect 53236 93604 53300 93618
rect 53300 93604 53386 93618
rect 53150 93382 53386 93604
rect 57980 93382 58216 93618
rect 59406 93382 59642 93618
rect 60878 94062 61114 94298
rect 60510 93382 60746 93618
rect 76702 94062 76938 94298
rect 77438 94062 77674 94298
rect 85986 165408 86222 165576
rect 85986 165344 86016 165408
rect 86016 165344 86032 165408
rect 86032 165344 86096 165408
rect 86096 165344 86112 165408
rect 86112 165344 86176 165408
rect 86176 165344 86192 165408
rect 86192 165344 86222 165408
rect 85986 165340 86222 165344
rect 84430 126022 84666 126258
rect 49286 93042 49522 93278
rect 4758 91342 4994 91578
rect 82982 90340 83218 90576
rect 5494 89302 5730 89538
rect 5126 88772 5362 88858
rect 5126 88708 5212 88772
rect 5212 88708 5276 88772
rect 5276 88708 5362 88772
rect 5126 88622 5362 88708
rect 5310 86732 5546 86818
rect 5310 86668 5396 86732
rect 5396 86668 5460 86732
rect 5460 86668 5546 86732
rect 5310 86582 5546 86668
rect 82536 85340 82772 85576
rect 82982 80340 83218 80576
rect 82536 75340 82772 75576
rect 82982 70340 83218 70576
rect 82536 65340 82772 65576
rect 82982 60340 83218 60576
rect 82536 55340 82772 55576
rect 82982 50340 83218 50576
rect 85986 155552 86016 155576
rect 86016 155552 86032 155576
rect 86032 155552 86096 155576
rect 86096 155552 86112 155576
rect 86112 155552 86176 155576
rect 86176 155552 86192 155576
rect 86192 155552 86222 155576
rect 85986 155340 86222 155552
rect 85986 145340 86222 145576
rect 85986 135340 86222 135576
rect 85986 125340 86222 125576
rect 85986 115360 86222 115576
rect 85986 115340 86016 115360
rect 86016 115340 86032 115360
rect 86032 115340 86096 115360
rect 86096 115340 86112 115360
rect 86112 115340 86176 115360
rect 86176 115340 86192 115360
rect 86192 115340 86222 115360
rect 85986 105568 86222 105576
rect 85986 105504 86016 105568
rect 86016 105504 86032 105568
rect 86032 105504 86096 105568
rect 86096 105504 86112 105568
rect 86112 105504 86176 105568
rect 86176 105504 86192 105568
rect 86192 105504 86222 105568
rect 85986 105340 86222 105504
rect 85986 95340 86222 95576
rect 87006 96782 87242 97018
rect 87986 180340 88222 180576
rect 87986 170340 88222 170576
rect 87986 160512 88222 160576
rect 87986 160448 88016 160512
rect 88016 160448 88032 160512
rect 88032 160448 88096 160512
rect 88096 160448 88112 160512
rect 88112 160448 88176 160512
rect 88176 160448 88192 160512
rect 88192 160448 88222 160512
rect 87986 160340 88222 160448
rect 87986 150340 88222 150576
rect 87986 140340 88222 140576
rect 87986 130340 88222 130576
rect 87986 120340 88222 120576
rect 87986 110464 88222 110576
rect 87986 110400 88016 110464
rect 88016 110400 88032 110464
rect 88032 110400 88096 110464
rect 88096 110400 88112 110464
rect 88112 110400 88176 110464
rect 88176 110400 88192 110464
rect 88192 110400 88222 110464
rect 87986 110340 88222 110400
rect 87986 100340 88222 100576
rect 89986 185340 90222 185576
rect 89986 175340 90222 175576
rect 89986 165408 90222 165576
rect 89986 165344 90016 165408
rect 90016 165344 90032 165408
rect 90032 165344 90096 165408
rect 90096 165344 90112 165408
rect 90112 165344 90176 165408
rect 90176 165344 90192 165408
rect 90192 165344 90222 165408
rect 89986 165340 90222 165344
rect 89986 155552 90016 155576
rect 90016 155552 90032 155576
rect 90032 155552 90096 155576
rect 90096 155552 90112 155576
rect 90112 155552 90176 155576
rect 90176 155552 90192 155576
rect 90192 155552 90222 155576
rect 89986 155340 90222 155552
rect 89986 145340 90222 145576
rect 89986 135340 90222 135576
rect 89986 125340 90222 125576
rect 90502 116502 90738 116738
rect 89986 115360 90222 115576
rect 89986 115340 90016 115360
rect 90016 115340 90032 115360
rect 90032 115340 90096 115360
rect 90096 115340 90112 115360
rect 90112 115340 90176 115360
rect 90176 115340 90192 115360
rect 90192 115340 90222 115360
rect 88662 96102 88898 96338
rect 88662 93382 88898 93618
rect 84614 92022 84850 92258
rect 86822 91342 87058 91578
rect 86822 89302 87058 89538
rect 86822 88622 87058 88858
rect 89986 105568 90222 105576
rect 89986 105504 90016 105568
rect 90016 105504 90032 105568
rect 90032 105504 90096 105568
rect 90096 105504 90112 105568
rect 90112 105504 90176 105568
rect 90176 105504 90192 105568
rect 90192 105504 90222 105568
rect 89986 105340 90222 105504
rect 90502 97462 90738 97698
rect 89986 95340 90222 95576
rect 89582 94062 89818 94298
rect 89030 92702 89266 92938
rect 87986 90340 88222 90576
rect 87190 86582 87426 86818
rect 85986 85340 86222 85576
rect 85986 75340 86222 75576
rect 85986 65340 86222 65576
rect 85986 55520 86222 55576
rect 85986 55456 86016 55520
rect 86016 55456 86032 55520
rect 86032 55456 86096 55520
rect 86096 55456 86112 55520
rect 86112 55456 86176 55520
rect 86176 55456 86192 55520
rect 86192 55456 86222 55520
rect 85986 55340 86222 55456
rect 82536 45340 82772 45576
rect 82982 40340 83218 40576
rect 82536 35340 82772 35576
rect 85986 45340 86222 45576
rect 82982 30340 83218 30576
rect 85986 35340 86222 35576
rect 82536 25340 82772 25576
rect 82982 20340 83218 20576
rect 82536 15340 82772 15576
rect 82982 10340 83218 10576
rect 82536 5340 82772 5576
rect 4758 3844 4844 3858
rect 4844 3844 4908 3858
rect 4908 3844 4994 3858
rect 4758 3622 4994 3844
rect 8070 2942 8306 3178
rect 36958 2942 37194 3178
rect 41374 2942 41610 3178
rect 85986 25340 86222 25576
rect 85986 15340 86222 15576
rect 85986 5472 86222 5576
rect 85986 5408 86016 5472
rect 86016 5408 86032 5472
rect 86032 5408 86096 5472
rect 86096 5408 86112 5472
rect 86112 5408 86176 5472
rect 86176 5408 86192 5472
rect 86192 5408 86222 5472
rect 85986 5340 86222 5408
rect 87986 80340 88222 80576
rect 87986 70340 88222 70576
rect 87986 60416 88222 60576
rect 87986 60352 88016 60416
rect 88016 60352 88032 60416
rect 88032 60352 88096 60416
rect 88096 60352 88112 60416
rect 88112 60352 88176 60416
rect 88176 60352 88192 60416
rect 88192 60352 88222 60416
rect 87986 60340 88222 60352
rect 87986 50560 88016 50576
rect 88016 50560 88032 50576
rect 88032 50560 88096 50576
rect 88096 50560 88112 50576
rect 88112 50560 88176 50576
rect 88176 50560 88192 50576
rect 88192 50560 88222 50576
rect 87986 50340 88222 50560
rect 87986 40340 88222 40576
rect 87986 30340 88222 30576
rect 87986 20340 88222 20576
rect 87986 10368 88222 10576
rect 87986 10340 88016 10368
rect 88016 10340 88032 10368
rect 88032 10340 88096 10368
rect 88096 10340 88112 10368
rect 88112 10340 88176 10368
rect 88176 10340 88192 10368
rect 88192 10340 88222 10368
rect 89986 85340 90222 85576
rect 89986 75340 90222 75576
rect 89986 65340 90222 65576
rect 89986 55520 90222 55576
rect 89986 55456 90016 55520
rect 90016 55456 90032 55520
rect 90032 55456 90096 55520
rect 90096 55456 90112 55520
rect 90112 55456 90176 55520
rect 90176 55456 90192 55520
rect 90192 55456 90222 55520
rect 89986 55340 90222 55456
rect 89986 45340 90222 45576
rect 89986 35340 90222 35576
rect 89986 25340 90222 25576
rect 89986 15340 90222 15576
rect 89986 5472 90222 5576
rect 89986 5408 90016 5472
rect 90016 5408 90032 5472
rect 90032 5408 90096 5472
rect 90096 5408 90112 5472
rect 90112 5408 90176 5472
rect 90176 5408 90192 5472
rect 90192 5408 90222 5472
rect 89986 5340 90222 5408
<< metal5 >>
rect 1104 185576 90896 185618
rect 1104 185340 1986 185576
rect 2222 185340 85986 185576
rect 86222 185340 89986 185576
rect 90222 185340 90896 185576
rect 1104 185298 90896 185340
rect 1104 180576 90896 180618
rect 1104 180340 3986 180576
rect 4222 180340 82982 180576
rect 83218 180340 87986 180576
rect 88222 180340 90896 180576
rect 1104 180298 90896 180340
rect 1104 175576 90896 175618
rect 1104 175340 1986 175576
rect 2222 175340 82536 175576
rect 82772 175340 85986 175576
rect 86222 175340 89986 175576
rect 90222 175340 90896 175576
rect 1104 175298 90896 175340
rect 1104 170576 90896 170618
rect 1104 170340 3986 170576
rect 4222 170340 82982 170576
rect 83218 170340 87986 170576
rect 88222 170340 90896 170576
rect 1104 170298 90896 170340
rect 1104 165576 90896 165618
rect 1104 165340 1986 165576
rect 2222 165340 82536 165576
rect 82772 165340 85986 165576
rect 86222 165340 89986 165576
rect 90222 165340 90896 165576
rect 1104 165298 90896 165340
rect 1104 160576 90896 160618
rect 1104 160340 3986 160576
rect 4222 160340 82982 160576
rect 83218 160340 87986 160576
rect 88222 160340 90896 160576
rect 1104 160298 90896 160340
rect 1104 155576 90896 155618
rect 1104 155340 1986 155576
rect 2222 155340 82536 155576
rect 82772 155340 85986 155576
rect 86222 155340 89986 155576
rect 90222 155340 90896 155576
rect 1104 155298 90896 155340
rect 1104 150576 90896 150618
rect 1104 150340 3986 150576
rect 4222 150340 82982 150576
rect 83218 150340 87986 150576
rect 88222 150340 90896 150576
rect 1104 150298 90896 150340
rect 1104 145576 90896 145618
rect 1104 145340 1986 145576
rect 2222 145340 82536 145576
rect 82772 145340 85986 145576
rect 86222 145340 89986 145576
rect 90222 145340 90896 145576
rect 1104 145298 90896 145340
rect 1104 140576 90896 140618
rect 1104 140340 3986 140576
rect 4222 140340 82982 140576
rect 83218 140340 87986 140576
rect 88222 140340 90896 140576
rect 1104 140298 90896 140340
rect 1104 135576 90896 135618
rect 1104 135340 1986 135576
rect 2222 135340 82536 135576
rect 82772 135340 85986 135576
rect 86222 135340 89986 135576
rect 90222 135340 90896 135576
rect 1104 135298 90896 135340
rect 1104 130576 90896 130618
rect 1104 130340 3986 130576
rect 4222 130340 82982 130576
rect 83218 130340 87986 130576
rect 88222 130340 90896 130576
rect 1104 130298 90896 130340
rect 6004 126258 84708 126300
rect 6004 126022 6046 126258
rect 6282 126022 84430 126258
rect 84666 126022 84708 126258
rect 6004 125980 84708 126022
rect 1104 125576 90896 125618
rect 1104 125340 1986 125576
rect 2222 125340 82536 125576
rect 82772 125340 85986 125576
rect 86222 125340 89986 125576
rect 90222 125340 90896 125576
rect 1104 125298 90896 125340
rect 1104 120576 90896 120618
rect 1104 120340 3986 120576
rect 4222 120340 82982 120576
rect 83218 120340 87986 120576
rect 88222 120340 90896 120576
rect 1104 120298 90896 120340
rect 5268 116738 90780 116780
rect 5268 116502 5310 116738
rect 5546 116502 90502 116738
rect 90738 116502 90780 116738
rect 5268 116460 90780 116502
rect 1104 115576 90896 115618
rect 1104 115340 1986 115576
rect 2222 115340 82536 115576
rect 82772 115340 85986 115576
rect 86222 115340 89986 115576
rect 90222 115340 90896 115576
rect 1104 115298 90896 115340
rect 1104 110576 90896 110618
rect 1104 110340 3986 110576
rect 4222 110340 82982 110576
rect 83218 110340 87986 110576
rect 88222 110340 90896 110576
rect 1104 110298 90896 110340
rect 1104 105576 90896 105618
rect 1104 105340 1986 105576
rect 2222 105340 82536 105576
rect 82772 105340 85986 105576
rect 86222 105340 89986 105576
rect 90222 105340 90896 105576
rect 1104 105298 90896 105340
rect 1104 100576 90896 100618
rect 1104 100340 3986 100576
rect 4222 100340 82982 100576
rect 83218 100340 87986 100576
rect 88222 100340 90896 100576
rect 1104 100298 90896 100340
rect 53108 97698 90780 97740
rect 53108 97462 90502 97698
rect 90738 97462 90780 97698
rect 53108 97420 90780 97462
rect 53108 97018 53428 97420
rect 53108 96782 53150 97018
rect 53386 96782 53428 97018
rect 53108 96740 53428 96782
rect 54028 97018 87284 97060
rect 54028 96782 54070 97018
rect 54306 96782 87006 97018
rect 87242 96782 87284 97018
rect 54028 96740 87284 96782
rect 50900 96338 88940 96380
rect 50900 96102 50942 96338
rect 51178 96102 88662 96338
rect 88898 96102 88940 96338
rect 50900 96060 88940 96102
rect 1104 95576 90896 95618
rect 1104 95340 1986 95576
rect 2222 95340 85986 95576
rect 86222 95340 89986 95576
rect 90222 95340 90896 95576
rect 1104 95298 90896 95340
rect 4348 94298 58948 94340
rect 4348 94062 4390 94298
rect 4626 94062 58948 94298
rect 4348 94020 58948 94062
rect 60836 94298 76980 94340
rect 60836 94062 60878 94298
rect 61114 94062 76702 94298
rect 76938 94062 76980 94298
rect 60836 94020 76980 94062
rect 77396 94298 89860 94340
rect 77396 94062 77438 94298
rect 77674 94062 89582 94298
rect 89818 94062 89860 94298
rect 77396 94020 89860 94062
rect 48140 93618 48460 93660
rect 48140 93382 48182 93618
rect 48418 93382 48460 93618
rect 48140 92300 48460 93382
rect 50900 93618 53428 93660
rect 50900 93382 53150 93618
rect 53386 93382 53428 93618
rect 50900 93340 53428 93382
rect 57123 93618 58258 93660
rect 57123 93382 57980 93618
rect 58216 93382 58258 93618
rect 57123 93340 58258 93382
rect 49244 93278 49564 93320
rect 49244 93042 49286 93278
rect 49522 93042 49564 93278
rect 49244 92980 49564 93042
rect 50900 92980 51220 93340
rect 49244 92660 51220 92980
rect 57123 92300 57443 93340
rect 58628 92980 58948 94020
rect 58444 92660 58948 92980
rect 59364 93618 59684 93660
rect 59364 93382 59406 93618
rect 59642 93382 59684 93618
rect 59364 92980 59684 93382
rect 60468 93618 88940 93660
rect 60468 93382 60510 93618
rect 60746 93382 88662 93618
rect 88898 93382 88940 93618
rect 60468 93340 88940 93382
rect 59364 92938 89308 92980
rect 59364 92702 89030 92938
rect 89266 92702 89308 92938
rect 59364 92660 89308 92702
rect 58444 92620 58764 92660
rect 48140 91980 57443 92300
rect 58260 92300 58764 92620
rect 58260 92258 84892 92300
rect 58260 92022 84614 92258
rect 84850 92022 84892 92258
rect 58260 91980 84892 92022
rect 4716 91578 87100 91620
rect 4716 91342 4758 91578
rect 4994 91342 86822 91578
rect 87058 91342 87100 91578
rect 4716 91300 87100 91342
rect 1104 90576 90896 90618
rect 1104 90340 3986 90576
rect 4222 90340 82982 90576
rect 83218 90340 87986 90576
rect 88222 90340 90896 90576
rect 1104 90298 90896 90340
rect 5452 89538 87100 89580
rect 5452 89302 5494 89538
rect 5730 89302 86822 89538
rect 87058 89302 87100 89538
rect 5452 89260 87100 89302
rect 5084 88858 87100 88900
rect 5084 88622 5126 88858
rect 5362 88622 86822 88858
rect 87058 88622 87100 88858
rect 5084 88580 87100 88622
rect 5268 86818 87468 86860
rect 5268 86582 5310 86818
rect 5546 86582 87190 86818
rect 87426 86582 87468 86818
rect 5268 86540 87468 86582
rect 1104 85576 90896 85618
rect 1104 85340 1986 85576
rect 2222 85340 82536 85576
rect 82772 85340 85986 85576
rect 86222 85340 89986 85576
rect 90222 85340 90896 85576
rect 1104 85298 90896 85340
rect 1104 80576 90896 80618
rect 1104 80340 3986 80576
rect 4222 80340 82982 80576
rect 83218 80340 87986 80576
rect 88222 80340 90896 80576
rect 1104 80298 90896 80340
rect 1104 75576 90896 75618
rect 1104 75340 1986 75576
rect 2222 75340 82536 75576
rect 82772 75340 85986 75576
rect 86222 75340 89986 75576
rect 90222 75340 90896 75576
rect 1104 75298 90896 75340
rect 1104 70576 90896 70618
rect 1104 70340 3986 70576
rect 4222 70340 82982 70576
rect 83218 70340 87986 70576
rect 88222 70340 90896 70576
rect 1104 70298 90896 70340
rect 1104 65576 90896 65618
rect 1104 65340 1986 65576
rect 2222 65340 82536 65576
rect 82772 65340 85986 65576
rect 86222 65340 89986 65576
rect 90222 65340 90896 65576
rect 1104 65298 90896 65340
rect 1104 60576 90896 60618
rect 1104 60340 3986 60576
rect 4222 60340 82982 60576
rect 83218 60340 87986 60576
rect 88222 60340 90896 60576
rect 1104 60298 90896 60340
rect 1104 55576 90896 55618
rect 1104 55340 1986 55576
rect 2222 55340 82536 55576
rect 82772 55340 85986 55576
rect 86222 55340 89986 55576
rect 90222 55340 90896 55576
rect 1104 55298 90896 55340
rect 1104 50576 90896 50618
rect 1104 50340 3986 50576
rect 4222 50340 82982 50576
rect 83218 50340 87986 50576
rect 88222 50340 90896 50576
rect 1104 50298 90896 50340
rect 1104 45576 90896 45618
rect 1104 45340 1986 45576
rect 2222 45340 82536 45576
rect 82772 45340 85986 45576
rect 86222 45340 89986 45576
rect 90222 45340 90896 45576
rect 1104 45298 90896 45340
rect 1104 40576 90896 40618
rect 1104 40340 3986 40576
rect 4222 40340 82982 40576
rect 83218 40340 87986 40576
rect 88222 40340 90896 40576
rect 1104 40298 90896 40340
rect 1104 35576 90896 35618
rect 1104 35340 1986 35576
rect 2222 35340 82536 35576
rect 82772 35340 85986 35576
rect 86222 35340 89986 35576
rect 90222 35340 90896 35576
rect 1104 35298 90896 35340
rect 1104 30576 90896 30618
rect 1104 30340 3986 30576
rect 4222 30340 82982 30576
rect 83218 30340 87986 30576
rect 88222 30340 90896 30576
rect 1104 30298 90896 30340
rect 1104 25576 90896 25618
rect 1104 25340 1986 25576
rect 2222 25340 82536 25576
rect 82772 25340 85986 25576
rect 86222 25340 89986 25576
rect 90222 25340 90896 25576
rect 1104 25298 90896 25340
rect 1104 20576 90896 20618
rect 1104 20340 3986 20576
rect 4222 20340 82982 20576
rect 83218 20340 87986 20576
rect 88222 20340 90896 20576
rect 1104 20298 90896 20340
rect 1104 15576 90896 15618
rect 1104 15340 1986 15576
rect 2222 15340 82536 15576
rect 82772 15340 85986 15576
rect 86222 15340 89986 15576
rect 90222 15340 90896 15576
rect 1104 15298 90896 15340
rect 1104 10576 90896 10618
rect 1104 10340 3986 10576
rect 4222 10340 82982 10576
rect 83218 10340 87986 10576
rect 88222 10340 90896 10576
rect 1104 10298 90896 10340
rect 1104 5576 90896 5618
rect 1104 5340 1986 5576
rect 2222 5340 82536 5576
rect 82772 5340 85986 5576
rect 86222 5340 89986 5576
rect 90222 5340 90896 5576
rect 1104 5298 90896 5340
rect 4716 3858 36868 3900
rect 4716 3622 4758 3858
rect 4994 3622 36868 3858
rect 4716 3580 36868 3622
rect 36548 3220 36868 3580
rect 8028 3178 36132 3220
rect 8028 2942 8070 3178
rect 8306 2942 36132 3178
rect 8028 2900 36132 2942
rect 36548 3178 37236 3220
rect 36548 2942 36958 3178
rect 37194 2942 37236 3178
rect 36548 2900 37236 2942
rect 37652 3178 41652 3220
rect 37652 2942 41374 3178
rect 41610 2942 41652 3178
rect 37652 2900 41652 2942
rect 35812 2540 36132 2900
rect 37652 2540 37972 2900
rect 35812 2220 37972 2540
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624015447
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_686
timestamp 1624015447
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624015447
transform 1 0 1380 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[5] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624015447
transform -1 0 2668 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_wmask0[0]
timestamp 1624015447
transform -1 0 2300 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_clk0
timestamp 1624015447
transform -1 0 2668 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624015447
transform 1 0 2668 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_13
timestamp 1624015447
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_17
timestamp 1624015447
transform 1 0 2668 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624015447
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_17
timestamp 1624015447
transform 1 0 2668 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1624015447
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_wmask0[2]
timestamp 1624015447
transform -1 0 2668 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1624015447
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_15
timestamp 1624015447
transform 1 0 2484 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1624015447
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1624015447
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_21
timestamp 1624015447
transform 1 0 3036 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21
timestamp 1624015447
transform 1 0 3036 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[9]
timestamp 1624015447
transform -1 0 3036 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[4]
timestamp 1624015447
transform -1 0 3404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[20]
timestamp 1624015447
transform -1 0 3036 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[18]
timestamp 1624015447
transform -1 0 3404 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_25
timestamp 1624015447
transform 1 0 3404 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25
timestamp 1624015447
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[1]
timestamp 1624015447
transform -1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[13]
timestamp 1624015447
transform -1 0 3772 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_29
timestamp 1624015447
transform 1 0 3772 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624015447
transform 1 0 3864 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[11]
timestamp 1624015447
transform -1 0 4140 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1548 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624015447
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_33
timestamp 1624015447
transform 1 0 4140 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624015447
transform 1 0 4232 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[15]
timestamp 1624015447
transform -1 0 4508 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[0]
timestamp 1624015447
transform -1 0 4508 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_21
timestamp 1624015447
transform 1 0 3036 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[7]
timestamp 1624015447
transform -1 0 3036 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[3]
timestamp 1624015447
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_25
timestamp 1624015447
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[17]
timestamp 1624015447
transform -1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_30
timestamp 1624015447
transform 1 0 3864 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1376
timestamp 1624015447
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_34
timestamp 1624015447
transform 1 0 4232 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[14]
timestamp 1624015447
transform -1 0 4508 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_wmask0[1]
timestamp 1624015447
transform -1 0 3404 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_25
timestamp 1624015447
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[6]
timestamp 1624015447
transform -1 0 3772 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_29
timestamp 1624015447
transform 1 0 3772 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[2]
timestamp 1624015447
transform 1 0 3956 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_33
timestamp 1624015447
transform 1 0 4140 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[19]
timestamp 1624015447
transform 1 0 4324 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_37
timestamp 1624015447
transform 1 0 4508 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37
timestamp 1624015447
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[12]
timestamp 1624015447
transform -1 0 4876 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr0[0]
timestamp 1624015447
transform -1 0 4876 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_687
timestamp 1624015447
transform -1 0 5152 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1624015447
transform -1 0 5152 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_37
timestamp 1624015447
transform 1 0 4508 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[10]
timestamp 1624015447
transform -1 0 4876 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1624015447
transform -1 0 5152 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_37
timestamp 1624015447
transform 1 0 4508 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[16]
timestamp 1624015447
transform -1 0 4876 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1624015447
transform -1 0 5152 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_690
timestamp 1624015447
transform 1 0 84180 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_688
timestamp 1624015447
transform 1 0 84180 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_906
timestamp 1624015447
transform 1 0 84456 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_906
timestamp 1624015447
transform 1 0 84456 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[26]
timestamp 1624015447
transform -1 0 84824 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[22]
timestamp 1624015447
transform 1 0 84640 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_692
timestamp 1624015447
transform 1 0 84180 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_906
timestamp 1624015447
transform 1 0 84456 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[23]
timestamp 1624015447
transform 1 0 84640 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_694
timestamp 1624015447
transform 1 0 84180 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_906
timestamp 1624015447
transform 1 0 84456 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[29]
timestamp 1624015447
transform 1 0 84640 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[24]
timestamp 1624015447
transform 1 0 85008 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[25]
timestamp 1624015447
transform 1 0 85376 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[28]
timestamp 1624015447
transform -1 0 85192 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_910
timestamp 1624015447
transform 1 0 84824 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_910
timestamp 1624015447
transform 1 0 84824 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_914
timestamp 1624015447
transform 1 0 85192 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_918
timestamp 1624015447
transform 1 0 85560 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[30]
timestamp 1624015447
transform 1 0 85744 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_926 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624015447
transform 1 0 86296 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_914
timestamp 1624015447
transform 1 0 85192 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_922
timestamp 1624015447
transform 1 0 85928 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_918
timestamp 1624015447
transform 1 0 85560 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_914
timestamp 1624015447
transform 1 0 85192 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_910
timestamp 1624015447
transform 1 0 84824 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[31]
timestamp 1624015447
transform 1 0 85376 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[27]
timestamp 1624015447
transform 1 0 85008 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_922
timestamp 1624015447
transform 1 0 85928 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_910
timestamp 1624015447
transform 1 0 84824 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_946
timestamp 1624015447
transform 1 0 88136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_934
timestamp 1624015447
transform 1 0 87032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_945
timestamp 1624015447
transform 1 0 88044 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_933
timestamp 1624015447
transform 1 0 86940 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1549
timestamp 1624015447
transform 1 0 86848 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_945
timestamp 1624015447
transform 1 0 88044 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_933
timestamp 1624015447
transform 1 0 86940 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_930
timestamp 1624015447
transform 1 0 86664 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1552
timestamp 1624015447
transform 1 0 86848 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_946
timestamp 1624015447
transform 1 0 88136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_934
timestamp 1624015447
transform 1 0 87032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_961
timestamp 1624015447
transform 1 0 89516 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_958
timestamp 1624015447
transform 1 0 89240 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_962
timestamp 1624015447
transform 1 0 89608 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_957
timestamp 1624015447
transform 1 0 89148 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1551
timestamp 1624015447
transform 1 0 89424 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1550
timestamp 1624015447
transform 1 0 89516 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_957
timestamp 1624015447
transform 1 0 89148 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_961
timestamp 1624015447
transform 1 0 89516 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_958
timestamp 1624015447
transform 1 0 89240 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1553
timestamp 1624015447
transform 1 0 89424 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_689
timestamp 1624015447
transform -1 0 90896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_691
timestamp 1624015447
transform -1 0 90896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_693
timestamp 1624015447
transform -1 0 90896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_695
timestamp 1624015447
transform -1 0 90896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_970
timestamp 1624015447
transform 1 0 90344 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_969
timestamp 1624015447
transform 1 0 90252 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1624015447
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1624015447
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1624015447
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1624015447
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1624015447
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1624015447
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1624015447
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1624015447
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1624015447
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1377
timestamp 1624015447
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1378
timestamp 1624015447
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[8]
timestamp 1624015447
transform 1 0 4324 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1624015447
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_30
timestamp 1624015447
transform 1 0 3864 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_34
timestamp 1624015447
transform 1 0 4232 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1624015447
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1624015447
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_30
timestamp 1624015447
transform 1 0 3864 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1624015447
transform -1 0 5152 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1624015447
transform -1 0 5152 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1624015447
transform -1 0 5152 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_din0[21]
timestamp 1624015447
transform 1 0 4692 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_wmask0[3]
timestamp 1624015447
transform -1 0 4876 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_37
timestamp 1624015447
transform 1 0 4508 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_38
timestamp 1624015447
transform 1 0 4600 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_696
timestamp 1624015447
transform 1 0 84180 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_698
timestamp 1624015447
transform 1 0 84180 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_700
timestamp 1624015447
transform 1 0 84180 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_906
timestamp 1624015447
transform 1 0 84456 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_906
timestamp 1624015447
transform 1 0 84456 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_906
timestamp 1624015447
transform 1 0 84456 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_918
timestamp 1624015447
transform 1 0 85560 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_918
timestamp 1624015447
transform 1 0 85560 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_918
timestamp 1624015447
transform 1 0 85560 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_945
timestamp 1624015447
transform 1 0 88044 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_933
timestamp 1624015447
transform 1 0 86940 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_930
timestamp 1624015447
transform 1 0 86664 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1554
timestamp 1624015447
transform 1 0 86848 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_942
timestamp 1624015447
transform 1 0 87768 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_930
timestamp 1624015447
transform 1 0 86664 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_945
timestamp 1624015447
transform 1 0 88044 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_933
timestamp 1624015447
transform 1 0 86940 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_930
timestamp 1624015447
transform 1 0 86664 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1556
timestamp 1624015447
transform 1 0 86848 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1555
timestamp 1624015447
transform 1 0 89424 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_957
timestamp 1624015447
transform 1 0 89148 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_954
timestamp 1624015447
transform 1 0 88872 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_961
timestamp 1624015447
transform 1 0 89516 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_957
timestamp 1624015447
transform 1 0 89148 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_697
timestamp 1624015447
transform -1 0 90896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_699
timestamp 1624015447
transform -1 0 90896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_701
timestamp 1624015447
transform -1 0 90896 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_969
timestamp 1624015447
transform 1 0 90252 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_969
timestamp 1624015447
transform 1 0 90252 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1624015447
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1624015447
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1624015447
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1624015447
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1624015447
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1624015447
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1624015447
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1624015447
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1624015447
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1379
timestamp 1624015447
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1624015447
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_27
timestamp 1624015447
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_30
timestamp 1624015447
transform 1 0 3864 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1624015447
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1624015447
transform -1 0 5152 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1624015447
transform -1 0 5152 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1624015447
transform -1 0 5152 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_39
timestamp 1624015447
transform 1 0 4692 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_38
timestamp 1624015447
transform 1 0 4600 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_39
timestamp 1624015447
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_702
timestamp 1624015447
transform 1 0 84180 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_704
timestamp 1624015447
transform 1 0 84180 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_706
timestamp 1624015447
transform 1 0 84180 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_906
timestamp 1624015447
transform 1 0 84456 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_906
timestamp 1624015447
transform 1 0 84456 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_906
timestamp 1624015447
transform 1 0 84456 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_918
timestamp 1624015447
transform 1 0 85560 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_918
timestamp 1624015447
transform 1 0 85560 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_918
timestamp 1624015447
transform 1 0 85560 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1558
timestamp 1624015447
transform 1 0 86848 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_930
timestamp 1624015447
transform 1 0 86664 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_942
timestamp 1624015447
transform 1 0 87768 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_930
timestamp 1624015447
transform 1 0 86664 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_933
timestamp 1624015447
transform 1 0 86940 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_945
timestamp 1624015447
transform 1 0 88044 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_930
timestamp 1624015447
transform 1 0 86664 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_942
timestamp 1624015447
transform 1 0 87768 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1557
timestamp 1624015447
transform 1 0 89424 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1559
timestamp 1624015447
transform 1 0 89424 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_954
timestamp 1624015447
transform 1 0 88872 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_961
timestamp 1624015447
transform 1 0 89516 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_957
timestamp 1624015447
transform 1 0 89148 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_954
timestamp 1624015447
transform 1 0 88872 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_961
timestamp 1624015447
transform 1 0 89516 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_703
timestamp 1624015447
transform -1 0 90896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_705
timestamp 1624015447
transform -1 0 90896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_707
timestamp 1624015447
transform -1 0 90896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_969
timestamp 1624015447
transform 1 0 90252 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1624015447
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1624015447
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1624015447
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1624015447
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1624015447
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1624015447
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1624015447
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1624015447
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1624015447
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1380
timestamp 1624015447
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1381
timestamp 1624015447
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1624015447
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_30
timestamp 1624015447
transform 1 0 3864 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1624015447
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1624015447
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_30
timestamp 1624015447
transform 1 0 3864 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1624015447
transform -1 0 5152 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1624015447
transform -1 0 5152 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1624015447
transform -1 0 5152 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_38
timestamp 1624015447
transform 1 0 4600 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_39
timestamp 1624015447
transform 1 0 4692 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_38
timestamp 1624015447
transform 1 0 4600 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_708
timestamp 1624015447
transform 1 0 84180 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_710
timestamp 1624015447
transform 1 0 84180 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_712
timestamp 1624015447
transform 1 0 84180 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_906
timestamp 1624015447
transform 1 0 84456 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_906
timestamp 1624015447
transform 1 0 84456 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_906
timestamp 1624015447
transform 1 0 84456 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_918
timestamp 1624015447
transform 1 0 85560 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_918
timestamp 1624015447
transform 1 0 85560 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_918
timestamp 1624015447
transform 1 0 85560 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_945
timestamp 1624015447
transform 1 0 88044 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_933
timestamp 1624015447
transform 1 0 86940 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_930
timestamp 1624015447
transform 1 0 86664 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1560
timestamp 1624015447
transform 1 0 86848 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_942
timestamp 1624015447
transform 1 0 87768 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_930
timestamp 1624015447
transform 1 0 86664 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_945
timestamp 1624015447
transform 1 0 88044 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_933
timestamp 1624015447
transform 1 0 86940 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_930
timestamp 1624015447
transform 1 0 86664 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1562
timestamp 1624015447
transform 1 0 86848 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1561
timestamp 1624015447
transform 1 0 89424 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_957
timestamp 1624015447
transform 1 0 89148 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_954
timestamp 1624015447
transform 1 0 88872 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_961
timestamp 1624015447
transform 1 0 89516 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_957
timestamp 1624015447
transform 1 0 89148 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_709
timestamp 1624015447
transform -1 0 90896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_711
timestamp 1624015447
transform -1 0 90896 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_713
timestamp 1624015447
transform -1 0 90896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_969
timestamp 1624015447
transform 1 0 90252 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_969
timestamp 1624015447
transform 1 0 90252 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1624015447
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1624015447
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1624015447
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1624015447
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1624015447
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1624015447
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1624015447
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1624015447
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1624015447
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _12_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624015447
transform 1 0 4232 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1382
timestamp 1624015447
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1624015447
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1624015447
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_30
timestamp 1624015447
transform 1 0 3864 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1624015447
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1624015447
transform -1 0 5152 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1624015447
transform -1 0 5152 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1624015447
transform -1 0 5152 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_39
timestamp 1624015447
transform 1 0 4692 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_37
timestamp 1624015447
transform 1 0 4508 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_39
timestamp 1624015447
transform 1 0 4692 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_714
timestamp 1624015447
transform 1 0 84180 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_716
timestamp 1624015447
transform 1 0 84180 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_718
timestamp 1624015447
transform 1 0 84180 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_906
timestamp 1624015447
transform 1 0 84456 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_906
timestamp 1624015447
transform 1 0 84456 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_906
timestamp 1624015447
transform 1 0 84456 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_918
timestamp 1624015447
transform 1 0 85560 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_918
timestamp 1624015447
transform 1 0 85560 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_918
timestamp 1624015447
transform 1 0 85560 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1564
timestamp 1624015447
transform 1 0 86848 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_930
timestamp 1624015447
transform 1 0 86664 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_942
timestamp 1624015447
transform 1 0 87768 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_930
timestamp 1624015447
transform 1 0 86664 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_933
timestamp 1624015447
transform 1 0 86940 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_945
timestamp 1624015447
transform 1 0 88044 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_930
timestamp 1624015447
transform 1 0 86664 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_942
timestamp 1624015447
transform 1 0 87768 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1563
timestamp 1624015447
transform 1 0 89424 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1565
timestamp 1624015447
transform 1 0 89424 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_954
timestamp 1624015447
transform 1 0 88872 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_961
timestamp 1624015447
transform 1 0 89516 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_957
timestamp 1624015447
transform 1 0 89148 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_954
timestamp 1624015447
transform 1 0 88872 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_961
timestamp 1624015447
transform 1 0 89516 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_715
timestamp 1624015447
transform -1 0 90896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_717
timestamp 1624015447
transform -1 0 90896 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_719
timestamp 1624015447
transform -1 0 90896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_969
timestamp 1624015447
transform 1 0 90252 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1624015447
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1624015447
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1624015447
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1624015447
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1624015447
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1624015447
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1624015447
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1624015447
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1624015447
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1383
timestamp 1624015447
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1384
timestamp 1624015447
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1624015447
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_30
timestamp 1624015447
transform 1 0 3864 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1624015447
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1624015447
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_30
timestamp 1624015447
transform 1 0 3864 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1624015447
transform -1 0 5152 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1624015447
transform -1 0 5152 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1624015447
transform -1 0 5152 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_38
timestamp 1624015447
transform 1 0 4600 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_39
timestamp 1624015447
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_38
timestamp 1624015447
transform 1 0 4600 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_720
timestamp 1624015447
transform 1 0 84180 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_722
timestamp 1624015447
transform 1 0 84180 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_724
timestamp 1624015447
transform 1 0 84180 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_906
timestamp 1624015447
transform 1 0 84456 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_906
timestamp 1624015447
transform 1 0 84456 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_906
timestamp 1624015447
transform 1 0 84456 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_918
timestamp 1624015447
transform 1 0 85560 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_918
timestamp 1624015447
transform 1 0 85560 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_918
timestamp 1624015447
transform 1 0 85560 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_945
timestamp 1624015447
transform 1 0 88044 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_933
timestamp 1624015447
transform 1 0 86940 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_930
timestamp 1624015447
transform 1 0 86664 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1566
timestamp 1624015447
transform 1 0 86848 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_942
timestamp 1624015447
transform 1 0 87768 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_930
timestamp 1624015447
transform 1 0 86664 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_945
timestamp 1624015447
transform 1 0 88044 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_933
timestamp 1624015447
transform 1 0 86940 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_930
timestamp 1624015447
transform 1 0 86664 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1568
timestamp 1624015447
transform 1 0 86848 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1567
timestamp 1624015447
transform 1 0 89424 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_957
timestamp 1624015447
transform 1 0 89148 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_954
timestamp 1624015447
transform 1 0 88872 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_961
timestamp 1624015447
transform 1 0 89516 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_957
timestamp 1624015447
transform 1 0 89148 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_721
timestamp 1624015447
transform -1 0 90896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_723
timestamp 1624015447
transform -1 0 90896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_725
timestamp 1624015447
transform -1 0 90896 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_969
timestamp 1624015447
transform 1 0 90252 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_969
timestamp 1624015447
transform 1 0 90252 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1624015447
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1624015447
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1624015447
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1624015447
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1624015447
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1624015447
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1624015447
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1624015447
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1624015447
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1385
timestamp 1624015447
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1624015447
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1624015447
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_30
timestamp 1624015447
transform 1 0 3864 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1624015447
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1624015447
transform -1 0 5152 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1624015447
transform -1 0 5152 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1624015447
transform -1 0 5152 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_39
timestamp 1624015447
transform 1 0 4692 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_38
timestamp 1624015447
transform 1 0 4600 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_39
timestamp 1624015447
transform 1 0 4692 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_8  BUF1_8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624015447
transform 1 0 84456 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_726
timestamp 1624015447
transform 1 0 84180 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_728
timestamp 1624015447
transform 1 0 84180 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_730
timestamp 1624015447
transform 1 0 84180 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_906
timestamp 1624015447
transform 1 0 84456 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_906
timestamp 1624015447
transform 1 0 84456 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_918
timestamp 1624015447
transform 1 0 85560 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_918
timestamp 1624015447
transform 1 0 85560 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_918
timestamp 1624015447
transform 1 0 85560 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1570
timestamp 1624015447
transform 1 0 86848 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_930
timestamp 1624015447
transform 1 0 86664 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_942
timestamp 1624015447
transform 1 0 87768 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_930
timestamp 1624015447
transform 1 0 86664 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_933
timestamp 1624015447
transform 1 0 86940 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_945
timestamp 1624015447
transform 1 0 88044 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_930
timestamp 1624015447
transform 1 0 86664 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_942
timestamp 1624015447
transform 1 0 87768 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1569
timestamp 1624015447
transform 1 0 89424 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1571
timestamp 1624015447
transform 1 0 89424 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_954
timestamp 1624015447
transform 1 0 88872 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_961
timestamp 1624015447
transform 1 0 89516 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_957
timestamp 1624015447
transform 1 0 89148 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_954
timestamp 1624015447
transform 1 0 88872 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_961
timestamp 1624015447
transform 1 0 89516 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_727
timestamp 1624015447
transform -1 0 90896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_729
timestamp 1624015447
transform -1 0 90896 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_731
timestamp 1624015447
transform -1 0 90896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_969
timestamp 1624015447
transform 1 0 90252 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1624015447
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1624015447
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1624015447
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1624015447
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1624015447
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1624015447
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1624015447
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1624015447
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1624015447
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1386
timestamp 1624015447
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1387
timestamp 1624015447
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1624015447
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_30
timestamp 1624015447
transform 1 0 3864 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1624015447
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1624015447
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_30
timestamp 1624015447
transform 1 0 3864 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1624015447
transform -1 0 5152 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1624015447
transform -1 0 5152 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1624015447
transform -1 0 5152 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_38
timestamp 1624015447
transform 1 0 4600 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_39
timestamp 1624015447
transform 1 0 4692 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_38
timestamp 1624015447
transform 1 0 4600 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_732
timestamp 1624015447
transform 1 0 84180 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_734
timestamp 1624015447
transform 1 0 84180 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_736
timestamp 1624015447
transform 1 0 84180 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF1_8_A
timestamp 1624015447
transform 1 0 84640 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_906
timestamp 1624015447
transform 1 0 84456 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_906
timestamp 1624015447
transform 1 0 84456 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_906
timestamp 1624015447
transform 1 0 84456 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_910
timestamp 1624015447
transform 1 0 84824 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_922
timestamp 1624015447
transform 1 0 85928 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_918
timestamp 1624015447
transform 1 0 85560 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_918
timestamp 1624015447
transform 1 0 85560 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_945
timestamp 1624015447
transform 1 0 88044 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_933
timestamp 1624015447
transform 1 0 86940 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_930
timestamp 1624015447
transform 1 0 86664 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1572
timestamp 1624015447
transform 1 0 86848 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_942
timestamp 1624015447
transform 1 0 87768 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_930
timestamp 1624015447
transform 1 0 86664 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_945
timestamp 1624015447
transform 1 0 88044 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_933
timestamp 1624015447
transform 1 0 86940 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_930
timestamp 1624015447
transform 1 0 86664 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1574
timestamp 1624015447
transform 1 0 86848 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1573
timestamp 1624015447
transform 1 0 89424 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_957
timestamp 1624015447
transform 1 0 89148 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_954
timestamp 1624015447
transform 1 0 88872 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_961
timestamp 1624015447
transform 1 0 89516 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_957
timestamp 1624015447
transform 1 0 89148 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_733
timestamp 1624015447
transform -1 0 90896 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_735
timestamp 1624015447
transform -1 0 90896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_737
timestamp 1624015447
transform -1 0 90896 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_969
timestamp 1624015447
transform 1 0 90252 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_969
timestamp 1624015447
transform 1 0 90252 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1624015447
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1624015447
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1624015447
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1624015447
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1624015447
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1624015447
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1624015447
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1624015447
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1624015447
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1388
timestamp 1624015447
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1624015447
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1624015447
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_30
timestamp 1624015447
transform 1 0 3864 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1624015447
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1624015447
transform -1 0 5152 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1624015447
transform -1 0 5152 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1624015447
transform -1 0 5152 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_39
timestamp 1624015447
transform 1 0 4692 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_38
timestamp 1624015447
transform 1 0 4600 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_39
timestamp 1624015447
transform 1 0 4692 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_738
timestamp 1624015447
transform 1 0 84180 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_740
timestamp 1624015447
transform 1 0 84180 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_742
timestamp 1624015447
transform 1 0 84180 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_906
timestamp 1624015447
transform 1 0 84456 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_906
timestamp 1624015447
transform 1 0 84456 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_906
timestamp 1624015447
transform 1 0 84456 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_918
timestamp 1624015447
transform 1 0 85560 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_918
timestamp 1624015447
transform 1 0 85560 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_918
timestamp 1624015447
transform 1 0 85560 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1576
timestamp 1624015447
transform 1 0 86848 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_930
timestamp 1624015447
transform 1 0 86664 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_942
timestamp 1624015447
transform 1 0 87768 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_930
timestamp 1624015447
transform 1 0 86664 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_933
timestamp 1624015447
transform 1 0 86940 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_945
timestamp 1624015447
transform 1 0 88044 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_930
timestamp 1624015447
transform 1 0 86664 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_942
timestamp 1624015447
transform 1 0 87768 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1575
timestamp 1624015447
transform 1 0 89424 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1577
timestamp 1624015447
transform 1 0 89424 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_954
timestamp 1624015447
transform 1 0 88872 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_961
timestamp 1624015447
transform 1 0 89516 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_957
timestamp 1624015447
transform 1 0 89148 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_954
timestamp 1624015447
transform 1 0 88872 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_961
timestamp 1624015447
transform 1 0 89516 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_739
timestamp 1624015447
transform -1 0 90896 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_741
timestamp 1624015447
transform -1 0 90896 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_743
timestamp 1624015447
transform -1 0 90896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_969
timestamp 1624015447
transform 1 0 90252 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1624015447
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1624015447
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1624015447
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1624015447
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1624015447
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1624015447
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1624015447
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1624015447
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1624015447
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1389
timestamp 1624015447
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1390
timestamp 1624015447
transform 1 0 3772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_27
timestamp 1624015447
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_30
timestamp 1624015447
transform 1 0 3864 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1624015447
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_27
timestamp 1624015447
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_30
timestamp 1624015447
transform 1 0 3864 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1624015447
transform -1 0 5152 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1624015447
transform -1 0 5152 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1624015447
transform -1 0 5152 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_38
timestamp 1624015447
transform 1 0 4600 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_39
timestamp 1624015447
transform 1 0 4692 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_38
timestamp 1624015447
transform 1 0 4600 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _15_
timestamp 1624015447
transform -1 0 84732 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_744
timestamp 1624015447
transform 1 0 84180 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_746
timestamp 1624015447
transform 1 0 84180 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_748
timestamp 1624015447
transform 1 0 84180 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_909
timestamp 1624015447
transform 1 0 84732 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_906
timestamp 1624015447
transform 1 0 84456 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_906
timestamp 1624015447
transform 1 0 84456 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_921
timestamp 1624015447
transform 1 0 85836 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_918
timestamp 1624015447
transform 1 0 85560 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_918
timestamp 1624015447
transform 1 0 85560 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_945
timestamp 1624015447
transform 1 0 88044 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_933
timestamp 1624015447
transform 1 0 86940 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_929
timestamp 1624015447
transform 1 0 86572 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1578
timestamp 1624015447
transform 1 0 86848 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_945
timestamp 1624015447
transform 1 0 88044 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_933
timestamp 1624015447
transform 1 0 86940 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_930
timestamp 1624015447
transform 1 0 86664 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_942
timestamp 1624015447
transform 1 0 87768 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_930
timestamp 1624015447
transform 1 0 86664 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1580
timestamp 1624015447
transform 1 0 86848 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1579
timestamp 1624015447
transform 1 0 89424 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_957
timestamp 1624015447
transform 1 0 89148 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_954
timestamp 1624015447
transform 1 0 88872 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_961
timestamp 1624015447
transform 1 0 89516 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_957
timestamp 1624015447
transform 1 0 89148 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_745
timestamp 1624015447
transform -1 0 90896 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_747
timestamp 1624015447
transform -1 0 90896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_749
timestamp 1624015447
transform -1 0 90896 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_969
timestamp 1624015447
transform 1 0 90252 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_969
timestamp 1624015447
transform 1 0 90252 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1624015447
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1624015447
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1624015447
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1624015447
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1624015447
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1624015447
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1624015447
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1624015447
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1624015447
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1391
timestamp 1624015447
transform 1 0 3772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1624015447
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_27
timestamp 1624015447
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_30
timestamp 1624015447
transform 1 0 3864 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1624015447
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1624015447
transform -1 0 5152 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1624015447
transform -1 0 5152 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1624015447
transform -1 0 5152 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_39
timestamp 1624015447
transform 1 0 4692 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_38
timestamp 1624015447
transform 1 0 4600 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_39
timestamp 1624015447
transform 1 0 4692 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_750
timestamp 1624015447
transform 1 0 84180 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_752
timestamp 1624015447
transform 1 0 84180 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_754
timestamp 1624015447
transform 1 0 84180 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_906
timestamp 1624015447
transform 1 0 84456 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_906
timestamp 1624015447
transform 1 0 84456 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_906
timestamp 1624015447
transform 1 0 84456 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_918
timestamp 1624015447
transform 1 0 85560 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_918
timestamp 1624015447
transform 1 0 85560 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_918
timestamp 1624015447
transform 1 0 85560 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1582
timestamp 1624015447
transform 1 0 86848 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_930
timestamp 1624015447
transform 1 0 86664 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_942
timestamp 1624015447
transform 1 0 87768 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_930
timestamp 1624015447
transform 1 0 86664 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_933
timestamp 1624015447
transform 1 0 86940 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_945
timestamp 1624015447
transform 1 0 88044 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_930
timestamp 1624015447
transform 1 0 86664 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_942
timestamp 1624015447
transform 1 0 87768 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1581
timestamp 1624015447
transform 1 0 89424 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1583
timestamp 1624015447
transform 1 0 89424 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_954
timestamp 1624015447
transform 1 0 88872 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_961
timestamp 1624015447
transform 1 0 89516 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_957
timestamp 1624015447
transform 1 0 89148 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_954
timestamp 1624015447
transform 1 0 88872 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_961
timestamp 1624015447
transform 1 0 89516 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_751
timestamp 1624015447
transform -1 0 90896 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_753
timestamp 1624015447
transform -1 0 90896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_755
timestamp 1624015447
transform -1 0 90896 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_969
timestamp 1624015447
transform 1 0 90252 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1624015447
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1624015447
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1624015447
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1624015447
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1624015447
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1624015447
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1624015447
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1624015447
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1624015447
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1392
timestamp 1624015447
transform 1 0 3772 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1393
timestamp 1624015447
transform 1 0 3772 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_27
timestamp 1624015447
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_30
timestamp 1624015447
transform 1 0 3864 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1624015447
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_27
timestamp 1624015447
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_30
timestamp 1624015447
transform 1 0 3864 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1624015447
transform -1 0 5152 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1624015447
transform -1 0 5152 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1624015447
transform -1 0 5152 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_csb0
timestamp 1624015447
transform -1 0 4876 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_38
timestamp 1624015447
transform 1 0 4600 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_39
timestamp 1624015447
transform 1 0 4692 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_38
timestamp 1624015447
transform 1 0 4600 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_756
timestamp 1624015447
transform 1 0 84180 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_758
timestamp 1624015447
transform 1 0 84180 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_760
timestamp 1624015447
transform 1 0 84180 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_906
timestamp 1624015447
transform 1 0 84456 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_906
timestamp 1624015447
transform 1 0 84456 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_906
timestamp 1624015447
transform 1 0 84456 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_918
timestamp 1624015447
transform 1 0 85560 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_918
timestamp 1624015447
transform 1 0 85560 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_918
timestamp 1624015447
transform 1 0 85560 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_942
timestamp 1624015447
transform 1 0 87768 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_930
timestamp 1624015447
transform 1 0 86664 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_945
timestamp 1624015447
transform 1 0 88044 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_933
timestamp 1624015447
transform 1 0 86940 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_930
timestamp 1624015447
transform 1 0 86664 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1584
timestamp 1624015447
transform 1 0 86848 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_945
timestamp 1624015447
transform 1 0 88044 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_933
timestamp 1624015447
transform 1 0 86940 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_930
timestamp 1624015447
transform 1 0 86664 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1586
timestamp 1624015447
transform 1 0 86848 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1585
timestamp 1624015447
transform 1 0 89424 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_957
timestamp 1624015447
transform 1 0 89148 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_954
timestamp 1624015447
transform 1 0 88872 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_961
timestamp 1624015447
transform 1 0 89516 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_957
timestamp 1624015447
transform 1 0 89148 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_757
timestamp 1624015447
transform -1 0 90896 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_759
timestamp 1624015447
transform -1 0 90896 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_761
timestamp 1624015447
transform -1 0 90896 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_969
timestamp 1624015447
transform 1 0 90252 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_969
timestamp 1624015447
transform 1 0 90252 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1624015447
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1624015447
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1624015447
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1624015447
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1624015447
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1624015447
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1624015447
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1624015447
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1624015447
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1624015447
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1624015447
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1624015447
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1394
timestamp 1624015447
transform 1 0 3772 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1395
timestamp 1624015447
transform 1 0 3772 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1624015447
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_27
timestamp 1624015447
transform 1 0 3588 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_30
timestamp 1624015447
transform 1 0 3864 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1624015447
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_27
timestamp 1624015447
transform 1 0 3588 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_30
timestamp 1624015447
transform 1 0 3864 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1624015447
transform -1 0 5152 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1624015447
transform -1 0 5152 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1624015447
transform -1 0 5152 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1624015447
transform -1 0 5152 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_web0
timestamp 1624015447
transform -1 0 4876 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_38
timestamp 1624015447
transform 1 0 4600 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_39
timestamp 1624015447
transform 1 0 4692 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_38
timestamp 1624015447
transform 1 0 4600 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_906
timestamp 1624015447
transform 1 0 84456 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_906
timestamp 1624015447
transform 1 0 84456 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr1[7]
timestamp 1624015447
transform -1 0 84824 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_764
timestamp 1624015447
transform 1 0 84180 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_762
timestamp 1624015447
transform 1 0 84180 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_906
timestamp 1624015447
transform 1 0 84456 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_766
timestamp 1624015447
transform 1 0 84180 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_906
timestamp 1624015447
transform 1 0 84456 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr1[6]
timestamp 1624015447
transform -1 0 84824 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_768
timestamp 1624015447
transform 1 0 84180 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_918
timestamp 1624015447
transform 1 0 85560 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_910
timestamp 1624015447
transform 1 0 84824 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_922
timestamp 1624015447
transform 1 0 85928 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_918
timestamp 1624015447
transform 1 0 85560 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_910
timestamp 1624015447
transform 1 0 84824 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_922
timestamp 1624015447
transform 1 0 85928 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_945
timestamp 1624015447
transform 1 0 88044 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_933
timestamp 1624015447
transform 1 0 86940 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_930
timestamp 1624015447
transform 1 0 86664 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_942
timestamp 1624015447
transform 1 0 87768 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_930
timestamp 1624015447
transform 1 0 86664 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1588
timestamp 1624015447
transform 1 0 86848 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_942
timestamp 1624015447
transform 1 0 87768 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_930
timestamp 1624015447
transform 1 0 86664 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_945
timestamp 1624015447
transform 1 0 88044 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_933
timestamp 1624015447
transform 1 0 86940 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_930
timestamp 1624015447
transform 1 0 86664 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1590
timestamp 1624015447
transform 1 0 86848 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1587
timestamp 1624015447
transform 1 0 89424 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1589
timestamp 1624015447
transform 1 0 89424 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_954
timestamp 1624015447
transform 1 0 88872 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_961
timestamp 1624015447
transform 1 0 89516 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_957
timestamp 1624015447
transform 1 0 89148 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_954
timestamp 1624015447
transform 1 0 88872 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_961
timestamp 1624015447
transform 1 0 89516 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_957
timestamp 1624015447
transform 1 0 89148 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_763
timestamp 1624015447
transform -1 0 90896 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_765
timestamp 1624015447
transform -1 0 90896 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_767
timestamp 1624015447
transform -1 0 90896 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_769
timestamp 1624015447
transform -1 0 90896 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_969
timestamp 1624015447
transform 1 0 90252 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_969
timestamp 1624015447
transform 1 0 90252 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1624015447
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1624015447
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1624015447
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1624015447
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1624015447
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1624015447
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1624015447
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1624015447
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1624015447
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1396
timestamp 1624015447
transform 1 0 3772 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1624015447
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_27
timestamp 1624015447
transform 1 0 3588 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_30
timestamp 1624015447
transform 1 0 3864 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1624015447
transform 1 0 3588 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1624015447
transform -1 0 5152 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1624015447
transform -1 0 5152 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1624015447
transform -1 0 5152 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_39
timestamp 1624015447
transform 1 0 4692 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_38
timestamp 1624015447
transform 1 0 4600 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_39
timestamp 1624015447
transform 1 0 4692 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_770
timestamp 1624015447
transform 1 0 84180 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_772
timestamp 1624015447
transform 1 0 84180 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_774
timestamp 1624015447
transform 1 0 84180 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_906
timestamp 1624015447
transform 1 0 84456 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_906
timestamp 1624015447
transform 1 0 84456 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_906
timestamp 1624015447
transform 1 0 84456 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_918
timestamp 1624015447
transform 1 0 85560 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_918
timestamp 1624015447
transform 1 0 85560 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_918
timestamp 1624015447
transform 1 0 85560 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1592
timestamp 1624015447
transform 1 0 86848 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_930
timestamp 1624015447
transform 1 0 86664 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_942
timestamp 1624015447
transform 1 0 87768 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_930
timestamp 1624015447
transform 1 0 86664 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_933
timestamp 1624015447
transform 1 0 86940 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_945
timestamp 1624015447
transform 1 0 88044 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_930
timestamp 1624015447
transform 1 0 86664 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_942
timestamp 1624015447
transform 1 0 87768 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1591
timestamp 1624015447
transform 1 0 89424 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1593
timestamp 1624015447
transform 1 0 89424 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_954
timestamp 1624015447
transform 1 0 88872 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_961
timestamp 1624015447
transform 1 0 89516 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_957
timestamp 1624015447
transform 1 0 89148 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_954
timestamp 1624015447
transform 1 0 88872 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_961
timestamp 1624015447
transform 1 0 89516 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_771
timestamp 1624015447
transform -1 0 90896 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_773
timestamp 1624015447
transform -1 0 90896 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_775
timestamp 1624015447
transform -1 0 90896 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_969
timestamp 1624015447
transform 1 0 90252 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1624015447
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1624015447
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1624015447
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1624015447
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1624015447
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1624015447
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1624015447
transform 1 0 2484 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1624015447
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1624015447
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1397
timestamp 1624015447
transform 1 0 3772 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1398
timestamp 1624015447
transform 1 0 3772 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_27
timestamp 1624015447
transform 1 0 3588 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_30
timestamp 1624015447
transform 1 0 3864 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1624015447
transform 1 0 3588 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_27
timestamp 1624015447
transform 1 0 3588 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_30
timestamp 1624015447
transform 1 0 3864 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1624015447
transform -1 0 5152 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1624015447
transform -1 0 5152 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1624015447
transform -1 0 5152 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_38
timestamp 1624015447
transform 1 0 4600 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_39
timestamp 1624015447
transform 1 0 4692 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_38
timestamp 1624015447
transform 1 0 4600 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_776
timestamp 1624015447
transform 1 0 84180 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_778
timestamp 1624015447
transform 1 0 84180 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_780
timestamp 1624015447
transform 1 0 84180 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr1[4]
timestamp 1624015447
transform 1 0 84640 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr1[5]
timestamp 1624015447
transform 1 0 84640 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_906
timestamp 1624015447
transform 1 0 84456 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_906
timestamp 1624015447
transform 1 0 84456 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_906
timestamp 1624015447
transform 1 0 84456 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_910
timestamp 1624015447
transform 1 0 84824 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_922
timestamp 1624015447
transform 1 0 85928 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_918
timestamp 1624015447
transform 1 0 85560 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_910
timestamp 1624015447
transform 1 0 84824 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_922
timestamp 1624015447
transform 1 0 85928 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_945
timestamp 1624015447
transform 1 0 88044 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_933
timestamp 1624015447
transform 1 0 86940 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_930
timestamp 1624015447
transform 1 0 86664 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1594
timestamp 1624015447
transform 1 0 86848 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_942
timestamp 1624015447
transform 1 0 87768 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_930
timestamp 1624015447
transform 1 0 86664 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_945
timestamp 1624015447
transform 1 0 88044 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_933
timestamp 1624015447
transform 1 0 86940 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_930
timestamp 1624015447
transform 1 0 86664 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1596
timestamp 1624015447
transform 1 0 86848 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1595
timestamp 1624015447
transform 1 0 89424 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_957
timestamp 1624015447
transform 1 0 89148 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_954
timestamp 1624015447
transform 1 0 88872 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_961
timestamp 1624015447
transform 1 0 89516 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_957
timestamp 1624015447
transform 1 0 89148 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_777
timestamp 1624015447
transform -1 0 90896 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_779
timestamp 1624015447
transform -1 0 90896 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_781
timestamp 1624015447
transform -1 0 90896 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_969
timestamp 1624015447
transform 1 0 90252 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_969
timestamp 1624015447
transform 1 0 90252 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1624015447
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1624015447
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1624015447
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1624015447
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1624015447
transform 1 0 2484 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1624015447
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1624015447
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1624015447
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1624015447
transform 1 0 2484 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1399
timestamp 1624015447
transform 1 0 3772 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1624015447
transform 1 0 3588 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_27
timestamp 1624015447
transform 1 0 3588 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_30
timestamp 1624015447
transform 1 0 3864 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1624015447
transform 1 0 3588 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1624015447
transform -1 0 5152 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1624015447
transform -1 0 5152 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1624015447
transform -1 0 5152 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_39
timestamp 1624015447
transform 1 0 4692 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_38
timestamp 1624015447
transform 1 0 4600 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_39
timestamp 1624015447
transform 1 0 4692 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_782
timestamp 1624015447
transform 1 0 84180 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_784
timestamp 1624015447
transform 1 0 84180 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_786
timestamp 1624015447
transform 1 0 84180 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr1[3]
timestamp 1624015447
transform 1 0 84640 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_906
timestamp 1624015447
transform 1 0 84456 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_906
timestamp 1624015447
transform 1 0 84456 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_906
timestamp 1624015447
transform 1 0 84456 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_918
timestamp 1624015447
transform 1 0 85560 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_918
timestamp 1624015447
transform 1 0 85560 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_910
timestamp 1624015447
transform 1 0 84824 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_922
timestamp 1624015447
transform 1 0 85928 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1598
timestamp 1624015447
transform 1 0 86848 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_930
timestamp 1624015447
transform 1 0 86664 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_942
timestamp 1624015447
transform 1 0 87768 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_930
timestamp 1624015447
transform 1 0 86664 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_933
timestamp 1624015447
transform 1 0 86940 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_945
timestamp 1624015447
transform 1 0 88044 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_934
timestamp 1624015447
transform 1 0 87032 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_946
timestamp 1624015447
transform 1 0 88136 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1597
timestamp 1624015447
transform 1 0 89424 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1599
timestamp 1624015447
transform 1 0 89424 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_954
timestamp 1624015447
transform 1 0 88872 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_961
timestamp 1624015447
transform 1 0 89516 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_957
timestamp 1624015447
transform 1 0 89148 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_958
timestamp 1624015447
transform 1 0 89240 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_961
timestamp 1624015447
transform 1 0 89516 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_783
timestamp 1624015447
transform -1 0 90896 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_785
timestamp 1624015447
transform -1 0 90896 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_787
timestamp 1624015447
transform -1 0 90896 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_969
timestamp 1624015447
transform 1 0 90252 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1624015447
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1624015447
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1624015447
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1624015447
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1624015447
transform 1 0 2484 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1624015447
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1624015447
transform 1 0 2484 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1624015447
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1624015447
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1400
timestamp 1624015447
transform 1 0 3772 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1401
timestamp 1624015447
transform 1 0 3772 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_27
timestamp 1624015447
transform 1 0 3588 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_30
timestamp 1624015447
transform 1 0 3864 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1624015447
transform 1 0 3588 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_27
timestamp 1624015447
transform 1 0 3588 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_30
timestamp 1624015447
transform 1 0 3864 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1624015447
transform -1 0 5152 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1624015447
transform -1 0 5152 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1624015447
transform -1 0 5152 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_38
timestamp 1624015447
transform 1 0 4600 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_39
timestamp 1624015447
transform 1 0 4692 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_38
timestamp 1624015447
transform 1 0 4600 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_788
timestamp 1624015447
transform 1 0 84180 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_790
timestamp 1624015447
transform 1 0 84180 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_792
timestamp 1624015447
transform 1 0 84180 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr1[2]
timestamp 1624015447
transform 1 0 84640 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_906
timestamp 1624015447
transform 1 0 84456 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_906
timestamp 1624015447
transform 1 0 84456 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_906
timestamp 1624015447
transform 1 0 84456 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_918
timestamp 1624015447
transform 1 0 85560 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_910
timestamp 1624015447
transform 1 0 84824 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_922
timestamp 1624015447
transform 1 0 85928 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_918
timestamp 1624015447
transform 1 0 85560 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_945
timestamp 1624015447
transform 1 0 88044 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_933
timestamp 1624015447
transform 1 0 86940 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_930
timestamp 1624015447
transform 1 0 86664 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1600
timestamp 1624015447
transform 1 0 86848 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_946
timestamp 1624015447
transform 1 0 88136 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_934
timestamp 1624015447
transform 1 0 87032 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_945
timestamp 1624015447
transform 1 0 88044 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_933
timestamp 1624015447
transform 1 0 86940 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_930
timestamp 1624015447
transform 1 0 86664 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1602
timestamp 1624015447
transform 1 0 86848 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1601
timestamp 1624015447
transform 1 0 89424 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_957
timestamp 1624015447
transform 1 0 89148 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_958
timestamp 1624015447
transform 1 0 89240 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_961
timestamp 1624015447
transform 1 0 89516 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_957
timestamp 1624015447
transform 1 0 89148 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_789
timestamp 1624015447
transform -1 0 90896 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_791
timestamp 1624015447
transform -1 0 90896 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_793
timestamp 1624015447
transform -1 0 90896 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_969
timestamp 1624015447
transform 1 0 90252 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_969
timestamp 1624015447
transform 1 0 90252 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1624015447
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1624015447
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1624015447
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1624015447
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1624015447
transform 1 0 2484 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1624015447
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1624015447
transform 1 0 2484 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1624015447
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1624015447
transform 1 0 2484 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1402
timestamp 1624015447
transform 1 0 3772 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1624015447
transform 1 0 3588 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_27
timestamp 1624015447
transform 1 0 3588 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_30
timestamp 1624015447
transform 1 0 3864 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1624015447
transform 1 0 3588 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1624015447
transform -1 0 5152 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1624015447
transform -1 0 5152 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1624015447
transform -1 0 5152 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_39
timestamp 1624015447
transform 1 0 4692 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_38
timestamp 1624015447
transform 1 0 4600 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_39
timestamp 1624015447
transform 1 0 4692 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_794
timestamp 1624015447
transform 1 0 84180 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_796
timestamp 1624015447
transform 1 0 84180 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_798
timestamp 1624015447
transform 1 0 84180 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr1[1]
timestamp 1624015447
transform 1 0 84640 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_906
timestamp 1624015447
transform 1 0 84456 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_906
timestamp 1624015447
transform 1 0 84456 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_906
timestamp 1624015447
transform 1 0 84456 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_918
timestamp 1624015447
transform 1 0 85560 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_910
timestamp 1624015447
transform 1 0 84824 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_922
timestamp 1624015447
transform 1 0 85928 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_918
timestamp 1624015447
transform 1 0 85560 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1604
timestamp 1624015447
transform 1 0 86848 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_930
timestamp 1624015447
transform 1 0 86664 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_942
timestamp 1624015447
transform 1 0 87768 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_930
timestamp 1624015447
transform 1 0 86664 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_933
timestamp 1624015447
transform 1 0 86940 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_945
timestamp 1624015447
transform 1 0 88044 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_930
timestamp 1624015447
transform 1 0 86664 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_942
timestamp 1624015447
transform 1 0 87768 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1603
timestamp 1624015447
transform 1 0 89424 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1605
timestamp 1624015447
transform 1 0 89424 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_954
timestamp 1624015447
transform 1 0 88872 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_961
timestamp 1624015447
transform 1 0 89516 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_957
timestamp 1624015447
transform 1 0 89148 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_954
timestamp 1624015447
transform 1 0 88872 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_961
timestamp 1624015447
transform 1 0 89516 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_795
timestamp 1624015447
transform -1 0 90896 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_797
timestamp 1624015447
transform -1 0 90896 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_799
timestamp 1624015447
transform -1 0 90896 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_969
timestamp 1624015447
transform 1 0 90252 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1624015447
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1624015447
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1624015447
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1624015447
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1624015447
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1624015447
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1624015447
transform 1 0 2484 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1624015447
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1624015447
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1403
timestamp 1624015447
transform 1 0 3772 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1404
timestamp 1624015447
transform 1 0 3772 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_27
timestamp 1624015447
transform 1 0 3588 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_30
timestamp 1624015447
transform 1 0 3864 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1624015447
transform 1 0 3588 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_27
timestamp 1624015447
transform 1 0 3588 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_30
timestamp 1624015447
transform 1 0 3864 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1624015447
transform -1 0 5152 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1624015447
transform -1 0 5152 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1624015447
transform -1 0 5152 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_38
timestamp 1624015447
transform 1 0 4600 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_39
timestamp 1624015447
transform 1 0 4692 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_38
timestamp 1624015447
transform 1 0 4600 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_800
timestamp 1624015447
transform 1 0 84180 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_802
timestamp 1624015447
transform 1 0 84180 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_804
timestamp 1624015447
transform 1 0 84180 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_906
timestamp 1624015447
transform 1 0 84456 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_906
timestamp 1624015447
transform 1 0 84456 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_906
timestamp 1624015447
transform 1 0 84456 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_918
timestamp 1624015447
transform 1 0 85560 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_918
timestamp 1624015447
transform 1 0 85560 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_918
timestamp 1624015447
transform 1 0 85560 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_945
timestamp 1624015447
transform 1 0 88044 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_933
timestamp 1624015447
transform 1 0 86940 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_930
timestamp 1624015447
transform 1 0 86664 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1606
timestamp 1624015447
transform 1 0 86848 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_942
timestamp 1624015447
transform 1 0 87768 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_930
timestamp 1624015447
transform 1 0 86664 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_945
timestamp 1624015447
transform 1 0 88044 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_933
timestamp 1624015447
transform 1 0 86940 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_930
timestamp 1624015447
transform 1 0 86664 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1608
timestamp 1624015447
transform 1 0 86848 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1607
timestamp 1624015447
transform 1 0 89424 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_957
timestamp 1624015447
transform 1 0 89148 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_954
timestamp 1624015447
transform 1 0 88872 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_961
timestamp 1624015447
transform 1 0 89516 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_957
timestamp 1624015447
transform 1 0 89148 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_801
timestamp 1624015447
transform -1 0 90896 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_803
timestamp 1624015447
transform -1 0 90896 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_805
timestamp 1624015447
transform -1 0 90896 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_969
timestamp 1624015447
transform 1 0 90252 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_969
timestamp 1624015447
transform 1 0 90252 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1624015447
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1624015447
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1624015447
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1624015447
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1624015447
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1624015447
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1624015447
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1624015447
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1624015447
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1405
timestamp 1624015447
transform 1 0 3772 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1624015447
transform 1 0 3588 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_27
timestamp 1624015447
transform 1 0 3588 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_30
timestamp 1624015447
transform 1 0 3864 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1624015447
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1624015447
transform -1 0 5152 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1624015447
transform -1 0 5152 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1624015447
transform -1 0 5152 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_39
timestamp 1624015447
transform 1 0 4692 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_38
timestamp 1624015447
transform 1 0 4600 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_39
timestamp 1624015447
transform 1 0 4692 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_806
timestamp 1624015447
transform 1 0 84180 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_808
timestamp 1624015447
transform 1 0 84180 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_810
timestamp 1624015447
transform 1 0 84180 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_906
timestamp 1624015447
transform 1 0 84456 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_906
timestamp 1624015447
transform 1 0 84456 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_906
timestamp 1624015447
transform 1 0 84456 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_918
timestamp 1624015447
transform 1 0 85560 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_918
timestamp 1624015447
transform 1 0 85560 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_918
timestamp 1624015447
transform 1 0 85560 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1610
timestamp 1624015447
transform 1 0 86848 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_930
timestamp 1624015447
transform 1 0 86664 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_942
timestamp 1624015447
transform 1 0 87768 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_930
timestamp 1624015447
transform 1 0 86664 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_933
timestamp 1624015447
transform 1 0 86940 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_945
timestamp 1624015447
transform 1 0 88044 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_930
timestamp 1624015447
transform 1 0 86664 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_942
timestamp 1624015447
transform 1 0 87768 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1609
timestamp 1624015447
transform 1 0 89424 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1611
timestamp 1624015447
transform 1 0 89424 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_954
timestamp 1624015447
transform 1 0 88872 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_961
timestamp 1624015447
transform 1 0 89516 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_957
timestamp 1624015447
transform 1 0 89148 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_954
timestamp 1624015447
transform 1 0 88872 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_961
timestamp 1624015447
transform 1 0 89516 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_807
timestamp 1624015447
transform -1 0 90896 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_809
timestamp 1624015447
transform -1 0 90896 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_811
timestamp 1624015447
transform -1 0 90896 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_969
timestamp 1624015447
transform 1 0 90252 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1624015447
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1624015447
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1624015447
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1624015447
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1624015447
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1624015447
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1624015447
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1624015447
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1624015447
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1406
timestamp 1624015447
transform 1 0 3772 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1407
timestamp 1624015447
transform 1 0 3772 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_27
timestamp 1624015447
transform 1 0 3588 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_30
timestamp 1624015447
transform 1 0 3864 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1624015447
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_27
timestamp 1624015447
transform 1 0 3588 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_30
timestamp 1624015447
transform 1 0 3864 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1624015447
transform -1 0 5152 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1624015447
transform -1 0 5152 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1624015447
transform -1 0 5152 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_62_38
timestamp 1624015447
transform 1 0 4600 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_39
timestamp 1624015447
transform 1 0 4692 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_38
timestamp 1624015447
transform 1 0 4600 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_812
timestamp 1624015447
transform 1 0 84180 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_814
timestamp 1624015447
transform 1 0 84180 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_816
timestamp 1624015447
transform 1 0 84180 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_906
timestamp 1624015447
transform 1 0 84456 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_906
timestamp 1624015447
transform 1 0 84456 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_906
timestamp 1624015447
transform 1 0 84456 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_918
timestamp 1624015447
transform 1 0 85560 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_918
timestamp 1624015447
transform 1 0 85560 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_918
timestamp 1624015447
transform 1 0 85560 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_945
timestamp 1624015447
transform 1 0 88044 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_933
timestamp 1624015447
transform 1 0 86940 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_930
timestamp 1624015447
transform 1 0 86664 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1612
timestamp 1624015447
transform 1 0 86848 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_942
timestamp 1624015447
transform 1 0 87768 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_930
timestamp 1624015447
transform 1 0 86664 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_945
timestamp 1624015447
transform 1 0 88044 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_933
timestamp 1624015447
transform 1 0 86940 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_930
timestamp 1624015447
transform 1 0 86664 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1614
timestamp 1624015447
transform 1 0 86848 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1613
timestamp 1624015447
transform 1 0 89424 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_957
timestamp 1624015447
transform 1 0 89148 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_954
timestamp 1624015447
transform 1 0 88872 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_961
timestamp 1624015447
transform 1 0 89516 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_957
timestamp 1624015447
transform 1 0 89148 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_813
timestamp 1624015447
transform -1 0 90896 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_815
timestamp 1624015447
transform -1 0 90896 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_817
timestamp 1624015447
transform -1 0 90896 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_969
timestamp 1624015447
transform 1 0 90252 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_969
timestamp 1624015447
transform 1 0 90252 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1624015447
transform 1 0 1104 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1624015447
transform 1 0 1104 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1624015447
transform 1 0 1104 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1624015447
transform 1 0 1380 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1624015447
transform 1 0 2484 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1624015447
transform 1 0 1380 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1624015447
transform 1 0 2484 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1624015447
transform 1 0 1380 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1624015447
transform 1 0 2484 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1408
timestamp 1624015447
transform 1 0 3772 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1624015447
transform 1 0 3588 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_27
timestamp 1624015447
transform 1 0 3588 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_30
timestamp 1624015447
transform 1 0 3864 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1624015447
transform 1 0 3588 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1624015447
transform -1 0 5152 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1624015447
transform -1 0 5152 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1624015447
transform -1 0 5152 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_39
timestamp 1624015447
transform 1 0 4692 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_66_38
timestamp 1624015447
transform 1 0 4600 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_39
timestamp 1624015447
transform 1 0 4692 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1624015447
transform -1 0 84732 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_818
timestamp 1624015447
transform 1 0 84180 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_820
timestamp 1624015447
transform 1 0 84180 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_822
timestamp 1624015447
transform 1 0 84180 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_906
timestamp 1624015447
transform 1 0 84456 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_906
timestamp 1624015447
transform 1 0 84456 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_909
timestamp 1624015447
transform 1 0 84732 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_918
timestamp 1624015447
transform 1 0 85560 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_918
timestamp 1624015447
transform 1 0 85560 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_921
timestamp 1624015447
transform 1 0 85836 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1616
timestamp 1624015447
transform 1 0 86848 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_930
timestamp 1624015447
transform 1 0 86664 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_942
timestamp 1624015447
transform 1 0 87768 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_930
timestamp 1624015447
transform 1 0 86664 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_933
timestamp 1624015447
transform 1 0 86940 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_945
timestamp 1624015447
transform 1 0 88044 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_933
timestamp 1624015447
transform 1 0 86940 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_945
timestamp 1624015447
transform 1 0 88044 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1615
timestamp 1624015447
transform 1 0 89424 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1617
timestamp 1624015447
transform 1 0 89424 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_954
timestamp 1624015447
transform 1 0 88872 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_961
timestamp 1624015447
transform 1 0 89516 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_957
timestamp 1624015447
transform 1 0 89148 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_957
timestamp 1624015447
transform 1 0 89148 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_961
timestamp 1624015447
transform 1 0 89516 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_819
timestamp 1624015447
transform -1 0 90896 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_821
timestamp 1624015447
transform -1 0 90896 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_823
timestamp 1624015447
transform -1 0 90896 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_969
timestamp 1624015447
transform 1 0 90252 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1624015447
transform 1 0 1104 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1624015447
transform 1 0 1104 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1624015447
transform 1 0 1104 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1624015447
transform 1 0 1380 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1624015447
transform 1 0 2484 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1624015447
transform 1 0 1380 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1624015447
transform 1 0 2484 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_3
timestamp 1624015447
transform 1 0 1380 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_15
timestamp 1624015447
transform 1 0 2484 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1409
timestamp 1624015447
transform 1 0 3772 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1410
timestamp 1624015447
transform 1 0 3772 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_27
timestamp 1624015447
transform 1 0 3588 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_30
timestamp 1624015447
transform 1 0 3864 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1624015447
transform 1 0 3588 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_27
timestamp 1624015447
transform 1 0 3588 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_30
timestamp 1624015447
transform 1 0 3864 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1624015447
transform -1 0 5152 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1624015447
transform -1 0 5152 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1624015447
transform -1 0 5152 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_68_38
timestamp 1624015447
transform 1 0 4600 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_39
timestamp 1624015447
transform 1 0 4692 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_70_38
timestamp 1624015447
transform 1 0 4600 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_824
timestamp 1624015447
transform 1 0 84180 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_826
timestamp 1624015447
transform 1 0 84180 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_828
timestamp 1624015447
transform 1 0 84180 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_906
timestamp 1624015447
transform 1 0 84456 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_906
timestamp 1624015447
transform 1 0 84456 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_906
timestamp 1624015447
transform 1 0 84456 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_918
timestamp 1624015447
transform 1 0 85560 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_918
timestamp 1624015447
transform 1 0 85560 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_918
timestamp 1624015447
transform 1 0 85560 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_945
timestamp 1624015447
transform 1 0 88044 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_933
timestamp 1624015447
transform 1 0 86940 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_930
timestamp 1624015447
transform 1 0 86664 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1618
timestamp 1624015447
transform 1 0 86848 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_945
timestamp 1624015447
transform 1 0 88044 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_933
timestamp 1624015447
transform 1 0 86940 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_930
timestamp 1624015447
transform 1 0 86664 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_942
timestamp 1624015447
transform 1 0 87768 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_930
timestamp 1624015447
transform 1 0 86664 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1620
timestamp 1624015447
transform 1 0 86848 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1619
timestamp 1624015447
transform 1 0 89424 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_957
timestamp 1624015447
transform 1 0 89148 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_954
timestamp 1624015447
transform 1 0 88872 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_69_961
timestamp 1624015447
transform 1 0 89516 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_957
timestamp 1624015447
transform 1 0 89148 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_825
timestamp 1624015447
transform -1 0 90896 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_827
timestamp 1624015447
transform -1 0 90896 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_829
timestamp 1624015447
transform -1 0 90896 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_969
timestamp 1624015447
transform 1 0 90252 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_969
timestamp 1624015447
transform 1 0 90252 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1624015447
transform 1 0 1104 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1624015447
transform 1 0 1104 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1624015447
transform 1 0 1104 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1624015447
transform 1 0 1380 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_15
timestamp 1624015447
transform 1 0 2484 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1624015447
transform 1 0 1380 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_15
timestamp 1624015447
transform 1 0 2484 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_3
timestamp 1624015447
transform 1 0 1380 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_15
timestamp 1624015447
transform 1 0 2484 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1411
timestamp 1624015447
transform 1 0 3772 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_27
timestamp 1624015447
transform 1 0 3588 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_27
timestamp 1624015447
transform 1 0 3588 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_30
timestamp 1624015447
transform 1 0 3864 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_27
timestamp 1624015447
transform 1 0 3588 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1624015447
transform -1 0 5152 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1624015447
transform -1 0 5152 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1624015447
transform -1 0 5152 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_39
timestamp 1624015447
transform 1 0 4692 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_72_38
timestamp 1624015447
transform 1 0 4600 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_73_39
timestamp 1624015447
transform 1 0 4692 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_830
timestamp 1624015447
transform 1 0 84180 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_832
timestamp 1624015447
transform 1 0 84180 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_834
timestamp 1624015447
transform 1 0 84180 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_906
timestamp 1624015447
transform 1 0 84456 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_906
timestamp 1624015447
transform 1 0 84456 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_906
timestamp 1624015447
transform 1 0 84456 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_918
timestamp 1624015447
transform 1 0 85560 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_918
timestamp 1624015447
transform 1 0 85560 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_918
timestamp 1624015447
transform 1 0 85560 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1622
timestamp 1624015447
transform 1 0 86848 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_930
timestamp 1624015447
transform 1 0 86664 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_942
timestamp 1624015447
transform 1 0 87768 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_930
timestamp 1624015447
transform 1 0 86664 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_933
timestamp 1624015447
transform 1 0 86940 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_945
timestamp 1624015447
transform 1 0 88044 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_930
timestamp 1624015447
transform 1 0 86664 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_942
timestamp 1624015447
transform 1 0 87768 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1621
timestamp 1624015447
transform 1 0 89424 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1623
timestamp 1624015447
transform 1 0 89424 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_954
timestamp 1624015447
transform 1 0 88872 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_961
timestamp 1624015447
transform 1 0 89516 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_957
timestamp 1624015447
transform 1 0 89148 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_954
timestamp 1624015447
transform 1 0 88872 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_73_961
timestamp 1624015447
transform 1 0 89516 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_831
timestamp 1624015447
transform -1 0 90896 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_833
timestamp 1624015447
transform -1 0 90896 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_835
timestamp 1624015447
transform -1 0 90896 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_969
timestamp 1624015447
transform 1 0 90252 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1624015447
transform 1 0 1104 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1624015447
transform 1 0 1104 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1624015447
transform 1 0 1104 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1624015447
transform 1 0 1380 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1624015447
transform 1 0 2484 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_3
timestamp 1624015447
transform 1 0 1380 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_15
timestamp 1624015447
transform 1 0 2484 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1624015447
transform 1 0 1380 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1624015447
transform 1 0 2484 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1412
timestamp 1624015447
transform 1 0 3772 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1413
timestamp 1624015447
transform 1 0 3772 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_27
timestamp 1624015447
transform 1 0 3588 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_30
timestamp 1624015447
transform 1 0 3864 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_27
timestamp 1624015447
transform 1 0 3588 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_27
timestamp 1624015447
transform 1 0 3588 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_76_30
timestamp 1624015447
transform 1 0 3864 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1624015447
transform -1 0 5152 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1624015447
transform -1 0 5152 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1624015447
transform -1 0 5152 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_74_38
timestamp 1624015447
transform 1 0 4600 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_39
timestamp 1624015447
transform 1 0 4692 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_76_38
timestamp 1624015447
transform 1 0 4600 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_836
timestamp 1624015447
transform 1 0 84180 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_838
timestamp 1624015447
transform 1 0 84180 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_840
timestamp 1624015447
transform 1 0 84180 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_906
timestamp 1624015447
transform 1 0 84456 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_906
timestamp 1624015447
transform 1 0 84456 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_906
timestamp 1624015447
transform 1 0 84456 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_918
timestamp 1624015447
transform 1 0 85560 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_918
timestamp 1624015447
transform 1 0 85560 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_918
timestamp 1624015447
transform 1 0 85560 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_942
timestamp 1624015447
transform 1 0 87768 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_930
timestamp 1624015447
transform 1 0 86664 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_945
timestamp 1624015447
transform 1 0 88044 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_933
timestamp 1624015447
transform 1 0 86940 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_930
timestamp 1624015447
transform 1 0 86664 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1624
timestamp 1624015447
transform 1 0 86848 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_945
timestamp 1624015447
transform 1 0 88044 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_933
timestamp 1624015447
transform 1 0 86940 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_930
timestamp 1624015447
transform 1 0 86664 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1626
timestamp 1624015447
transform 1 0 86848 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1625
timestamp 1624015447
transform 1 0 89424 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_957
timestamp 1624015447
transform 1 0 89148 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_954
timestamp 1624015447
transform 1 0 88872 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_961
timestamp 1624015447
transform 1 0 89516 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_957
timestamp 1624015447
transform 1 0 89148 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_837
timestamp 1624015447
transform -1 0 90896 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_839
timestamp 1624015447
transform -1 0 90896 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_841
timestamp 1624015447
transform -1 0 90896 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_969
timestamp 1624015447
transform 1 0 90252 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_969
timestamp 1624015447
transform 1 0 90252 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1624015447
transform 1 0 2484 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_3
timestamp 1624015447
transform 1 0 1380 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1624015447
transform 1 0 2484 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1624015447
transform 1 0 1380 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1624015447
transform 1 0 1104 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1624015447
transform 1 0 1104 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_15
timestamp 1624015447
transform 1 0 2484 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_3
timestamp 1624015447
transform 1 0 1380 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1624015447
transform 1 0 1104 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_15
timestamp 1624015447
transform 1 0 2484 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_3
timestamp 1624015447
transform 1 0 1380 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1624015447
transform 1 0 1104 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1414
timestamp 1624015447
transform 1 0 3772 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1415
timestamp 1624015447
transform 1 0 3772 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1624015447
transform 1 0 3588 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_27
timestamp 1624015447
transform 1 0 3588 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_78_30
timestamp 1624015447
transform 1 0 3864 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_27
timestamp 1624015447
transform 1 0 3588 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_27
timestamp 1624015447
transform 1 0 3588 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_30
timestamp 1624015447
transform 1 0 3864 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1624015447
transform -1 0 5152 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1624015447
transform -1 0 5152 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1624015447
transform -1 0 5152 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1624015447
transform -1 0 5152 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_77_39
timestamp 1624015447
transform 1 0 4692 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_78_38
timestamp 1624015447
transform 1 0 4600 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_39
timestamp 1624015447
transform 1 0 4692 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_80_38
timestamp 1624015447
transform 1 0 4600 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_842
timestamp 1624015447
transform 1 0 84180 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_844
timestamp 1624015447
transform 1 0 84180 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_846
timestamp 1624015447
transform 1 0 84180 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_848
timestamp 1624015447
transform 1 0 84180 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_906
timestamp 1624015447
transform 1 0 84456 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_906
timestamp 1624015447
transform 1 0 84456 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_906
timestamp 1624015447
transform 1 0 84456 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_906
timestamp 1624015447
transform 1 0 84456 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_918
timestamp 1624015447
transform 1 0 85560 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_918
timestamp 1624015447
transform 1 0 85560 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_918
timestamp 1624015447
transform 1 0 85560 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_918
timestamp 1624015447
transform 1 0 85560 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_945
timestamp 1624015447
transform 1 0 88044 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_933
timestamp 1624015447
transform 1 0 86940 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_930
timestamp 1624015447
transform 1 0 86664 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_77_942
timestamp 1624015447
transform 1 0 87768 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_930
timestamp 1624015447
transform 1 0 86664 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1628
timestamp 1624015447
transform 1 0 86848 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_942
timestamp 1624015447
transform 1 0 87768 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_930
timestamp 1624015447
transform 1 0 86664 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_945
timestamp 1624015447
transform 1 0 88044 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_933
timestamp 1624015447
transform 1 0 86940 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_930
timestamp 1624015447
transform 1 0 86664 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1630
timestamp 1624015447
transform 1 0 86848 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1627
timestamp 1624015447
transform 1 0 89424 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1629
timestamp 1624015447
transform 1 0 89424 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_954
timestamp 1624015447
transform 1 0 88872 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_77_961
timestamp 1624015447
transform 1 0 89516 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_957
timestamp 1624015447
transform 1 0 89148 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_954
timestamp 1624015447
transform 1 0 88872 0 1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_79_961
timestamp 1624015447
transform 1 0 89516 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_957
timestamp 1624015447
transform 1 0 89148 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_843
timestamp 1624015447
transform -1 0 90896 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_845
timestamp 1624015447
transform -1 0 90896 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_847
timestamp 1624015447
transform -1 0 90896 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_849
timestamp 1624015447
transform -1 0 90896 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_969
timestamp 1624015447
transform 1 0 90252 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_969
timestamp 1624015447
transform 1 0 90252 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1624015447
transform 1 0 1104 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1624015447
transform 1 0 1104 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1624015447
transform 1 0 1104 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_3
timestamp 1624015447
transform 1 0 1380 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_15
timestamp 1624015447
transform 1 0 2484 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_3
timestamp 1624015447
transform 1 0 1380 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_15
timestamp 1624015447
transform 1 0 2484 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_3
timestamp 1624015447
transform 1 0 1380 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_15
timestamp 1624015447
transform 1 0 2484 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1416
timestamp 1624015447
transform 1 0 3772 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_27
timestamp 1624015447
transform 1 0 3588 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_27
timestamp 1624015447
transform 1 0 3588 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_30
timestamp 1624015447
transform 1 0 3864 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_27
timestamp 1624015447
transform 1 0 3588 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1624015447
transform -1 0 5152 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1624015447
transform -1 0 5152 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1624015447
transform -1 0 5152 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_81_39
timestamp 1624015447
transform 1 0 4692 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_82_38
timestamp 1624015447
transform 1 0 4600 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_83_39
timestamp 1624015447
transform 1 0 4692 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_850
timestamp 1624015447
transform 1 0 84180 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_852
timestamp 1624015447
transform 1 0 84180 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_854
timestamp 1624015447
transform 1 0 84180 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_906
timestamp 1624015447
transform 1 0 84456 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_906
timestamp 1624015447
transform 1 0 84456 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_906
timestamp 1624015447
transform 1 0 84456 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_918
timestamp 1624015447
transform 1 0 85560 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_918
timestamp 1624015447
transform 1 0 85560 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_918
timestamp 1624015447
transform 1 0 85560 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1632
timestamp 1624015447
transform 1 0 86848 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_930
timestamp 1624015447
transform 1 0 86664 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_942
timestamp 1624015447
transform 1 0 87768 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_930
timestamp 1624015447
transform 1 0 86664 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_933
timestamp 1624015447
transform 1 0 86940 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_945
timestamp 1624015447
transform 1 0 88044 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_930
timestamp 1624015447
transform 1 0 86664 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_942
timestamp 1624015447
transform 1 0 87768 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1631
timestamp 1624015447
transform 1 0 89424 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1633
timestamp 1624015447
transform 1 0 89424 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_954
timestamp 1624015447
transform 1 0 88872 0 1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_81_961
timestamp 1624015447
transform 1 0 89516 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_957
timestamp 1624015447
transform 1 0 89148 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_954
timestamp 1624015447
transform 1 0 88872 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_83_961
timestamp 1624015447
transform 1 0 89516 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_851
timestamp 1624015447
transform -1 0 90896 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_853
timestamp 1624015447
transform -1 0 90896 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_855
timestamp 1624015447
transform -1 0 90896 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_969
timestamp 1624015447
transform 1 0 90252 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_15
timestamp 1624015447
transform 1 0 2484 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_3
timestamp 1624015447
transform 1 0 1380 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_15
timestamp 1624015447
transform 1 0 2484 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_3
timestamp 1624015447
transform 1 0 1380 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1624015447
transform 1 0 1104 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1624015447
transform 1 0 1104 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_86_15
timestamp 1624015447
transform 1 0 2484 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_3
timestamp 1624015447
transform 1 0 1380 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1624015447
transform 1 0 1104 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_87_15
timestamp 1624015447
transform 1 0 2484 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_3
timestamp 1624015447
transform 1 0 1380 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1624015447
transform 1 0 1104 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_85_27
timestamp 1624015447
transform 1 0 3588 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_30
timestamp 1624015447
transform 1 0 3864 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_27
timestamp 1624015447
transform 1 0 3588 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1417
timestamp 1624015447
transform 1 0 3772 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_30
timestamp 1624015447
transform 1 0 3864 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_27
timestamp 1624015447
transform 1 0 3588 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1418
timestamp 1624015447
transform 1 0 3772 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_37
timestamp 1624015447
transform 1 0 4508 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_33
timestamp 1624015447
transform 1 0 4140 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_87_27
timestamp 1624015447
transform 1 0 3588 0 1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _16_
timestamp 1624015447
transform 1 0 4232 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1624015447
transform -1 0 5152 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1624015447
transform -1 0 5152 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1624015447
transform -1 0 5152 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1624015447
transform -1 0 5152 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_84_38
timestamp 1624015447
transform 1 0 4600 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_85_39
timestamp 1624015447
transform 1 0 4692 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_86_38
timestamp 1624015447
transform 1 0 4600 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_856
timestamp 1624015447
transform 1 0 84180 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_858
timestamp 1624015447
transform 1 0 84180 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_860
timestamp 1624015447
transform 1 0 84180 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_862
timestamp 1624015447
transform 1 0 84180 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_906
timestamp 1624015447
transform 1 0 84456 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_906
timestamp 1624015447
transform 1 0 84456 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_906
timestamp 1624015447
transform 1 0 84456 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_906
timestamp 1624015447
transform 1 0 84456 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_918
timestamp 1624015447
transform 1 0 85560 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_84_930
timestamp 1624015447
transform 1 0 86664 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_85_918
timestamp 1624015447
transform 1 0 85560 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_930
timestamp 1624015447
transform 1 0 86664 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_918
timestamp 1624015447
transform 1 0 85560 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_86_930
timestamp 1624015447
transform 1 0 86664 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_87_918
timestamp 1624015447
transform 1 0 85560 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_930
timestamp 1624015447
transform 1 0 86664 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1634
timestamp 1624015447
transform 1 0 86848 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1636
timestamp 1624015447
transform 1 0 86848 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_933
timestamp 1624015447
transform 1 0 86940 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_945
timestamp 1624015447
transform 1 0 88044 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_942
timestamp 1624015447
transform 1 0 87768 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_933
timestamp 1624015447
transform 1 0 86940 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_945
timestamp 1624015447
transform 1 0 88044 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_942
timestamp 1624015447
transform 1 0 87768 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1635
timestamp 1624015447
transform 1 0 89424 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1637
timestamp 1624015447
transform 1 0 89424 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_957
timestamp 1624015447
transform 1 0 89148 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_954
timestamp 1624015447
transform 1 0 88872 0 1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_85_961
timestamp 1624015447
transform 1 0 89516 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_957
timestamp 1624015447
transform 1 0 89148 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_954
timestamp 1624015447
transform 1 0 88872 0 1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_87_961
timestamp 1624015447
transform 1 0 89516 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_857
timestamp 1624015447
transform -1 0 90896 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_859
timestamp 1624015447
transform -1 0 90896 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_861
timestamp 1624015447
transform -1 0 90896 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_863
timestamp 1624015447
transform -1 0 90896 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_84_969
timestamp 1624015447
transform 1 0 90252 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_969
timestamp 1624015447
transform 1 0 90252 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1624015447
transform 1 0 1104 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1624015447
transform 1 0 1104 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1624015447
transform 1 0 1104 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_88_3
timestamp 1624015447
transform 1 0 1380 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_15
timestamp 1624015447
transform 1 0 2484 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_3
timestamp 1624015447
transform 1 0 1380 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_15
timestamp 1624015447
transform 1 0 2484 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_3
timestamp 1624015447
transform 1 0 1380 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_15
timestamp 1624015447
transform 1 0 2484 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1419
timestamp 1624015447
transform 1 0 3772 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1420
timestamp 1624015447
transform 1 0 3772 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_88_27
timestamp 1624015447
transform 1 0 3588 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_88_30
timestamp 1624015447
transform 1 0 3864 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_89_27
timestamp 1624015447
transform 1 0 3588 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_90_27
timestamp 1624015447
transform 1 0 3588 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_90_30
timestamp 1624015447
transform 1 0 3864 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1624015447
transform -1 0 5152 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1624015447
transform -1 0 5152 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1624015447
transform -1 0 5152 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_88_38
timestamp 1624015447
transform 1 0 4600 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_89_39
timestamp 1624015447
transform 1 0 4692 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_90_38
timestamp 1624015447
transform 1 0 4600 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_864
timestamp 1624015447
transform 1 0 84180 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_866
timestamp 1624015447
transform 1 0 84180 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_868
timestamp 1624015447
transform 1 0 84180 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_88_906
timestamp 1624015447
transform 1 0 84456 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_906
timestamp 1624015447
transform 1 0 84456 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_906
timestamp 1624015447
transform 1 0 84456 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_918
timestamp 1624015447
transform 1 0 85560 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_88_930
timestamp 1624015447
transform 1 0 86664 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_89_918
timestamp 1624015447
transform 1 0 85560 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_930
timestamp 1624015447
transform 1 0 86664 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_918
timestamp 1624015447
transform 1 0 85560 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_90_930
timestamp 1624015447
transform 1 0 86664 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1638
timestamp 1624015447
transform 1 0 86848 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1640
timestamp 1624015447
transform 1 0 86848 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_933
timestamp 1624015447
transform 1 0 86940 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_945
timestamp 1624015447
transform 1 0 88044 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_942
timestamp 1624015447
transform 1 0 87768 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_933
timestamp 1624015447
transform 1 0 86940 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_945
timestamp 1624015447
transform 1 0 88044 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1639
timestamp 1624015447
transform 1 0 89424 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_957
timestamp 1624015447
transform 1 0 89148 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_954
timestamp 1624015447
transform 1 0 88872 0 1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_89_961
timestamp 1624015447
transform 1 0 89516 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_957
timestamp 1624015447
transform 1 0 89148 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_865
timestamp 1624015447
transform -1 0 90896 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_867
timestamp 1624015447
transform -1 0 90896 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_869
timestamp 1624015447
transform -1 0 90896 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_88_969
timestamp 1624015447
transform 1 0 90252 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_969
timestamp 1624015447
transform 1 0 90252 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1624015447
transform 1 0 1104 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1624015447
transform 1 0 1104 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1624015447
transform 1 0 1104 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_3
timestamp 1624015447
transform 1 0 1380 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_15
timestamp 1624015447
transform 1 0 2484 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_3
timestamp 1624015447
transform 1 0 1380 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_15
timestamp 1624015447
transform 1 0 2484 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_3
timestamp 1624015447
transform 1 0 1380 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_15
timestamp 1624015447
transform 1 0 2484 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1421
timestamp 1624015447
transform 1 0 3772 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_27
timestamp 1624015447
transform 1 0 3588 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_92_27
timestamp 1624015447
transform 1 0 3588 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_92_30
timestamp 1624015447
transform 1 0 3864 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_27
timestamp 1624015447
transform 1 0 3588 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1624015447
transform -1 0 5152 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1624015447
transform -1 0 5152 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1624015447
transform -1 0 5152 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_91_39
timestamp 1624015447
transform 1 0 4692 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_92_38
timestamp 1624015447
transform 1 0 4600 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_93_39
timestamp 1624015447
transform 1 0 4692 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_870
timestamp 1624015447
transform 1 0 84180 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_872
timestamp 1624015447
transform 1 0 84180 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_874
timestamp 1624015447
transform 1 0 84180 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_906
timestamp 1624015447
transform 1 0 84456 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_906
timestamp 1624015447
transform 1 0 84456 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_906
timestamp 1624015447
transform 1 0 84456 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_918
timestamp 1624015447
transform 1 0 85560 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_930
timestamp 1624015447
transform 1 0 86664 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_918
timestamp 1624015447
transform 1 0 85560 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_92_930
timestamp 1624015447
transform 1 0 86664 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_93_918
timestamp 1624015447
transform 1 0 85560 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_930
timestamp 1624015447
transform 1 0 86664 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1642
timestamp 1624015447
transform 1 0 86848 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_942
timestamp 1624015447
transform 1 0 87768 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_933
timestamp 1624015447
transform 1 0 86940 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_945
timestamp 1624015447
transform 1 0 88044 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_942
timestamp 1624015447
transform 1 0 87768 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1641
timestamp 1624015447
transform 1 0 89424 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1643
timestamp 1624015447
transform 1 0 89424 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_91_954
timestamp 1624015447
transform 1 0 88872 0 1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_91_961
timestamp 1624015447
transform 1 0 89516 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_957
timestamp 1624015447
transform 1 0 89148 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_954
timestamp 1624015447
transform 1 0 88872 0 1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_93_961
timestamp 1624015447
transform 1 0 89516 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_871
timestamp 1624015447
transform -1 0 90896 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_873
timestamp 1624015447
transform -1 0 90896 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_875
timestamp 1624015447
transform -1 0 90896 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_92_969
timestamp 1624015447
transform 1 0 90252 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1624015447
transform 1 0 1104 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1624015447
transform 1 0 1104 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1624015447
transform 1 0 1104 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_94_3
timestamp 1624015447
transform 1 0 1380 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_15
timestamp 1624015447
transform 1 0 2484 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_3
timestamp 1624015447
transform 1 0 1380 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_15
timestamp 1624015447
transform 1 0 2484 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_3
timestamp 1624015447
transform 1 0 1380 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_15
timestamp 1624015447
transform 1 0 2484 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1422
timestamp 1624015447
transform 1 0 3772 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1423
timestamp 1624015447
transform 1 0 3772 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_27
timestamp 1624015447
transform 1 0 3588 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_94_30
timestamp 1624015447
transform 1 0 3864 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_27
timestamp 1624015447
transform 1 0 3588 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_96_27
timestamp 1624015447
transform 1 0 3588 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_96_30
timestamp 1624015447
transform 1 0 3864 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1624015447
transform -1 0 5152 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1624015447
transform -1 0 5152 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1624015447
transform -1 0 5152 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_94_38
timestamp 1624015447
transform 1 0 4600 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_39
timestamp 1624015447
transform 1 0 4692 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_96_38
timestamp 1624015447
transform 1 0 4600 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_876
timestamp 1624015447
transform 1 0 84180 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_878
timestamp 1624015447
transform 1 0 84180 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_880
timestamp 1624015447
transform 1 0 84180 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_94_906
timestamp 1624015447
transform 1 0 84456 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_906
timestamp 1624015447
transform 1 0 84456 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_906
timestamp 1624015447
transform 1 0 84456 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_918
timestamp 1624015447
transform 1 0 85560 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_94_930
timestamp 1624015447
transform 1 0 86664 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_95_918
timestamp 1624015447
transform 1 0 85560 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_930
timestamp 1624015447
transform 1 0 86664 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_918
timestamp 1624015447
transform 1 0 85560 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_96_930
timestamp 1624015447
transform 1 0 86664 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1644
timestamp 1624015447
transform 1 0 86848 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1646
timestamp 1624015447
transform 1 0 86848 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_933
timestamp 1624015447
transform 1 0 86940 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_945
timestamp 1624015447
transform 1 0 88044 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_942
timestamp 1624015447
transform 1 0 87768 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_933
timestamp 1624015447
transform 1 0 86940 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_945
timestamp 1624015447
transform 1 0 88044 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1645
timestamp 1624015447
transform 1 0 89424 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_957
timestamp 1624015447
transform 1 0 89148 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_954
timestamp 1624015447
transform 1 0 88872 0 1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_95_961
timestamp 1624015447
transform 1 0 89516 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_957
timestamp 1624015447
transform 1 0 89148 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_877
timestamp 1624015447
transform -1 0 90896 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_879
timestamp 1624015447
transform -1 0 90896 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_881
timestamp 1624015447
transform -1 0 90896 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_94_969
timestamp 1624015447
transform 1 0 90252 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_969
timestamp 1624015447
transform 1 0 90252 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1624015447
transform 1 0 1104 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1624015447
transform 1 0 1104 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1624015447
transform 1 0 1104 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_3
timestamp 1624015447
transform 1 0 1380 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_15
timestamp 1624015447
transform 1 0 2484 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_3
timestamp 1624015447
transform 1 0 1380 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_15
timestamp 1624015447
transform 1 0 2484 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_3
timestamp 1624015447
transform 1 0 1380 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_15
timestamp 1624015447
transform 1 0 2484 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1424
timestamp 1624015447
transform 1 0 3772 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_27
timestamp 1624015447
transform 1 0 3588 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_98_27
timestamp 1624015447
transform 1 0 3588 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_98_30
timestamp 1624015447
transform 1 0 3864 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_99_27
timestamp 1624015447
transform 1 0 3588 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1624015447
transform -1 0 5152 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1624015447
transform -1 0 5152 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1624015447
transform -1 0 5152 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_97_39
timestamp 1624015447
transform 1 0 4692 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_98_38
timestamp 1624015447
transform 1 0 4600 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_99_39
timestamp 1624015447
transform 1 0 4692 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_882
timestamp 1624015447
transform 1 0 84180 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_884
timestamp 1624015447
transform 1 0 84180 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_886
timestamp 1624015447
transform 1 0 84180 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_906
timestamp 1624015447
transform 1 0 84456 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_906
timestamp 1624015447
transform 1 0 84456 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_906
timestamp 1624015447
transform 1 0 84456 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_918
timestamp 1624015447
transform 1 0 85560 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_930
timestamp 1624015447
transform 1 0 86664 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_918
timestamp 1624015447
transform 1 0 85560 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_98_930
timestamp 1624015447
transform 1 0 86664 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_99_918
timestamp 1624015447
transform 1 0 85560 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_930
timestamp 1624015447
transform 1 0 86664 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1648
timestamp 1624015447
transform 1 0 86848 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_942
timestamp 1624015447
transform 1 0 87768 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_933
timestamp 1624015447
transform 1 0 86940 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_945
timestamp 1624015447
transform 1 0 88044 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_942
timestamp 1624015447
transform 1 0 87768 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1647
timestamp 1624015447
transform 1 0 89424 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1649
timestamp 1624015447
transform 1 0 89424 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_97_954
timestamp 1624015447
transform 1 0 88872 0 1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_97_961
timestamp 1624015447
transform 1 0 89516 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_957
timestamp 1624015447
transform 1 0 89148 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_954
timestamp 1624015447
transform 1 0 88872 0 1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_99_961
timestamp 1624015447
transform 1 0 89516 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_883
timestamp 1624015447
transform -1 0 90896 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_885
timestamp 1624015447
transform -1 0 90896 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_887
timestamp 1624015447
transform -1 0 90896 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_98_969
timestamp 1624015447
transform 1 0 90252 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1624015447
transform 1 0 1104 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1624015447
transform 1 0 1104 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1624015447
transform 1 0 1104 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_3
timestamp 1624015447
transform 1 0 1380 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_15
timestamp 1624015447
transform 1 0 2484 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_3
timestamp 1624015447
transform 1 0 1380 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_15
timestamp 1624015447
transform 1 0 2484 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_3
timestamp 1624015447
transform 1 0 1380 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_15
timestamp 1624015447
transform 1 0 2484 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1624015447
transform 1 0 4232 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1425
timestamp 1624015447
transform 1 0 3772 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1426
timestamp 1624015447
transform 1 0 3772 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_100_27
timestamp 1624015447
transform 1 0 3588 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_100_30
timestamp 1624015447
transform 1 0 3864 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_101_27
timestamp 1624015447
transform 1 0 3588 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_102_27
timestamp 1624015447
transform 1 0 3588 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_102_30
timestamp 1624015447
transform 1 0 3864 0 -1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_102_37
timestamp 1624015447
transform 1 0 4508 0 -1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1624015447
transform -1 0 5152 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1624015447
transform -1 0 5152 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1624015447
transform -1 0 5152 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_100_38
timestamp 1624015447
transform 1 0 4600 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_39
timestamp 1624015447
transform 1 0 4692 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_888
timestamp 1624015447
transform 1 0 84180 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_890
timestamp 1624015447
transform 1 0 84180 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_892
timestamp 1624015447
transform 1 0 84180 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_906
timestamp 1624015447
transform 1 0 84456 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_906
timestamp 1624015447
transform 1 0 84456 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_906
timestamp 1624015447
transform 1 0 84456 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_918
timestamp 1624015447
transform 1 0 85560 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_930
timestamp 1624015447
transform 1 0 86664 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_101_918
timestamp 1624015447
transform 1 0 85560 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_930
timestamp 1624015447
transform 1 0 86664 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_918
timestamp 1624015447
transform 1 0 85560 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_102_930
timestamp 1624015447
transform 1 0 86664 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1650
timestamp 1624015447
transform 1 0 86848 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1652
timestamp 1624015447
transform 1 0 86848 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_933
timestamp 1624015447
transform 1 0 86940 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_945
timestamp 1624015447
transform 1 0 88044 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_942
timestamp 1624015447
transform 1 0 87768 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_933
timestamp 1624015447
transform 1 0 86940 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_945
timestamp 1624015447
transform 1 0 88044 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1651
timestamp 1624015447
transform 1 0 89424 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_957
timestamp 1624015447
transform 1 0 89148 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_954
timestamp 1624015447
transform 1 0 88872 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_101_961
timestamp 1624015447
transform 1 0 89516 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_957
timestamp 1624015447
transform 1 0 89148 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_889
timestamp 1624015447
transform -1 0 90896 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_891
timestamp 1624015447
transform -1 0 90896 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_893
timestamp 1624015447
transform -1 0 90896 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_100_969
timestamp 1624015447
transform 1 0 90252 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_102_969
timestamp 1624015447
transform 1 0 90252 0 -1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1624015447
transform 1 0 1104 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1624015447
transform 1 0 1104 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1624015447
transform 1 0 1104 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_3
timestamp 1624015447
transform 1 0 1380 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_15
timestamp 1624015447
transform 1 0 2484 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_3
timestamp 1624015447
transform 1 0 1380 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_15
timestamp 1624015447
transform 1 0 2484 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_3
timestamp 1624015447
transform 1 0 1380 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_15
timestamp 1624015447
transform 1 0 2484 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1427
timestamp 1624015447
transform 1 0 3772 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_27
timestamp 1624015447
transform 1 0 3588 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_104_27
timestamp 1624015447
transform 1 0 3588 0 -1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_104_30
timestamp 1624015447
transform 1 0 3864 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_105_27
timestamp 1624015447
transform 1 0 3588 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1624015447
transform -1 0 5152 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1624015447
transform -1 0 5152 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1624015447
transform -1 0 5152 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_103_39
timestamp 1624015447
transform 1 0 4692 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_104_38
timestamp 1624015447
transform 1 0 4600 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_105_39
timestamp 1624015447
transform 1 0 4692 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_894
timestamp 1624015447
transform 1 0 84180 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_896
timestamp 1624015447
transform 1 0 84180 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_898
timestamp 1624015447
transform 1 0 84180 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_906
timestamp 1624015447
transform 1 0 84456 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_906
timestamp 1624015447
transform 1 0 84456 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_906
timestamp 1624015447
transform 1 0 84456 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_918
timestamp 1624015447
transform 1 0 85560 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_930
timestamp 1624015447
transform 1 0 86664 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_918
timestamp 1624015447
transform 1 0 85560 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_104_930
timestamp 1624015447
transform 1 0 86664 0 -1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_105_918
timestamp 1624015447
transform 1 0 85560 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_930
timestamp 1624015447
transform 1 0 86664 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1654
timestamp 1624015447
transform 1 0 86848 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_942
timestamp 1624015447
transform 1 0 87768 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_933
timestamp 1624015447
transform 1 0 86940 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_945
timestamp 1624015447
transform 1 0 88044 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_942
timestamp 1624015447
transform 1 0 87768 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1653
timestamp 1624015447
transform 1 0 89424 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1655
timestamp 1624015447
transform 1 0 89424 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_103_954
timestamp 1624015447
transform 1 0 88872 0 1 58208
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_103_961
timestamp 1624015447
transform 1 0 89516 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_957
timestamp 1624015447
transform 1 0 89148 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_954
timestamp 1624015447
transform 1 0 88872 0 1 59296
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_105_961
timestamp 1624015447
transform 1 0 89516 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_895
timestamp 1624015447
transform -1 0 90896 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_897
timestamp 1624015447
transform -1 0 90896 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_899
timestamp 1624015447
transform -1 0 90896 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_104_969
timestamp 1624015447
transform 1 0 90252 0 -1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_107_15
timestamp 1624015447
transform 1 0 2484 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_3
timestamp 1624015447
transform 1 0 1380 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_15
timestamp 1624015447
transform 1 0 2484 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_3
timestamp 1624015447
transform 1 0 1380 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1624015447
transform 1 0 1104 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1624015447
transform 1 0 1104 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_108_15
timestamp 1624015447
transform 1 0 2484 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_3
timestamp 1624015447
transform 1 0 1380 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1624015447
transform 1 0 1104 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_109_15
timestamp 1624015447
transform 1 0 2484 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_3
timestamp 1624015447
transform 1 0 1380 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1624015447
transform 1 0 1104 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1428
timestamp 1624015447
transform 1 0 3772 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1429
timestamp 1624015447
transform 1 0 3772 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_106_27
timestamp 1624015447
transform 1 0 3588 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_106_30
timestamp 1624015447
transform 1 0 3864 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_107_27
timestamp 1624015447
transform 1 0 3588 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_108_27
timestamp 1624015447
transform 1 0 3588 0 -1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_108_30
timestamp 1624015447
transform 1 0 3864 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_109_27
timestamp 1624015447
transform 1 0 3588 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1624015447
transform -1 0 5152 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1624015447
transform -1 0 5152 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1624015447
transform -1 0 5152 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1624015447
transform -1 0 5152 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_106_38
timestamp 1624015447
transform 1 0 4600 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_107_39
timestamp 1624015447
transform 1 0 4692 0 1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_108_38
timestamp 1624015447
transform 1 0 4600 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_109_39
timestamp 1624015447
transform 1 0 4692 0 1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_900
timestamp 1624015447
transform 1 0 84180 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_902
timestamp 1624015447
transform 1 0 84180 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_904
timestamp 1624015447
transform 1 0 84180 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_906
timestamp 1624015447
transform 1 0 84180 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_106_906
timestamp 1624015447
transform 1 0 84456 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_906
timestamp 1624015447
transform 1 0 84456 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_906
timestamp 1624015447
transform 1 0 84456 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_906
timestamp 1624015447
transform 1 0 84456 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_918
timestamp 1624015447
transform 1 0 85560 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_106_930
timestamp 1624015447
transform 1 0 86664 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_107_918
timestamp 1624015447
transform 1 0 85560 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_930
timestamp 1624015447
transform 1 0 86664 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_918
timestamp 1624015447
transform 1 0 85560 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_108_930
timestamp 1624015447
transform 1 0 86664 0 -1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_109_918
timestamp 1624015447
transform 1 0 85560 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_930
timestamp 1624015447
transform 1 0 86664 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1656
timestamp 1624015447
transform 1 0 86848 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1658
timestamp 1624015447
transform 1 0 86848 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_933
timestamp 1624015447
transform 1 0 86940 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_945
timestamp 1624015447
transform 1 0 88044 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_942
timestamp 1624015447
transform 1 0 87768 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_933
timestamp 1624015447
transform 1 0 86940 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_945
timestamp 1624015447
transform 1 0 88044 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_942
timestamp 1624015447
transform 1 0 87768 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1657
timestamp 1624015447
transform 1 0 89424 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1659
timestamp 1624015447
transform 1 0 89424 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_957
timestamp 1624015447
transform 1 0 89148 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_954
timestamp 1624015447
transform 1 0 88872 0 1 60384
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_107_961
timestamp 1624015447
transform 1 0 89516 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_957
timestamp 1624015447
transform 1 0 89148 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_954
timestamp 1624015447
transform 1 0 88872 0 1 61472
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_109_961
timestamp 1624015447
transform 1 0 89516 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_901
timestamp 1624015447
transform -1 0 90896 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_903
timestamp 1624015447
transform -1 0 90896 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_905
timestamp 1624015447
transform -1 0 90896 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_907
timestamp 1624015447
transform -1 0 90896 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_106_969
timestamp 1624015447
transform 1 0 90252 0 -1 60384
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_969
timestamp 1624015447
transform 1 0 90252 0 -1 61472
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1624015447
transform 1 0 1104 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1624015447
transform 1 0 1104 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1624015447
transform 1 0 1104 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_110_3
timestamp 1624015447
transform 1 0 1380 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_15
timestamp 1624015447
transform 1 0 2484 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_3
timestamp 1624015447
transform 1 0 1380 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_15
timestamp 1624015447
transform 1 0 2484 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_3
timestamp 1624015447
transform 1 0 1380 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_15
timestamp 1624015447
transform 1 0 2484 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1430
timestamp 1624015447
transform 1 0 3772 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1431
timestamp 1624015447
transform 1 0 3772 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_110_27
timestamp 1624015447
transform 1 0 3588 0 -1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_110_30
timestamp 1624015447
transform 1 0 3864 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_111_27
timestamp 1624015447
transform 1 0 3588 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_112_27
timestamp 1624015447
transform 1 0 3588 0 -1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_112_30
timestamp 1624015447
transform 1 0 3864 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1624015447
transform -1 0 5152 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1624015447
transform -1 0 5152 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1624015447
transform -1 0 5152 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_110_38
timestamp 1624015447
transform 1 0 4600 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_111_39
timestamp 1624015447
transform 1 0 4692 0 1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_112_38
timestamp 1624015447
transform 1 0 4600 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_908
timestamp 1624015447
transform 1 0 84180 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_910
timestamp 1624015447
transform 1 0 84180 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_912
timestamp 1624015447
transform 1 0 84180 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_110_906
timestamp 1624015447
transform 1 0 84456 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_906
timestamp 1624015447
transform 1 0 84456 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_906
timestamp 1624015447
transform 1 0 84456 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_918
timestamp 1624015447
transform 1 0 85560 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_110_930
timestamp 1624015447
transform 1 0 86664 0 -1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_111_918
timestamp 1624015447
transform 1 0 85560 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_930
timestamp 1624015447
transform 1 0 86664 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_918
timestamp 1624015447
transform 1 0 85560 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_112_930
timestamp 1624015447
transform 1 0 86664 0 -1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1660
timestamp 1624015447
transform 1 0 86848 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1662
timestamp 1624015447
transform 1 0 86848 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_933
timestamp 1624015447
transform 1 0 86940 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_945
timestamp 1624015447
transform 1 0 88044 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_942
timestamp 1624015447
transform 1 0 87768 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_933
timestamp 1624015447
transform 1 0 86940 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_945
timestamp 1624015447
transform 1 0 88044 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1661
timestamp 1624015447
transform 1 0 89424 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_957
timestamp 1624015447
transform 1 0 89148 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_954
timestamp 1624015447
transform 1 0 88872 0 1 62560
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_111_961
timestamp 1624015447
transform 1 0 89516 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_957
timestamp 1624015447
transform 1 0 89148 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_909
timestamp 1624015447
transform -1 0 90896 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_911
timestamp 1624015447
transform -1 0 90896 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_913
timestamp 1624015447
transform -1 0 90896 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_110_969
timestamp 1624015447
transform 1 0 90252 0 -1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_112_969
timestamp 1624015447
transform 1 0 90252 0 -1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1624015447
transform 1 0 1104 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1624015447
transform 1 0 1104 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1624015447
transform 1 0 1104 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_113_3
timestamp 1624015447
transform 1 0 1380 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_15
timestamp 1624015447
transform 1 0 2484 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_3
timestamp 1624015447
transform 1 0 1380 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_15
timestamp 1624015447
transform 1 0 2484 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_3
timestamp 1624015447
transform 1 0 1380 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_15
timestamp 1624015447
transform 1 0 2484 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1432
timestamp 1624015447
transform 1 0 3772 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_27
timestamp 1624015447
transform 1 0 3588 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_114_27
timestamp 1624015447
transform 1 0 3588 0 -1 64736
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_114_30
timestamp 1624015447
transform 1 0 3864 0 -1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_115_27
timestamp 1624015447
transform 1 0 3588 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1624015447
transform -1 0 5152 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1624015447
transform -1 0 5152 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1624015447
transform -1 0 5152 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_113_39
timestamp 1624015447
transform 1 0 4692 0 1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_114_38
timestamp 1624015447
transform 1 0 4600 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_115_39
timestamp 1624015447
transform 1 0 4692 0 1 64736
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_914
timestamp 1624015447
transform 1 0 84180 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_916
timestamp 1624015447
transform 1 0 84180 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_918
timestamp 1624015447
transform 1 0 84180 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_113_906
timestamp 1624015447
transform 1 0 84456 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_906
timestamp 1624015447
transform 1 0 84456 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_906
timestamp 1624015447
transform 1 0 84456 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_918
timestamp 1624015447
transform 1 0 85560 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_930
timestamp 1624015447
transform 1 0 86664 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_918
timestamp 1624015447
transform 1 0 85560 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_114_930
timestamp 1624015447
transform 1 0 86664 0 -1 64736
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_115_918
timestamp 1624015447
transform 1 0 85560 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_930
timestamp 1624015447
transform 1 0 86664 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1664
timestamp 1624015447
transform 1 0 86848 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_942
timestamp 1624015447
transform 1 0 87768 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_933
timestamp 1624015447
transform 1 0 86940 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_945
timestamp 1624015447
transform 1 0 88044 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_942
timestamp 1624015447
transform 1 0 87768 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1663
timestamp 1624015447
transform 1 0 89424 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1665
timestamp 1624015447
transform 1 0 89424 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_113_954
timestamp 1624015447
transform 1 0 88872 0 1 63648
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_113_961
timestamp 1624015447
transform 1 0 89516 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_957
timestamp 1624015447
transform 1 0 89148 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_954
timestamp 1624015447
transform 1 0 88872 0 1 64736
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_115_961
timestamp 1624015447
transform 1 0 89516 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_915
timestamp 1624015447
transform -1 0 90896 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_917
timestamp 1624015447
transform -1 0 90896 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_919
timestamp 1624015447
transform -1 0 90896 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_114_969
timestamp 1624015447
transform 1 0 90252 0 -1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_230
timestamp 1624015447
transform 1 0 1104 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_232
timestamp 1624015447
transform 1 0 1104 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_234
timestamp 1624015447
transform 1 0 1104 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_116_3
timestamp 1624015447
transform 1 0 1380 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_15
timestamp 1624015447
transform 1 0 2484 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_3
timestamp 1624015447
transform 1 0 1380 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_15
timestamp 1624015447
transform 1 0 2484 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_3
timestamp 1624015447
transform 1 0 1380 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_15
timestamp 1624015447
transform 1 0 2484 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1433
timestamp 1624015447
transform 1 0 3772 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1434
timestamp 1624015447
transform 1 0 3772 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_116_27
timestamp 1624015447
transform 1 0 3588 0 -1 65824
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_116_30
timestamp 1624015447
transform 1 0 3864 0 -1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_117_27
timestamp 1624015447
transform 1 0 3588 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_118_27
timestamp 1624015447
transform 1 0 3588 0 -1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_118_30
timestamp 1624015447
transform 1 0 3864 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_231
timestamp 1624015447
transform -1 0 5152 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_233
timestamp 1624015447
transform -1 0 5152 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_235
timestamp 1624015447
transform -1 0 5152 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_116_38
timestamp 1624015447
transform 1 0 4600 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_117_39
timestamp 1624015447
transform 1 0 4692 0 1 65824
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_118_38
timestamp 1624015447
transform 1 0 4600 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_920
timestamp 1624015447
transform 1 0 84180 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_922
timestamp 1624015447
transform 1 0 84180 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_924
timestamp 1624015447
transform 1 0 84180 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_116_906
timestamp 1624015447
transform 1 0 84456 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_906
timestamp 1624015447
transform 1 0 84456 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_906
timestamp 1624015447
transform 1 0 84456 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_918
timestamp 1624015447
transform 1 0 85560 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_116_930
timestamp 1624015447
transform 1 0 86664 0 -1 65824
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_117_918
timestamp 1624015447
transform 1 0 85560 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_930
timestamp 1624015447
transform 1 0 86664 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_918
timestamp 1624015447
transform 1 0 85560 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_118_930
timestamp 1624015447
transform 1 0 86664 0 -1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1666
timestamp 1624015447
transform 1 0 86848 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1668
timestamp 1624015447
transform 1 0 86848 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_933
timestamp 1624015447
transform 1 0 86940 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_945
timestamp 1624015447
transform 1 0 88044 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_942
timestamp 1624015447
transform 1 0 87768 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_933
timestamp 1624015447
transform 1 0 86940 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_945
timestamp 1624015447
transform 1 0 88044 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1667
timestamp 1624015447
transform 1 0 89424 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_957
timestamp 1624015447
transform 1 0 89148 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_954
timestamp 1624015447
transform 1 0 88872 0 1 65824
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_117_961
timestamp 1624015447
transform 1 0 89516 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_957
timestamp 1624015447
transform 1 0 89148 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_921
timestamp 1624015447
transform -1 0 90896 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_923
timestamp 1624015447
transform -1 0 90896 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_925
timestamp 1624015447
transform -1 0 90896 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_116_969
timestamp 1624015447
transform 1 0 90252 0 -1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_118_969
timestamp 1624015447
transform 1 0 90252 0 -1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_236
timestamp 1624015447
transform 1 0 1104 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_238
timestamp 1624015447
transform 1 0 1104 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_240
timestamp 1624015447
transform 1 0 1104 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_119_3
timestamp 1624015447
transform 1 0 1380 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_15
timestamp 1624015447
transform 1 0 2484 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_3
timestamp 1624015447
transform 1 0 1380 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_15
timestamp 1624015447
transform 1 0 2484 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_3
timestamp 1624015447
transform 1 0 1380 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_15
timestamp 1624015447
transform 1 0 2484 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1435
timestamp 1624015447
transform 1 0 3772 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_27
timestamp 1624015447
transform 1 0 3588 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_120_27
timestamp 1624015447
transform 1 0 3588 0 -1 68000
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_120_30
timestamp 1624015447
transform 1 0 3864 0 -1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_121_27
timestamp 1624015447
transform 1 0 3588 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_237
timestamp 1624015447
transform -1 0 5152 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_239
timestamp 1624015447
transform -1 0 5152 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_241
timestamp 1624015447
transform -1 0 5152 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_119_39
timestamp 1624015447
transform 1 0 4692 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_120_38
timestamp 1624015447
transform 1 0 4600 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_121_39
timestamp 1624015447
transform 1 0 4692 0 1 68000
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_926
timestamp 1624015447
transform 1 0 84180 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_928
timestamp 1624015447
transform 1 0 84180 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_930
timestamp 1624015447
transform 1 0 84180 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_119_906
timestamp 1624015447
transform 1 0 84456 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_906
timestamp 1624015447
transform 1 0 84456 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_906
timestamp 1624015447
transform 1 0 84456 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_918
timestamp 1624015447
transform 1 0 85560 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_930
timestamp 1624015447
transform 1 0 86664 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_918
timestamp 1624015447
transform 1 0 85560 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_120_930
timestamp 1624015447
transform 1 0 86664 0 -1 68000
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_121_918
timestamp 1624015447
transform 1 0 85560 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_930
timestamp 1624015447
transform 1 0 86664 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1670
timestamp 1624015447
transform 1 0 86848 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_942
timestamp 1624015447
transform 1 0 87768 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_933
timestamp 1624015447
transform 1 0 86940 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_945
timestamp 1624015447
transform 1 0 88044 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_942
timestamp 1624015447
transform 1 0 87768 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1669
timestamp 1624015447
transform 1 0 89424 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1671
timestamp 1624015447
transform 1 0 89424 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_119_954
timestamp 1624015447
transform 1 0 88872 0 1 66912
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_119_961
timestamp 1624015447
transform 1 0 89516 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_957
timestamp 1624015447
transform 1 0 89148 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_954
timestamp 1624015447
transform 1 0 88872 0 1 68000
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_121_961
timestamp 1624015447
transform 1 0 89516 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_927
timestamp 1624015447
transform -1 0 90896 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_929
timestamp 1624015447
transform -1 0 90896 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_931
timestamp 1624015447
transform -1 0 90896 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_120_969
timestamp 1624015447
transform 1 0 90252 0 -1 68000
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_242
timestamp 1624015447
transform 1 0 1104 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_244
timestamp 1624015447
transform 1 0 1104 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_246
timestamp 1624015447
transform 1 0 1104 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_122_3
timestamp 1624015447
transform 1 0 1380 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_15
timestamp 1624015447
transform 1 0 2484 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_3
timestamp 1624015447
transform 1 0 1380 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_15
timestamp 1624015447
transform 1 0 2484 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_3
timestamp 1624015447
transform 1 0 1380 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_15
timestamp 1624015447
transform 1 0 2484 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1436
timestamp 1624015447
transform 1 0 3772 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1437
timestamp 1624015447
transform 1 0 3772 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_122_27
timestamp 1624015447
transform 1 0 3588 0 -1 69088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_122_30
timestamp 1624015447
transform 1 0 3864 0 -1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_123_27
timestamp 1624015447
transform 1 0 3588 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_124_27
timestamp 1624015447
transform 1 0 3588 0 -1 70176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_124_30
timestamp 1624015447
transform 1 0 3864 0 -1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_243
timestamp 1624015447
transform -1 0 5152 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_245
timestamp 1624015447
transform -1 0 5152 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_247
timestamp 1624015447
transform -1 0 5152 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_122_38
timestamp 1624015447
transform 1 0 4600 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_123_39
timestamp 1624015447
transform 1 0 4692 0 1 69088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_124_38
timestamp 1624015447
transform 1 0 4600 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_932
timestamp 1624015447
transform 1 0 84180 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_934
timestamp 1624015447
transform 1 0 84180 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_936
timestamp 1624015447
transform 1 0 84180 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_122_906
timestamp 1624015447
transform 1 0 84456 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_906
timestamp 1624015447
transform 1 0 84456 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_906
timestamp 1624015447
transform 1 0 84456 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_918
timestamp 1624015447
transform 1 0 85560 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_122_930
timestamp 1624015447
transform 1 0 86664 0 -1 69088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_123_918
timestamp 1624015447
transform 1 0 85560 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_930
timestamp 1624015447
transform 1 0 86664 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_918
timestamp 1624015447
transform 1 0 85560 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_124_930
timestamp 1624015447
transform 1 0 86664 0 -1 70176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1672
timestamp 1624015447
transform 1 0 86848 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1674
timestamp 1624015447
transform 1 0 86848 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_933
timestamp 1624015447
transform 1 0 86940 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_945
timestamp 1624015447
transform 1 0 88044 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_942
timestamp 1624015447
transform 1 0 87768 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_933
timestamp 1624015447
transform 1 0 86940 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_945
timestamp 1624015447
transform 1 0 88044 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1673
timestamp 1624015447
transform 1 0 89424 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_957
timestamp 1624015447
transform 1 0 89148 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_954
timestamp 1624015447
transform 1 0 88872 0 1 69088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_123_961
timestamp 1624015447
transform 1 0 89516 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_957
timestamp 1624015447
transform 1 0 89148 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_933
timestamp 1624015447
transform -1 0 90896 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_935
timestamp 1624015447
transform -1 0 90896 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_937
timestamp 1624015447
transform -1 0 90896 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_122_969
timestamp 1624015447
transform 1 0 90252 0 -1 69088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_124_969
timestamp 1624015447
transform 1 0 90252 0 -1 70176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_248
timestamp 1624015447
transform 1 0 1104 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_250
timestamp 1624015447
transform 1 0 1104 0 -1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_252
timestamp 1624015447
transform 1 0 1104 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_125_3
timestamp 1624015447
transform 1 0 1380 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_15
timestamp 1624015447
transform 1 0 2484 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_3
timestamp 1624015447
transform 1 0 1380 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_15
timestamp 1624015447
transform 1 0 2484 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_3
timestamp 1624015447
transform 1 0 1380 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_15
timestamp 1624015447
transform 1 0 2484 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1438
timestamp 1624015447
transform 1 0 3772 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_27
timestamp 1624015447
transform 1 0 3588 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_126_27
timestamp 1624015447
transform 1 0 3588 0 -1 71264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_126_30
timestamp 1624015447
transform 1 0 3864 0 -1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_127_27
timestamp 1624015447
transform 1 0 3588 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_249
timestamp 1624015447
transform -1 0 5152 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_251
timestamp 1624015447
transform -1 0 5152 0 -1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_253
timestamp 1624015447
transform -1 0 5152 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_125_39
timestamp 1624015447
transform 1 0 4692 0 1 70176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_126_38
timestamp 1624015447
transform 1 0 4600 0 -1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_127_39
timestamp 1624015447
transform 1 0 4692 0 1 71264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_938
timestamp 1624015447
transform 1 0 84180 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_940
timestamp 1624015447
transform 1 0 84180 0 -1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_942
timestamp 1624015447
transform 1 0 84180 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_125_906
timestamp 1624015447
transform 1 0 84456 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_906
timestamp 1624015447
transform 1 0 84456 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_906
timestamp 1624015447
transform 1 0 84456 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_918
timestamp 1624015447
transform 1 0 85560 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_930
timestamp 1624015447
transform 1 0 86664 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_918
timestamp 1624015447
transform 1 0 85560 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_126_930
timestamp 1624015447
transform 1 0 86664 0 -1 71264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_127_918
timestamp 1624015447
transform 1 0 85560 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_930
timestamp 1624015447
transform 1 0 86664 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1676
timestamp 1624015447
transform 1 0 86848 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_942
timestamp 1624015447
transform 1 0 87768 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_933
timestamp 1624015447
transform 1 0 86940 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_945
timestamp 1624015447
transform 1 0 88044 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_942
timestamp 1624015447
transform 1 0 87768 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1675
timestamp 1624015447
transform 1 0 89424 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1677
timestamp 1624015447
transform 1 0 89424 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_125_954
timestamp 1624015447
transform 1 0 88872 0 1 70176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_125_961
timestamp 1624015447
transform 1 0 89516 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_957
timestamp 1624015447
transform 1 0 89148 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_954
timestamp 1624015447
transform 1 0 88872 0 1 71264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_127_961
timestamp 1624015447
transform 1 0 89516 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_939
timestamp 1624015447
transform -1 0 90896 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_941
timestamp 1624015447
transform -1 0 90896 0 -1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_943
timestamp 1624015447
transform -1 0 90896 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_126_969
timestamp 1624015447
transform 1 0 90252 0 -1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_129_15
timestamp 1624015447
transform 1 0 2484 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_3
timestamp 1624015447
transform 1 0 1380 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_15
timestamp 1624015447
transform 1 0 2484 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_3
timestamp 1624015447
transform 1 0 1380 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_256
timestamp 1624015447
transform 1 0 1104 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_254
timestamp 1624015447
transform 1 0 1104 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_130_15
timestamp 1624015447
transform 1 0 2484 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_3
timestamp 1624015447
transform 1 0 1380 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_258
timestamp 1624015447
transform 1 0 1104 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_131_15
timestamp 1624015447
transform 1 0 2484 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_3
timestamp 1624015447
transform 1 0 1380 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_260
timestamp 1624015447
transform 1 0 1104 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1439
timestamp 1624015447
transform 1 0 3772 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1440
timestamp 1624015447
transform 1 0 3772 0 -1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_128_27
timestamp 1624015447
transform 1 0 3588 0 -1 72352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_128_30
timestamp 1624015447
transform 1 0 3864 0 -1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_129_27
timestamp 1624015447
transform 1 0 3588 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_130_27
timestamp 1624015447
transform 1 0 3588 0 -1 73440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_130_30
timestamp 1624015447
transform 1 0 3864 0 -1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_131_27
timestamp 1624015447
transform 1 0 3588 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_255
timestamp 1624015447
transform -1 0 5152 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_257
timestamp 1624015447
transform -1 0 5152 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_259
timestamp 1624015447
transform -1 0 5152 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_261
timestamp 1624015447
transform -1 0 5152 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_128_38
timestamp 1624015447
transform 1 0 4600 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_129_39
timestamp 1624015447
transform 1 0 4692 0 1 72352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_130_38
timestamp 1624015447
transform 1 0 4600 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_131_39
timestamp 1624015447
transform 1 0 4692 0 1 73440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_944
timestamp 1624015447
transform 1 0 84180 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_946
timestamp 1624015447
transform 1 0 84180 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_948
timestamp 1624015447
transform 1 0 84180 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_950
timestamp 1624015447
transform 1 0 84180 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_128_906
timestamp 1624015447
transform 1 0 84456 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_906
timestamp 1624015447
transform 1 0 84456 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_906
timestamp 1624015447
transform 1 0 84456 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_906
timestamp 1624015447
transform 1 0 84456 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_918
timestamp 1624015447
transform 1 0 85560 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_128_930
timestamp 1624015447
transform 1 0 86664 0 -1 72352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_129_918
timestamp 1624015447
transform 1 0 85560 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_930
timestamp 1624015447
transform 1 0 86664 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_918
timestamp 1624015447
transform 1 0 85560 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_130_930
timestamp 1624015447
transform 1 0 86664 0 -1 73440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_131_918
timestamp 1624015447
transform 1 0 85560 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_930
timestamp 1624015447
transform 1 0 86664 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1678
timestamp 1624015447
transform 1 0 86848 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1680
timestamp 1624015447
transform 1 0 86848 0 -1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_933
timestamp 1624015447
transform 1 0 86940 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_945
timestamp 1624015447
transform 1 0 88044 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_942
timestamp 1624015447
transform 1 0 87768 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_933
timestamp 1624015447
transform 1 0 86940 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_945
timestamp 1624015447
transform 1 0 88044 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_942
timestamp 1624015447
transform 1 0 87768 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1679
timestamp 1624015447
transform 1 0 89424 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1681
timestamp 1624015447
transform 1 0 89424 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_957
timestamp 1624015447
transform 1 0 89148 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_954
timestamp 1624015447
transform 1 0 88872 0 1 72352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_129_961
timestamp 1624015447
transform 1 0 89516 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_957
timestamp 1624015447
transform 1 0 89148 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_954
timestamp 1624015447
transform 1 0 88872 0 1 73440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_131_961
timestamp 1624015447
transform 1 0 89516 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_945
timestamp 1624015447
transform -1 0 90896 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_947
timestamp 1624015447
transform -1 0 90896 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_949
timestamp 1624015447
transform -1 0 90896 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_951
timestamp 1624015447
transform -1 0 90896 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_128_969
timestamp 1624015447
transform 1 0 90252 0 -1 72352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_130_969
timestamp 1624015447
transform 1 0 90252 0 -1 73440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_262
timestamp 1624015447
transform 1 0 1104 0 -1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_264
timestamp 1624015447
transform 1 0 1104 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_266
timestamp 1624015447
transform 1 0 1104 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_132_3
timestamp 1624015447
transform 1 0 1380 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_15
timestamp 1624015447
transform 1 0 2484 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_3
timestamp 1624015447
transform 1 0 1380 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_15
timestamp 1624015447
transform 1 0 2484 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_3
timestamp 1624015447
transform 1 0 1380 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_15
timestamp 1624015447
transform 1 0 2484 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1441
timestamp 1624015447
transform 1 0 3772 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1442
timestamp 1624015447
transform 1 0 3772 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_132_27
timestamp 1624015447
transform 1 0 3588 0 -1 74528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_132_30
timestamp 1624015447
transform 1 0 3864 0 -1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_133_27
timestamp 1624015447
transform 1 0 3588 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_134_27
timestamp 1624015447
transform 1 0 3588 0 -1 75616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_134_30
timestamp 1624015447
transform 1 0 3864 0 -1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_263
timestamp 1624015447
transform -1 0 5152 0 -1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_265
timestamp 1624015447
transform -1 0 5152 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_267
timestamp 1624015447
transform -1 0 5152 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_132_38
timestamp 1624015447
transform 1 0 4600 0 -1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_133_39
timestamp 1624015447
transform 1 0 4692 0 1 74528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_134_38
timestamp 1624015447
transform 1 0 4600 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_952
timestamp 1624015447
transform 1 0 84180 0 -1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_954
timestamp 1624015447
transform 1 0 84180 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_956
timestamp 1624015447
transform 1 0 84180 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_132_906
timestamp 1624015447
transform 1 0 84456 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_906
timestamp 1624015447
transform 1 0 84456 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_906
timestamp 1624015447
transform 1 0 84456 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_918
timestamp 1624015447
transform 1 0 85560 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_132_930
timestamp 1624015447
transform 1 0 86664 0 -1 74528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_133_918
timestamp 1624015447
transform 1 0 85560 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_930
timestamp 1624015447
transform 1 0 86664 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_918
timestamp 1624015447
transform 1 0 85560 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_134_930
timestamp 1624015447
transform 1 0 86664 0 -1 75616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1682
timestamp 1624015447
transform 1 0 86848 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1684
timestamp 1624015447
transform 1 0 86848 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_933
timestamp 1624015447
transform 1 0 86940 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_945
timestamp 1624015447
transform 1 0 88044 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_942
timestamp 1624015447
transform 1 0 87768 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_933
timestamp 1624015447
transform 1 0 86940 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_945
timestamp 1624015447
transform 1 0 88044 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1683
timestamp 1624015447
transform 1 0 89424 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_957
timestamp 1624015447
transform 1 0 89148 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_954
timestamp 1624015447
transform 1 0 88872 0 1 74528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_133_961
timestamp 1624015447
transform 1 0 89516 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_957
timestamp 1624015447
transform 1 0 89148 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_953
timestamp 1624015447
transform -1 0 90896 0 -1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_955
timestamp 1624015447
transform -1 0 90896 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_957
timestamp 1624015447
transform -1 0 90896 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_132_969
timestamp 1624015447
transform 1 0 90252 0 -1 74528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_134_969
timestamp 1624015447
transform 1 0 90252 0 -1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_268
timestamp 1624015447
transform 1 0 1104 0 1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_270
timestamp 1624015447
transform 1 0 1104 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_272
timestamp 1624015447
transform 1 0 1104 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_135_3
timestamp 1624015447
transform 1 0 1380 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_15
timestamp 1624015447
transform 1 0 2484 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_3
timestamp 1624015447
transform 1 0 1380 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_15
timestamp 1624015447
transform 1 0 2484 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_3
timestamp 1624015447
transform 1 0 1380 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_15
timestamp 1624015447
transform 1 0 2484 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1443
timestamp 1624015447
transform 1 0 3772 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_27
timestamp 1624015447
transform 1 0 3588 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_136_27
timestamp 1624015447
transform 1 0 3588 0 -1 76704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_136_30
timestamp 1624015447
transform 1 0 3864 0 -1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_137_27
timestamp 1624015447
transform 1 0 3588 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_269
timestamp 1624015447
transform -1 0 5152 0 1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_271
timestamp 1624015447
transform -1 0 5152 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_273
timestamp 1624015447
transform -1 0 5152 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_135_39
timestamp 1624015447
transform 1 0 4692 0 1 75616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_136_38
timestamp 1624015447
transform 1 0 4600 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_137_39
timestamp 1624015447
transform 1 0 4692 0 1 76704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_958
timestamp 1624015447
transform 1 0 84180 0 1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_960
timestamp 1624015447
transform 1 0 84180 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_962
timestamp 1624015447
transform 1 0 84180 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_135_906
timestamp 1624015447
transform 1 0 84456 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_906
timestamp 1624015447
transform 1 0 84456 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_906
timestamp 1624015447
transform 1 0 84456 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_918
timestamp 1624015447
transform 1 0 85560 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_930
timestamp 1624015447
transform 1 0 86664 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_918
timestamp 1624015447
transform 1 0 85560 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_136_930
timestamp 1624015447
transform 1 0 86664 0 -1 76704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_137_918
timestamp 1624015447
transform 1 0 85560 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_930
timestamp 1624015447
transform 1 0 86664 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1686
timestamp 1624015447
transform 1 0 86848 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_942
timestamp 1624015447
transform 1 0 87768 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_933
timestamp 1624015447
transform 1 0 86940 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_945
timestamp 1624015447
transform 1 0 88044 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_942
timestamp 1624015447
transform 1 0 87768 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1685
timestamp 1624015447
transform 1 0 89424 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1687
timestamp 1624015447
transform 1 0 89424 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_135_954
timestamp 1624015447
transform 1 0 88872 0 1 75616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_135_961
timestamp 1624015447
transform 1 0 89516 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_957
timestamp 1624015447
transform 1 0 89148 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_954
timestamp 1624015447
transform 1 0 88872 0 1 76704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_137_961
timestamp 1624015447
transform 1 0 89516 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_959
timestamp 1624015447
transform -1 0 90896 0 1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_961
timestamp 1624015447
transform -1 0 90896 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_963
timestamp 1624015447
transform -1 0 90896 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_136_969
timestamp 1624015447
transform 1 0 90252 0 -1 76704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_274
timestamp 1624015447
transform 1 0 1104 0 -1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_276
timestamp 1624015447
transform 1 0 1104 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_278
timestamp 1624015447
transform 1 0 1104 0 -1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_138_3
timestamp 1624015447
transform 1 0 1380 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_15
timestamp 1624015447
transform 1 0 2484 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_3
timestamp 1624015447
transform 1 0 1380 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_15
timestamp 1624015447
transform 1 0 2484 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_3
timestamp 1624015447
transform 1 0 1380 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_15
timestamp 1624015447
transform 1 0 2484 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1444
timestamp 1624015447
transform 1 0 3772 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1445
timestamp 1624015447
transform 1 0 3772 0 -1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_138_27
timestamp 1624015447
transform 1 0 3588 0 -1 77792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_138_30
timestamp 1624015447
transform 1 0 3864 0 -1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_139_27
timestamp 1624015447
transform 1 0 3588 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_140_27
timestamp 1624015447
transform 1 0 3588 0 -1 78880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_140_30
timestamp 1624015447
transform 1 0 3864 0 -1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_275
timestamp 1624015447
transform -1 0 5152 0 -1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_277
timestamp 1624015447
transform -1 0 5152 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_279
timestamp 1624015447
transform -1 0 5152 0 -1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_138_38
timestamp 1624015447
transform 1 0 4600 0 -1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_139_39
timestamp 1624015447
transform 1 0 4692 0 1 77792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_140_38
timestamp 1624015447
transform 1 0 4600 0 -1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_964
timestamp 1624015447
transform 1 0 84180 0 -1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_966
timestamp 1624015447
transform 1 0 84180 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_968
timestamp 1624015447
transform 1 0 84180 0 -1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_138_906
timestamp 1624015447
transform 1 0 84456 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_906
timestamp 1624015447
transform 1 0 84456 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_906
timestamp 1624015447
transform 1 0 84456 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_918
timestamp 1624015447
transform 1 0 85560 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_138_930
timestamp 1624015447
transform 1 0 86664 0 -1 77792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_139_918
timestamp 1624015447
transform 1 0 85560 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_930
timestamp 1624015447
transform 1 0 86664 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_918
timestamp 1624015447
transform 1 0 85560 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_140_930
timestamp 1624015447
transform 1 0 86664 0 -1 78880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1688
timestamp 1624015447
transform 1 0 86848 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1690
timestamp 1624015447
transform 1 0 86848 0 -1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_933
timestamp 1624015447
transform 1 0 86940 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_945
timestamp 1624015447
transform 1 0 88044 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_942
timestamp 1624015447
transform 1 0 87768 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_933
timestamp 1624015447
transform 1 0 86940 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_945
timestamp 1624015447
transform 1 0 88044 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1689
timestamp 1624015447
transform 1 0 89424 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_957
timestamp 1624015447
transform 1 0 89148 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_954
timestamp 1624015447
transform 1 0 88872 0 1 77792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_139_961
timestamp 1624015447
transform 1 0 89516 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_957
timestamp 1624015447
transform 1 0 89148 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_965
timestamp 1624015447
transform -1 0 90896 0 -1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_967
timestamp 1624015447
transform -1 0 90896 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_969
timestamp 1624015447
transform -1 0 90896 0 -1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_138_969
timestamp 1624015447
transform 1 0 90252 0 -1 77792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_140_969
timestamp 1624015447
transform 1 0 90252 0 -1 78880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_280
timestamp 1624015447
transform 1 0 1104 0 1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_282
timestamp 1624015447
transform 1 0 1104 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_284
timestamp 1624015447
transform 1 0 1104 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_141_3
timestamp 1624015447
transform 1 0 1380 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_15
timestamp 1624015447
transform 1 0 2484 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_3
timestamp 1624015447
transform 1 0 1380 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_15
timestamp 1624015447
transform 1 0 2484 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_3
timestamp 1624015447
transform 1 0 1380 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_15
timestamp 1624015447
transform 1 0 2484 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1446
timestamp 1624015447
transform 1 0 3772 0 -1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_141_27
timestamp 1624015447
transform 1 0 3588 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_142_27
timestamp 1624015447
transform 1 0 3588 0 -1 79968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_142_30
timestamp 1624015447
transform 1 0 3864 0 -1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_143_27
timestamp 1624015447
transform 1 0 3588 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_281
timestamp 1624015447
transform -1 0 5152 0 1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_283
timestamp 1624015447
transform -1 0 5152 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_285
timestamp 1624015447
transform -1 0 5152 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr0[1]
timestamp 1624015447
transform -1 0 4876 0 1 79968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_141_39
timestamp 1624015447
transform 1 0 4692 0 1 78880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_142_38
timestamp 1624015447
transform 1 0 4600 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_970
timestamp 1624015447
transform 1 0 84180 0 1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_972
timestamp 1624015447
transform 1 0 84180 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_974
timestamp 1624015447
transform 1 0 84180 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_141_906
timestamp 1624015447
transform 1 0 84456 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_906
timestamp 1624015447
transform 1 0 84456 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_906
timestamp 1624015447
transform 1 0 84456 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_918
timestamp 1624015447
transform 1 0 85560 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_930
timestamp 1624015447
transform 1 0 86664 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_918
timestamp 1624015447
transform 1 0 85560 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_142_930
timestamp 1624015447
transform 1 0 86664 0 -1 79968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_143_918
timestamp 1624015447
transform 1 0 85560 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_930
timestamp 1624015447
transform 1 0 86664 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1692
timestamp 1624015447
transform 1 0 86848 0 -1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_141_942
timestamp 1624015447
transform 1 0 87768 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_933
timestamp 1624015447
transform 1 0 86940 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_945
timestamp 1624015447
transform 1 0 88044 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_942
timestamp 1624015447
transform 1 0 87768 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1691
timestamp 1624015447
transform 1 0 89424 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1693
timestamp 1624015447
transform 1 0 89424 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_141_954
timestamp 1624015447
transform 1 0 88872 0 1 78880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_141_961
timestamp 1624015447
transform 1 0 89516 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_957
timestamp 1624015447
transform 1 0 89148 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_954
timestamp 1624015447
transform 1 0 88872 0 1 79968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_143_961
timestamp 1624015447
transform 1 0 89516 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_971
timestamp 1624015447
transform -1 0 90896 0 1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_973
timestamp 1624015447
transform -1 0 90896 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_975
timestamp 1624015447
transform -1 0 90896 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_142_969
timestamp 1624015447
transform 1 0 90252 0 -1 79968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_286
timestamp 1624015447
transform 1 0 1104 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_288
timestamp 1624015447
transform 1 0 1104 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_290
timestamp 1624015447
transform 1 0 1104 0 -1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_144_3
timestamp 1624015447
transform 1 0 1380 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_15
timestamp 1624015447
transform 1 0 2484 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_3
timestamp 1624015447
transform 1 0 1380 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_15
timestamp 1624015447
transform 1 0 2484 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_3
timestamp 1624015447
transform 1 0 1380 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_15
timestamp 1624015447
transform 1 0 2484 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1447
timestamp 1624015447
transform 1 0 3772 0 -1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1448
timestamp 1624015447
transform 1 0 3772 0 -1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_144_27
timestamp 1624015447
transform 1 0 3588 0 -1 81056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_144_30
timestamp 1624015447
transform 1 0 3864 0 -1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_145_27
timestamp 1624015447
transform 1 0 3588 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_146_27
timestamp 1624015447
transform 1 0 3588 0 -1 82144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_146_30
timestamp 1624015447
transform 1 0 3864 0 -1 82144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_287
timestamp 1624015447
transform -1 0 5152 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_289
timestamp 1624015447
transform -1 0 5152 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_291
timestamp 1624015447
transform -1 0 5152 0 -1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_144_38
timestamp 1624015447
transform 1 0 4600 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_145_39
timestamp 1624015447
transform 1 0 4692 0 1 81056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_146_38
timestamp 1624015447
transform 1 0 4600 0 -1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_976
timestamp 1624015447
transform 1 0 84180 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_978
timestamp 1624015447
transform 1 0 84180 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_980
timestamp 1624015447
transform 1 0 84180 0 -1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_144_906
timestamp 1624015447
transform 1 0 84456 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_906
timestamp 1624015447
transform 1 0 84456 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_906
timestamp 1624015447
transform 1 0 84456 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_918
timestamp 1624015447
transform 1 0 85560 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_144_930
timestamp 1624015447
transform 1 0 86664 0 -1 81056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_145_918
timestamp 1624015447
transform 1 0 85560 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_930
timestamp 1624015447
transform 1 0 86664 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_918
timestamp 1624015447
transform 1 0 85560 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_146_930
timestamp 1624015447
transform 1 0 86664 0 -1 82144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1694
timestamp 1624015447
transform 1 0 86848 0 -1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1696
timestamp 1624015447
transform 1 0 86848 0 -1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_144_933
timestamp 1624015447
transform 1 0 86940 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_945
timestamp 1624015447
transform 1 0 88044 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_942
timestamp 1624015447
transform 1 0 87768 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_933
timestamp 1624015447
transform 1 0 86940 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_945
timestamp 1624015447
transform 1 0 88044 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1695
timestamp 1624015447
transform 1 0 89424 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_144_957
timestamp 1624015447
transform 1 0 89148 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_954
timestamp 1624015447
transform 1 0 88872 0 1 81056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_145_961
timestamp 1624015447
transform 1 0 89516 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_957
timestamp 1624015447
transform 1 0 89148 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_977
timestamp 1624015447
transform -1 0 90896 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_979
timestamp 1624015447
transform -1 0 90896 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_981
timestamp 1624015447
transform -1 0 90896 0 -1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_144_969
timestamp 1624015447
transform 1 0 90252 0 -1 81056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_146_969
timestamp 1624015447
transform 1 0 90252 0 -1 82144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_292
timestamp 1624015447
transform 1 0 1104 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_294
timestamp 1624015447
transform 1 0 1104 0 -1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_296
timestamp 1624015447
transform 1 0 1104 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_147_3
timestamp 1624015447
transform 1 0 1380 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_15
timestamp 1624015447
transform 1 0 2484 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_3
timestamp 1624015447
transform 1 0 1380 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_15
timestamp 1624015447
transform 1 0 2484 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_3
timestamp 1624015447
transform 1 0 1380 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_15
timestamp 1624015447
transform 1 0 2484 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1449
timestamp 1624015447
transform 1 0 3772 0 -1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_147_27
timestamp 1624015447
transform 1 0 3588 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_148_27
timestamp 1624015447
transform 1 0 3588 0 -1 83232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_148_30
timestamp 1624015447
transform 1 0 3864 0 -1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_149_27
timestamp 1624015447
transform 1 0 3588 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_293
timestamp 1624015447
transform -1 0 5152 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_295
timestamp 1624015447
transform -1 0 5152 0 -1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_297
timestamp 1624015447
transform -1 0 5152 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr0[2]
timestamp 1624015447
transform -1 0 4876 0 1 82144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr0[3]
timestamp 1624015447
transform -1 0 4876 0 1 83232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_148_38
timestamp 1624015447
transform 1 0 4600 0 -1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_982
timestamp 1624015447
transform 1 0 84180 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_984
timestamp 1624015447
transform 1 0 84180 0 -1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_986
timestamp 1624015447
transform 1 0 84180 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_147_906
timestamp 1624015447
transform 1 0 84456 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_906
timestamp 1624015447
transform 1 0 84456 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_906
timestamp 1624015447
transform 1 0 84456 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_918
timestamp 1624015447
transform 1 0 85560 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_930
timestamp 1624015447
transform 1 0 86664 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_918
timestamp 1624015447
transform 1 0 85560 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_148_930
timestamp 1624015447
transform 1 0 86664 0 -1 83232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_149_918
timestamp 1624015447
transform 1 0 85560 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_930
timestamp 1624015447
transform 1 0 86664 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1698
timestamp 1624015447
transform 1 0 86848 0 -1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_147_942
timestamp 1624015447
transform 1 0 87768 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_933
timestamp 1624015447
transform 1 0 86940 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_945
timestamp 1624015447
transform 1 0 88044 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_942
timestamp 1624015447
transform 1 0 87768 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1697
timestamp 1624015447
transform 1 0 89424 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1699
timestamp 1624015447
transform 1 0 89424 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_147_954
timestamp 1624015447
transform 1 0 88872 0 1 82144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_147_961
timestamp 1624015447
transform 1 0 89516 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_957
timestamp 1624015447
transform 1 0 89148 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_954
timestamp 1624015447
transform 1 0 88872 0 1 83232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_149_961
timestamp 1624015447
transform 1 0 89516 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_983
timestamp 1624015447
transform -1 0 90896 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_985
timestamp 1624015447
transform -1 0 90896 0 -1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_987
timestamp 1624015447
transform -1 0 90896 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_148_969
timestamp 1624015447
transform 1 0 90252 0 -1 83232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_151_15
timestamp 1624015447
transform 1 0 2484 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_3
timestamp 1624015447
transform 1 0 1380 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_15
timestamp 1624015447
transform 1 0 2484 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_3
timestamp 1624015447
transform 1 0 1380 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_300
timestamp 1624015447
transform 1 0 1104 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_298
timestamp 1624015447
transform 1 0 1104 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_152_15
timestamp 1624015447
transform 1 0 2484 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_3
timestamp 1624015447
transform 1 0 1380 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_302
timestamp 1624015447
transform 1 0 1104 0 -1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_153_15
timestamp 1624015447
transform 1 0 2484 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_3
timestamp 1624015447
transform 1 0 1380 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_304
timestamp 1624015447
transform 1 0 1104 0 1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1450
timestamp 1624015447
transform 1 0 3772 0 -1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1451
timestamp 1624015447
transform 1 0 3772 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_150_27
timestamp 1624015447
transform 1 0 3588 0 -1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_150_30
timestamp 1624015447
transform 1 0 3864 0 -1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_151_27
timestamp 1624015447
transform 1 0 3588 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_152_27
timestamp 1624015447
transform 1 0 3588 0 -1 85408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_152_30
timestamp 1624015447
transform 1 0 3864 0 -1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_153_27
timestamp 1624015447
transform 1 0 3588 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_299
timestamp 1624015447
transform -1 0 5152 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_301
timestamp 1624015447
transform -1 0 5152 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_303
timestamp 1624015447
transform -1 0 5152 0 -1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_305
timestamp 1624015447
transform -1 0 5152 0 1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr0[4]
timestamp 1624015447
transform -1 0 4876 0 -1 85408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_150_38
timestamp 1624015447
transform 1 0 4600 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_151_39
timestamp 1624015447
transform 1 0 4692 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_152_38
timestamp 1624015447
transform 1 0 4600 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_153_39
timestamp 1624015447
transform 1 0 4692 0 1 85408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_988
timestamp 1624015447
transform 1 0 84180 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_990
timestamp 1624015447
transform 1 0 84180 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_992
timestamp 1624015447
transform 1 0 84180 0 -1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_994
timestamp 1624015447
transform 1 0 84180 0 1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_150_906
timestamp 1624015447
transform 1 0 84456 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_906
timestamp 1624015447
transform 1 0 84456 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_906
timestamp 1624015447
transform 1 0 84456 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_906
timestamp 1624015447
transform 1 0 84456 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_918
timestamp 1624015447
transform 1 0 85560 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_150_930
timestamp 1624015447
transform 1 0 86664 0 -1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_151_918
timestamp 1624015447
transform 1 0 85560 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_930
timestamp 1624015447
transform 1 0 86664 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_918
timestamp 1624015447
transform 1 0 85560 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_152_930
timestamp 1624015447
transform 1 0 86664 0 -1 85408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_153_918
timestamp 1624015447
transform 1 0 85560 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_930
timestamp 1624015447
transform 1 0 86664 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1700
timestamp 1624015447
transform 1 0 86848 0 -1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1702
timestamp 1624015447
transform 1 0 86848 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_150_933
timestamp 1624015447
transform 1 0 86940 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_945
timestamp 1624015447
transform 1 0 88044 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_942
timestamp 1624015447
transform 1 0 87768 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_933
timestamp 1624015447
transform 1 0 86940 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_945
timestamp 1624015447
transform 1 0 88044 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_942
timestamp 1624015447
transform 1 0 87768 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1701
timestamp 1624015447
transform 1 0 89424 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1703
timestamp 1624015447
transform 1 0 89424 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_150_957
timestamp 1624015447
transform 1 0 89148 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_954
timestamp 1624015447
transform 1 0 88872 0 1 84320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_151_961
timestamp 1624015447
transform 1 0 89516 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_957
timestamp 1624015447
transform 1 0 89148 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_954
timestamp 1624015447
transform 1 0 88872 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_153_961
timestamp 1624015447
transform 1 0 89516 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_989
timestamp 1624015447
transform -1 0 90896 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_991
timestamp 1624015447
transform -1 0 90896 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_993
timestamp 1624015447
transform -1 0 90896 0 -1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_995
timestamp 1624015447
transform -1 0 90896 0 1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_150_969
timestamp 1624015447
transform 1 0 90252 0 -1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_152_969
timestamp 1624015447
transform 1 0 90252 0 -1 85408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_306
timestamp 1624015447
transform 1 0 1104 0 -1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_308
timestamp 1624015447
transform 1 0 1104 0 1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_310
timestamp 1624015447
transform 1 0 1104 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_154_3
timestamp 1624015447
transform 1 0 1380 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_15
timestamp 1624015447
transform 1 0 2484 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_3
timestamp 1624015447
transform 1 0 1380 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_15
timestamp 1624015447
transform 1 0 2484 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_3
timestamp 1624015447
transform 1 0 1380 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_15
timestamp 1624015447
transform 1 0 2484 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1452
timestamp 1624015447
transform 1 0 3772 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1453
timestamp 1624015447
transform 1 0 3772 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_154_27
timestamp 1624015447
transform 1 0 3588 0 -1 86496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_154_30
timestamp 1624015447
transform 1 0 3864 0 -1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_155_27
timestamp 1624015447
transform 1 0 3588 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_156_27
timestamp 1624015447
transform 1 0 3588 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_156_30
timestamp 1624015447
transform 1 0 3864 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_307
timestamp 1624015447
transform -1 0 5152 0 -1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_309
timestamp 1624015447
transform -1 0 5152 0 1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_311
timestamp 1624015447
transform -1 0 5152 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr0[5]
timestamp 1624015447
transform -1 0 4876 0 -1 86496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_154_38
timestamp 1624015447
transform 1 0 4600 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_155_39
timestamp 1624015447
transform 1 0 4692 0 1 86496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_156_38
timestamp 1624015447
transform 1 0 4600 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_996
timestamp 1624015447
transform 1 0 84180 0 -1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_998
timestamp 1624015447
transform 1 0 84180 0 1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1000
timestamp 1624015447
transform 1 0 84180 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_154_906
timestamp 1624015447
transform 1 0 84456 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_906
timestamp 1624015447
transform 1 0 84456 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_906
timestamp 1624015447
transform 1 0 84456 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_918
timestamp 1624015447
transform 1 0 85560 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_154_930
timestamp 1624015447
transform 1 0 86664 0 -1 86496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_155_918
timestamp 1624015447
transform 1 0 85560 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_930
timestamp 1624015447
transform 1 0 86664 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_918
timestamp 1624015447
transform 1 0 85560 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_156_930
timestamp 1624015447
transform 1 0 86664 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1704
timestamp 1624015447
transform 1 0 86848 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1706
timestamp 1624015447
transform 1 0 86848 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_154_933
timestamp 1624015447
transform 1 0 86940 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_945
timestamp 1624015447
transform 1 0 88044 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_942
timestamp 1624015447
transform 1 0 87768 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_933
timestamp 1624015447
transform 1 0 86940 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_945
timestamp 1624015447
transform 1 0 88044 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1705
timestamp 1624015447
transform 1 0 89424 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_154_957
timestamp 1624015447
transform 1 0 89148 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_954
timestamp 1624015447
transform 1 0 88872 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_155_961
timestamp 1624015447
transform 1 0 89516 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_957
timestamp 1624015447
transform 1 0 89148 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_997
timestamp 1624015447
transform -1 0 90896 0 -1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_999
timestamp 1624015447
transform -1 0 90896 0 1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1001
timestamp 1624015447
transform -1 0 90896 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_154_969
timestamp 1624015447
transform 1 0 90252 0 -1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_156_969
timestamp 1624015447
transform 1 0 90252 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_312
timestamp 1624015447
transform 1 0 1104 0 1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_314
timestamp 1624015447
transform 1 0 1104 0 -1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_316
timestamp 1624015447
transform 1 0 1104 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_157_3
timestamp 1624015447
transform 1 0 1380 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_15
timestamp 1624015447
transform 1 0 2484 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_3
timestamp 1624015447
transform 1 0 1380 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_15
timestamp 1624015447
transform 1 0 2484 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_3
timestamp 1624015447
transform 1 0 1380 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_15
timestamp 1624015447
transform 1 0 2484 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1454
timestamp 1624015447
transform 1 0 3772 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_157_27
timestamp 1624015447
transform 1 0 3588 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_158_27
timestamp 1624015447
transform 1 0 3588 0 -1 88672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_158_30
timestamp 1624015447
transform 1 0 3864 0 -1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_159_27
timestamp 1624015447
transform 1 0 3588 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_313
timestamp 1624015447
transform -1 0 5152 0 1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_315
timestamp 1624015447
transform -1 0 5152 0 -1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_317
timestamp 1624015447
transform -1 0 5152 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr0[6]
timestamp 1624015447
transform -1 0 4876 0 1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr0[7]
timestamp 1624015447
transform -1 0 4876 0 1 88672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_158_38
timestamp 1624015447
transform 1 0 4600 0 -1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1002
timestamp 1624015447
transform 1 0 84180 0 1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1004
timestamp 1624015447
transform 1 0 84180 0 -1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1006
timestamp 1624015447
transform 1 0 84180 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_157_906
timestamp 1624015447
transform 1 0 84456 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_906
timestamp 1624015447
transform 1 0 84456 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_906
timestamp 1624015447
transform 1 0 84456 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_918
timestamp 1624015447
transform 1 0 85560 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_930
timestamp 1624015447
transform 1 0 86664 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_918
timestamp 1624015447
transform 1 0 85560 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_158_930
timestamp 1624015447
transform 1 0 86664 0 -1 88672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_159_918
timestamp 1624015447
transform 1 0 85560 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_930
timestamp 1624015447
transform 1 0 86664 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1708
timestamp 1624015447
transform 1 0 86848 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_157_942
timestamp 1624015447
transform 1 0 87768 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_933
timestamp 1624015447
transform 1 0 86940 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_945
timestamp 1624015447
transform 1 0 88044 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_942
timestamp 1624015447
transform 1 0 87768 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1707
timestamp 1624015447
transform 1 0 89424 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1709
timestamp 1624015447
transform 1 0 89424 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_157_954
timestamp 1624015447
transform 1 0 88872 0 1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_157_961
timestamp 1624015447
transform 1 0 89516 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_957
timestamp 1624015447
transform 1 0 89148 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_954
timestamp 1624015447
transform 1 0 88872 0 1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_159_961
timestamp 1624015447
transform 1 0 89516 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1003
timestamp 1624015447
transform -1 0 90896 0 1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1005
timestamp 1624015447
transform -1 0 90896 0 -1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1007
timestamp 1624015447
transform -1 0 90896 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_158_969
timestamp 1624015447
transform 1 0 90252 0 -1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_318
timestamp 1624015447
transform 1 0 1104 0 -1 89760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_320
timestamp 1624015447
transform 1 0 1104 0 1 89760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_322
timestamp 1624015447
transform 1 0 1104 0 -1 90848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_160_3
timestamp 1624015447
transform 1 0 1380 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_15
timestamp 1624015447
transform 1 0 2484 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_3
timestamp 1624015447
transform 1 0 1380 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_15
timestamp 1624015447
transform 1 0 2484 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_3
timestamp 1624015447
transform 1 0 1380 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_15
timestamp 1624015447
transform 1 0 2484 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1455
timestamp 1624015447
transform 1 0 3772 0 -1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1456
timestamp 1624015447
transform 1 0 3772 0 -1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_160_27
timestamp 1624015447
transform 1 0 3588 0 -1 89760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_160_30
timestamp 1624015447
transform 1 0 3864 0 -1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_161_27
timestamp 1624015447
transform 1 0 3588 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_162_27
timestamp 1624015447
transform 1 0 3588 0 -1 90848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_162_30
timestamp 1624015447
transform 1 0 3864 0 -1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_319
timestamp 1624015447
transform -1 0 5152 0 -1 89760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_321
timestamp 1624015447
transform -1 0 5152 0 1 89760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_323
timestamp 1624015447
transform -1 0 5152 0 -1 90848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_160_38
timestamp 1624015447
transform 1 0 4600 0 -1 89760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_161_39
timestamp 1624015447
transform 1 0 4692 0 1 89760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_162_38
timestamp 1624015447
transform 1 0 4600 0 -1 90848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1008
timestamp 1624015447
transform 1 0 84180 0 -1 89760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1010
timestamp 1624015447
transform 1 0 84180 0 1 89760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1012
timestamp 1624015447
transform 1 0 84180 0 -1 90848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_160_906
timestamp 1624015447
transform 1 0 84456 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_906
timestamp 1624015447
transform 1 0 84456 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_906
timestamp 1624015447
transform 1 0 84456 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_918
timestamp 1624015447
transform 1 0 85560 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_160_930
timestamp 1624015447
transform 1 0 86664 0 -1 89760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_161_918
timestamp 1624015447
transform 1 0 85560 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_930
timestamp 1624015447
transform 1 0 86664 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_918
timestamp 1624015447
transform 1 0 85560 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_162_930
timestamp 1624015447
transform 1 0 86664 0 -1 90848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1710
timestamp 1624015447
transform 1 0 86848 0 -1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1712
timestamp 1624015447
transform 1 0 86848 0 -1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_160_933
timestamp 1624015447
transform 1 0 86940 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_945
timestamp 1624015447
transform 1 0 88044 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_942
timestamp 1624015447
transform 1 0 87768 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_933
timestamp 1624015447
transform 1 0 86940 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_945
timestamp 1624015447
transform 1 0 88044 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1711
timestamp 1624015447
transform 1 0 89424 0 1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_160_957
timestamp 1624015447
transform 1 0 89148 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_954
timestamp 1624015447
transform 1 0 88872 0 1 89760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_161_961
timestamp 1624015447
transform 1 0 89516 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_957
timestamp 1624015447
transform 1 0 89148 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1009
timestamp 1624015447
transform -1 0 90896 0 -1 89760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1011
timestamp 1624015447
transform -1 0 90896 0 1 89760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1013
timestamp 1624015447
transform -1 0 90896 0 -1 90848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_160_969
timestamp 1624015447
transform 1 0 90252 0 -1 89760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_162_969
timestamp 1624015447
transform 1 0 90252 0 -1 90848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_324
timestamp 1624015447
transform 1 0 1104 0 1 90848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_326
timestamp 1624015447
transform 1 0 1104 0 -1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_328
timestamp 1624015447
transform 1 0 1104 0 1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_163_3
timestamp 1624015447
transform 1 0 1380 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_15
timestamp 1624015447
transform 1 0 2484 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_3
timestamp 1624015447
transform 1 0 1380 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_15
timestamp 1624015447
transform 1 0 2484 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_3
timestamp 1624015447
transform 1 0 1380 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_15
timestamp 1624015447
transform 1 0 2484 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1457
timestamp 1624015447
transform 1 0 3772 0 -1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_163_27
timestamp 1624015447
transform 1 0 3588 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_164_27
timestamp 1624015447
transform 1 0 3588 0 -1 91936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_164_30
timestamp 1624015447
transform 1 0 3864 0 -1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_165_27
timestamp 1624015447
transform 1 0 3588 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_325
timestamp 1624015447
transform -1 0 5152 0 1 90848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_327
timestamp 1624015447
transform -1 0 5152 0 -1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_329
timestamp 1624015447
transform -1 0 5152 0 1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_163_39
timestamp 1624015447
transform 1 0 4692 0 1 90848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_164_38
timestamp 1624015447
transform 1 0 4600 0 -1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_165_39
timestamp 1624015447
transform 1 0 4692 0 1 91936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1014
timestamp 1624015447
transform 1 0 84180 0 1 90848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1016
timestamp 1624015447
transform 1 0 84180 0 -1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1018
timestamp 1624015447
transform 1 0 84180 0 1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_csb1
timestamp 1624015447
transform -1 0 84824 0 1 91936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_163_906
timestamp 1624015447
transform 1 0 84456 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_906
timestamp 1624015447
transform 1 0 84456 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_165_906
timestamp 1624015447
transform 1 0 84456 0 1 91936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_165_910
timestamp 1624015447
transform 1 0 84824 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_918
timestamp 1624015447
transform 1 0 85560 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_930
timestamp 1624015447
transform 1 0 86664 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_918
timestamp 1624015447
transform 1 0 85560 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_164_930
timestamp 1624015447
transform 1 0 86664 0 -1 91936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_165_922
timestamp 1624015447
transform 1 0 85928 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1714
timestamp 1624015447
transform 1 0 86848 0 -1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_163_942
timestamp 1624015447
transform 1 0 87768 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_933
timestamp 1624015447
transform 1 0 86940 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_945
timestamp 1624015447
transform 1 0 88044 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_934
timestamp 1624015447
transform 1 0 87032 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_946
timestamp 1624015447
transform 1 0 88136 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1713
timestamp 1624015447
transform 1 0 89424 0 1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1715
timestamp 1624015447
transform 1 0 89424 0 1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_163_954
timestamp 1624015447
transform 1 0 88872 0 1 90848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_163_961
timestamp 1624015447
transform 1 0 89516 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_957
timestamp 1624015447
transform 1 0 89148 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_165_958
timestamp 1624015447
transform 1 0 89240 0 1 91936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_165_961
timestamp 1624015447
transform 1 0 89516 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1015
timestamp 1624015447
transform -1 0 90896 0 1 90848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1017
timestamp 1624015447
transform -1 0 90896 0 -1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1019
timestamp 1624015447
transform -1 0 90896 0 1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_164_969
timestamp 1624015447
transform 1 0 90252 0 -1 91936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_330
timestamp 1624015447
transform 1 0 1104 0 -1 93024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_332
timestamp 1624015447
transform 1 0 1104 0 1 93024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_166_3
timestamp 1624015447
transform 1 0 1380 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_15
timestamp 1624015447
transform 1 0 2484 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_3
timestamp 1624015447
transform 1 0 1380 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_15
timestamp 1624015447
transform 1 0 2484 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1458
timestamp 1624015447
transform 1 0 3772 0 -1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_166_27
timestamp 1624015447
transform 1 0 3588 0 -1 93024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_166_30
timestamp 1624015447
transform 1 0 3864 0 -1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_167_27
timestamp 1624015447
transform 1 0 3588 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_331
timestamp 1624015447
transform -1 0 5152 0 -1 93024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_333
timestamp 1624015447
transform -1 0 5152 0 1 93024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_166_38
timestamp 1624015447
transform 1 0 4600 0 -1 93024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_167_39
timestamp 1624015447
transform 1 0 4692 0 1 93024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1020
timestamp 1624015447
transform 1 0 84180 0 -1 93024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1022
timestamp 1624015447
transform 1 0 84180 0 1 93024
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_addr1[0]
timestamp 1624015447
transform 1 0 84640 0 1 93024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_0_clk1
timestamp 1624015447
transform 1 0 85008 0 1 93024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_166_906
timestamp 1624015447
transform 1 0 84456 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_167_906
timestamp 1624015447
transform 1 0 84456 0 1 93024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_167_910
timestamp 1624015447
transform 1 0 84824 0 1 93024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_166_918
timestamp 1624015447
transform 1 0 85560 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_166_930
timestamp 1624015447
transform 1 0 86664 0 -1 93024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_167_914
timestamp 1624015447
transform 1 0 85192 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_926
timestamp 1624015447
transform 1 0 86296 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1716
timestamp 1624015447
transform 1 0 86848 0 -1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_166_933
timestamp 1624015447
transform 1 0 86940 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_945
timestamp 1624015447
transform 1 0 88044 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_938
timestamp 1624015447
transform 1 0 87400 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1717
timestamp 1624015447
transform 1 0 89424 0 1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_166_957
timestamp 1624015447
transform 1 0 89148 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_167_950
timestamp 1624015447
transform 1 0 88504 0 1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_167_958
timestamp 1624015447
transform 1 0 89240 0 1 93024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_167_961
timestamp 1624015447
transform 1 0 89516 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1021
timestamp 1624015447
transform -1 0 90896 0 -1 93024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1023
timestamp 1624015447
transform -1 0 90896 0 1 93024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_166_969
timestamp 1624015447
transform 1 0 90252 0 -1 93024
box -38 -48 406 592
use sram_1rw1r_32_256_8_sky130  SRAM_0
timestamp 1624446551
transform 1 0 6000 0 1 2361
box 0 0 77296 91247
use sky130_fd_sc_hd__decap_3  PHY_334
timestamp 1624015447
transform 1 0 1104 0 -1 94112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_336
timestamp 1624015447
transform 1 0 1104 0 1 94112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_338
timestamp 1624015447
transform 1 0 1104 0 -1 95200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_168_3
timestamp 1624015447
transform 1 0 1380 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_15
timestamp 1624015447
transform 1 0 2484 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_3
timestamp 1624015447
transform 1 0 1380 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_15
timestamp 1624015447
transform 1 0 2484 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_3
timestamp 1624015447
transform 1 0 1380 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_15
timestamp 1624015447
transform 1 0 2484 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1459
timestamp 1624015447
transform 1 0 3772 0 -1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1460
timestamp 1624015447
transform 1 0 3772 0 -1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_168_27
timestamp 1624015447
transform 1 0 3588 0 -1 94112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_168_30
timestamp 1624015447
transform 1 0 3864 0 -1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_169_27
timestamp 1624015447
transform 1 0 3588 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_170_27
timestamp 1624015447
transform 1 0 3588 0 -1 95200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_170_30
timestamp 1624015447
transform 1 0 3864 0 -1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_335
timestamp 1624015447
transform -1 0 5152 0 -1 94112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_337
timestamp 1624015447
transform -1 0 5152 0 1 94112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_339
timestamp 1624015447
transform -1 0 5152 0 -1 95200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_168_38
timestamp 1624015447
transform 1 0 4600 0 -1 94112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_169_39
timestamp 1624015447
transform 1 0 4692 0 1 94112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_170_38
timestamp 1624015447
transform 1 0 4600 0 -1 95200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1024
timestamp 1624015447
transform 1 0 84180 0 -1 94112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1026
timestamp 1624015447
transform 1 0 84180 0 1 94112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1028
timestamp 1624015447
transform 1 0 84180 0 -1 95200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_168_906
timestamp 1624015447
transform 1 0 84456 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_906
timestamp 1624015447
transform 1 0 84456 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_906
timestamp 1624015447
transform 1 0 84456 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_918
timestamp 1624015447
transform 1 0 85560 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_918
timestamp 1624015447
transform 1 0 85560 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_918
timestamp 1624015447
transform 1 0 85560 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_945
timestamp 1624015447
transform 1 0 88044 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_933
timestamp 1624015447
transform 1 0 86940 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_168_930
timestamp 1624015447
transform 1 0 86664 0 -1 94112
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1718
timestamp 1624015447
transform 1 0 86848 0 -1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_170_945
timestamp 1624015447
transform 1 0 88044 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_933
timestamp 1624015447
transform 1 0 86940 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_170_930
timestamp 1624015447
transform 1 0 86664 0 -1 95200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_169_942
timestamp 1624015447
transform 1 0 87768 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_930
timestamp 1624015447
transform 1 0 86664 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1720
timestamp 1624015447
transform 1 0 86848 0 -1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1719
timestamp 1624015447
transform 1 0 89424 0 1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_168_957
timestamp 1624015447
transform 1 0 89148 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_954
timestamp 1624015447
transform 1 0 88872 0 1 94112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_169_961
timestamp 1624015447
transform 1 0 89516 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_957
timestamp 1624015447
transform 1 0 89148 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1025
timestamp 1624015447
transform -1 0 90896 0 -1 94112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1027
timestamp 1624015447
transform -1 0 90896 0 1 94112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1029
timestamp 1624015447
transform -1 0 90896 0 -1 95200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_168_969
timestamp 1624015447
transform 1 0 90252 0 -1 94112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_170_969
timestamp 1624015447
transform 1 0 90252 0 -1 95200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_340
timestamp 1624015447
transform 1 0 1104 0 1 95200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_342
timestamp 1624015447
transform 1 0 1104 0 -1 96288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_344
timestamp 1624015447
transform 1 0 1104 0 1 96288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_171_3
timestamp 1624015447
transform 1 0 1380 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_15
timestamp 1624015447
transform 1 0 2484 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_3
timestamp 1624015447
transform 1 0 1380 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_15
timestamp 1624015447
transform 1 0 2484 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_3
timestamp 1624015447
transform 1 0 1380 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_173_15
timestamp 1624015447
transform 1 0 2484 0 1 96288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_171_27
timestamp 1624015447
transform 1 0 3588 0 1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_wmask0[1]
timestamp 1624015447
transform -1 0 4508 0 1 95200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_173_25
timestamp 1624015447
transform 1 0 3404 0 1 96288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_clk0
timestamp 1624015447
transform -1 0 3772 0 -1 96288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[8]
timestamp 1624015447
transform -1 0 3404 0 1 96288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[2]
timestamp 1624015447
transform -1 0 3772 0 1 96288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_173_33
timestamp 1624015447
transform 1 0 4140 0 1 96288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_173_29
timestamp 1624015447
transform 1 0 3772 0 1 96288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_172_34
timestamp 1624015447
transform 1 0 4232 0 -1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_172_30
timestamp 1624015447
transform 1 0 3864 0 -1 96288
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[20]
timestamp 1624015447
transform 1 0 4324 0 -1 96288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[18]
timestamp 1624015447
transform 1 0 3956 0 1 96288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[14]
timestamp 1624015447
transform -1 0 4508 0 1 96288
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1461
timestamp 1624015447
transform 1 0 3772 0 -1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_341
timestamp 1624015447
transform -1 0 5152 0 1 95200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_343
timestamp 1624015447
transform -1 0 5152 0 -1 96288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_345
timestamp 1624015447
transform -1 0 5152 0 1 96288
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[11]
timestamp 1624015447
transform 1 0 4692 0 1 96288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[17]
timestamp 1624015447
transform 1 0 4692 0 -1 96288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[7]
timestamp 1624015447
transform 1 0 4692 0 1 95200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_171_37
timestamp 1624015447
transform 1 0 4508 0 1 95200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_172_37
timestamp 1624015447
transform 1 0 4508 0 -1 96288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_173_37
timestamp 1624015447
transform 1 0 4508 0 1 96288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_171_906
timestamp 1624015447
transform 1 0 84456 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1030
timestamp 1624015447
transform 1 0 84180 0 1 95200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_173_910
timestamp 1624015447
transform 1 0 84824 0 1 96288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_173_906
timestamp 1624015447
transform 1 0 84456 0 1 96288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_172_910
timestamp 1624015447
transform 1 0 84824 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_172_906
timestamp 1624015447
transform 1 0 84456 0 -1 96288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[31]
timestamp 1624015447
transform 1 0 84640 0 -1 96288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[26]
timestamp 1624015447
transform 1 0 84640 0 1 96288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1034
timestamp 1624015447
transform 1 0 84180 0 1 96288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1032
timestamp 1624015447
transform 1 0 84180 0 -1 96288
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[28]
timestamp 1624015447
transform 1 0 85008 0 1 96288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_171_918
timestamp 1624015447
transform 1 0 85560 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_172_922
timestamp 1624015447
transform 1 0 85928 0 -1 96288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_173_914
timestamp 1624015447
transform 1 0 85192 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_926
timestamp 1624015447
transform 1 0 86296 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1722
timestamp 1624015447
transform 1 0 86848 0 -1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_930
timestamp 1624015447
transform 1 0 86664 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_942
timestamp 1624015447
transform 1 0 87768 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_172_930
timestamp 1624015447
transform 1 0 86664 0 -1 96288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_172_933
timestamp 1624015447
transform 1 0 86940 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_945
timestamp 1624015447
transform 1 0 88044 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_938
timestamp 1624015447
transform 1 0 87400 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1721
timestamp 1624015447
transform 1 0 89424 0 1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1723
timestamp 1624015447
transform 1 0 89424 0 1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_171_954
timestamp 1624015447
transform 1 0 88872 0 1 95200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_171_961
timestamp 1624015447
transform 1 0 89516 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_957
timestamp 1624015447
transform 1 0 89148 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_173_950
timestamp 1624015447
transform 1 0 88504 0 1 96288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_173_958
timestamp 1624015447
transform 1 0 89240 0 1 96288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_173_961
timestamp 1624015447
transform 1 0 89516 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1031
timestamp 1624015447
transform -1 0 90896 0 1 95200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1033
timestamp 1624015447
transform -1 0 90896 0 -1 96288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1035
timestamp 1624015447
transform -1 0 90896 0 1 96288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_172_969
timestamp 1624015447
transform 1 0 90252 0 -1 96288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_175_15
timestamp 1624015447
transform 1 0 2484 0 1 97376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_175_3
timestamp 1624015447
transform 1 0 1380 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_174_17
timestamp 1624015447
transform 1 0 2668 0 -1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_174_13
timestamp 1624015447
transform 1 0 2300 0 -1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_174_3
timestamp 1624015447
transform 1 0 1380 0 -1 97376
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_wmask0[0]
timestamp 1624015447
transform -1 0 2300 0 -1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[5]
timestamp 1624015447
transform -1 0 2668 0 -1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_348
timestamp 1624015447
transform 1 0 1104 0 1 97376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_346
timestamp 1624015447
transform 1 0 1104 0 -1 97376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_176_15
timestamp 1624015447
transform 1 0 2484 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_3
timestamp 1624015447
transform 1 0 1380 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_350
timestamp 1624015447
transform 1 0 1104 0 -1 98464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_175_21
timestamp 1624015447
transform 1 0 3036 0 1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_174_21
timestamp 1624015447
transform 1 0 3036 0 -1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_wmask0[3]
timestamp 1624015447
transform -1 0 3036 0 1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[4]
timestamp 1624015447
transform -1 0 3404 0 1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[3]
timestamp 1624015447
transform -1 0 3036 0 -1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[19]
timestamp 1624015447
transform -1 0 3404 0 -1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_175_25
timestamp 1624015447
transform 1 0 3404 0 1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_174_25
timestamp 1624015447
transform 1 0 3404 0 -1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[21]
timestamp 1624015447
transform -1 0 3772 0 1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[13]
timestamp 1624015447
transform -1 0 3772 0 -1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_175_29
timestamp 1624015447
transform 1 0 3772 0 1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_174_30
timestamp 1624015447
transform 1 0 3864 0 -1 97376
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[15]
timestamp 1624015447
transform -1 0 4140 0 1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1462
timestamp 1624015447
transform 1 0 3772 0 -1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_175_33
timestamp 1624015447
transform 1 0 4140 0 1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_174_34
timestamp 1624015447
transform 1 0 4232 0 -1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[12]
timestamp 1624015447
transform -1 0 4508 0 1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[0]
timestamp 1624015447
transform -1 0 4508 0 -1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_wmask0[2]
timestamp 1624015447
transform -1 0 3772 0 -1 98464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_176_30
timestamp 1624015447
transform 1 0 3864 0 -1 98464
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1463
timestamp 1624015447
transform 1 0 3772 0 -1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_176_34
timestamp 1624015447
transform 1 0 4232 0 -1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[1]
timestamp 1624015447
transform 1 0 4324 0 -1 98464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_347
timestamp 1624015447
transform -1 0 5152 0 -1 97376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_349
timestamp 1624015447
transform -1 0 5152 0 1 97376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_351
timestamp 1624015447
transform -1 0 5152 0 -1 98464
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_addr0[0]
timestamp 1624015447
transform -1 0 4876 0 -1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[10]
timestamp 1624015447
transform -1 0 4876 0 1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[16]
timestamp 1624015447
transform -1 0 4876 0 -1 98464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_174_37
timestamp 1624015447
transform 1 0 4508 0 -1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_175_37
timestamp 1624015447
transform 1 0 4508 0 1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_176_37
timestamp 1624015447
transform 1 0 4508 0 -1 98464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_175_910
timestamp 1624015447
transform 1 0 84824 0 1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_175_906
timestamp 1624015447
transform 1 0 84456 0 1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_174_910
timestamp 1624015447
transform 1 0 84824 0 -1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_174_906
timestamp 1624015447
transform 1 0 84456 0 -1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[24]
timestamp 1624015447
transform 1 0 84640 0 1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[22]
timestamp 1624015447
transform 1 0 84640 0 -1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1038
timestamp 1624015447
transform 1 0 84180 0 1 97376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1036
timestamp 1624015447
transform 1 0 84180 0 -1 97376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_176_910
timestamp 1624015447
transform 1 0 84824 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_176_906
timestamp 1624015447
transform 1 0 84456 0 -1 98464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[29]
timestamp 1624015447
transform 1 0 84640 0 -1 98464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1040
timestamp 1624015447
transform 1 0 84180 0 -1 98464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_175_926
timestamp 1624015447
transform 1 0 86296 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_914
timestamp 1624015447
transform 1 0 85192 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_174_922
timestamp 1624015447
transform 1 0 85928 0 -1 97376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_174_918
timestamp 1624015447
transform 1 0 85560 0 -1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_174_914
timestamp 1624015447
transform 1 0 85192 0 -1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[30]
timestamp 1624015447
transform 1 0 85744 0 -1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[27]
timestamp 1624015447
transform 1 0 85008 0 1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[25]
timestamp 1624015447
transform 1 0 85376 0 -1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[23]
timestamp 1624015447
transform 1 0 85008 0 -1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_176_922
timestamp 1624015447
transform 1 0 85928 0 -1 98464
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1724
timestamp 1624015447
transform 1 0 86848 0 -1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1726
timestamp 1624015447
transform 1 0 86848 0 -1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_174_930
timestamp 1624015447
transform 1 0 86664 0 -1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_174_933
timestamp 1624015447
transform 1 0 86940 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_945
timestamp 1624015447
transform 1 0 88044 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_938
timestamp 1624015447
transform 1 0 87400 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_176_930
timestamp 1624015447
transform 1 0 86664 0 -1 98464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_176_933
timestamp 1624015447
transform 1 0 86940 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_945
timestamp 1624015447
transform 1 0 88044 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1725
timestamp 1624015447
transform 1 0 89424 0 1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_174_957
timestamp 1624015447
transform 1 0 89148 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_175_950
timestamp 1624015447
transform 1 0 88504 0 1 97376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_175_958
timestamp 1624015447
transform 1 0 89240 0 1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_175_961
timestamp 1624015447
transform 1 0 89516 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_957
timestamp 1624015447
transform 1 0 89148 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1037
timestamp 1624015447
transform -1 0 90896 0 -1 97376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1039
timestamp 1624015447
transform -1 0 90896 0 1 97376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1041
timestamp 1624015447
transform -1 0 90896 0 -1 98464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_174_969
timestamp 1624015447
transform 1 0 90252 0 -1 97376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_176_969
timestamp 1624015447
transform 1 0 90252 0 -1 98464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_178_15
timestamp 1624015447
transform 1 0 2484 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_3
timestamp 1624015447
transform 1 0 1380 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_15
timestamp 1624015447
transform 1 0 2484 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_3
timestamp 1624015447
transform 1 0 1380 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_354
timestamp 1624015447
transform 1 0 1104 0 -1 99552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_352
timestamp 1624015447
transform 1 0 1104 0 1 98464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_179_15
timestamp 1624015447
transform 1 0 2484 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_3
timestamp 1624015447
transform 1 0 1380 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_356
timestamp 1624015447
transform 1 0 1104 0 1 99552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_180_15
timestamp 1624015447
transform 1 0 2484 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_3
timestamp 1624015447
transform 1 0 1380 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_358
timestamp 1624015447
transform 1 0 1104 0 -1 100640
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1464
timestamp 1624015447
transform 1 0 3772 0 -1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1465
timestamp 1624015447
transform 1 0 3772 0 -1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[9]
timestamp 1624015447
transform 1 0 4324 0 1 98464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_177_27
timestamp 1624015447
transform 1 0 3588 0 1 98464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_178_27
timestamp 1624015447
transform 1 0 3588 0 -1 99552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_178_30
timestamp 1624015447
transform 1 0 3864 0 -1 99552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_179_27
timestamp 1624015447
transform 1 0 3588 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_180_27
timestamp 1624015447
transform 1 0 3588 0 -1 100640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_180_30
timestamp 1624015447
transform 1 0 3864 0 -1 100640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_353
timestamp 1624015447
transform -1 0 5152 0 1 98464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_355
timestamp 1624015447
transform -1 0 5152 0 -1 99552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_357
timestamp 1624015447
transform -1 0 5152 0 1 99552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_359
timestamp 1624015447
transform -1 0 5152 0 -1 100640
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_din0[6]
timestamp 1624015447
transform 1 0 4692 0 1 98464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_177_37
timestamp 1624015447
transform 1 0 4508 0 1 98464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_178_38
timestamp 1624015447
transform 1 0 4600 0 -1 99552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_179_39
timestamp 1624015447
transform 1 0 4692 0 1 99552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_180_38
timestamp 1624015447
transform 1 0 4600 0 -1 100640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1042
timestamp 1624015447
transform 1 0 84180 0 1 98464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1044
timestamp 1624015447
transform 1 0 84180 0 -1 99552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1046
timestamp 1624015447
transform 1 0 84180 0 1 99552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1048
timestamp 1624015447
transform 1 0 84180 0 -1 100640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_177_906
timestamp 1624015447
transform 1 0 84456 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_906
timestamp 1624015447
transform 1 0 84456 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_906
timestamp 1624015447
transform 1 0 84456 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_906
timestamp 1624015447
transform 1 0 84456 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_918
timestamp 1624015447
transform 1 0 85560 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_918
timestamp 1624015447
transform 1 0 85560 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_918
timestamp 1624015447
transform 1 0 85560 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_918
timestamp 1624015447
transform 1 0 85560 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_945
timestamp 1624015447
transform 1 0 88044 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_933
timestamp 1624015447
transform 1 0 86940 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_178_930
timestamp 1624015447
transform 1 0 86664 0 -1 99552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_177_942
timestamp 1624015447
transform 1 0 87768 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_930
timestamp 1624015447
transform 1 0 86664 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1728
timestamp 1624015447
transform 1 0 86848 0 -1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_179_942
timestamp 1624015447
transform 1 0 87768 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_930
timestamp 1624015447
transform 1 0 86664 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_945
timestamp 1624015447
transform 1 0 88044 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_933
timestamp 1624015447
transform 1 0 86940 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_180_930
timestamp 1624015447
transform 1 0 86664 0 -1 100640
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1730
timestamp 1624015447
transform 1 0 86848 0 -1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1727
timestamp 1624015447
transform 1 0 89424 0 1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1729
timestamp 1624015447
transform 1 0 89424 0 1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_177_954
timestamp 1624015447
transform 1 0 88872 0 1 98464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_177_961
timestamp 1624015447
transform 1 0 89516 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_957
timestamp 1624015447
transform 1 0 89148 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_954
timestamp 1624015447
transform 1 0 88872 0 1 99552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_179_961
timestamp 1624015447
transform 1 0 89516 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_957
timestamp 1624015447
transform 1 0 89148 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1043
timestamp 1624015447
transform -1 0 90896 0 1 98464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1045
timestamp 1624015447
transform -1 0 90896 0 -1 99552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1047
timestamp 1624015447
transform -1 0 90896 0 1 99552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1049
timestamp 1624015447
transform -1 0 90896 0 -1 100640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_178_969
timestamp 1624015447
transform 1 0 90252 0 -1 99552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_180_969
timestamp 1624015447
transform 1 0 90252 0 -1 100640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_360
timestamp 1624015447
transform 1 0 1104 0 1 100640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_362
timestamp 1624015447
transform 1 0 1104 0 -1 101728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_364
timestamp 1624015447
transform 1 0 1104 0 1 101728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_181_3
timestamp 1624015447
transform 1 0 1380 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_15
timestamp 1624015447
transform 1 0 2484 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_3
timestamp 1624015447
transform 1 0 1380 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_15
timestamp 1624015447
transform 1 0 2484 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_3
timestamp 1624015447
transform 1 0 1380 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_15
timestamp 1624015447
transform 1 0 2484 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1466
timestamp 1624015447
transform 1 0 3772 0 -1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_181_27
timestamp 1624015447
transform 1 0 3588 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_182_27
timestamp 1624015447
transform 1 0 3588 0 -1 101728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_182_30
timestamp 1624015447
transform 1 0 3864 0 -1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_183_27
timestamp 1624015447
transform 1 0 3588 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_361
timestamp 1624015447
transform -1 0 5152 0 1 100640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_363
timestamp 1624015447
transform -1 0 5152 0 -1 101728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_365
timestamp 1624015447
transform -1 0 5152 0 1 101728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_181_39
timestamp 1624015447
transform 1 0 4692 0 1 100640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_182_38
timestamp 1624015447
transform 1 0 4600 0 -1 101728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_183_39
timestamp 1624015447
transform 1 0 4692 0 1 101728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1050
timestamp 1624015447
transform 1 0 84180 0 1 100640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1052
timestamp 1624015447
transform 1 0 84180 0 -1 101728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1054
timestamp 1624015447
transform 1 0 84180 0 1 101728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_181_906
timestamp 1624015447
transform 1 0 84456 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_906
timestamp 1624015447
transform 1 0 84456 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_906
timestamp 1624015447
transform 1 0 84456 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_918
timestamp 1624015447
transform 1 0 85560 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_918
timestamp 1624015447
transform 1 0 85560 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_918
timestamp 1624015447
transform 1 0 85560 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1732
timestamp 1624015447
transform 1 0 86848 0 -1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_181_930
timestamp 1624015447
transform 1 0 86664 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_942
timestamp 1624015447
transform 1 0 87768 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_182_930
timestamp 1624015447
transform 1 0 86664 0 -1 101728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_182_933
timestamp 1624015447
transform 1 0 86940 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_945
timestamp 1624015447
transform 1 0 88044 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_930
timestamp 1624015447
transform 1 0 86664 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_942
timestamp 1624015447
transform 1 0 87768 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1731
timestamp 1624015447
transform 1 0 89424 0 1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1733
timestamp 1624015447
transform 1 0 89424 0 1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_181_954
timestamp 1624015447
transform 1 0 88872 0 1 100640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_181_961
timestamp 1624015447
transform 1 0 89516 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_957
timestamp 1624015447
transform 1 0 89148 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_183_954
timestamp 1624015447
transform 1 0 88872 0 1 101728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_183_961
timestamp 1624015447
transform 1 0 89516 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1051
timestamp 1624015447
transform -1 0 90896 0 1 100640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1053
timestamp 1624015447
transform -1 0 90896 0 -1 101728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1055
timestamp 1624015447
transform -1 0 90896 0 1 101728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_182_969
timestamp 1624015447
transform 1 0 90252 0 -1 101728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_366
timestamp 1624015447
transform 1 0 1104 0 -1 102816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_368
timestamp 1624015447
transform 1 0 1104 0 1 102816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_370
timestamp 1624015447
transform 1 0 1104 0 -1 103904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_184_3
timestamp 1624015447
transform 1 0 1380 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_15
timestamp 1624015447
transform 1 0 2484 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_3
timestamp 1624015447
transform 1 0 1380 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_15
timestamp 1624015447
transform 1 0 2484 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_3
timestamp 1624015447
transform 1 0 1380 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_15
timestamp 1624015447
transform 1 0 2484 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1467
timestamp 1624015447
transform 1 0 3772 0 -1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1468
timestamp 1624015447
transform 1 0 3772 0 -1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_184_27
timestamp 1624015447
transform 1 0 3588 0 -1 102816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_184_30
timestamp 1624015447
transform 1 0 3864 0 -1 102816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_185_27
timestamp 1624015447
transform 1 0 3588 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_186_27
timestamp 1624015447
transform 1 0 3588 0 -1 103904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_186_30
timestamp 1624015447
transform 1 0 3864 0 -1 103904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_367
timestamp 1624015447
transform -1 0 5152 0 -1 102816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_369
timestamp 1624015447
transform -1 0 5152 0 1 102816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_371
timestamp 1624015447
transform -1 0 5152 0 -1 103904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_184_38
timestamp 1624015447
transform 1 0 4600 0 -1 102816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_185_39
timestamp 1624015447
transform 1 0 4692 0 1 102816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_186_38
timestamp 1624015447
transform 1 0 4600 0 -1 103904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1056
timestamp 1624015447
transform 1 0 84180 0 -1 102816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1058
timestamp 1624015447
transform 1 0 84180 0 1 102816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1060
timestamp 1624015447
transform 1 0 84180 0 -1 103904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_184_906
timestamp 1624015447
transform 1 0 84456 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_906
timestamp 1624015447
transform 1 0 84456 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_906
timestamp 1624015447
transform 1 0 84456 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_918
timestamp 1624015447
transform 1 0 85560 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_918
timestamp 1624015447
transform 1 0 85560 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_918
timestamp 1624015447
transform 1 0 85560 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_945
timestamp 1624015447
transform 1 0 88044 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_933
timestamp 1624015447
transform 1 0 86940 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_184_930
timestamp 1624015447
transform 1 0 86664 0 -1 102816
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1734
timestamp 1624015447
transform 1 0 86848 0 -1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_942
timestamp 1624015447
transform 1 0 87768 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_930
timestamp 1624015447
transform 1 0 86664 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_945
timestamp 1624015447
transform 1 0 88044 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_933
timestamp 1624015447
transform 1 0 86940 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_186_930
timestamp 1624015447
transform 1 0 86664 0 -1 103904
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1736
timestamp 1624015447
transform 1 0 86848 0 -1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1735
timestamp 1624015447
transform 1 0 89424 0 1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_184_957
timestamp 1624015447
transform 1 0 89148 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_185_954
timestamp 1624015447
transform 1 0 88872 0 1 102816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_185_961
timestamp 1624015447
transform 1 0 89516 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_957
timestamp 1624015447
transform 1 0 89148 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1057
timestamp 1624015447
transform -1 0 90896 0 -1 102816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1059
timestamp 1624015447
transform -1 0 90896 0 1 102816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1061
timestamp 1624015447
transform -1 0 90896 0 -1 103904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_184_969
timestamp 1624015447
transform 1 0 90252 0 -1 102816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_186_969
timestamp 1624015447
transform 1 0 90252 0 -1 103904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_372
timestamp 1624015447
transform 1 0 1104 0 1 103904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_374
timestamp 1624015447
transform 1 0 1104 0 -1 104992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_376
timestamp 1624015447
transform 1 0 1104 0 1 104992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_187_3
timestamp 1624015447
transform 1 0 1380 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_15
timestamp 1624015447
transform 1 0 2484 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_3
timestamp 1624015447
transform 1 0 1380 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_15
timestamp 1624015447
transform 1 0 2484 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_3
timestamp 1624015447
transform 1 0 1380 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_15
timestamp 1624015447
transform 1 0 2484 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1469
timestamp 1624015447
transform 1 0 3772 0 -1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_187_27
timestamp 1624015447
transform 1 0 3588 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_188_27
timestamp 1624015447
transform 1 0 3588 0 -1 104992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_188_30
timestamp 1624015447
transform 1 0 3864 0 -1 104992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_189_27
timestamp 1624015447
transform 1 0 3588 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_373
timestamp 1624015447
transform -1 0 5152 0 1 103904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_375
timestamp 1624015447
transform -1 0 5152 0 -1 104992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_377
timestamp 1624015447
transform -1 0 5152 0 1 104992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_187_39
timestamp 1624015447
transform 1 0 4692 0 1 103904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_188_38
timestamp 1624015447
transform 1 0 4600 0 -1 104992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_189_39
timestamp 1624015447
transform 1 0 4692 0 1 104992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1062
timestamp 1624015447
transform 1 0 84180 0 1 103904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1064
timestamp 1624015447
transform 1 0 84180 0 -1 104992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1066
timestamp 1624015447
transform 1 0 84180 0 1 104992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_187_906
timestamp 1624015447
transform 1 0 84456 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_906
timestamp 1624015447
transform 1 0 84456 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_906
timestamp 1624015447
transform 1 0 84456 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_918
timestamp 1624015447
transform 1 0 85560 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_918
timestamp 1624015447
transform 1 0 85560 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_918
timestamp 1624015447
transform 1 0 85560 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1738
timestamp 1624015447
transform 1 0 86848 0 -1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_187_930
timestamp 1624015447
transform 1 0 86664 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_942
timestamp 1624015447
transform 1 0 87768 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_188_930
timestamp 1624015447
transform 1 0 86664 0 -1 104992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_188_933
timestamp 1624015447
transform 1 0 86940 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_945
timestamp 1624015447
transform 1 0 88044 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_930
timestamp 1624015447
transform 1 0 86664 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_942
timestamp 1624015447
transform 1 0 87768 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1737
timestamp 1624015447
transform 1 0 89424 0 1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1739
timestamp 1624015447
transform 1 0 89424 0 1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_187_954
timestamp 1624015447
transform 1 0 88872 0 1 103904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_187_961
timestamp 1624015447
transform 1 0 89516 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_957
timestamp 1624015447
transform 1 0 89148 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_189_954
timestamp 1624015447
transform 1 0 88872 0 1 104992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_189_961
timestamp 1624015447
transform 1 0 89516 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1063
timestamp 1624015447
transform -1 0 90896 0 1 103904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1065
timestamp 1624015447
transform -1 0 90896 0 -1 104992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1067
timestamp 1624015447
transform -1 0 90896 0 1 104992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_188_969
timestamp 1624015447
transform 1 0 90252 0 -1 104992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_378
timestamp 1624015447
transform 1 0 1104 0 -1 106080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_380
timestamp 1624015447
transform 1 0 1104 0 1 106080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_382
timestamp 1624015447
transform 1 0 1104 0 -1 107168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_190_3
timestamp 1624015447
transform 1 0 1380 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_15
timestamp 1624015447
transform 1 0 2484 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_3
timestamp 1624015447
transform 1 0 1380 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_15
timestamp 1624015447
transform 1 0 2484 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_3
timestamp 1624015447
transform 1 0 1380 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_15
timestamp 1624015447
transform 1 0 2484 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1624015447
transform 1 0 4232 0 -1 106080
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1470
timestamp 1624015447
transform 1 0 3772 0 -1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1471
timestamp 1624015447
transform 1 0 3772 0 -1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_190_27
timestamp 1624015447
transform 1 0 3588 0 -1 106080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_190_30
timestamp 1624015447
transform 1 0 3864 0 -1 106080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_191_27
timestamp 1624015447
transform 1 0 3588 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_192_27
timestamp 1624015447
transform 1 0 3588 0 -1 107168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_192_30
timestamp 1624015447
transform 1 0 3864 0 -1 107168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_379
timestamp 1624015447
transform -1 0 5152 0 -1 106080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_381
timestamp 1624015447
transform -1 0 5152 0 1 106080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_383
timestamp 1624015447
transform -1 0 5152 0 -1 107168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_190_37
timestamp 1624015447
transform 1 0 4508 0 -1 106080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_191_39
timestamp 1624015447
transform 1 0 4692 0 1 106080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_192_38
timestamp 1624015447
transform 1 0 4600 0 -1 107168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1068
timestamp 1624015447
transform 1 0 84180 0 -1 106080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1070
timestamp 1624015447
transform 1 0 84180 0 1 106080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1072
timestamp 1624015447
transform 1 0 84180 0 -1 107168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_190_906
timestamp 1624015447
transform 1 0 84456 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_906
timestamp 1624015447
transform 1 0 84456 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_906
timestamp 1624015447
transform 1 0 84456 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_918
timestamp 1624015447
transform 1 0 85560 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_918
timestamp 1624015447
transform 1 0 85560 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_918
timestamp 1624015447
transform 1 0 85560 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_945
timestamp 1624015447
transform 1 0 88044 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_933
timestamp 1624015447
transform 1 0 86940 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_190_930
timestamp 1624015447
transform 1 0 86664 0 -1 106080
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1740
timestamp 1624015447
transform 1 0 86848 0 -1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_942
timestamp 1624015447
transform 1 0 87768 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_930
timestamp 1624015447
transform 1 0 86664 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_945
timestamp 1624015447
transform 1 0 88044 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_933
timestamp 1624015447
transform 1 0 86940 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_192_930
timestamp 1624015447
transform 1 0 86664 0 -1 107168
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1742
timestamp 1624015447
transform 1 0 86848 0 -1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1741
timestamp 1624015447
transform 1 0 89424 0 1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_190_957
timestamp 1624015447
transform 1 0 89148 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_191_954
timestamp 1624015447
transform 1 0 88872 0 1 106080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_191_961
timestamp 1624015447
transform 1 0 89516 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_957
timestamp 1624015447
transform 1 0 89148 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1069
timestamp 1624015447
transform -1 0 90896 0 -1 106080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1071
timestamp 1624015447
transform -1 0 90896 0 1 106080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1073
timestamp 1624015447
transform -1 0 90896 0 -1 107168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_190_969
timestamp 1624015447
transform 1 0 90252 0 -1 106080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_192_969
timestamp 1624015447
transform 1 0 90252 0 -1 107168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_384
timestamp 1624015447
transform 1 0 1104 0 1 107168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_386
timestamp 1624015447
transform 1 0 1104 0 -1 108256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_388
timestamp 1624015447
transform 1 0 1104 0 1 108256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_193_3
timestamp 1624015447
transform 1 0 1380 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_15
timestamp 1624015447
transform 1 0 2484 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_3
timestamp 1624015447
transform 1 0 1380 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_15
timestamp 1624015447
transform 1 0 2484 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_3
timestamp 1624015447
transform 1 0 1380 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_15
timestamp 1624015447
transform 1 0 2484 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1472
timestamp 1624015447
transform 1 0 3772 0 -1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_193_27
timestamp 1624015447
transform 1 0 3588 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_194_27
timestamp 1624015447
transform 1 0 3588 0 -1 108256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_194_30
timestamp 1624015447
transform 1 0 3864 0 -1 108256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_195_27
timestamp 1624015447
transform 1 0 3588 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_385
timestamp 1624015447
transform -1 0 5152 0 1 107168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_387
timestamp 1624015447
transform -1 0 5152 0 -1 108256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_389
timestamp 1624015447
transform -1 0 5152 0 1 108256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_193_39
timestamp 1624015447
transform 1 0 4692 0 1 107168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_194_38
timestamp 1624015447
transform 1 0 4600 0 -1 108256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_195_39
timestamp 1624015447
transform 1 0 4692 0 1 108256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1074
timestamp 1624015447
transform 1 0 84180 0 1 107168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1076
timestamp 1624015447
transform 1 0 84180 0 -1 108256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1078
timestamp 1624015447
transform 1 0 84180 0 1 108256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_193_906
timestamp 1624015447
transform 1 0 84456 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_906
timestamp 1624015447
transform 1 0 84456 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_906
timestamp 1624015447
transform 1 0 84456 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_918
timestamp 1624015447
transform 1 0 85560 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_918
timestamp 1624015447
transform 1 0 85560 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_918
timestamp 1624015447
transform 1 0 85560 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1744
timestamp 1624015447
transform 1 0 86848 0 -1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_193_930
timestamp 1624015447
transform 1 0 86664 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_942
timestamp 1624015447
transform 1 0 87768 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_194_930
timestamp 1624015447
transform 1 0 86664 0 -1 108256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_194_933
timestamp 1624015447
transform 1 0 86940 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_945
timestamp 1624015447
transform 1 0 88044 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_930
timestamp 1624015447
transform 1 0 86664 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_942
timestamp 1624015447
transform 1 0 87768 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1743
timestamp 1624015447
transform 1 0 89424 0 1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1745
timestamp 1624015447
transform 1 0 89424 0 1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_193_954
timestamp 1624015447
transform 1 0 88872 0 1 107168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_193_961
timestamp 1624015447
transform 1 0 89516 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_957
timestamp 1624015447
transform 1 0 89148 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_195_954
timestamp 1624015447
transform 1 0 88872 0 1 108256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_195_961
timestamp 1624015447
transform 1 0 89516 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1075
timestamp 1624015447
transform -1 0 90896 0 1 107168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1077
timestamp 1624015447
transform -1 0 90896 0 -1 108256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1079
timestamp 1624015447
transform -1 0 90896 0 1 108256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_194_969
timestamp 1624015447
transform 1 0 90252 0 -1 108256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_390
timestamp 1624015447
transform 1 0 1104 0 -1 109344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_392
timestamp 1624015447
transform 1 0 1104 0 1 109344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_394
timestamp 1624015447
transform 1 0 1104 0 -1 110432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_196_3
timestamp 1624015447
transform 1 0 1380 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_15
timestamp 1624015447
transform 1 0 2484 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_3
timestamp 1624015447
transform 1 0 1380 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_15
timestamp 1624015447
transform 1 0 2484 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_3
timestamp 1624015447
transform 1 0 1380 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_15
timestamp 1624015447
transform 1 0 2484 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1473
timestamp 1624015447
transform 1 0 3772 0 -1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1474
timestamp 1624015447
transform 1 0 3772 0 -1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_196_27
timestamp 1624015447
transform 1 0 3588 0 -1 109344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_196_30
timestamp 1624015447
transform 1 0 3864 0 -1 109344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_197_27
timestamp 1624015447
transform 1 0 3588 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_198_27
timestamp 1624015447
transform 1 0 3588 0 -1 110432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_198_30
timestamp 1624015447
transform 1 0 3864 0 -1 110432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_391
timestamp 1624015447
transform -1 0 5152 0 -1 109344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_393
timestamp 1624015447
transform -1 0 5152 0 1 109344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_395
timestamp 1624015447
transform -1 0 5152 0 -1 110432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_196_38
timestamp 1624015447
transform 1 0 4600 0 -1 109344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_197_39
timestamp 1624015447
transform 1 0 4692 0 1 109344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_198_38
timestamp 1624015447
transform 1 0 4600 0 -1 110432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1080
timestamp 1624015447
transform 1 0 84180 0 -1 109344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1082
timestamp 1624015447
transform 1 0 84180 0 1 109344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1084
timestamp 1624015447
transform 1 0 84180 0 -1 110432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_196_906
timestamp 1624015447
transform 1 0 84456 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_906
timestamp 1624015447
transform 1 0 84456 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_906
timestamp 1624015447
transform 1 0 84456 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_918
timestamp 1624015447
transform 1 0 85560 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_918
timestamp 1624015447
transform 1 0 85560 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_918
timestamp 1624015447
transform 1 0 85560 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_945
timestamp 1624015447
transform 1 0 88044 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_933
timestamp 1624015447
transform 1 0 86940 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_196_930
timestamp 1624015447
transform 1 0 86664 0 -1 109344
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1746
timestamp 1624015447
transform 1 0 86848 0 -1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_197_942
timestamp 1624015447
transform 1 0 87768 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_930
timestamp 1624015447
transform 1 0 86664 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_945
timestamp 1624015447
transform 1 0 88044 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_933
timestamp 1624015447
transform 1 0 86940 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_198_930
timestamp 1624015447
transform 1 0 86664 0 -1 110432
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1748
timestamp 1624015447
transform 1 0 86848 0 -1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1747
timestamp 1624015447
transform 1 0 89424 0 1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_196_957
timestamp 1624015447
transform 1 0 89148 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_197_954
timestamp 1624015447
transform 1 0 88872 0 1 109344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_197_961
timestamp 1624015447
transform 1 0 89516 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_957
timestamp 1624015447
transform 1 0 89148 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1081
timestamp 1624015447
transform -1 0 90896 0 -1 109344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1083
timestamp 1624015447
transform -1 0 90896 0 1 109344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1085
timestamp 1624015447
transform -1 0 90896 0 -1 110432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_196_969
timestamp 1624015447
transform 1 0 90252 0 -1 109344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_198_969
timestamp 1624015447
transform 1 0 90252 0 -1 110432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_396
timestamp 1624015447
transform 1 0 1104 0 1 110432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_398
timestamp 1624015447
transform 1 0 1104 0 -1 111520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_400
timestamp 1624015447
transform 1 0 1104 0 1 111520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_199_3
timestamp 1624015447
transform 1 0 1380 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_15
timestamp 1624015447
transform 1 0 2484 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_3
timestamp 1624015447
transform 1 0 1380 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_15
timestamp 1624015447
transform 1 0 2484 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_3
timestamp 1624015447
transform 1 0 1380 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_15
timestamp 1624015447
transform 1 0 2484 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1475
timestamp 1624015447
transform 1 0 3772 0 -1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_199_27
timestamp 1624015447
transform 1 0 3588 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_200_27
timestamp 1624015447
transform 1 0 3588 0 -1 111520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_200_30
timestamp 1624015447
transform 1 0 3864 0 -1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_201_27
timestamp 1624015447
transform 1 0 3588 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_397
timestamp 1624015447
transform -1 0 5152 0 1 110432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_399
timestamp 1624015447
transform -1 0 5152 0 -1 111520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_401
timestamp 1624015447
transform -1 0 5152 0 1 111520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_199_39
timestamp 1624015447
transform 1 0 4692 0 1 110432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_200_38
timestamp 1624015447
transform 1 0 4600 0 -1 111520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_201_39
timestamp 1624015447
transform 1 0 4692 0 1 111520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1086
timestamp 1624015447
transform 1 0 84180 0 1 110432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1088
timestamp 1624015447
transform 1 0 84180 0 -1 111520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1090
timestamp 1624015447
transform 1 0 84180 0 1 111520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_199_906
timestamp 1624015447
transform 1 0 84456 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_906
timestamp 1624015447
transform 1 0 84456 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_906
timestamp 1624015447
transform 1 0 84456 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_918
timestamp 1624015447
transform 1 0 85560 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_918
timestamp 1624015447
transform 1 0 85560 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_918
timestamp 1624015447
transform 1 0 85560 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1750
timestamp 1624015447
transform 1 0 86848 0 -1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_199_930
timestamp 1624015447
transform 1 0 86664 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_942
timestamp 1624015447
transform 1 0 87768 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_200_930
timestamp 1624015447
transform 1 0 86664 0 -1 111520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_200_933
timestamp 1624015447
transform 1 0 86940 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_945
timestamp 1624015447
transform 1 0 88044 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_930
timestamp 1624015447
transform 1 0 86664 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_942
timestamp 1624015447
transform 1 0 87768 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1749
timestamp 1624015447
transform 1 0 89424 0 1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1751
timestamp 1624015447
transform 1 0 89424 0 1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_199_954
timestamp 1624015447
transform 1 0 88872 0 1 110432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_199_961
timestamp 1624015447
transform 1 0 89516 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_957
timestamp 1624015447
transform 1 0 89148 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_201_954
timestamp 1624015447
transform 1 0 88872 0 1 111520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_201_961
timestamp 1624015447
transform 1 0 89516 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1087
timestamp 1624015447
transform -1 0 90896 0 1 110432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1089
timestamp 1624015447
transform -1 0 90896 0 -1 111520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1091
timestamp 1624015447
transform -1 0 90896 0 1 111520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_200_969
timestamp 1624015447
transform 1 0 90252 0 -1 111520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_402
timestamp 1624015447
transform 1 0 1104 0 -1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_404
timestamp 1624015447
transform 1 0 1104 0 1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_406
timestamp 1624015447
transform 1 0 1104 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_202_3
timestamp 1624015447
transform 1 0 1380 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_15
timestamp 1624015447
transform 1 0 2484 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_3
timestamp 1624015447
transform 1 0 1380 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_15
timestamp 1624015447
transform 1 0 2484 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_3
timestamp 1624015447
transform 1 0 1380 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_15
timestamp 1624015447
transform 1 0 2484 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1476
timestamp 1624015447
transform 1 0 3772 0 -1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1477
timestamp 1624015447
transform 1 0 3772 0 -1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_202_27
timestamp 1624015447
transform 1 0 3588 0 -1 112608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_202_30
timestamp 1624015447
transform 1 0 3864 0 -1 112608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_203_27
timestamp 1624015447
transform 1 0 3588 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_204_27
timestamp 1624015447
transform 1 0 3588 0 -1 113696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_204_30
timestamp 1624015447
transform 1 0 3864 0 -1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_403
timestamp 1624015447
transform -1 0 5152 0 -1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_405
timestamp 1624015447
transform -1 0 5152 0 1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_407
timestamp 1624015447
transform -1 0 5152 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_202_38
timestamp 1624015447
transform 1 0 4600 0 -1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_203_39
timestamp 1624015447
transform 1 0 4692 0 1 112608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_204_38
timestamp 1624015447
transform 1 0 4600 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1092
timestamp 1624015447
transform 1 0 84180 0 -1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1094
timestamp 1624015447
transform 1 0 84180 0 1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1096
timestamp 1624015447
transform 1 0 84180 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_202_906
timestamp 1624015447
transform 1 0 84456 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_906
timestamp 1624015447
transform 1 0 84456 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_906
timestamp 1624015447
transform 1 0 84456 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_918
timestamp 1624015447
transform 1 0 85560 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_918
timestamp 1624015447
transform 1 0 85560 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_918
timestamp 1624015447
transform 1 0 85560 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_945
timestamp 1624015447
transform 1 0 88044 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_933
timestamp 1624015447
transform 1 0 86940 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_202_930
timestamp 1624015447
transform 1 0 86664 0 -1 112608
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1752
timestamp 1624015447
transform 1 0 86848 0 -1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_204_945
timestamp 1624015447
transform 1 0 88044 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_933
timestamp 1624015447
transform 1 0 86940 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_204_930
timestamp 1624015447
transform 1 0 86664 0 -1 113696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_203_942
timestamp 1624015447
transform 1 0 87768 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_930
timestamp 1624015447
transform 1 0 86664 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1754
timestamp 1624015447
transform 1 0 86848 0 -1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1753
timestamp 1624015447
transform 1 0 89424 0 1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_202_957
timestamp 1624015447
transform 1 0 89148 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_203_954
timestamp 1624015447
transform 1 0 88872 0 1 112608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_203_961
timestamp 1624015447
transform 1 0 89516 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_957
timestamp 1624015447
transform 1 0 89148 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1093
timestamp 1624015447
transform -1 0 90896 0 -1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1095
timestamp 1624015447
transform -1 0 90896 0 1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1097
timestamp 1624015447
transform -1 0 90896 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_202_969
timestamp 1624015447
transform 1 0 90252 0 -1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_204_969
timestamp 1624015447
transform 1 0 90252 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_408
timestamp 1624015447
transform 1 0 1104 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_410
timestamp 1624015447
transform 1 0 1104 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_412
timestamp 1624015447
transform 1 0 1104 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_205_3
timestamp 1624015447
transform 1 0 1380 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_15
timestamp 1624015447
transform 1 0 2484 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_3
timestamp 1624015447
transform 1 0 1380 0 -1 114784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_15
timestamp 1624015447
transform 1 0 2484 0 -1 114784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_3
timestamp 1624015447
transform 1 0 1380 0 1 114784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_15
timestamp 1624015447
transform 1 0 2484 0 1 114784
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1478
timestamp 1624015447
transform 1 0 3772 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_205_27
timestamp 1624015447
transform 1 0 3588 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_206_27
timestamp 1624015447
transform 1 0 3588 0 -1 114784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_206_30
timestamp 1624015447
transform 1 0 3864 0 -1 114784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_207_27
timestamp 1624015447
transform 1 0 3588 0 1 114784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_409
timestamp 1624015447
transform -1 0 5152 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_411
timestamp 1624015447
transform -1 0 5152 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_413
timestamp 1624015447
transform -1 0 5152 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_csb0
timestamp 1624015447
transform -1 0 4876 0 1 114784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_205_39
timestamp 1624015447
transform 1 0 4692 0 1 113696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_206_38
timestamp 1624015447
transform 1 0 4600 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1098
timestamp 1624015447
transform 1 0 84180 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1100
timestamp 1624015447
transform 1 0 84180 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1102
timestamp 1624015447
transform 1 0 84180 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_205_906
timestamp 1624015447
transform 1 0 84456 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_906
timestamp 1624015447
transform 1 0 84456 0 -1 114784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_906
timestamp 1624015447
transform 1 0 84456 0 1 114784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_918
timestamp 1624015447
transform 1 0 85560 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_918
timestamp 1624015447
transform 1 0 85560 0 -1 114784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_918
timestamp 1624015447
transform 1 0 85560 0 1 114784
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1756
timestamp 1624015447
transform 1 0 86848 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_205_930
timestamp 1624015447
transform 1 0 86664 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_942
timestamp 1624015447
transform 1 0 87768 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_206_930
timestamp 1624015447
transform 1 0 86664 0 -1 114784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_206_933
timestamp 1624015447
transform 1 0 86940 0 -1 114784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_945
timestamp 1624015447
transform 1 0 88044 0 -1 114784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_930
timestamp 1624015447
transform 1 0 86664 0 1 114784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_942
timestamp 1624015447
transform 1 0 87768 0 1 114784
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1755
timestamp 1624015447
transform 1 0 89424 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1757
timestamp 1624015447
transform 1 0 89424 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_205_954
timestamp 1624015447
transform 1 0 88872 0 1 113696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_205_961
timestamp 1624015447
transform 1 0 89516 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_957
timestamp 1624015447
transform 1 0 89148 0 -1 114784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_207_954
timestamp 1624015447
transform 1 0 88872 0 1 114784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_207_961
timestamp 1624015447
transform 1 0 89516 0 1 114784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1099
timestamp 1624015447
transform -1 0 90896 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1101
timestamp 1624015447
transform -1 0 90896 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1103
timestamp 1624015447
transform -1 0 90896 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_206_969
timestamp 1624015447
transform 1 0 90252 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_414
timestamp 1624015447
transform 1 0 1104 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_416
timestamp 1624015447
transform 1 0 1104 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_418
timestamp 1624015447
transform 1 0 1104 0 -1 116960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_208_3
timestamp 1624015447
transform 1 0 1380 0 -1 115872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_15
timestamp 1624015447
transform 1 0 2484 0 -1 115872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_3
timestamp 1624015447
transform 1 0 1380 0 1 115872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_15
timestamp 1624015447
transform 1 0 2484 0 1 115872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_3
timestamp 1624015447
transform 1 0 1380 0 -1 116960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_15
timestamp 1624015447
transform 1 0 2484 0 -1 116960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1479
timestamp 1624015447
transform 1 0 3772 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1480
timestamp 1624015447
transform 1 0 3772 0 -1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_208_27
timestamp 1624015447
transform 1 0 3588 0 -1 115872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_208_30
timestamp 1624015447
transform 1 0 3864 0 -1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_209_27
timestamp 1624015447
transform 1 0 3588 0 1 115872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_210_27
timestamp 1624015447
transform 1 0 3588 0 -1 116960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_210_30
timestamp 1624015447
transform 1 0 3864 0 -1 116960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_415
timestamp 1624015447
transform -1 0 5152 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_417
timestamp 1624015447
transform -1 0 5152 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_419
timestamp 1624015447
transform -1 0 5152 0 -1 116960
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_web0
timestamp 1624015447
transform -1 0 4876 0 -1 116960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_208_38
timestamp 1624015447
transform 1 0 4600 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_209_39
timestamp 1624015447
transform 1 0 4692 0 1 115872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_210_38
timestamp 1624015447
transform 1 0 4600 0 -1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1104
timestamp 1624015447
transform 1 0 84180 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1106
timestamp 1624015447
transform 1 0 84180 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1108
timestamp 1624015447
transform 1 0 84180 0 -1 116960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_208_906
timestamp 1624015447
transform 1 0 84456 0 -1 115872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_906
timestamp 1624015447
transform 1 0 84456 0 1 115872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_906
timestamp 1624015447
transform 1 0 84456 0 -1 116960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_918
timestamp 1624015447
transform 1 0 85560 0 -1 115872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_918
timestamp 1624015447
transform 1 0 85560 0 1 115872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_918
timestamp 1624015447
transform 1 0 85560 0 -1 116960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_945
timestamp 1624015447
transform 1 0 88044 0 -1 115872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_933
timestamp 1624015447
transform 1 0 86940 0 -1 115872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_208_930
timestamp 1624015447
transform 1 0 86664 0 -1 115872
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1758
timestamp 1624015447
transform 1 0 86848 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_210_945
timestamp 1624015447
transform 1 0 88044 0 -1 116960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_933
timestamp 1624015447
transform 1 0 86940 0 -1 116960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_210_930
timestamp 1624015447
transform 1 0 86664 0 -1 116960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_209_942
timestamp 1624015447
transform 1 0 87768 0 1 115872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_930
timestamp 1624015447
transform 1 0 86664 0 1 115872
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1760
timestamp 1624015447
transform 1 0 86848 0 -1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1759
timestamp 1624015447
transform 1 0 89424 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_208_957
timestamp 1624015447
transform 1 0 89148 0 -1 115872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_209_954
timestamp 1624015447
transform 1 0 88872 0 1 115872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_209_961
timestamp 1624015447
transform 1 0 89516 0 1 115872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_957
timestamp 1624015447
transform 1 0 89148 0 -1 116960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1105
timestamp 1624015447
transform -1 0 90896 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1107
timestamp 1624015447
transform -1 0 90896 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1109
timestamp 1624015447
transform -1 0 90896 0 -1 116960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_208_969
timestamp 1624015447
transform 1 0 90252 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_969
timestamp 1624015447
transform 1 0 90252 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_420
timestamp 1624015447
transform 1 0 1104 0 1 116960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_422
timestamp 1624015447
transform 1 0 1104 0 -1 118048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_424
timestamp 1624015447
transform 1 0 1104 0 1 118048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_211_3
timestamp 1624015447
transform 1 0 1380 0 1 116960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_211_15
timestamp 1624015447
transform 1 0 2484 0 1 116960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_212_3
timestamp 1624015447
transform 1 0 1380 0 -1 118048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_212_15
timestamp 1624015447
transform 1 0 2484 0 -1 118048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_213_3
timestamp 1624015447
transform 1 0 1380 0 1 118048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_213_15
timestamp 1624015447
transform 1 0 2484 0 1 118048
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1481
timestamp 1624015447
transform 1 0 3772 0 -1 118048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_211_27
timestamp 1624015447
transform 1 0 3588 0 1 116960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_212_27
timestamp 1624015447
transform 1 0 3588 0 -1 118048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_212_30
timestamp 1624015447
transform 1 0 3864 0 -1 118048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_213_27
timestamp 1624015447
transform 1 0 3588 0 1 118048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_421
timestamp 1624015447
transform -1 0 5152 0 1 116960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_423
timestamp 1624015447
transform -1 0 5152 0 -1 118048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_425
timestamp 1624015447
transform -1 0 5152 0 1 118048
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_211_39
timestamp 1624015447
transform 1 0 4692 0 1 116960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_212_38
timestamp 1624015447
transform 1 0 4600 0 -1 118048
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_213_39
timestamp 1624015447
transform 1 0 4692 0 1 118048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_212_906
timestamp 1624015447
transform 1 0 84456 0 -1 118048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_211_910
timestamp 1624015447
transform 1 0 84824 0 1 116960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_211_906
timestamp 1624015447
transform 1 0 84456 0 1 116960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_addr1[7]
timestamp 1624015447
transform -1 0 84824 0 1 116960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1112
timestamp 1624015447
transform 1 0 84180 0 -1 118048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1110
timestamp 1624015447
transform 1 0 84180 0 1 116960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_213_910
timestamp 1624015447
transform 1 0 84824 0 1 118048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_213_906
timestamp 1624015447
transform 1 0 84456 0 1 118048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_addr1[6]
timestamp 1624015447
transform -1 0 84824 0 1 118048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1114
timestamp 1624015447
transform 1 0 84180 0 1 118048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_211_922
timestamp 1624015447
transform 1 0 85928 0 1 116960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_212_918
timestamp 1624015447
transform 1 0 85560 0 -1 118048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_213_922
timestamp 1624015447
transform 1 0 85928 0 1 118048
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1762
timestamp 1624015447
transform 1 0 86848 0 -1 118048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_211_934
timestamp 1624015447
transform 1 0 87032 0 1 116960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_211_946
timestamp 1624015447
transform 1 0 88136 0 1 116960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_212_930
timestamp 1624015447
transform 1 0 86664 0 -1 118048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_212_933
timestamp 1624015447
transform 1 0 86940 0 -1 118048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_212_945
timestamp 1624015447
transform 1 0 88044 0 -1 118048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_213_934
timestamp 1624015447
transform 1 0 87032 0 1 118048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_213_946
timestamp 1624015447
transform 1 0 88136 0 1 118048
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1761
timestamp 1624015447
transform 1 0 89424 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1763
timestamp 1624015447
transform 1 0 89424 0 1 118048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_211_958
timestamp 1624015447
transform 1 0 89240 0 1 116960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_211_961
timestamp 1624015447
transform 1 0 89516 0 1 116960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_212_957
timestamp 1624015447
transform 1 0 89148 0 -1 118048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_213_958
timestamp 1624015447
transform 1 0 89240 0 1 118048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_213_961
timestamp 1624015447
transform 1 0 89516 0 1 118048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1111
timestamp 1624015447
transform -1 0 90896 0 1 116960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1113
timestamp 1624015447
transform -1 0 90896 0 -1 118048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1115
timestamp 1624015447
transform -1 0 90896 0 1 118048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_212_969
timestamp 1624015447
transform 1 0 90252 0 -1 118048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_215_15
timestamp 1624015447
transform 1 0 2484 0 1 119136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_215_3
timestamp 1624015447
transform 1 0 1380 0 1 119136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_214_15
timestamp 1624015447
transform 1 0 2484 0 -1 119136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_214_3
timestamp 1624015447
transform 1 0 1380 0 -1 119136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_428
timestamp 1624015447
transform 1 0 1104 0 1 119136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_426
timestamp 1624015447
transform 1 0 1104 0 -1 119136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_216_15
timestamp 1624015447
transform 1 0 2484 0 -1 120224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_216_3
timestamp 1624015447
transform 1 0 1380 0 -1 120224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_430
timestamp 1624015447
transform 1 0 1104 0 -1 120224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_217_15
timestamp 1624015447
transform 1 0 2484 0 1 120224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_217_3
timestamp 1624015447
transform 1 0 1380 0 1 120224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_432
timestamp 1624015447
transform 1 0 1104 0 1 120224
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1482
timestamp 1624015447
transform 1 0 3772 0 -1 119136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1483
timestamp 1624015447
transform 1 0 3772 0 -1 120224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_214_27
timestamp 1624015447
transform 1 0 3588 0 -1 119136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_214_30
timestamp 1624015447
transform 1 0 3864 0 -1 119136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_215_27
timestamp 1624015447
transform 1 0 3588 0 1 119136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_216_27
timestamp 1624015447
transform 1 0 3588 0 -1 120224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_216_30
timestamp 1624015447
transform 1 0 3864 0 -1 120224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_217_27
timestamp 1624015447
transform 1 0 3588 0 1 120224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_427
timestamp 1624015447
transform -1 0 5152 0 -1 119136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_429
timestamp 1624015447
transform -1 0 5152 0 1 119136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_431
timestamp 1624015447
transform -1 0 5152 0 -1 120224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_433
timestamp 1624015447
transform -1 0 5152 0 1 120224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_214_38
timestamp 1624015447
transform 1 0 4600 0 -1 119136
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_215_39
timestamp 1624015447
transform 1 0 4692 0 1 119136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_216_38
timestamp 1624015447
transform 1 0 4600 0 -1 120224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_217_39
timestamp 1624015447
transform 1 0 4692 0 1 120224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_215_906
timestamp 1624015447
transform 1 0 84456 0 1 119136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_214_906
timestamp 1624015447
transform 1 0 84456 0 -1 119136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1118
timestamp 1624015447
transform 1 0 84180 0 1 119136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1116
timestamp 1624015447
transform 1 0 84180 0 -1 119136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_216_910
timestamp 1624015447
transform 1 0 84824 0 -1 120224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_216_906
timestamp 1624015447
transform 1 0 84456 0 -1 120224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_addr1[5]
timestamp 1624015447
transform -1 0 84824 0 -1 120224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1120
timestamp 1624015447
transform 1 0 84180 0 -1 120224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_217_906
timestamp 1624015447
transform 1 0 84456 0 1 120224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1122
timestamp 1624015447
transform 1 0 84180 0 1 120224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_214_918
timestamp 1624015447
transform 1 0 85560 0 -1 119136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_215_918
timestamp 1624015447
transform 1 0 85560 0 1 119136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_216_922
timestamp 1624015447
transform 1 0 85928 0 -1 120224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_217_918
timestamp 1624015447
transform 1 0 85560 0 1 120224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_215_942
timestamp 1624015447
transform 1 0 87768 0 1 119136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_215_930
timestamp 1624015447
transform 1 0 86664 0 1 119136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_214_945
timestamp 1624015447
transform 1 0 88044 0 -1 119136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_214_933
timestamp 1624015447
transform 1 0 86940 0 -1 119136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_214_930
timestamp 1624015447
transform 1 0 86664 0 -1 119136
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1764
timestamp 1624015447
transform 1 0 86848 0 -1 119136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_216_945
timestamp 1624015447
transform 1 0 88044 0 -1 120224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_216_933
timestamp 1624015447
transform 1 0 86940 0 -1 120224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_216_930
timestamp 1624015447
transform 1 0 86664 0 -1 120224
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1766
timestamp 1624015447
transform 1 0 86848 0 -1 120224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_217_942
timestamp 1624015447
transform 1 0 87768 0 1 120224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_217_930
timestamp 1624015447
transform 1 0 86664 0 1 120224
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1765
timestamp 1624015447
transform 1 0 89424 0 1 119136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1767
timestamp 1624015447
transform 1 0 89424 0 1 120224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_214_957
timestamp 1624015447
transform 1 0 89148 0 -1 119136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_215_954
timestamp 1624015447
transform 1 0 88872 0 1 119136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_215_961
timestamp 1624015447
transform 1 0 89516 0 1 119136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_216_957
timestamp 1624015447
transform 1 0 89148 0 -1 120224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_217_954
timestamp 1624015447
transform 1 0 88872 0 1 120224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_217_961
timestamp 1624015447
transform 1 0 89516 0 1 120224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1117
timestamp 1624015447
transform -1 0 90896 0 -1 119136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1119
timestamp 1624015447
transform -1 0 90896 0 1 119136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1121
timestamp 1624015447
transform -1 0 90896 0 -1 120224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1123
timestamp 1624015447
transform -1 0 90896 0 1 120224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_214_969
timestamp 1624015447
transform 1 0 90252 0 -1 119136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_216_969
timestamp 1624015447
transform 1 0 90252 0 -1 120224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_434
timestamp 1624015447
transform 1 0 1104 0 -1 121312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_436
timestamp 1624015447
transform 1 0 1104 0 1 121312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_438
timestamp 1624015447
transform 1 0 1104 0 -1 122400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_218_3
timestamp 1624015447
transform 1 0 1380 0 -1 121312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_218_15
timestamp 1624015447
transform 1 0 2484 0 -1 121312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_219_3
timestamp 1624015447
transform 1 0 1380 0 1 121312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_219_15
timestamp 1624015447
transform 1 0 2484 0 1 121312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_220_3
timestamp 1624015447
transform 1 0 1380 0 -1 122400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_220_15
timestamp 1624015447
transform 1 0 2484 0 -1 122400
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1484
timestamp 1624015447
transform 1 0 3772 0 -1 121312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1485
timestamp 1624015447
transform 1 0 3772 0 -1 122400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_218_27
timestamp 1624015447
transform 1 0 3588 0 -1 121312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_218_30
timestamp 1624015447
transform 1 0 3864 0 -1 121312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_219_27
timestamp 1624015447
transform 1 0 3588 0 1 121312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_220_27
timestamp 1624015447
transform 1 0 3588 0 -1 122400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_220_30
timestamp 1624015447
transform 1 0 3864 0 -1 122400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_435
timestamp 1624015447
transform -1 0 5152 0 -1 121312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_437
timestamp 1624015447
transform -1 0 5152 0 1 121312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_439
timestamp 1624015447
transform -1 0 5152 0 -1 122400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_218_38
timestamp 1624015447
transform 1 0 4600 0 -1 121312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_219_39
timestamp 1624015447
transform 1 0 4692 0 1 121312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_220_38
timestamp 1624015447
transform 1 0 4600 0 -1 122400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1124
timestamp 1624015447
transform 1 0 84180 0 -1 121312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1126
timestamp 1624015447
transform 1 0 84180 0 1 121312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1128
timestamp 1624015447
transform 1 0 84180 0 -1 122400
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_addr1[4]
timestamp 1624015447
transform -1 0 84824 0 -1 121312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_218_906
timestamp 1624015447
transform 1 0 84456 0 -1 121312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_218_910
timestamp 1624015447
transform 1 0 84824 0 -1 121312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_219_906
timestamp 1624015447
transform 1 0 84456 0 1 121312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_220_906
timestamp 1624015447
transform 1 0 84456 0 -1 122400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_218_922
timestamp 1624015447
transform 1 0 85928 0 -1 121312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_219_918
timestamp 1624015447
transform 1 0 85560 0 1 121312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_220_918
timestamp 1624015447
transform 1 0 85560 0 -1 122400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_218_945
timestamp 1624015447
transform 1 0 88044 0 -1 121312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_218_933
timestamp 1624015447
transform 1 0 86940 0 -1 121312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_218_930
timestamp 1624015447
transform 1 0 86664 0 -1 121312
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1768
timestamp 1624015447
transform 1 0 86848 0 -1 121312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_219_942
timestamp 1624015447
transform 1 0 87768 0 1 121312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_219_930
timestamp 1624015447
transform 1 0 86664 0 1 121312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_220_945
timestamp 1624015447
transform 1 0 88044 0 -1 122400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_220_933
timestamp 1624015447
transform 1 0 86940 0 -1 122400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_220_930
timestamp 1624015447
transform 1 0 86664 0 -1 122400
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1770
timestamp 1624015447
transform 1 0 86848 0 -1 122400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1769
timestamp 1624015447
transform 1 0 89424 0 1 121312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_218_957
timestamp 1624015447
transform 1 0 89148 0 -1 121312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_219_954
timestamp 1624015447
transform 1 0 88872 0 1 121312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_219_961
timestamp 1624015447
transform 1 0 89516 0 1 121312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_220_957
timestamp 1624015447
transform 1 0 89148 0 -1 122400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1125
timestamp 1624015447
transform -1 0 90896 0 -1 121312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1127
timestamp 1624015447
transform -1 0 90896 0 1 121312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1129
timestamp 1624015447
transform -1 0 90896 0 -1 122400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_218_969
timestamp 1624015447
transform 1 0 90252 0 -1 121312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_220_969
timestamp 1624015447
transform 1 0 90252 0 -1 122400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_440
timestamp 1624015447
transform 1 0 1104 0 1 122400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_442
timestamp 1624015447
transform 1 0 1104 0 -1 123488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_444
timestamp 1624015447
transform 1 0 1104 0 1 123488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_221_3
timestamp 1624015447
transform 1 0 1380 0 1 122400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_221_15
timestamp 1624015447
transform 1 0 2484 0 1 122400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_222_3
timestamp 1624015447
transform 1 0 1380 0 -1 123488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_222_15
timestamp 1624015447
transform 1 0 2484 0 -1 123488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_223_3
timestamp 1624015447
transform 1 0 1380 0 1 123488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_223_15
timestamp 1624015447
transform 1 0 2484 0 1 123488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1486
timestamp 1624015447
transform 1 0 3772 0 -1 123488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_221_27
timestamp 1624015447
transform 1 0 3588 0 1 122400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_222_27
timestamp 1624015447
transform 1 0 3588 0 -1 123488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_222_30
timestamp 1624015447
transform 1 0 3864 0 -1 123488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_223_27
timestamp 1624015447
transform 1 0 3588 0 1 123488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_441
timestamp 1624015447
transform -1 0 5152 0 1 122400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_443
timestamp 1624015447
transform -1 0 5152 0 -1 123488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_445
timestamp 1624015447
transform -1 0 5152 0 1 123488
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_221_39
timestamp 1624015447
transform 1 0 4692 0 1 122400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_222_38
timestamp 1624015447
transform 1 0 4600 0 -1 123488
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_223_39
timestamp 1624015447
transform 1 0 4692 0 1 123488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1130
timestamp 1624015447
transform 1 0 84180 0 1 122400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1132
timestamp 1624015447
transform 1 0 84180 0 -1 123488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1134
timestamp 1624015447
transform 1 0 84180 0 1 123488
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_addr1[3]
timestamp 1624015447
transform -1 0 84824 0 -1 123488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_221_906
timestamp 1624015447
transform 1 0 84456 0 1 122400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_222_906
timestamp 1624015447
transform 1 0 84456 0 -1 123488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_222_910
timestamp 1624015447
transform 1 0 84824 0 -1 123488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_223_906
timestamp 1624015447
transform 1 0 84456 0 1 123488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_221_918
timestamp 1624015447
transform 1 0 85560 0 1 122400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_222_922
timestamp 1624015447
transform 1 0 85928 0 -1 123488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_223_918
timestamp 1624015447
transform 1 0 85560 0 1 123488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1772
timestamp 1624015447
transform 1 0 86848 0 -1 123488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_221_930
timestamp 1624015447
transform 1 0 86664 0 1 122400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_221_942
timestamp 1624015447
transform 1 0 87768 0 1 122400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_222_930
timestamp 1624015447
transform 1 0 86664 0 -1 123488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_222_933
timestamp 1624015447
transform 1 0 86940 0 -1 123488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_222_945
timestamp 1624015447
transform 1 0 88044 0 -1 123488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_223_930
timestamp 1624015447
transform 1 0 86664 0 1 123488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_223_942
timestamp 1624015447
transform 1 0 87768 0 1 123488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1771
timestamp 1624015447
transform 1 0 89424 0 1 122400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1773
timestamp 1624015447
transform 1 0 89424 0 1 123488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_221_954
timestamp 1624015447
transform 1 0 88872 0 1 122400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_221_961
timestamp 1624015447
transform 1 0 89516 0 1 122400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_222_957
timestamp 1624015447
transform 1 0 89148 0 -1 123488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_223_954
timestamp 1624015447
transform 1 0 88872 0 1 123488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_223_961
timestamp 1624015447
transform 1 0 89516 0 1 123488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1131
timestamp 1624015447
transform -1 0 90896 0 1 122400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1133
timestamp 1624015447
transform -1 0 90896 0 -1 123488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1135
timestamp 1624015447
transform -1 0 90896 0 1 123488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_222_969
timestamp 1624015447
transform 1 0 90252 0 -1 123488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_446
timestamp 1624015447
transform 1 0 1104 0 -1 124576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_448
timestamp 1624015447
transform 1 0 1104 0 1 124576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_450
timestamp 1624015447
transform 1 0 1104 0 -1 125664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_224_3
timestamp 1624015447
transform 1 0 1380 0 -1 124576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_224_15
timestamp 1624015447
transform 1 0 2484 0 -1 124576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_225_3
timestamp 1624015447
transform 1 0 1380 0 1 124576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_225_15
timestamp 1624015447
transform 1 0 2484 0 1 124576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_226_3
timestamp 1624015447
transform 1 0 1380 0 -1 125664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_226_15
timestamp 1624015447
transform 1 0 2484 0 -1 125664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1487
timestamp 1624015447
transform 1 0 3772 0 -1 124576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1488
timestamp 1624015447
transform 1 0 3772 0 -1 125664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_224_27
timestamp 1624015447
transform 1 0 3588 0 -1 124576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_224_30
timestamp 1624015447
transform 1 0 3864 0 -1 124576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_225_27
timestamp 1624015447
transform 1 0 3588 0 1 124576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_226_27
timestamp 1624015447
transform 1 0 3588 0 -1 125664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_226_30
timestamp 1624015447
transform 1 0 3864 0 -1 125664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_447
timestamp 1624015447
transform -1 0 5152 0 -1 124576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_449
timestamp 1624015447
transform -1 0 5152 0 1 124576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_451
timestamp 1624015447
transform -1 0 5152 0 -1 125664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_224_38
timestamp 1624015447
transform 1 0 4600 0 -1 124576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_225_39
timestamp 1624015447
transform 1 0 4692 0 1 124576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_226_38
timestamp 1624015447
transform 1 0 4600 0 -1 125664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1136
timestamp 1624015447
transform 1 0 84180 0 -1 124576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1138
timestamp 1624015447
transform 1 0 84180 0 1 124576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1140
timestamp 1624015447
transform 1 0 84180 0 -1 125664
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_addr1[2]
timestamp 1624015447
transform -1 0 84824 0 -1 124576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_224_906
timestamp 1624015447
transform 1 0 84456 0 -1 124576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_224_910
timestamp 1624015447
transform 1 0 84824 0 -1 124576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_225_906
timestamp 1624015447
transform 1 0 84456 0 1 124576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_226_906
timestamp 1624015447
transform 1 0 84456 0 -1 125664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_224_922
timestamp 1624015447
transform 1 0 85928 0 -1 124576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_225_918
timestamp 1624015447
transform 1 0 85560 0 1 124576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_226_918
timestamp 1624015447
transform 1 0 85560 0 -1 125664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_224_945
timestamp 1624015447
transform 1 0 88044 0 -1 124576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_224_933
timestamp 1624015447
transform 1 0 86940 0 -1 124576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_224_930
timestamp 1624015447
transform 1 0 86664 0 -1 124576
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1774
timestamp 1624015447
transform 1 0 86848 0 -1 124576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_225_942
timestamp 1624015447
transform 1 0 87768 0 1 124576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_225_930
timestamp 1624015447
transform 1 0 86664 0 1 124576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_226_945
timestamp 1624015447
transform 1 0 88044 0 -1 125664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_226_933
timestamp 1624015447
transform 1 0 86940 0 -1 125664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_226_930
timestamp 1624015447
transform 1 0 86664 0 -1 125664
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1776
timestamp 1624015447
transform 1 0 86848 0 -1 125664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1775
timestamp 1624015447
transform 1 0 89424 0 1 124576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_224_957
timestamp 1624015447
transform 1 0 89148 0 -1 124576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_225_954
timestamp 1624015447
transform 1 0 88872 0 1 124576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_225_961
timestamp 1624015447
transform 1 0 89516 0 1 124576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_226_957
timestamp 1624015447
transform 1 0 89148 0 -1 125664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1137
timestamp 1624015447
transform -1 0 90896 0 -1 124576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1139
timestamp 1624015447
transform -1 0 90896 0 1 124576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1141
timestamp 1624015447
transform -1 0 90896 0 -1 125664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_224_969
timestamp 1624015447
transform 1 0 90252 0 -1 124576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_226_969
timestamp 1624015447
transform 1 0 90252 0 -1 125664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_452
timestamp 1624015447
transform 1 0 1104 0 1 125664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_454
timestamp 1624015447
transform 1 0 1104 0 -1 126752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_456
timestamp 1624015447
transform 1 0 1104 0 1 126752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_227_3
timestamp 1624015447
transform 1 0 1380 0 1 125664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_227_15
timestamp 1624015447
transform 1 0 2484 0 1 125664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_228_3
timestamp 1624015447
transform 1 0 1380 0 -1 126752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_228_15
timestamp 1624015447
transform 1 0 2484 0 -1 126752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_229_3
timestamp 1624015447
transform 1 0 1380 0 1 126752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_229_15
timestamp 1624015447
transform 1 0 2484 0 1 126752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1489
timestamp 1624015447
transform 1 0 3772 0 -1 126752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_227_27
timestamp 1624015447
transform 1 0 3588 0 1 125664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_228_27
timestamp 1624015447
transform 1 0 3588 0 -1 126752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_228_30
timestamp 1624015447
transform 1 0 3864 0 -1 126752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_229_27
timestamp 1624015447
transform 1 0 3588 0 1 126752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_453
timestamp 1624015447
transform -1 0 5152 0 1 125664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_455
timestamp 1624015447
transform -1 0 5152 0 -1 126752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_457
timestamp 1624015447
transform -1 0 5152 0 1 126752
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_227_39
timestamp 1624015447
transform 1 0 4692 0 1 125664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_228_38
timestamp 1624015447
transform 1 0 4600 0 -1 126752
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_229_39
timestamp 1624015447
transform 1 0 4692 0 1 126752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1142
timestamp 1624015447
transform 1 0 84180 0 1 125664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1144
timestamp 1624015447
transform 1 0 84180 0 -1 126752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1146
timestamp 1624015447
transform 1 0 84180 0 1 126752
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_addr1[1]
timestamp 1624015447
transform -1 0 84824 0 1 125664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_227_906
timestamp 1624015447
transform 1 0 84456 0 1 125664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_227_910
timestamp 1624015447
transform 1 0 84824 0 1 125664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_228_906
timestamp 1624015447
transform 1 0 84456 0 -1 126752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_229_906
timestamp 1624015447
transform 1 0 84456 0 1 126752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_227_922
timestamp 1624015447
transform 1 0 85928 0 1 125664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_228_918
timestamp 1624015447
transform 1 0 85560 0 -1 126752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_229_918
timestamp 1624015447
transform 1 0 85560 0 1 126752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1778
timestamp 1624015447
transform 1 0 86848 0 -1 126752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_227_934
timestamp 1624015447
transform 1 0 87032 0 1 125664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_227_946
timestamp 1624015447
transform 1 0 88136 0 1 125664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_228_930
timestamp 1624015447
transform 1 0 86664 0 -1 126752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_228_933
timestamp 1624015447
transform 1 0 86940 0 -1 126752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_228_945
timestamp 1624015447
transform 1 0 88044 0 -1 126752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_229_930
timestamp 1624015447
transform 1 0 86664 0 1 126752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_229_942
timestamp 1624015447
transform 1 0 87768 0 1 126752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1777
timestamp 1624015447
transform 1 0 89424 0 1 125664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1779
timestamp 1624015447
transform 1 0 89424 0 1 126752
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_227_958
timestamp 1624015447
transform 1 0 89240 0 1 125664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_227_961
timestamp 1624015447
transform 1 0 89516 0 1 125664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_228_957
timestamp 1624015447
transform 1 0 89148 0 -1 126752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_229_954
timestamp 1624015447
transform 1 0 88872 0 1 126752
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_229_961
timestamp 1624015447
transform 1 0 89516 0 1 126752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1143
timestamp 1624015447
transform -1 0 90896 0 1 125664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1145
timestamp 1624015447
transform -1 0 90896 0 -1 126752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1147
timestamp 1624015447
transform -1 0 90896 0 1 126752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_228_969
timestamp 1624015447
transform 1 0 90252 0 -1 126752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_458
timestamp 1624015447
transform 1 0 1104 0 -1 127840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_460
timestamp 1624015447
transform 1 0 1104 0 1 127840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_462
timestamp 1624015447
transform 1 0 1104 0 -1 128928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_230_3
timestamp 1624015447
transform 1 0 1380 0 -1 127840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_230_15
timestamp 1624015447
transform 1 0 2484 0 -1 127840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_231_3
timestamp 1624015447
transform 1 0 1380 0 1 127840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_231_15
timestamp 1624015447
transform 1 0 2484 0 1 127840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_232_3
timestamp 1624015447
transform 1 0 1380 0 -1 128928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_232_15
timestamp 1624015447
transform 1 0 2484 0 -1 128928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1490
timestamp 1624015447
transform 1 0 3772 0 -1 127840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1491
timestamp 1624015447
transform 1 0 3772 0 -1 128928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_230_27
timestamp 1624015447
transform 1 0 3588 0 -1 127840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_230_30
timestamp 1624015447
transform 1 0 3864 0 -1 127840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_231_27
timestamp 1624015447
transform 1 0 3588 0 1 127840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_232_27
timestamp 1624015447
transform 1 0 3588 0 -1 128928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_232_30
timestamp 1624015447
transform 1 0 3864 0 -1 128928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_459
timestamp 1624015447
transform -1 0 5152 0 -1 127840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_461
timestamp 1624015447
transform -1 0 5152 0 1 127840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_463
timestamp 1624015447
transform -1 0 5152 0 -1 128928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_230_38
timestamp 1624015447
transform 1 0 4600 0 -1 127840
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_231_39
timestamp 1624015447
transform 1 0 4692 0 1 127840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_232_38
timestamp 1624015447
transform 1 0 4600 0 -1 128928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1148
timestamp 1624015447
transform 1 0 84180 0 -1 127840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1150
timestamp 1624015447
transform 1 0 84180 0 1 127840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1152
timestamp 1624015447
transform 1 0 84180 0 -1 128928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_230_906
timestamp 1624015447
transform 1 0 84456 0 -1 127840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_231_906
timestamp 1624015447
transform 1 0 84456 0 1 127840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_232_906
timestamp 1624015447
transform 1 0 84456 0 -1 128928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_230_918
timestamp 1624015447
transform 1 0 85560 0 -1 127840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_231_918
timestamp 1624015447
transform 1 0 85560 0 1 127840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_232_918
timestamp 1624015447
transform 1 0 85560 0 -1 128928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_230_945
timestamp 1624015447
transform 1 0 88044 0 -1 127840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_230_933
timestamp 1624015447
transform 1 0 86940 0 -1 127840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_230_930
timestamp 1624015447
transform 1 0 86664 0 -1 127840
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1780
timestamp 1624015447
transform 1 0 86848 0 -1 127840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_231_942
timestamp 1624015447
transform 1 0 87768 0 1 127840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_231_930
timestamp 1624015447
transform 1 0 86664 0 1 127840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_232_945
timestamp 1624015447
transform 1 0 88044 0 -1 128928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_232_933
timestamp 1624015447
transform 1 0 86940 0 -1 128928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_232_930
timestamp 1624015447
transform 1 0 86664 0 -1 128928
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1782
timestamp 1624015447
transform 1 0 86848 0 -1 128928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1781
timestamp 1624015447
transform 1 0 89424 0 1 127840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_230_957
timestamp 1624015447
transform 1 0 89148 0 -1 127840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_231_954
timestamp 1624015447
transform 1 0 88872 0 1 127840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_231_961
timestamp 1624015447
transform 1 0 89516 0 1 127840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_232_957
timestamp 1624015447
transform 1 0 89148 0 -1 128928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1149
timestamp 1624015447
transform -1 0 90896 0 -1 127840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1151
timestamp 1624015447
transform -1 0 90896 0 1 127840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1153
timestamp 1624015447
transform -1 0 90896 0 -1 128928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_230_969
timestamp 1624015447
transform 1 0 90252 0 -1 127840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_232_969
timestamp 1624015447
transform 1 0 90252 0 -1 128928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_464
timestamp 1624015447
transform 1 0 1104 0 1 128928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_466
timestamp 1624015447
transform 1 0 1104 0 -1 130016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_468
timestamp 1624015447
transform 1 0 1104 0 1 130016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_233_3
timestamp 1624015447
transform 1 0 1380 0 1 128928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_233_15
timestamp 1624015447
transform 1 0 2484 0 1 128928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_234_3
timestamp 1624015447
transform 1 0 1380 0 -1 130016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_234_15
timestamp 1624015447
transform 1 0 2484 0 -1 130016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_235_3
timestamp 1624015447
transform 1 0 1380 0 1 130016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_235_15
timestamp 1624015447
transform 1 0 2484 0 1 130016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1492
timestamp 1624015447
transform 1 0 3772 0 -1 130016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_233_27
timestamp 1624015447
transform 1 0 3588 0 1 128928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_234_27
timestamp 1624015447
transform 1 0 3588 0 -1 130016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_234_30
timestamp 1624015447
transform 1 0 3864 0 -1 130016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_235_27
timestamp 1624015447
transform 1 0 3588 0 1 130016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_465
timestamp 1624015447
transform -1 0 5152 0 1 128928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_467
timestamp 1624015447
transform -1 0 5152 0 -1 130016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_469
timestamp 1624015447
transform -1 0 5152 0 1 130016
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_233_39
timestamp 1624015447
transform 1 0 4692 0 1 128928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_234_38
timestamp 1624015447
transform 1 0 4600 0 -1 130016
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_235_39
timestamp 1624015447
transform 1 0 4692 0 1 130016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1154
timestamp 1624015447
transform 1 0 84180 0 1 128928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1156
timestamp 1624015447
transform 1 0 84180 0 -1 130016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1158
timestamp 1624015447
transform 1 0 84180 0 1 130016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_233_906
timestamp 1624015447
transform 1 0 84456 0 1 128928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_234_906
timestamp 1624015447
transform 1 0 84456 0 -1 130016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_235_906
timestamp 1624015447
transform 1 0 84456 0 1 130016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_233_918
timestamp 1624015447
transform 1 0 85560 0 1 128928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_234_918
timestamp 1624015447
transform 1 0 85560 0 -1 130016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_235_918
timestamp 1624015447
transform 1 0 85560 0 1 130016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1784
timestamp 1624015447
transform 1 0 86848 0 -1 130016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_233_930
timestamp 1624015447
transform 1 0 86664 0 1 128928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_233_942
timestamp 1624015447
transform 1 0 87768 0 1 128928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_234_930
timestamp 1624015447
transform 1 0 86664 0 -1 130016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_234_933
timestamp 1624015447
transform 1 0 86940 0 -1 130016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_234_945
timestamp 1624015447
transform 1 0 88044 0 -1 130016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_235_930
timestamp 1624015447
transform 1 0 86664 0 1 130016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_235_942
timestamp 1624015447
transform 1 0 87768 0 1 130016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1783
timestamp 1624015447
transform 1 0 89424 0 1 128928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1785
timestamp 1624015447
transform 1 0 89424 0 1 130016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_233_954
timestamp 1624015447
transform 1 0 88872 0 1 128928
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_233_961
timestamp 1624015447
transform 1 0 89516 0 1 128928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_234_957
timestamp 1624015447
transform 1 0 89148 0 -1 130016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_235_954
timestamp 1624015447
transform 1 0 88872 0 1 130016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_235_961
timestamp 1624015447
transform 1 0 89516 0 1 130016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1155
timestamp 1624015447
transform -1 0 90896 0 1 128928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1157
timestamp 1624015447
transform -1 0 90896 0 -1 130016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1159
timestamp 1624015447
transform -1 0 90896 0 1 130016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_234_969
timestamp 1624015447
transform 1 0 90252 0 -1 130016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_470
timestamp 1624015447
transform 1 0 1104 0 -1 131104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_472
timestamp 1624015447
transform 1 0 1104 0 1 131104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_474
timestamp 1624015447
transform 1 0 1104 0 -1 132192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_236_3
timestamp 1624015447
transform 1 0 1380 0 -1 131104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_236_15
timestamp 1624015447
transform 1 0 2484 0 -1 131104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_237_3
timestamp 1624015447
transform 1 0 1380 0 1 131104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_237_15
timestamp 1624015447
transform 1 0 2484 0 1 131104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_238_3
timestamp 1624015447
transform 1 0 1380 0 -1 132192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_238_15
timestamp 1624015447
transform 1 0 2484 0 -1 132192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1493
timestamp 1624015447
transform 1 0 3772 0 -1 131104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1494
timestamp 1624015447
transform 1 0 3772 0 -1 132192
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_236_27
timestamp 1624015447
transform 1 0 3588 0 -1 131104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_236_30
timestamp 1624015447
transform 1 0 3864 0 -1 131104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_237_27
timestamp 1624015447
transform 1 0 3588 0 1 131104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_238_27
timestamp 1624015447
transform 1 0 3588 0 -1 132192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_238_30
timestamp 1624015447
transform 1 0 3864 0 -1 132192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_471
timestamp 1624015447
transform -1 0 5152 0 -1 131104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_473
timestamp 1624015447
transform -1 0 5152 0 1 131104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_475
timestamp 1624015447
transform -1 0 5152 0 -1 132192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_236_38
timestamp 1624015447
transform 1 0 4600 0 -1 131104
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_237_39
timestamp 1624015447
transform 1 0 4692 0 1 131104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_238_38
timestamp 1624015447
transform 1 0 4600 0 -1 132192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1160
timestamp 1624015447
transform 1 0 84180 0 -1 131104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1162
timestamp 1624015447
transform 1 0 84180 0 1 131104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1164
timestamp 1624015447
transform 1 0 84180 0 -1 132192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_236_906
timestamp 1624015447
transform 1 0 84456 0 -1 131104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_237_906
timestamp 1624015447
transform 1 0 84456 0 1 131104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_238_906
timestamp 1624015447
transform 1 0 84456 0 -1 132192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_236_918
timestamp 1624015447
transform 1 0 85560 0 -1 131104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_237_918
timestamp 1624015447
transform 1 0 85560 0 1 131104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_238_918
timestamp 1624015447
transform 1 0 85560 0 -1 132192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_236_945
timestamp 1624015447
transform 1 0 88044 0 -1 131104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_236_933
timestamp 1624015447
transform 1 0 86940 0 -1 131104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_236_930
timestamp 1624015447
transform 1 0 86664 0 -1 131104
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1786
timestamp 1624015447
transform 1 0 86848 0 -1 131104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_237_942
timestamp 1624015447
transform 1 0 87768 0 1 131104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_237_930
timestamp 1624015447
transform 1 0 86664 0 1 131104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_238_945
timestamp 1624015447
transform 1 0 88044 0 -1 132192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_238_933
timestamp 1624015447
transform 1 0 86940 0 -1 132192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_238_930
timestamp 1624015447
transform 1 0 86664 0 -1 132192
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1788
timestamp 1624015447
transform 1 0 86848 0 -1 132192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1787
timestamp 1624015447
transform 1 0 89424 0 1 131104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_236_957
timestamp 1624015447
transform 1 0 89148 0 -1 131104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_237_954
timestamp 1624015447
transform 1 0 88872 0 1 131104
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_237_961
timestamp 1624015447
transform 1 0 89516 0 1 131104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_238_957
timestamp 1624015447
transform 1 0 89148 0 -1 132192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1161
timestamp 1624015447
transform -1 0 90896 0 -1 131104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1163
timestamp 1624015447
transform -1 0 90896 0 1 131104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1165
timestamp 1624015447
transform -1 0 90896 0 -1 132192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_236_969
timestamp 1624015447
transform 1 0 90252 0 -1 131104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_238_969
timestamp 1624015447
transform 1 0 90252 0 -1 132192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_476
timestamp 1624015447
transform 1 0 1104 0 1 132192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_478
timestamp 1624015447
transform 1 0 1104 0 -1 133280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_480
timestamp 1624015447
transform 1 0 1104 0 1 133280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_239_3
timestamp 1624015447
transform 1 0 1380 0 1 132192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_239_15
timestamp 1624015447
transform 1 0 2484 0 1 132192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_240_3
timestamp 1624015447
transform 1 0 1380 0 -1 133280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_240_15
timestamp 1624015447
transform 1 0 2484 0 -1 133280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_241_3
timestamp 1624015447
transform 1 0 1380 0 1 133280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_241_15
timestamp 1624015447
transform 1 0 2484 0 1 133280
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1495
timestamp 1624015447
transform 1 0 3772 0 -1 133280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_239_27
timestamp 1624015447
transform 1 0 3588 0 1 132192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_240_27
timestamp 1624015447
transform 1 0 3588 0 -1 133280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_240_30
timestamp 1624015447
transform 1 0 3864 0 -1 133280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_241_27
timestamp 1624015447
transform 1 0 3588 0 1 133280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_477
timestamp 1624015447
transform -1 0 5152 0 1 132192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_479
timestamp 1624015447
transform -1 0 5152 0 -1 133280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_481
timestamp 1624015447
transform -1 0 5152 0 1 133280
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_239_39
timestamp 1624015447
transform 1 0 4692 0 1 132192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_240_38
timestamp 1624015447
transform 1 0 4600 0 -1 133280
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_241_39
timestamp 1624015447
transform 1 0 4692 0 1 133280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1166
timestamp 1624015447
transform 1 0 84180 0 1 132192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1168
timestamp 1624015447
transform 1 0 84180 0 -1 133280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1170
timestamp 1624015447
transform 1 0 84180 0 1 133280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_239_906
timestamp 1624015447
transform 1 0 84456 0 1 132192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_240_906
timestamp 1624015447
transform 1 0 84456 0 -1 133280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_241_906
timestamp 1624015447
transform 1 0 84456 0 1 133280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_239_918
timestamp 1624015447
transform 1 0 85560 0 1 132192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_240_918
timestamp 1624015447
transform 1 0 85560 0 -1 133280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_241_918
timestamp 1624015447
transform 1 0 85560 0 1 133280
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1790
timestamp 1624015447
transform 1 0 86848 0 -1 133280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_239_930
timestamp 1624015447
transform 1 0 86664 0 1 132192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_239_942
timestamp 1624015447
transform 1 0 87768 0 1 132192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_240_930
timestamp 1624015447
transform 1 0 86664 0 -1 133280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_240_933
timestamp 1624015447
transform 1 0 86940 0 -1 133280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_240_945
timestamp 1624015447
transform 1 0 88044 0 -1 133280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_241_930
timestamp 1624015447
transform 1 0 86664 0 1 133280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_241_942
timestamp 1624015447
transform 1 0 87768 0 1 133280
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1789
timestamp 1624015447
transform 1 0 89424 0 1 132192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1791
timestamp 1624015447
transform 1 0 89424 0 1 133280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_239_954
timestamp 1624015447
transform 1 0 88872 0 1 132192
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_239_961
timestamp 1624015447
transform 1 0 89516 0 1 132192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_240_957
timestamp 1624015447
transform 1 0 89148 0 -1 133280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_241_954
timestamp 1624015447
transform 1 0 88872 0 1 133280
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_241_961
timestamp 1624015447
transform 1 0 89516 0 1 133280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1167
timestamp 1624015447
transform -1 0 90896 0 1 132192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1169
timestamp 1624015447
transform -1 0 90896 0 -1 133280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1171
timestamp 1624015447
transform -1 0 90896 0 1 133280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_240_969
timestamp 1624015447
transform 1 0 90252 0 -1 133280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_482
timestamp 1624015447
transform 1 0 1104 0 -1 134368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_484
timestamp 1624015447
transform 1 0 1104 0 1 134368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_486
timestamp 1624015447
transform 1 0 1104 0 -1 135456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_242_3
timestamp 1624015447
transform 1 0 1380 0 -1 134368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_242_15
timestamp 1624015447
transform 1 0 2484 0 -1 134368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_243_3
timestamp 1624015447
transform 1 0 1380 0 1 134368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_243_15
timestamp 1624015447
transform 1 0 2484 0 1 134368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_244_3
timestamp 1624015447
transform 1 0 1380 0 -1 135456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_244_15
timestamp 1624015447
transform 1 0 2484 0 -1 135456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1496
timestamp 1624015447
transform 1 0 3772 0 -1 134368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1497
timestamp 1624015447
transform 1 0 3772 0 -1 135456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_242_27
timestamp 1624015447
transform 1 0 3588 0 -1 134368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_242_30
timestamp 1624015447
transform 1 0 3864 0 -1 134368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_243_27
timestamp 1624015447
transform 1 0 3588 0 1 134368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_244_27
timestamp 1624015447
transform 1 0 3588 0 -1 135456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_244_30
timestamp 1624015447
transform 1 0 3864 0 -1 135456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_483
timestamp 1624015447
transform -1 0 5152 0 -1 134368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_485
timestamp 1624015447
transform -1 0 5152 0 1 134368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_487
timestamp 1624015447
transform -1 0 5152 0 -1 135456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_242_38
timestamp 1624015447
transform 1 0 4600 0 -1 134368
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_243_39
timestamp 1624015447
transform 1 0 4692 0 1 134368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_244_38
timestamp 1624015447
transform 1 0 4600 0 -1 135456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1172
timestamp 1624015447
transform 1 0 84180 0 -1 134368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1174
timestamp 1624015447
transform 1 0 84180 0 1 134368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1176
timestamp 1624015447
transform 1 0 84180 0 -1 135456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_242_906
timestamp 1624015447
transform 1 0 84456 0 -1 134368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_243_906
timestamp 1624015447
transform 1 0 84456 0 1 134368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_244_906
timestamp 1624015447
transform 1 0 84456 0 -1 135456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_242_918
timestamp 1624015447
transform 1 0 85560 0 -1 134368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_243_918
timestamp 1624015447
transform 1 0 85560 0 1 134368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_244_918
timestamp 1624015447
transform 1 0 85560 0 -1 135456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_242_945
timestamp 1624015447
transform 1 0 88044 0 -1 134368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_242_933
timestamp 1624015447
transform 1 0 86940 0 -1 134368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_242_930
timestamp 1624015447
transform 1 0 86664 0 -1 134368
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1792
timestamp 1624015447
transform 1 0 86848 0 -1 134368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_244_945
timestamp 1624015447
transform 1 0 88044 0 -1 135456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_244_933
timestamp 1624015447
transform 1 0 86940 0 -1 135456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_244_930
timestamp 1624015447
transform 1 0 86664 0 -1 135456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_243_942
timestamp 1624015447
transform 1 0 87768 0 1 134368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_243_930
timestamp 1624015447
transform 1 0 86664 0 1 134368
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1794
timestamp 1624015447
transform 1 0 86848 0 -1 135456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1793
timestamp 1624015447
transform 1 0 89424 0 1 134368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_242_957
timestamp 1624015447
transform 1 0 89148 0 -1 134368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_243_954
timestamp 1624015447
transform 1 0 88872 0 1 134368
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_243_961
timestamp 1624015447
transform 1 0 89516 0 1 134368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_244_957
timestamp 1624015447
transform 1 0 89148 0 -1 135456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1173
timestamp 1624015447
transform -1 0 90896 0 -1 134368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1175
timestamp 1624015447
transform -1 0 90896 0 1 134368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1177
timestamp 1624015447
transform -1 0 90896 0 -1 135456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_242_969
timestamp 1624015447
transform 1 0 90252 0 -1 134368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_244_969
timestamp 1624015447
transform 1 0 90252 0 -1 135456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_488
timestamp 1624015447
transform 1 0 1104 0 1 135456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_490
timestamp 1624015447
transform 1 0 1104 0 -1 136544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_492
timestamp 1624015447
transform 1 0 1104 0 1 136544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_245_3
timestamp 1624015447
transform 1 0 1380 0 1 135456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_245_15
timestamp 1624015447
transform 1 0 2484 0 1 135456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_246_3
timestamp 1624015447
transform 1 0 1380 0 -1 136544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_246_15
timestamp 1624015447
transform 1 0 2484 0 -1 136544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_247_3
timestamp 1624015447
transform 1 0 1380 0 1 136544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_247_15
timestamp 1624015447
transform 1 0 2484 0 1 136544
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1498
timestamp 1624015447
transform 1 0 3772 0 -1 136544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_245_27
timestamp 1624015447
transform 1 0 3588 0 1 135456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_246_27
timestamp 1624015447
transform 1 0 3588 0 -1 136544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_246_30
timestamp 1624015447
transform 1 0 3864 0 -1 136544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_247_27
timestamp 1624015447
transform 1 0 3588 0 1 136544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_489
timestamp 1624015447
transform -1 0 5152 0 1 135456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_491
timestamp 1624015447
transform -1 0 5152 0 -1 136544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_493
timestamp 1624015447
transform -1 0 5152 0 1 136544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_245_39
timestamp 1624015447
transform 1 0 4692 0 1 135456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_246_38
timestamp 1624015447
transform 1 0 4600 0 -1 136544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_247_39
timestamp 1624015447
transform 1 0 4692 0 1 136544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1178
timestamp 1624015447
transform 1 0 84180 0 1 135456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1180
timestamp 1624015447
transform 1 0 84180 0 -1 136544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1182
timestamp 1624015447
transform 1 0 84180 0 1 136544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_245_906
timestamp 1624015447
transform 1 0 84456 0 1 135456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_246_906
timestamp 1624015447
transform 1 0 84456 0 -1 136544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_247_906
timestamp 1624015447
transform 1 0 84456 0 1 136544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_245_918
timestamp 1624015447
transform 1 0 85560 0 1 135456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_246_918
timestamp 1624015447
transform 1 0 85560 0 -1 136544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_247_918
timestamp 1624015447
transform 1 0 85560 0 1 136544
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1796
timestamp 1624015447
transform 1 0 86848 0 -1 136544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_245_930
timestamp 1624015447
transform 1 0 86664 0 1 135456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_245_942
timestamp 1624015447
transform 1 0 87768 0 1 135456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_246_930
timestamp 1624015447
transform 1 0 86664 0 -1 136544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_246_933
timestamp 1624015447
transform 1 0 86940 0 -1 136544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_246_945
timestamp 1624015447
transform 1 0 88044 0 -1 136544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_247_930
timestamp 1624015447
transform 1 0 86664 0 1 136544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_247_942
timestamp 1624015447
transform 1 0 87768 0 1 136544
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1795
timestamp 1624015447
transform 1 0 89424 0 1 135456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1797
timestamp 1624015447
transform 1 0 89424 0 1 136544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_245_954
timestamp 1624015447
transform 1 0 88872 0 1 135456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_245_961
timestamp 1624015447
transform 1 0 89516 0 1 135456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_246_957
timestamp 1624015447
transform 1 0 89148 0 -1 136544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_954
timestamp 1624015447
transform 1 0 88872 0 1 136544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_247_961
timestamp 1624015447
transform 1 0 89516 0 1 136544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1179
timestamp 1624015447
transform -1 0 90896 0 1 135456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1181
timestamp 1624015447
transform -1 0 90896 0 -1 136544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1183
timestamp 1624015447
transform -1 0 90896 0 1 136544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_246_969
timestamp 1624015447
transform 1 0 90252 0 -1 136544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_494
timestamp 1624015447
transform 1 0 1104 0 -1 137632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_496
timestamp 1624015447
transform 1 0 1104 0 1 137632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_498
timestamp 1624015447
transform 1 0 1104 0 -1 138720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_248_3
timestamp 1624015447
transform 1 0 1380 0 -1 137632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_248_15
timestamp 1624015447
transform 1 0 2484 0 -1 137632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_249_3
timestamp 1624015447
transform 1 0 1380 0 1 137632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_249_15
timestamp 1624015447
transform 1 0 2484 0 1 137632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_250_3
timestamp 1624015447
transform 1 0 1380 0 -1 138720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_250_15
timestamp 1624015447
transform 1 0 2484 0 -1 138720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1499
timestamp 1624015447
transform 1 0 3772 0 -1 137632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1500
timestamp 1624015447
transform 1 0 3772 0 -1 138720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_248_27
timestamp 1624015447
transform 1 0 3588 0 -1 137632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_248_30
timestamp 1624015447
transform 1 0 3864 0 -1 137632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_249_27
timestamp 1624015447
transform 1 0 3588 0 1 137632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_250_27
timestamp 1624015447
transform 1 0 3588 0 -1 138720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_250_30
timestamp 1624015447
transform 1 0 3864 0 -1 138720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_495
timestamp 1624015447
transform -1 0 5152 0 -1 137632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_497
timestamp 1624015447
transform -1 0 5152 0 1 137632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_499
timestamp 1624015447
transform -1 0 5152 0 -1 138720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_248_38
timestamp 1624015447
transform 1 0 4600 0 -1 137632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_249_39
timestamp 1624015447
transform 1 0 4692 0 1 137632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_250_38
timestamp 1624015447
transform 1 0 4600 0 -1 138720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1184
timestamp 1624015447
transform 1 0 84180 0 -1 137632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1186
timestamp 1624015447
transform 1 0 84180 0 1 137632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1188
timestamp 1624015447
transform 1 0 84180 0 -1 138720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_248_906
timestamp 1624015447
transform 1 0 84456 0 -1 137632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_249_906
timestamp 1624015447
transform 1 0 84456 0 1 137632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_250_906
timestamp 1624015447
transform 1 0 84456 0 -1 138720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_248_918
timestamp 1624015447
transform 1 0 85560 0 -1 137632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_249_918
timestamp 1624015447
transform 1 0 85560 0 1 137632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_250_918
timestamp 1624015447
transform 1 0 85560 0 -1 138720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_249_942
timestamp 1624015447
transform 1 0 87768 0 1 137632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_249_930
timestamp 1624015447
transform 1 0 86664 0 1 137632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_248_945
timestamp 1624015447
transform 1 0 88044 0 -1 137632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_248_933
timestamp 1624015447
transform 1 0 86940 0 -1 137632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_248_930
timestamp 1624015447
transform 1 0 86664 0 -1 137632
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1798
timestamp 1624015447
transform 1 0 86848 0 -1 137632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_250_945
timestamp 1624015447
transform 1 0 88044 0 -1 138720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_250_933
timestamp 1624015447
transform 1 0 86940 0 -1 138720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_250_930
timestamp 1624015447
transform 1 0 86664 0 -1 138720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1800
timestamp 1624015447
transform 1 0 86848 0 -1 138720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1799
timestamp 1624015447
transform 1 0 89424 0 1 137632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_248_957
timestamp 1624015447
transform 1 0 89148 0 -1 137632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_954
timestamp 1624015447
transform 1 0 88872 0 1 137632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_249_961
timestamp 1624015447
transform 1 0 89516 0 1 137632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_250_957
timestamp 1624015447
transform 1 0 89148 0 -1 138720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1185
timestamp 1624015447
transform -1 0 90896 0 -1 137632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1187
timestamp 1624015447
transform -1 0 90896 0 1 137632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1189
timestamp 1624015447
transform -1 0 90896 0 -1 138720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_248_969
timestamp 1624015447
transform 1 0 90252 0 -1 137632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_250_969
timestamp 1624015447
transform 1 0 90252 0 -1 138720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_500
timestamp 1624015447
transform 1 0 1104 0 1 138720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_251_3
timestamp 1624015447
transform 1 0 1380 0 1 138720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_251_15
timestamp 1624015447
transform 1 0 2484 0 1 138720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_251_27
timestamp 1624015447
transform 1 0 3588 0 1 138720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_501
timestamp 1624015447
transform -1 0 5152 0 1 138720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_251_39
timestamp 1624015447
transform 1 0 4692 0 1 138720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1190
timestamp 1624015447
transform 1 0 84180 0 1 138720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_251_906
timestamp 1624015447
transform 1 0 84456 0 1 138720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_251_918
timestamp 1624015447
transform 1 0 85560 0 1 138720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_251_930
timestamp 1624015447
transform 1 0 86664 0 1 138720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_251_942
timestamp 1624015447
transform 1 0 87768 0 1 138720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1801
timestamp 1624015447
transform 1 0 89424 0 1 138720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_251_954
timestamp 1624015447
transform 1 0 88872 0 1 138720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_251_961
timestamp 1624015447
transform 1 0 89516 0 1 138720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1191
timestamp 1624015447
transform -1 0 90896 0 1 138720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_502
timestamp 1624015447
transform 1 0 1104 0 -1 139808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_504
timestamp 1624015447
transform 1 0 1104 0 1 139808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_506
timestamp 1624015447
transform 1 0 1104 0 -1 140896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_252_3
timestamp 1624015447
transform 1 0 1380 0 -1 139808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_252_15
timestamp 1624015447
transform 1 0 2484 0 -1 139808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_253_3
timestamp 1624015447
transform 1 0 1380 0 1 139808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_253_15
timestamp 1624015447
transform 1 0 2484 0 1 139808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_254_3
timestamp 1624015447
transform 1 0 1380 0 -1 140896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_254_15
timestamp 1624015447
transform 1 0 2484 0 -1 140896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1501
timestamp 1624015447
transform 1 0 3772 0 -1 139808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1502
timestamp 1624015447
transform 1 0 3772 0 -1 140896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_252_27
timestamp 1624015447
transform 1 0 3588 0 -1 139808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_252_30
timestamp 1624015447
transform 1 0 3864 0 -1 139808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_253_27
timestamp 1624015447
transform 1 0 3588 0 1 139808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_254_27
timestamp 1624015447
transform 1 0 3588 0 -1 140896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_254_30
timestamp 1624015447
transform 1 0 3864 0 -1 140896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_503
timestamp 1624015447
transform -1 0 5152 0 -1 139808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_505
timestamp 1624015447
transform -1 0 5152 0 1 139808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_507
timestamp 1624015447
transform -1 0 5152 0 -1 140896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_252_38
timestamp 1624015447
transform 1 0 4600 0 -1 139808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_253_39
timestamp 1624015447
transform 1 0 4692 0 1 139808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_254_38
timestamp 1624015447
transform 1 0 4600 0 -1 140896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1192
timestamp 1624015447
transform 1 0 84180 0 -1 139808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1194
timestamp 1624015447
transform 1 0 84180 0 1 139808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1196
timestamp 1624015447
transform 1 0 84180 0 -1 140896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_252_906
timestamp 1624015447
transform 1 0 84456 0 -1 139808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_253_906
timestamp 1624015447
transform 1 0 84456 0 1 139808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_254_906
timestamp 1624015447
transform 1 0 84456 0 -1 140896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_252_918
timestamp 1624015447
transform 1 0 85560 0 -1 139808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_252_930
timestamp 1624015447
transform 1 0 86664 0 -1 139808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_253_918
timestamp 1624015447
transform 1 0 85560 0 1 139808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_253_930
timestamp 1624015447
transform 1 0 86664 0 1 139808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_254_918
timestamp 1624015447
transform 1 0 85560 0 -1 140896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_254_930
timestamp 1624015447
transform 1 0 86664 0 -1 140896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1802
timestamp 1624015447
transform 1 0 86848 0 -1 139808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1804
timestamp 1624015447
transform 1 0 86848 0 -1 140896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_252_933
timestamp 1624015447
transform 1 0 86940 0 -1 139808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_252_945
timestamp 1624015447
transform 1 0 88044 0 -1 139808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_253_942
timestamp 1624015447
transform 1 0 87768 0 1 139808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_254_933
timestamp 1624015447
transform 1 0 86940 0 -1 140896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_254_945
timestamp 1624015447
transform 1 0 88044 0 -1 140896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1803
timestamp 1624015447
transform 1 0 89424 0 1 139808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_252_957
timestamp 1624015447
transform 1 0 89148 0 -1 139808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_954
timestamp 1624015447
transform 1 0 88872 0 1 139808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_253_961
timestamp 1624015447
transform 1 0 89516 0 1 139808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_254_957
timestamp 1624015447
transform 1 0 89148 0 -1 140896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1193
timestamp 1624015447
transform -1 0 90896 0 -1 139808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1195
timestamp 1624015447
transform -1 0 90896 0 1 139808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1197
timestamp 1624015447
transform -1 0 90896 0 -1 140896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_252_969
timestamp 1624015447
transform 1 0 90252 0 -1 139808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_254_969
timestamp 1624015447
transform 1 0 90252 0 -1 140896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_508
timestamp 1624015447
transform 1 0 1104 0 1 140896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_510
timestamp 1624015447
transform 1 0 1104 0 -1 141984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_512
timestamp 1624015447
transform 1 0 1104 0 1 141984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_255_3
timestamp 1624015447
transform 1 0 1380 0 1 140896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_255_15
timestamp 1624015447
transform 1 0 2484 0 1 140896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_256_3
timestamp 1624015447
transform 1 0 1380 0 -1 141984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_256_15
timestamp 1624015447
transform 1 0 2484 0 -1 141984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_257_3
timestamp 1624015447
transform 1 0 1380 0 1 141984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_257_15
timestamp 1624015447
transform 1 0 2484 0 1 141984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1503
timestamp 1624015447
transform 1 0 3772 0 -1 141984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_255_27
timestamp 1624015447
transform 1 0 3588 0 1 140896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_256_27
timestamp 1624015447
transform 1 0 3588 0 -1 141984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_256_30
timestamp 1624015447
transform 1 0 3864 0 -1 141984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_257_27
timestamp 1624015447
transform 1 0 3588 0 1 141984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_509
timestamp 1624015447
transform -1 0 5152 0 1 140896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_511
timestamp 1624015447
transform -1 0 5152 0 -1 141984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_513
timestamp 1624015447
transform -1 0 5152 0 1 141984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_255_39
timestamp 1624015447
transform 1 0 4692 0 1 140896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_256_38
timestamp 1624015447
transform 1 0 4600 0 -1 141984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_257_39
timestamp 1624015447
transform 1 0 4692 0 1 141984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  BUF_4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624015447
transform -1 0 85008 0 1 140896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_1198
timestamp 1624015447
transform 1 0 84180 0 1 140896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1200
timestamp 1624015447
transform 1 0 84180 0 -1 141984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1202
timestamp 1624015447
transform 1 0 84180 0 1 141984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_256_906
timestamp 1624015447
transform 1 0 84456 0 -1 141984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_257_906
timestamp 1624015447
transform 1 0 84456 0 1 141984
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF_4_A
timestamp 1624015447
transform -1 0 85376 0 1 140896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_255_912
timestamp 1624015447
transform 1 0 85008 0 1 140896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_255_916
timestamp 1624015447
transform 1 0 85376 0 1 140896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_255_928
timestamp 1624015447
transform 1 0 86480 0 1 140896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_256_918
timestamp 1624015447
transform 1 0 85560 0 -1 141984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_256_930
timestamp 1624015447
transform 1 0 86664 0 -1 141984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_257_918
timestamp 1624015447
transform 1 0 85560 0 1 141984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_257_930
timestamp 1624015447
transform 1 0 86664 0 1 141984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1806
timestamp 1624015447
transform 1 0 86848 0 -1 141984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_255_940
timestamp 1624015447
transform 1 0 87584 0 1 140896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_256_933
timestamp 1624015447
transform 1 0 86940 0 -1 141984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_256_945
timestamp 1624015447
transform 1 0 88044 0 -1 141984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_257_942
timestamp 1624015447
transform 1 0 87768 0 1 141984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1805
timestamp 1624015447
transform 1 0 89424 0 1 140896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1807
timestamp 1624015447
transform 1 0 89424 0 1 141984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_255_952
timestamp 1624015447
transform 1 0 88688 0 1 140896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_255_961
timestamp 1624015447
transform 1 0 89516 0 1 140896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_256_957
timestamp 1624015447
transform 1 0 89148 0 -1 141984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_954
timestamp 1624015447
transform 1 0 88872 0 1 141984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_257_961
timestamp 1624015447
transform 1 0 89516 0 1 141984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1199
timestamp 1624015447
transform -1 0 90896 0 1 140896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1201
timestamp 1624015447
transform -1 0 90896 0 -1 141984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1203
timestamp 1624015447
transform -1 0 90896 0 1 141984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_256_969
timestamp 1624015447
transform 1 0 90252 0 -1 141984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_259_15
timestamp 1624015447
transform 1 0 2484 0 1 143072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_259_3
timestamp 1624015447
transform 1 0 1380 0 1 143072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_258_15
timestamp 1624015447
transform 1 0 2484 0 -1 143072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_258_3
timestamp 1624015447
transform 1 0 1380 0 -1 143072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_516
timestamp 1624015447
transform 1 0 1104 0 1 143072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_514
timestamp 1624015447
transform 1 0 1104 0 -1 143072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_260_15
timestamp 1624015447
transform 1 0 2484 0 -1 144160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_260_3
timestamp 1624015447
transform 1 0 1380 0 -1 144160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_518
timestamp 1624015447
transform 1 0 1104 0 -1 144160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_261_15
timestamp 1624015447
transform 1 0 2484 0 1 144160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_261_3
timestamp 1624015447
transform 1 0 1380 0 1 144160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_520
timestamp 1624015447
transform 1 0 1104 0 1 144160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1504
timestamp 1624015447
transform 1 0 3772 0 -1 143072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1505
timestamp 1624015447
transform 1 0 3772 0 -1 144160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_258_27
timestamp 1624015447
transform 1 0 3588 0 -1 143072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_258_30
timestamp 1624015447
transform 1 0 3864 0 -1 143072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_259_27
timestamp 1624015447
transform 1 0 3588 0 1 143072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_260_27
timestamp 1624015447
transform 1 0 3588 0 -1 144160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_260_30
timestamp 1624015447
transform 1 0 3864 0 -1 144160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_261_27
timestamp 1624015447
transform 1 0 3588 0 1 144160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_515
timestamp 1624015447
transform -1 0 5152 0 -1 143072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_517
timestamp 1624015447
transform -1 0 5152 0 1 143072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_519
timestamp 1624015447
transform -1 0 5152 0 -1 144160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_521
timestamp 1624015447
transform -1 0 5152 0 1 144160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_258_38
timestamp 1624015447
transform 1 0 4600 0 -1 143072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_259_39
timestamp 1624015447
transform 1 0 4692 0 1 143072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_260_38
timestamp 1624015447
transform 1 0 4600 0 -1 144160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_261_39
timestamp 1624015447
transform 1 0 4692 0 1 144160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1204
timestamp 1624015447
transform 1 0 84180 0 -1 143072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1206
timestamp 1624015447
transform 1 0 84180 0 1 143072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1208
timestamp 1624015447
transform 1 0 84180 0 -1 144160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1210
timestamp 1624015447
transform 1 0 84180 0 1 144160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_258_906
timestamp 1624015447
transform 1 0 84456 0 -1 143072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_259_906
timestamp 1624015447
transform 1 0 84456 0 1 143072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_260_906
timestamp 1624015447
transform 1 0 84456 0 -1 144160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_261_906
timestamp 1624015447
transform 1 0 84456 0 1 144160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_258_918
timestamp 1624015447
transform 1 0 85560 0 -1 143072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_258_930
timestamp 1624015447
transform 1 0 86664 0 -1 143072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_259_918
timestamp 1624015447
transform 1 0 85560 0 1 143072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_259_930
timestamp 1624015447
transform 1 0 86664 0 1 143072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_260_918
timestamp 1624015447
transform 1 0 85560 0 -1 144160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_260_930
timestamp 1624015447
transform 1 0 86664 0 -1 144160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_261_918
timestamp 1624015447
transform 1 0 85560 0 1 144160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_261_930
timestamp 1624015447
transform 1 0 86664 0 1 144160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1808
timestamp 1624015447
transform 1 0 86848 0 -1 143072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1810
timestamp 1624015447
transform 1 0 86848 0 -1 144160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_258_933
timestamp 1624015447
transform 1 0 86940 0 -1 143072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_258_945
timestamp 1624015447
transform 1 0 88044 0 -1 143072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_259_942
timestamp 1624015447
transform 1 0 87768 0 1 143072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_260_933
timestamp 1624015447
transform 1 0 86940 0 -1 144160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_260_945
timestamp 1624015447
transform 1 0 88044 0 -1 144160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_261_942
timestamp 1624015447
transform 1 0 87768 0 1 144160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1809
timestamp 1624015447
transform 1 0 89424 0 1 143072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1811
timestamp 1624015447
transform 1 0 89424 0 1 144160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_258_957
timestamp 1624015447
transform 1 0 89148 0 -1 143072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_954
timestamp 1624015447
transform 1 0 88872 0 1 143072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_259_961
timestamp 1624015447
transform 1 0 89516 0 1 143072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_260_957
timestamp 1624015447
transform 1 0 89148 0 -1 144160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_954
timestamp 1624015447
transform 1 0 88872 0 1 144160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_261_961
timestamp 1624015447
transform 1 0 89516 0 1 144160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1205
timestamp 1624015447
transform -1 0 90896 0 -1 143072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1207
timestamp 1624015447
transform -1 0 90896 0 1 143072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1209
timestamp 1624015447
transform -1 0 90896 0 -1 144160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1211
timestamp 1624015447
transform -1 0 90896 0 1 144160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_258_969
timestamp 1624015447
transform 1 0 90252 0 -1 143072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_260_969
timestamp 1624015447
transform 1 0 90252 0 -1 144160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_522
timestamp 1624015447
transform 1 0 1104 0 -1 145248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_524
timestamp 1624015447
transform 1 0 1104 0 1 145248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_526
timestamp 1624015447
transform 1 0 1104 0 -1 146336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_262_3
timestamp 1624015447
transform 1 0 1380 0 -1 145248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_262_15
timestamp 1624015447
transform 1 0 2484 0 -1 145248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_263_3
timestamp 1624015447
transform 1 0 1380 0 1 145248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_263_15
timestamp 1624015447
transform 1 0 2484 0 1 145248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_264_3
timestamp 1624015447
transform 1 0 1380 0 -1 146336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_264_15
timestamp 1624015447
transform 1 0 2484 0 -1 146336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1506
timestamp 1624015447
transform 1 0 3772 0 -1 145248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1507
timestamp 1624015447
transform 1 0 3772 0 -1 146336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_262_27
timestamp 1624015447
transform 1 0 3588 0 -1 145248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_262_30
timestamp 1624015447
transform 1 0 3864 0 -1 145248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_263_27
timestamp 1624015447
transform 1 0 3588 0 1 145248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_264_27
timestamp 1624015447
transform 1 0 3588 0 -1 146336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_264_30
timestamp 1624015447
transform 1 0 3864 0 -1 146336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_523
timestamp 1624015447
transform -1 0 5152 0 -1 145248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_525
timestamp 1624015447
transform -1 0 5152 0 1 145248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_527
timestamp 1624015447
transform -1 0 5152 0 -1 146336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_262_38
timestamp 1624015447
transform 1 0 4600 0 -1 145248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_263_39
timestamp 1624015447
transform 1 0 4692 0 1 145248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_264_38
timestamp 1624015447
transform 1 0 4600 0 -1 146336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1212
timestamp 1624015447
transform 1 0 84180 0 -1 145248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1214
timestamp 1624015447
transform 1 0 84180 0 1 145248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1216
timestamp 1624015447
transform 1 0 84180 0 -1 146336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_262_906
timestamp 1624015447
transform 1 0 84456 0 -1 145248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_263_906
timestamp 1624015447
transform 1 0 84456 0 1 145248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_264_906
timestamp 1624015447
transform 1 0 84456 0 -1 146336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_262_918
timestamp 1624015447
transform 1 0 85560 0 -1 145248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_262_930
timestamp 1624015447
transform 1 0 86664 0 -1 145248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_263_918
timestamp 1624015447
transform 1 0 85560 0 1 145248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_263_930
timestamp 1624015447
transform 1 0 86664 0 1 145248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_264_918
timestamp 1624015447
transform 1 0 85560 0 -1 146336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_264_930
timestamp 1624015447
transform 1 0 86664 0 -1 146336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1812
timestamp 1624015447
transform 1 0 86848 0 -1 145248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1814
timestamp 1624015447
transform 1 0 86848 0 -1 146336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_262_933
timestamp 1624015447
transform 1 0 86940 0 -1 145248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_262_945
timestamp 1624015447
transform 1 0 88044 0 -1 145248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_263_942
timestamp 1624015447
transform 1 0 87768 0 1 145248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_264_933
timestamp 1624015447
transform 1 0 86940 0 -1 146336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_264_945
timestamp 1624015447
transform 1 0 88044 0 -1 146336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1813
timestamp 1624015447
transform 1 0 89424 0 1 145248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_262_957
timestamp 1624015447
transform 1 0 89148 0 -1 145248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_954
timestamp 1624015447
transform 1 0 88872 0 1 145248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_263_961
timestamp 1624015447
transform 1 0 89516 0 1 145248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_264_957
timestamp 1624015447
transform 1 0 89148 0 -1 146336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1213
timestamp 1624015447
transform -1 0 90896 0 -1 145248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1215
timestamp 1624015447
transform -1 0 90896 0 1 145248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1217
timestamp 1624015447
transform -1 0 90896 0 -1 146336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_262_969
timestamp 1624015447
transform 1 0 90252 0 -1 145248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_264_969
timestamp 1624015447
transform 1 0 90252 0 -1 146336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_528
timestamp 1624015447
transform 1 0 1104 0 1 146336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_530
timestamp 1624015447
transform 1 0 1104 0 -1 147424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_532
timestamp 1624015447
transform 1 0 1104 0 1 147424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_265_3
timestamp 1624015447
transform 1 0 1380 0 1 146336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_265_15
timestamp 1624015447
transform 1 0 2484 0 1 146336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_266_3
timestamp 1624015447
transform 1 0 1380 0 -1 147424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_266_15
timestamp 1624015447
transform 1 0 2484 0 -1 147424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_267_3
timestamp 1624015447
transform 1 0 1380 0 1 147424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_267_15
timestamp 1624015447
transform 1 0 2484 0 1 147424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1508
timestamp 1624015447
transform 1 0 3772 0 -1 147424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_265_27
timestamp 1624015447
transform 1 0 3588 0 1 146336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_266_27
timestamp 1624015447
transform 1 0 3588 0 -1 147424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_266_30
timestamp 1624015447
transform 1 0 3864 0 -1 147424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_267_27
timestamp 1624015447
transform 1 0 3588 0 1 147424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_529
timestamp 1624015447
transform -1 0 5152 0 1 146336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_531
timestamp 1624015447
transform -1 0 5152 0 -1 147424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_533
timestamp 1624015447
transform -1 0 5152 0 1 147424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_265_39
timestamp 1624015447
transform 1 0 4692 0 1 146336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_266_38
timestamp 1624015447
transform 1 0 4600 0 -1 147424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_267_39
timestamp 1624015447
transform 1 0 4692 0 1 147424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1218
timestamp 1624015447
transform 1 0 84180 0 1 146336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1220
timestamp 1624015447
transform 1 0 84180 0 -1 147424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1222
timestamp 1624015447
transform 1 0 84180 0 1 147424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_265_906
timestamp 1624015447
transform 1 0 84456 0 1 146336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_266_906
timestamp 1624015447
transform 1 0 84456 0 -1 147424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_267_906
timestamp 1624015447
transform 1 0 84456 0 1 147424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_265_918
timestamp 1624015447
transform 1 0 85560 0 1 146336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_265_930
timestamp 1624015447
transform 1 0 86664 0 1 146336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_266_918
timestamp 1624015447
transform 1 0 85560 0 -1 147424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_266_930
timestamp 1624015447
transform 1 0 86664 0 -1 147424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_267_918
timestamp 1624015447
transform 1 0 85560 0 1 147424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_267_930
timestamp 1624015447
transform 1 0 86664 0 1 147424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1816
timestamp 1624015447
transform 1 0 86848 0 -1 147424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_265_942
timestamp 1624015447
transform 1 0 87768 0 1 146336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_266_933
timestamp 1624015447
transform 1 0 86940 0 -1 147424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_266_945
timestamp 1624015447
transform 1 0 88044 0 -1 147424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_267_942
timestamp 1624015447
transform 1 0 87768 0 1 147424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1815
timestamp 1624015447
transform 1 0 89424 0 1 146336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1817
timestamp 1624015447
transform 1 0 89424 0 1 147424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_265_954
timestamp 1624015447
transform 1 0 88872 0 1 146336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_265_961
timestamp 1624015447
transform 1 0 89516 0 1 146336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_266_957
timestamp 1624015447
transform 1 0 89148 0 -1 147424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_267_954
timestamp 1624015447
transform 1 0 88872 0 1 147424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_267_961
timestamp 1624015447
transform 1 0 89516 0 1 147424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1219
timestamp 1624015447
transform -1 0 90896 0 1 146336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1221
timestamp 1624015447
transform -1 0 90896 0 -1 147424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1223
timestamp 1624015447
transform -1 0 90896 0 1 147424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_266_969
timestamp 1624015447
transform 1 0 90252 0 -1 147424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_534
timestamp 1624015447
transform 1 0 1104 0 -1 148512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_536
timestamp 1624015447
transform 1 0 1104 0 1 148512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_538
timestamp 1624015447
transform 1 0 1104 0 -1 149600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_268_3
timestamp 1624015447
transform 1 0 1380 0 -1 148512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_268_15
timestamp 1624015447
transform 1 0 2484 0 -1 148512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_269_3
timestamp 1624015447
transform 1 0 1380 0 1 148512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_269_15
timestamp 1624015447
transform 1 0 2484 0 1 148512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_270_3
timestamp 1624015447
transform 1 0 1380 0 -1 149600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_270_15
timestamp 1624015447
transform 1 0 2484 0 -1 149600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1509
timestamp 1624015447
transform 1 0 3772 0 -1 148512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1510
timestamp 1624015447
transform 1 0 3772 0 -1 149600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_268_27
timestamp 1624015447
transform 1 0 3588 0 -1 148512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_268_30
timestamp 1624015447
transform 1 0 3864 0 -1 148512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_269_27
timestamp 1624015447
transform 1 0 3588 0 1 148512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_270_27
timestamp 1624015447
transform 1 0 3588 0 -1 149600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_270_30
timestamp 1624015447
transform 1 0 3864 0 -1 149600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_535
timestamp 1624015447
transform -1 0 5152 0 -1 148512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_537
timestamp 1624015447
transform -1 0 5152 0 1 148512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_539
timestamp 1624015447
transform -1 0 5152 0 -1 149600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_268_38
timestamp 1624015447
transform 1 0 4600 0 -1 148512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_269_39
timestamp 1624015447
transform 1 0 4692 0 1 148512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_270_38
timestamp 1624015447
transform 1 0 4600 0 -1 149600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1224
timestamp 1624015447
transform 1 0 84180 0 -1 148512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1226
timestamp 1624015447
transform 1 0 84180 0 1 148512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1228
timestamp 1624015447
transform 1 0 84180 0 -1 149600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_268_906
timestamp 1624015447
transform 1 0 84456 0 -1 148512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_269_906
timestamp 1624015447
transform 1 0 84456 0 1 148512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_270_906
timestamp 1624015447
transform 1 0 84456 0 -1 149600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_268_918
timestamp 1624015447
transform 1 0 85560 0 -1 148512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_268_930
timestamp 1624015447
transform 1 0 86664 0 -1 148512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_269_918
timestamp 1624015447
transform 1 0 85560 0 1 148512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_269_930
timestamp 1624015447
transform 1 0 86664 0 1 148512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_270_918
timestamp 1624015447
transform 1 0 85560 0 -1 149600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_270_930
timestamp 1624015447
transform 1 0 86664 0 -1 149600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1818
timestamp 1624015447
transform 1 0 86848 0 -1 148512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1820
timestamp 1624015447
transform 1 0 86848 0 -1 149600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_268_933
timestamp 1624015447
transform 1 0 86940 0 -1 148512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_268_945
timestamp 1624015447
transform 1 0 88044 0 -1 148512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_269_942
timestamp 1624015447
transform 1 0 87768 0 1 148512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_270_933
timestamp 1624015447
transform 1 0 86940 0 -1 149600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_270_945
timestamp 1624015447
transform 1 0 88044 0 -1 149600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1819
timestamp 1624015447
transform 1 0 89424 0 1 148512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_268_957
timestamp 1624015447
transform 1 0 89148 0 -1 148512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_269_954
timestamp 1624015447
transform 1 0 88872 0 1 148512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_269_961
timestamp 1624015447
transform 1 0 89516 0 1 148512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_270_957
timestamp 1624015447
transform 1 0 89148 0 -1 149600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1225
timestamp 1624015447
transform -1 0 90896 0 -1 148512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1227
timestamp 1624015447
transform -1 0 90896 0 1 148512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1229
timestamp 1624015447
transform -1 0 90896 0 -1 149600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_268_969
timestamp 1624015447
transform 1 0 90252 0 -1 148512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_270_969
timestamp 1624015447
transform 1 0 90252 0 -1 149600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_540
timestamp 1624015447
transform 1 0 1104 0 1 149600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_542
timestamp 1624015447
transform 1 0 1104 0 -1 150688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_544
timestamp 1624015447
transform 1 0 1104 0 1 150688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_271_3
timestamp 1624015447
transform 1 0 1380 0 1 149600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_271_15
timestamp 1624015447
transform 1 0 2484 0 1 149600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_272_3
timestamp 1624015447
transform 1 0 1380 0 -1 150688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_272_15
timestamp 1624015447
transform 1 0 2484 0 -1 150688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_273_3
timestamp 1624015447
transform 1 0 1380 0 1 150688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_273_15
timestamp 1624015447
transform 1 0 2484 0 1 150688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1511
timestamp 1624015447
transform 1 0 3772 0 -1 150688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_271_27
timestamp 1624015447
transform 1 0 3588 0 1 149600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_272_27
timestamp 1624015447
transform 1 0 3588 0 -1 150688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_272_30
timestamp 1624015447
transform 1 0 3864 0 -1 150688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_273_27
timestamp 1624015447
transform 1 0 3588 0 1 150688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_541
timestamp 1624015447
transform -1 0 5152 0 1 149600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_543
timestamp 1624015447
transform -1 0 5152 0 -1 150688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_545
timestamp 1624015447
transform -1 0 5152 0 1 150688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_271_39
timestamp 1624015447
transform 1 0 4692 0 1 149600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_272_38
timestamp 1624015447
transform 1 0 4600 0 -1 150688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_273_39
timestamp 1624015447
transform 1 0 4692 0 1 150688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1230
timestamp 1624015447
transform 1 0 84180 0 1 149600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1232
timestamp 1624015447
transform 1 0 84180 0 -1 150688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1234
timestamp 1624015447
transform 1 0 84180 0 1 150688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_271_906
timestamp 1624015447
transform 1 0 84456 0 1 149600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_272_906
timestamp 1624015447
transform 1 0 84456 0 -1 150688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_273_906
timestamp 1624015447
transform 1 0 84456 0 1 150688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_271_918
timestamp 1624015447
transform 1 0 85560 0 1 149600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_271_930
timestamp 1624015447
transform 1 0 86664 0 1 149600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_272_918
timestamp 1624015447
transform 1 0 85560 0 -1 150688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_272_930
timestamp 1624015447
transform 1 0 86664 0 -1 150688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_273_918
timestamp 1624015447
transform 1 0 85560 0 1 150688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_273_930
timestamp 1624015447
transform 1 0 86664 0 1 150688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1822
timestamp 1624015447
transform 1 0 86848 0 -1 150688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_271_942
timestamp 1624015447
transform 1 0 87768 0 1 149600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_272_933
timestamp 1624015447
transform 1 0 86940 0 -1 150688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_272_945
timestamp 1624015447
transform 1 0 88044 0 -1 150688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_273_942
timestamp 1624015447
transform 1 0 87768 0 1 150688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1821
timestamp 1624015447
transform 1 0 89424 0 1 149600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1823
timestamp 1624015447
transform 1 0 89424 0 1 150688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_271_954
timestamp 1624015447
transform 1 0 88872 0 1 149600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_271_961
timestamp 1624015447
transform 1 0 89516 0 1 149600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_272_957
timestamp 1624015447
transform 1 0 89148 0 -1 150688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_273_954
timestamp 1624015447
transform 1 0 88872 0 1 150688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_273_961
timestamp 1624015447
transform 1 0 89516 0 1 150688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1231
timestamp 1624015447
transform -1 0 90896 0 1 149600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1233
timestamp 1624015447
transform -1 0 90896 0 -1 150688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1235
timestamp 1624015447
transform -1 0 90896 0 1 150688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_272_969
timestamp 1624015447
transform 1 0 90252 0 -1 150688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_546
timestamp 1624015447
transform 1 0 1104 0 -1 151776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_548
timestamp 1624015447
transform 1 0 1104 0 1 151776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_550
timestamp 1624015447
transform 1 0 1104 0 -1 152864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_274_3
timestamp 1624015447
transform 1 0 1380 0 -1 151776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_274_15
timestamp 1624015447
transform 1 0 2484 0 -1 151776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_275_3
timestamp 1624015447
transform 1 0 1380 0 1 151776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_275_15
timestamp 1624015447
transform 1 0 2484 0 1 151776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_276_3
timestamp 1624015447
transform 1 0 1380 0 -1 152864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_276_15
timestamp 1624015447
transform 1 0 2484 0 -1 152864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1512
timestamp 1624015447
transform 1 0 3772 0 -1 151776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1513
timestamp 1624015447
transform 1 0 3772 0 -1 152864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_274_27
timestamp 1624015447
transform 1 0 3588 0 -1 151776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_274_30
timestamp 1624015447
transform 1 0 3864 0 -1 151776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_275_27
timestamp 1624015447
transform 1 0 3588 0 1 151776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_276_27
timestamp 1624015447
transform 1 0 3588 0 -1 152864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_276_30
timestamp 1624015447
transform 1 0 3864 0 -1 152864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_547
timestamp 1624015447
transform -1 0 5152 0 -1 151776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_549
timestamp 1624015447
transform -1 0 5152 0 1 151776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_551
timestamp 1624015447
transform -1 0 5152 0 -1 152864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_274_38
timestamp 1624015447
transform 1 0 4600 0 -1 151776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_275_39
timestamp 1624015447
transform 1 0 4692 0 1 151776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_276_38
timestamp 1624015447
transform 1 0 4600 0 -1 152864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1236
timestamp 1624015447
transform 1 0 84180 0 -1 151776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1238
timestamp 1624015447
transform 1 0 84180 0 1 151776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1240
timestamp 1624015447
transform 1 0 84180 0 -1 152864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_274_906
timestamp 1624015447
transform 1 0 84456 0 -1 151776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_275_906
timestamp 1624015447
transform 1 0 84456 0 1 151776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_276_906
timestamp 1624015447
transform 1 0 84456 0 -1 152864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_274_918
timestamp 1624015447
transform 1 0 85560 0 -1 151776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_274_930
timestamp 1624015447
transform 1 0 86664 0 -1 151776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_275_918
timestamp 1624015447
transform 1 0 85560 0 1 151776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_275_930
timestamp 1624015447
transform 1 0 86664 0 1 151776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_276_918
timestamp 1624015447
transform 1 0 85560 0 -1 152864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_276_930
timestamp 1624015447
transform 1 0 86664 0 -1 152864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1824
timestamp 1624015447
transform 1 0 86848 0 -1 151776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1826
timestamp 1624015447
transform 1 0 86848 0 -1 152864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_274_933
timestamp 1624015447
transform 1 0 86940 0 -1 151776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_274_945
timestamp 1624015447
transform 1 0 88044 0 -1 151776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_275_942
timestamp 1624015447
transform 1 0 87768 0 1 151776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_276_933
timestamp 1624015447
transform 1 0 86940 0 -1 152864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_276_945
timestamp 1624015447
transform 1 0 88044 0 -1 152864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1825
timestamp 1624015447
transform 1 0 89424 0 1 151776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_274_957
timestamp 1624015447
transform 1 0 89148 0 -1 151776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_275_954
timestamp 1624015447
transform 1 0 88872 0 1 151776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_275_961
timestamp 1624015447
transform 1 0 89516 0 1 151776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_276_957
timestamp 1624015447
transform 1 0 89148 0 -1 152864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1237
timestamp 1624015447
transform -1 0 90896 0 -1 151776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1239
timestamp 1624015447
transform -1 0 90896 0 1 151776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1241
timestamp 1624015447
transform -1 0 90896 0 -1 152864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_274_969
timestamp 1624015447
transform 1 0 90252 0 -1 151776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_276_969
timestamp 1624015447
transform 1 0 90252 0 -1 152864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_552
timestamp 1624015447
transform 1 0 1104 0 1 152864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_554
timestamp 1624015447
transform 1 0 1104 0 -1 153952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_556
timestamp 1624015447
transform 1 0 1104 0 1 153952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_277_3
timestamp 1624015447
transform 1 0 1380 0 1 152864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_277_15
timestamp 1624015447
transform 1 0 2484 0 1 152864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_278_3
timestamp 1624015447
transform 1 0 1380 0 -1 153952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_278_15
timestamp 1624015447
transform 1 0 2484 0 -1 153952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_279_3
timestamp 1624015447
transform 1 0 1380 0 1 153952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_279_15
timestamp 1624015447
transform 1 0 2484 0 1 153952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1514
timestamp 1624015447
transform 1 0 3772 0 -1 153952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_277_27
timestamp 1624015447
transform 1 0 3588 0 1 152864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_278_27
timestamp 1624015447
transform 1 0 3588 0 -1 153952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_278_30
timestamp 1624015447
transform 1 0 3864 0 -1 153952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_279_27
timestamp 1624015447
transform 1 0 3588 0 1 153952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_553
timestamp 1624015447
transform -1 0 5152 0 1 152864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_555
timestamp 1624015447
transform -1 0 5152 0 -1 153952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_557
timestamp 1624015447
transform -1 0 5152 0 1 153952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_277_39
timestamp 1624015447
transform 1 0 4692 0 1 152864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_278_38
timestamp 1624015447
transform 1 0 4600 0 -1 153952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_279_39
timestamp 1624015447
transform 1 0 4692 0 1 153952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _10_
timestamp 1624015447
transform 1 0 84640 0 -1 153952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1242
timestamp 1624015447
transform 1 0 84180 0 1 152864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1244
timestamp 1624015447
transform 1 0 84180 0 -1 153952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1246
timestamp 1624015447
transform 1 0 84180 0 1 153952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_277_906
timestamp 1624015447
transform 1 0 84456 0 1 152864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_278_906
timestamp 1624015447
transform 1 0 84456 0 -1 153952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_278_911
timestamp 1624015447
transform 1 0 84916 0 -1 153952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_279_906
timestamp 1624015447
transform 1 0 84456 0 1 153952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_277_918
timestamp 1624015447
transform 1 0 85560 0 1 152864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_277_930
timestamp 1624015447
transform 1 0 86664 0 1 152864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_278_923
timestamp 1624015447
transform 1 0 86020 0 -1 153952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_279_918
timestamp 1624015447
transform 1 0 85560 0 1 153952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_279_930
timestamp 1624015447
transform 1 0 86664 0 1 153952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1828
timestamp 1624015447
transform 1 0 86848 0 -1 153952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_277_942
timestamp 1624015447
transform 1 0 87768 0 1 152864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_278_931
timestamp 1624015447
transform 1 0 86756 0 -1 153952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_278_933
timestamp 1624015447
transform 1 0 86940 0 -1 153952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_278_945
timestamp 1624015447
transform 1 0 88044 0 -1 153952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_279_942
timestamp 1624015447
transform 1 0 87768 0 1 153952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1827
timestamp 1624015447
transform 1 0 89424 0 1 152864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1829
timestamp 1624015447
transform 1 0 89424 0 1 153952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_277_954
timestamp 1624015447
transform 1 0 88872 0 1 152864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_277_961
timestamp 1624015447
transform 1 0 89516 0 1 152864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_278_957
timestamp 1624015447
transform 1 0 89148 0 -1 153952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_279_954
timestamp 1624015447
transform 1 0 88872 0 1 153952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_279_961
timestamp 1624015447
transform 1 0 89516 0 1 153952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1243
timestamp 1624015447
transform -1 0 90896 0 1 152864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1245
timestamp 1624015447
transform -1 0 90896 0 -1 153952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1247
timestamp 1624015447
transform -1 0 90896 0 1 153952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_278_969
timestamp 1624015447
transform 1 0 90252 0 -1 153952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_281_15
timestamp 1624015447
transform 1 0 2484 0 1 155040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_281_3
timestamp 1624015447
transform 1 0 1380 0 1 155040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_280_15
timestamp 1624015447
transform 1 0 2484 0 -1 155040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_280_3
timestamp 1624015447
transform 1 0 1380 0 -1 155040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_560
timestamp 1624015447
transform 1 0 1104 0 1 155040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_558
timestamp 1624015447
transform 1 0 1104 0 -1 155040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_282_15
timestamp 1624015447
transform 1 0 2484 0 -1 156128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_282_3
timestamp 1624015447
transform 1 0 1380 0 -1 156128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_562
timestamp 1624015447
transform 1 0 1104 0 -1 156128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_283_15
timestamp 1624015447
transform 1 0 2484 0 1 156128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_283_3
timestamp 1624015447
transform 1 0 1380 0 1 156128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_564
timestamp 1624015447
transform 1 0 1104 0 1 156128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1515
timestamp 1624015447
transform 1 0 3772 0 -1 155040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1516
timestamp 1624015447
transform 1 0 3772 0 -1 156128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_280_27
timestamp 1624015447
transform 1 0 3588 0 -1 155040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_280_30
timestamp 1624015447
transform 1 0 3864 0 -1 155040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_281_27
timestamp 1624015447
transform 1 0 3588 0 1 155040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_282_27
timestamp 1624015447
transform 1 0 3588 0 -1 156128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_282_30
timestamp 1624015447
transform 1 0 3864 0 -1 156128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_283_27
timestamp 1624015447
transform 1 0 3588 0 1 156128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_559
timestamp 1624015447
transform -1 0 5152 0 -1 155040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_561
timestamp 1624015447
transform -1 0 5152 0 1 155040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_563
timestamp 1624015447
transform -1 0 5152 0 -1 156128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_565
timestamp 1624015447
transform -1 0 5152 0 1 156128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_280_38
timestamp 1624015447
transform 1 0 4600 0 -1 155040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_281_39
timestamp 1624015447
transform 1 0 4692 0 1 155040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_282_38
timestamp 1624015447
transform 1 0 4600 0 -1 156128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_283_39
timestamp 1624015447
transform 1 0 4692 0 1 156128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1248
timestamp 1624015447
transform 1 0 84180 0 -1 155040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1250
timestamp 1624015447
transform 1 0 84180 0 1 155040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1252
timestamp 1624015447
transform 1 0 84180 0 -1 156128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1254
timestamp 1624015447
transform 1 0 84180 0 1 156128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_280_906
timestamp 1624015447
transform 1 0 84456 0 -1 155040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_281_906
timestamp 1624015447
transform 1 0 84456 0 1 155040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_282_906
timestamp 1624015447
transform 1 0 84456 0 -1 156128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_283_906
timestamp 1624015447
transform 1 0 84456 0 1 156128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_280_918
timestamp 1624015447
transform 1 0 85560 0 -1 155040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_280_930
timestamp 1624015447
transform 1 0 86664 0 -1 155040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_281_918
timestamp 1624015447
transform 1 0 85560 0 1 155040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_281_930
timestamp 1624015447
transform 1 0 86664 0 1 155040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_282_918
timestamp 1624015447
transform 1 0 85560 0 -1 156128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_282_930
timestamp 1624015447
transform 1 0 86664 0 -1 156128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_283_918
timestamp 1624015447
transform 1 0 85560 0 1 156128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_283_930
timestamp 1624015447
transform 1 0 86664 0 1 156128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1830
timestamp 1624015447
transform 1 0 86848 0 -1 155040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1832
timestamp 1624015447
transform 1 0 86848 0 -1 156128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_280_933
timestamp 1624015447
transform 1 0 86940 0 -1 155040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_280_945
timestamp 1624015447
transform 1 0 88044 0 -1 155040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_281_942
timestamp 1624015447
transform 1 0 87768 0 1 155040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_282_933
timestamp 1624015447
transform 1 0 86940 0 -1 156128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_282_945
timestamp 1624015447
transform 1 0 88044 0 -1 156128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_283_942
timestamp 1624015447
transform 1 0 87768 0 1 156128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1831
timestamp 1624015447
transform 1 0 89424 0 1 155040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1833
timestamp 1624015447
transform 1 0 89424 0 1 156128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_280_957
timestamp 1624015447
transform 1 0 89148 0 -1 155040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_281_954
timestamp 1624015447
transform 1 0 88872 0 1 155040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_281_961
timestamp 1624015447
transform 1 0 89516 0 1 155040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_282_957
timestamp 1624015447
transform 1 0 89148 0 -1 156128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_283_954
timestamp 1624015447
transform 1 0 88872 0 1 156128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_283_961
timestamp 1624015447
transform 1 0 89516 0 1 156128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1249
timestamp 1624015447
transform -1 0 90896 0 -1 155040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1251
timestamp 1624015447
transform -1 0 90896 0 1 155040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1253
timestamp 1624015447
transform -1 0 90896 0 -1 156128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1255
timestamp 1624015447
transform -1 0 90896 0 1 156128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_280_969
timestamp 1624015447
transform 1 0 90252 0 -1 155040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_282_969
timestamp 1624015447
transform 1 0 90252 0 -1 156128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_566
timestamp 1624015447
transform 1 0 1104 0 -1 157216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_568
timestamp 1624015447
transform 1 0 1104 0 1 157216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_570
timestamp 1624015447
transform 1 0 1104 0 -1 158304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_284_3
timestamp 1624015447
transform 1 0 1380 0 -1 157216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_284_15
timestamp 1624015447
transform 1 0 2484 0 -1 157216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_285_3
timestamp 1624015447
transform 1 0 1380 0 1 157216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_285_15
timestamp 1624015447
transform 1 0 2484 0 1 157216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_286_3
timestamp 1624015447
transform 1 0 1380 0 -1 158304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_286_15
timestamp 1624015447
transform 1 0 2484 0 -1 158304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1517
timestamp 1624015447
transform 1 0 3772 0 -1 157216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1518
timestamp 1624015447
transform 1 0 3772 0 -1 158304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_284_27
timestamp 1624015447
transform 1 0 3588 0 -1 157216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_284_30
timestamp 1624015447
transform 1 0 3864 0 -1 157216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_285_27
timestamp 1624015447
transform 1 0 3588 0 1 157216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_286_27
timestamp 1624015447
transform 1 0 3588 0 -1 158304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_286_30
timestamp 1624015447
transform 1 0 3864 0 -1 158304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_567
timestamp 1624015447
transform -1 0 5152 0 -1 157216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_569
timestamp 1624015447
transform -1 0 5152 0 1 157216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_571
timestamp 1624015447
transform -1 0 5152 0 -1 158304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_284_38
timestamp 1624015447
transform 1 0 4600 0 -1 157216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_285_39
timestamp 1624015447
transform 1 0 4692 0 1 157216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_286_38
timestamp 1624015447
transform 1 0 4600 0 -1 158304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1256
timestamp 1624015447
transform 1 0 84180 0 -1 157216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1258
timestamp 1624015447
transform 1 0 84180 0 1 157216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1260
timestamp 1624015447
transform 1 0 84180 0 -1 158304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_284_906
timestamp 1624015447
transform 1 0 84456 0 -1 157216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_285_906
timestamp 1624015447
transform 1 0 84456 0 1 157216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_286_906
timestamp 1624015447
transform 1 0 84456 0 -1 158304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_284_918
timestamp 1624015447
transform 1 0 85560 0 -1 157216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_284_930
timestamp 1624015447
transform 1 0 86664 0 -1 157216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_285_918
timestamp 1624015447
transform 1 0 85560 0 1 157216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_285_930
timestamp 1624015447
transform 1 0 86664 0 1 157216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_286_918
timestamp 1624015447
transform 1 0 85560 0 -1 158304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_286_930
timestamp 1624015447
transform 1 0 86664 0 -1 158304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1834
timestamp 1624015447
transform 1 0 86848 0 -1 157216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1836
timestamp 1624015447
transform 1 0 86848 0 -1 158304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_284_933
timestamp 1624015447
transform 1 0 86940 0 -1 157216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_284_945
timestamp 1624015447
transform 1 0 88044 0 -1 157216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_285_942
timestamp 1624015447
transform 1 0 87768 0 1 157216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_286_933
timestamp 1624015447
transform 1 0 86940 0 -1 158304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_286_945
timestamp 1624015447
transform 1 0 88044 0 -1 158304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1835
timestamp 1624015447
transform 1 0 89424 0 1 157216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_284_957
timestamp 1624015447
transform 1 0 89148 0 -1 157216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_285_954
timestamp 1624015447
transform 1 0 88872 0 1 157216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_285_961
timestamp 1624015447
transform 1 0 89516 0 1 157216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_286_957
timestamp 1624015447
transform 1 0 89148 0 -1 158304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1257
timestamp 1624015447
transform -1 0 90896 0 -1 157216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1259
timestamp 1624015447
transform -1 0 90896 0 1 157216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1261
timestamp 1624015447
transform -1 0 90896 0 -1 158304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_284_969
timestamp 1624015447
transform 1 0 90252 0 -1 157216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_286_969
timestamp 1624015447
transform 1 0 90252 0 -1 158304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_572
timestamp 1624015447
transform 1 0 1104 0 1 158304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_574
timestamp 1624015447
transform 1 0 1104 0 -1 159392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_576
timestamp 1624015447
transform 1 0 1104 0 1 159392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_287_3
timestamp 1624015447
transform 1 0 1380 0 1 158304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_287_15
timestamp 1624015447
transform 1 0 2484 0 1 158304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_288_3
timestamp 1624015447
transform 1 0 1380 0 -1 159392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_288_15
timestamp 1624015447
transform 1 0 2484 0 -1 159392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_289_3
timestamp 1624015447
transform 1 0 1380 0 1 159392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_289_15
timestamp 1624015447
transform 1 0 2484 0 1 159392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1519
timestamp 1624015447
transform 1 0 3772 0 -1 159392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_287_27
timestamp 1624015447
transform 1 0 3588 0 1 158304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_288_27
timestamp 1624015447
transform 1 0 3588 0 -1 159392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_288_30
timestamp 1624015447
transform 1 0 3864 0 -1 159392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_289_27
timestamp 1624015447
transform 1 0 3588 0 1 159392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_573
timestamp 1624015447
transform -1 0 5152 0 1 158304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_575
timestamp 1624015447
transform -1 0 5152 0 -1 159392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_577
timestamp 1624015447
transform -1 0 5152 0 1 159392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_287_39
timestamp 1624015447
transform 1 0 4692 0 1 158304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_288_38
timestamp 1624015447
transform 1 0 4600 0 -1 159392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_289_39
timestamp 1624015447
transform 1 0 4692 0 1 159392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1262
timestamp 1624015447
transform 1 0 84180 0 1 158304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1264
timestamp 1624015447
transform 1 0 84180 0 -1 159392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1266
timestamp 1624015447
transform 1 0 84180 0 1 159392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_287_906
timestamp 1624015447
transform 1 0 84456 0 1 158304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_288_906
timestamp 1624015447
transform 1 0 84456 0 -1 159392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_289_906
timestamp 1624015447
transform 1 0 84456 0 1 159392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_287_918
timestamp 1624015447
transform 1 0 85560 0 1 158304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_287_930
timestamp 1624015447
transform 1 0 86664 0 1 158304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_288_918
timestamp 1624015447
transform 1 0 85560 0 -1 159392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_288_930
timestamp 1624015447
transform 1 0 86664 0 -1 159392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_289_918
timestamp 1624015447
transform 1 0 85560 0 1 159392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_289_930
timestamp 1624015447
transform 1 0 86664 0 1 159392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1838
timestamp 1624015447
transform 1 0 86848 0 -1 159392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_287_942
timestamp 1624015447
transform 1 0 87768 0 1 158304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_288_933
timestamp 1624015447
transform 1 0 86940 0 -1 159392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_288_945
timestamp 1624015447
transform 1 0 88044 0 -1 159392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_289_942
timestamp 1624015447
transform 1 0 87768 0 1 159392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1837
timestamp 1624015447
transform 1 0 89424 0 1 158304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1839
timestamp 1624015447
transform 1 0 89424 0 1 159392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_287_954
timestamp 1624015447
transform 1 0 88872 0 1 158304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_287_961
timestamp 1624015447
transform 1 0 89516 0 1 158304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_288_957
timestamp 1624015447
transform 1 0 89148 0 -1 159392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_289_954
timestamp 1624015447
transform 1 0 88872 0 1 159392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_289_961
timestamp 1624015447
transform 1 0 89516 0 1 159392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1263
timestamp 1624015447
transform -1 0 90896 0 1 158304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1265
timestamp 1624015447
transform -1 0 90896 0 -1 159392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1267
timestamp 1624015447
transform -1 0 90896 0 1 159392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_288_969
timestamp 1624015447
transform 1 0 90252 0 -1 159392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_578
timestamp 1624015447
transform 1 0 1104 0 -1 160480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_580
timestamp 1624015447
transform 1 0 1104 0 1 160480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_582
timestamp 1624015447
transform 1 0 1104 0 -1 161568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_290_3
timestamp 1624015447
transform 1 0 1380 0 -1 160480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_290_15
timestamp 1624015447
transform 1 0 2484 0 -1 160480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_291_3
timestamp 1624015447
transform 1 0 1380 0 1 160480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_291_15
timestamp 1624015447
transform 1 0 2484 0 1 160480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_292_3
timestamp 1624015447
transform 1 0 1380 0 -1 161568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_292_15
timestamp 1624015447
transform 1 0 2484 0 -1 161568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1520
timestamp 1624015447
transform 1 0 3772 0 -1 160480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1521
timestamp 1624015447
transform 1 0 3772 0 -1 161568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_290_27
timestamp 1624015447
transform 1 0 3588 0 -1 160480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_290_30
timestamp 1624015447
transform 1 0 3864 0 -1 160480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_291_27
timestamp 1624015447
transform 1 0 3588 0 1 160480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_292_27
timestamp 1624015447
transform 1 0 3588 0 -1 161568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_292_30
timestamp 1624015447
transform 1 0 3864 0 -1 161568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_579
timestamp 1624015447
transform -1 0 5152 0 -1 160480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_581
timestamp 1624015447
transform -1 0 5152 0 1 160480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_583
timestamp 1624015447
transform -1 0 5152 0 -1 161568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_290_38
timestamp 1624015447
transform 1 0 4600 0 -1 160480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_291_39
timestamp 1624015447
transform 1 0 4692 0 1 160480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_292_38
timestamp 1624015447
transform 1 0 4600 0 -1 161568
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _14_
timestamp 1624015447
transform -1 0 84732 0 -1 160480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1268
timestamp 1624015447
transform 1 0 84180 0 -1 160480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1270
timestamp 1624015447
transform 1 0 84180 0 1 160480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1272
timestamp 1624015447
transform 1 0 84180 0 -1 161568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_290_909
timestamp 1624015447
transform 1 0 84732 0 -1 160480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_291_906
timestamp 1624015447
transform 1 0 84456 0 1 160480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_292_906
timestamp 1624015447
transform 1 0 84456 0 -1 161568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_290_921
timestamp 1624015447
transform 1 0 85836 0 -1 160480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_290_929
timestamp 1624015447
transform 1 0 86572 0 -1 160480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_291_918
timestamp 1624015447
transform 1 0 85560 0 1 160480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_291_930
timestamp 1624015447
transform 1 0 86664 0 1 160480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_292_918
timestamp 1624015447
transform 1 0 85560 0 -1 161568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_292_930
timestamp 1624015447
transform 1 0 86664 0 -1 161568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1840
timestamp 1624015447
transform 1 0 86848 0 -1 160480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1842
timestamp 1624015447
transform 1 0 86848 0 -1 161568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_290_933
timestamp 1624015447
transform 1 0 86940 0 -1 160480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_290_945
timestamp 1624015447
transform 1 0 88044 0 -1 160480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_291_942
timestamp 1624015447
transform 1 0 87768 0 1 160480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_292_933
timestamp 1624015447
transform 1 0 86940 0 -1 161568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_292_945
timestamp 1624015447
transform 1 0 88044 0 -1 161568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1841
timestamp 1624015447
transform 1 0 89424 0 1 160480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_290_957
timestamp 1624015447
transform 1 0 89148 0 -1 160480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_291_954
timestamp 1624015447
transform 1 0 88872 0 1 160480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_291_961
timestamp 1624015447
transform 1 0 89516 0 1 160480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_292_957
timestamp 1624015447
transform 1 0 89148 0 -1 161568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1269
timestamp 1624015447
transform -1 0 90896 0 -1 160480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1271
timestamp 1624015447
transform -1 0 90896 0 1 160480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1273
timestamp 1624015447
transform -1 0 90896 0 -1 161568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_290_969
timestamp 1624015447
transform 1 0 90252 0 -1 160480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_292_969
timestamp 1624015447
transform 1 0 90252 0 -1 161568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_584
timestamp 1624015447
transform 1 0 1104 0 1 161568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_586
timestamp 1624015447
transform 1 0 1104 0 -1 162656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_588
timestamp 1624015447
transform 1 0 1104 0 1 162656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_293_3
timestamp 1624015447
transform 1 0 1380 0 1 161568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_293_15
timestamp 1624015447
transform 1 0 2484 0 1 161568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_294_3
timestamp 1624015447
transform 1 0 1380 0 -1 162656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_294_15
timestamp 1624015447
transform 1 0 2484 0 -1 162656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_295_3
timestamp 1624015447
transform 1 0 1380 0 1 162656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_295_15
timestamp 1624015447
transform 1 0 2484 0 1 162656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1522
timestamp 1624015447
transform 1 0 3772 0 -1 162656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_293_27
timestamp 1624015447
transform 1 0 3588 0 1 161568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_294_27
timestamp 1624015447
transform 1 0 3588 0 -1 162656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_294_30
timestamp 1624015447
transform 1 0 3864 0 -1 162656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_295_27
timestamp 1624015447
transform 1 0 3588 0 1 162656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_585
timestamp 1624015447
transform -1 0 5152 0 1 161568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_587
timestamp 1624015447
transform -1 0 5152 0 -1 162656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_589
timestamp 1624015447
transform -1 0 5152 0 1 162656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_293_39
timestamp 1624015447
transform 1 0 4692 0 1 161568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_294_38
timestamp 1624015447
transform 1 0 4600 0 -1 162656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_295_39
timestamp 1624015447
transform 1 0 4692 0 1 162656
box -38 -48 222 592
use sky130_fd_sc_hd__buf_8  BUF0_8
timestamp 1624015447
transform 1 0 84456 0 -1 162656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1274
timestamp 1624015447
transform 1 0 84180 0 1 161568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1276
timestamp 1624015447
transform 1 0 84180 0 -1 162656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1278
timestamp 1624015447
transform 1 0 84180 0 1 162656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF0_8_A
timestamp 1624015447
transform 1 0 84640 0 1 161568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_293_906
timestamp 1624015447
transform 1 0 84456 0 1 161568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_293_910
timestamp 1624015447
transform 1 0 84824 0 1 161568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_295_906
timestamp 1624015447
transform 1 0 84456 0 1 162656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_293_922
timestamp 1624015447
transform 1 0 85928 0 1 161568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_294_918
timestamp 1624015447
transform 1 0 85560 0 -1 162656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_294_930
timestamp 1624015447
transform 1 0 86664 0 -1 162656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_295_918
timestamp 1624015447
transform 1 0 85560 0 1 162656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_295_930
timestamp 1624015447
transform 1 0 86664 0 1 162656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1844
timestamp 1624015447
transform 1 0 86848 0 -1 162656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_293_934
timestamp 1624015447
transform 1 0 87032 0 1 161568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_293_946
timestamp 1624015447
transform 1 0 88136 0 1 161568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_294_933
timestamp 1624015447
transform 1 0 86940 0 -1 162656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_294_945
timestamp 1624015447
transform 1 0 88044 0 -1 162656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_295_942
timestamp 1624015447
transform 1 0 87768 0 1 162656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1843
timestamp 1624015447
transform 1 0 89424 0 1 161568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1845
timestamp 1624015447
transform 1 0 89424 0 1 162656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_293_958
timestamp 1624015447
transform 1 0 89240 0 1 161568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_293_961
timestamp 1624015447
transform 1 0 89516 0 1 161568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_294_957
timestamp 1624015447
transform 1 0 89148 0 -1 162656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_295_954
timestamp 1624015447
transform 1 0 88872 0 1 162656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_295_961
timestamp 1624015447
transform 1 0 89516 0 1 162656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1275
timestamp 1624015447
transform -1 0 90896 0 1 161568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1277
timestamp 1624015447
transform -1 0 90896 0 -1 162656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1279
timestamp 1624015447
transform -1 0 90896 0 1 162656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_294_969
timestamp 1624015447
transform 1 0 90252 0 -1 162656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_590
timestamp 1624015447
transform 1 0 1104 0 -1 163744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_592
timestamp 1624015447
transform 1 0 1104 0 1 163744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_594
timestamp 1624015447
transform 1 0 1104 0 -1 164832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_296_3
timestamp 1624015447
transform 1 0 1380 0 -1 163744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_296_15
timestamp 1624015447
transform 1 0 2484 0 -1 163744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_297_3
timestamp 1624015447
transform 1 0 1380 0 1 163744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_297_15
timestamp 1624015447
transform 1 0 2484 0 1 163744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_298_3
timestamp 1624015447
transform 1 0 1380 0 -1 164832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_298_15
timestamp 1624015447
transform 1 0 2484 0 -1 164832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1523
timestamp 1624015447
transform 1 0 3772 0 -1 163744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1524
timestamp 1624015447
transform 1 0 3772 0 -1 164832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_296_27
timestamp 1624015447
transform 1 0 3588 0 -1 163744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_296_30
timestamp 1624015447
transform 1 0 3864 0 -1 163744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_297_27
timestamp 1624015447
transform 1 0 3588 0 1 163744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_298_27
timestamp 1624015447
transform 1 0 3588 0 -1 164832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_298_30
timestamp 1624015447
transform 1 0 3864 0 -1 164832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_591
timestamp 1624015447
transform -1 0 5152 0 -1 163744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_593
timestamp 1624015447
transform -1 0 5152 0 1 163744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_595
timestamp 1624015447
transform -1 0 5152 0 -1 164832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_296_38
timestamp 1624015447
transform 1 0 4600 0 -1 163744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_297_39
timestamp 1624015447
transform 1 0 4692 0 1 163744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_298_38
timestamp 1624015447
transform 1 0 4600 0 -1 164832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1280
timestamp 1624015447
transform 1 0 84180 0 -1 163744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1282
timestamp 1624015447
transform 1 0 84180 0 1 163744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1284
timestamp 1624015447
transform 1 0 84180 0 -1 164832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_296_906
timestamp 1624015447
transform 1 0 84456 0 -1 163744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_297_906
timestamp 1624015447
transform 1 0 84456 0 1 163744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_298_906
timestamp 1624015447
transform 1 0 84456 0 -1 164832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_296_918
timestamp 1624015447
transform 1 0 85560 0 -1 163744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_296_930
timestamp 1624015447
transform 1 0 86664 0 -1 163744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_297_918
timestamp 1624015447
transform 1 0 85560 0 1 163744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_297_930
timestamp 1624015447
transform 1 0 86664 0 1 163744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_298_918
timestamp 1624015447
transform 1 0 85560 0 -1 164832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_298_930
timestamp 1624015447
transform 1 0 86664 0 -1 164832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1846
timestamp 1624015447
transform 1 0 86848 0 -1 163744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1848
timestamp 1624015447
transform 1 0 86848 0 -1 164832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_296_933
timestamp 1624015447
transform 1 0 86940 0 -1 163744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_296_945
timestamp 1624015447
transform 1 0 88044 0 -1 163744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_297_942
timestamp 1624015447
transform 1 0 87768 0 1 163744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_298_933
timestamp 1624015447
transform 1 0 86940 0 -1 164832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_298_945
timestamp 1624015447
transform 1 0 88044 0 -1 164832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1847
timestamp 1624015447
transform 1 0 89424 0 1 163744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_296_957
timestamp 1624015447
transform 1 0 89148 0 -1 163744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_297_954
timestamp 1624015447
transform 1 0 88872 0 1 163744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_297_961
timestamp 1624015447
transform 1 0 89516 0 1 163744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_298_957
timestamp 1624015447
transform 1 0 89148 0 -1 164832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1281
timestamp 1624015447
transform -1 0 90896 0 -1 163744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1283
timestamp 1624015447
transform -1 0 90896 0 1 163744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1285
timestamp 1624015447
transform -1 0 90896 0 -1 164832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_296_969
timestamp 1624015447
transform 1 0 90252 0 -1 163744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_298_969
timestamp 1624015447
transform 1 0 90252 0 -1 164832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_596
timestamp 1624015447
transform 1 0 1104 0 1 164832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_598
timestamp 1624015447
transform 1 0 1104 0 -1 165920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_600
timestamp 1624015447
transform 1 0 1104 0 1 165920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_299_3
timestamp 1624015447
transform 1 0 1380 0 1 164832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_299_15
timestamp 1624015447
transform 1 0 2484 0 1 164832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_300_3
timestamp 1624015447
transform 1 0 1380 0 -1 165920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_300_15
timestamp 1624015447
transform 1 0 2484 0 -1 165920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_301_3
timestamp 1624015447
transform 1 0 1380 0 1 165920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_301_15
timestamp 1624015447
transform 1 0 2484 0 1 165920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1525
timestamp 1624015447
transform 1 0 3772 0 -1 165920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_299_27
timestamp 1624015447
transform 1 0 3588 0 1 164832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_300_27
timestamp 1624015447
transform 1 0 3588 0 -1 165920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_300_30
timestamp 1624015447
transform 1 0 3864 0 -1 165920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_301_27
timestamp 1624015447
transform 1 0 3588 0 1 165920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_597
timestamp 1624015447
transform -1 0 5152 0 1 164832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_599
timestamp 1624015447
transform -1 0 5152 0 -1 165920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_601
timestamp 1624015447
transform -1 0 5152 0 1 165920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_299_39
timestamp 1624015447
transform 1 0 4692 0 1 164832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_300_38
timestamp 1624015447
transform 1 0 4600 0 -1 165920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_301_39
timestamp 1624015447
transform 1 0 4692 0 1 165920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1286
timestamp 1624015447
transform 1 0 84180 0 1 164832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1288
timestamp 1624015447
transform 1 0 84180 0 -1 165920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1290
timestamp 1624015447
transform 1 0 84180 0 1 165920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_299_906
timestamp 1624015447
transform 1 0 84456 0 1 164832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_300_906
timestamp 1624015447
transform 1 0 84456 0 -1 165920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_301_906
timestamp 1624015447
transform 1 0 84456 0 1 165920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_299_918
timestamp 1624015447
transform 1 0 85560 0 1 164832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_299_930
timestamp 1624015447
transform 1 0 86664 0 1 164832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_300_918
timestamp 1624015447
transform 1 0 85560 0 -1 165920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_300_930
timestamp 1624015447
transform 1 0 86664 0 -1 165920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_301_918
timestamp 1624015447
transform 1 0 85560 0 1 165920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_301_930
timestamp 1624015447
transform 1 0 86664 0 1 165920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1850
timestamp 1624015447
transform 1 0 86848 0 -1 165920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_299_942
timestamp 1624015447
transform 1 0 87768 0 1 164832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_300_933
timestamp 1624015447
transform 1 0 86940 0 -1 165920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_300_945
timestamp 1624015447
transform 1 0 88044 0 -1 165920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_301_942
timestamp 1624015447
transform 1 0 87768 0 1 165920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1849
timestamp 1624015447
transform 1 0 89424 0 1 164832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1851
timestamp 1624015447
transform 1 0 89424 0 1 165920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_299_954
timestamp 1624015447
transform 1 0 88872 0 1 164832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_299_961
timestamp 1624015447
transform 1 0 89516 0 1 164832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_300_957
timestamp 1624015447
transform 1 0 89148 0 -1 165920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_301_954
timestamp 1624015447
transform 1 0 88872 0 1 165920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_301_961
timestamp 1624015447
transform 1 0 89516 0 1 165920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1287
timestamp 1624015447
transform -1 0 90896 0 1 164832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1289
timestamp 1624015447
transform -1 0 90896 0 -1 165920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1291
timestamp 1624015447
transform -1 0 90896 0 1 165920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_300_969
timestamp 1624015447
transform 1 0 90252 0 -1 165920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_303_15
timestamp 1624015447
transform 1 0 2484 0 1 167008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_303_3
timestamp 1624015447
transform 1 0 1380 0 1 167008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_302_15
timestamp 1624015447
transform 1 0 2484 0 -1 167008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_302_3
timestamp 1624015447
transform 1 0 1380 0 -1 167008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_604
timestamp 1624015447
transform 1 0 1104 0 1 167008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_602
timestamp 1624015447
transform 1 0 1104 0 -1 167008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_304_15
timestamp 1624015447
transform 1 0 2484 0 -1 168096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_304_3
timestamp 1624015447
transform 1 0 1380 0 -1 168096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_606
timestamp 1624015447
transform 1 0 1104 0 -1 168096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_305_15
timestamp 1624015447
transform 1 0 2484 0 1 168096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_305_3
timestamp 1624015447
transform 1 0 1380 0 1 168096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_608
timestamp 1624015447
transform 1 0 1104 0 1 168096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1526
timestamp 1624015447
transform 1 0 3772 0 -1 167008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1527
timestamp 1624015447
transform 1 0 3772 0 -1 168096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_302_27
timestamp 1624015447
transform 1 0 3588 0 -1 167008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_302_30
timestamp 1624015447
transform 1 0 3864 0 -1 167008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_303_27
timestamp 1624015447
transform 1 0 3588 0 1 167008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_304_27
timestamp 1624015447
transform 1 0 3588 0 -1 168096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_304_30
timestamp 1624015447
transform 1 0 3864 0 -1 168096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_305_27
timestamp 1624015447
transform 1 0 3588 0 1 168096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_603
timestamp 1624015447
transform -1 0 5152 0 -1 167008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_605
timestamp 1624015447
transform -1 0 5152 0 1 167008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_607
timestamp 1624015447
transform -1 0 5152 0 -1 168096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_609
timestamp 1624015447
transform -1 0 5152 0 1 168096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_302_38
timestamp 1624015447
transform 1 0 4600 0 -1 167008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_303_39
timestamp 1624015447
transform 1 0 4692 0 1 167008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_304_38
timestamp 1624015447
transform 1 0 4600 0 -1 168096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_305_39
timestamp 1624015447
transform 1 0 4692 0 1 168096
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _11_
timestamp 1624015447
transform -1 0 84732 0 1 167008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1292
timestamp 1624015447
transform 1 0 84180 0 -1 167008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1294
timestamp 1624015447
transform 1 0 84180 0 1 167008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1296
timestamp 1624015447
transform 1 0 84180 0 -1 168096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1298
timestamp 1624015447
transform 1 0 84180 0 1 168096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_302_906
timestamp 1624015447
transform 1 0 84456 0 -1 167008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_303_909
timestamp 1624015447
transform 1 0 84732 0 1 167008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_304_906
timestamp 1624015447
transform 1 0 84456 0 -1 168096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_305_906
timestamp 1624015447
transform 1 0 84456 0 1 168096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_302_918
timestamp 1624015447
transform 1 0 85560 0 -1 167008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_302_930
timestamp 1624015447
transform 1 0 86664 0 -1 167008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_303_921
timestamp 1624015447
transform 1 0 85836 0 1 167008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_304_918
timestamp 1624015447
transform 1 0 85560 0 -1 168096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_304_930
timestamp 1624015447
transform 1 0 86664 0 -1 168096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_305_918
timestamp 1624015447
transform 1 0 85560 0 1 168096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_305_930
timestamp 1624015447
transform 1 0 86664 0 1 168096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1852
timestamp 1624015447
transform 1 0 86848 0 -1 167008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1854
timestamp 1624015447
transform 1 0 86848 0 -1 168096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_302_933
timestamp 1624015447
transform 1 0 86940 0 -1 167008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_302_945
timestamp 1624015447
transform 1 0 88044 0 -1 167008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_303_933
timestamp 1624015447
transform 1 0 86940 0 1 167008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_303_945
timestamp 1624015447
transform 1 0 88044 0 1 167008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_304_933
timestamp 1624015447
transform 1 0 86940 0 -1 168096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_304_945
timestamp 1624015447
transform 1 0 88044 0 -1 168096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_305_942
timestamp 1624015447
transform 1 0 87768 0 1 168096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1853
timestamp 1624015447
transform 1 0 89424 0 1 167008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1855
timestamp 1624015447
transform 1 0 89424 0 1 168096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_302_957
timestamp 1624015447
transform 1 0 89148 0 -1 167008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_303_957
timestamp 1624015447
transform 1 0 89148 0 1 167008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_303_961
timestamp 1624015447
transform 1 0 89516 0 1 167008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_304_957
timestamp 1624015447
transform 1 0 89148 0 -1 168096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_305_954
timestamp 1624015447
transform 1 0 88872 0 1 168096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_305_961
timestamp 1624015447
transform 1 0 89516 0 1 168096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1293
timestamp 1624015447
transform -1 0 90896 0 -1 167008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1295
timestamp 1624015447
transform -1 0 90896 0 1 167008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1297
timestamp 1624015447
transform -1 0 90896 0 -1 168096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1299
timestamp 1624015447
transform -1 0 90896 0 1 168096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_302_969
timestamp 1624015447
transform 1 0 90252 0 -1 167008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_304_969
timestamp 1624015447
transform 1 0 90252 0 -1 168096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_610
timestamp 1624015447
transform 1 0 1104 0 -1 169184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_612
timestamp 1624015447
transform 1 0 1104 0 1 169184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_614
timestamp 1624015447
transform 1 0 1104 0 -1 170272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_306_3
timestamp 1624015447
transform 1 0 1380 0 -1 169184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_306_15
timestamp 1624015447
transform 1 0 2484 0 -1 169184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_307_3
timestamp 1624015447
transform 1 0 1380 0 1 169184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_307_15
timestamp 1624015447
transform 1 0 2484 0 1 169184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_308_3
timestamp 1624015447
transform 1 0 1380 0 -1 170272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_308_15
timestamp 1624015447
transform 1 0 2484 0 -1 170272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1528
timestamp 1624015447
transform 1 0 3772 0 -1 169184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1529
timestamp 1624015447
transform 1 0 3772 0 -1 170272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_306_27
timestamp 1624015447
transform 1 0 3588 0 -1 169184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_306_30
timestamp 1624015447
transform 1 0 3864 0 -1 169184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_307_27
timestamp 1624015447
transform 1 0 3588 0 1 169184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_308_27
timestamp 1624015447
transform 1 0 3588 0 -1 170272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_308_30
timestamp 1624015447
transform 1 0 3864 0 -1 170272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_611
timestamp 1624015447
transform -1 0 5152 0 -1 169184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_613
timestamp 1624015447
transform -1 0 5152 0 1 169184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_615
timestamp 1624015447
transform -1 0 5152 0 -1 170272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_306_38
timestamp 1624015447
transform 1 0 4600 0 -1 169184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_307_39
timestamp 1624015447
transform 1 0 4692 0 1 169184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_308_38
timestamp 1624015447
transform 1 0 4600 0 -1 170272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1300
timestamp 1624015447
transform 1 0 84180 0 -1 169184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1302
timestamp 1624015447
transform 1 0 84180 0 1 169184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1304
timestamp 1624015447
transform 1 0 84180 0 -1 170272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_306_906
timestamp 1624015447
transform 1 0 84456 0 -1 169184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_307_906
timestamp 1624015447
transform 1 0 84456 0 1 169184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_308_906
timestamp 1624015447
transform 1 0 84456 0 -1 170272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_306_918
timestamp 1624015447
transform 1 0 85560 0 -1 169184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_306_930
timestamp 1624015447
transform 1 0 86664 0 -1 169184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_307_918
timestamp 1624015447
transform 1 0 85560 0 1 169184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_307_930
timestamp 1624015447
transform 1 0 86664 0 1 169184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_308_918
timestamp 1624015447
transform 1 0 85560 0 -1 170272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_308_930
timestamp 1624015447
transform 1 0 86664 0 -1 170272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1856
timestamp 1624015447
transform 1 0 86848 0 -1 169184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1858
timestamp 1624015447
transform 1 0 86848 0 -1 170272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_306_933
timestamp 1624015447
transform 1 0 86940 0 -1 169184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_306_945
timestamp 1624015447
transform 1 0 88044 0 -1 169184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_307_942
timestamp 1624015447
transform 1 0 87768 0 1 169184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_308_933
timestamp 1624015447
transform 1 0 86940 0 -1 170272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_308_945
timestamp 1624015447
transform 1 0 88044 0 -1 170272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1857
timestamp 1624015447
transform 1 0 89424 0 1 169184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_306_957
timestamp 1624015447
transform 1 0 89148 0 -1 169184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_307_954
timestamp 1624015447
transform 1 0 88872 0 1 169184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_307_961
timestamp 1624015447
transform 1 0 89516 0 1 169184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_308_957
timestamp 1624015447
transform 1 0 89148 0 -1 170272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1301
timestamp 1624015447
transform -1 0 90896 0 -1 169184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1303
timestamp 1624015447
transform -1 0 90896 0 1 169184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1305
timestamp 1624015447
transform -1 0 90896 0 -1 170272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_306_969
timestamp 1624015447
transform 1 0 90252 0 -1 169184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_308_969
timestamp 1624015447
transform 1 0 90252 0 -1 170272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_616
timestamp 1624015447
transform 1 0 1104 0 1 170272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_618
timestamp 1624015447
transform 1 0 1104 0 -1 171360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_620
timestamp 1624015447
transform 1 0 1104 0 1 171360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_309_3
timestamp 1624015447
transform 1 0 1380 0 1 170272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_309_15
timestamp 1624015447
transform 1 0 2484 0 1 170272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_310_3
timestamp 1624015447
transform 1 0 1380 0 -1 171360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_310_15
timestamp 1624015447
transform 1 0 2484 0 -1 171360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_311_3
timestamp 1624015447
transform 1 0 1380 0 1 171360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_311_15
timestamp 1624015447
transform 1 0 2484 0 1 171360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1530
timestamp 1624015447
transform 1 0 3772 0 -1 171360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_309_27
timestamp 1624015447
transform 1 0 3588 0 1 170272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_310_27
timestamp 1624015447
transform 1 0 3588 0 -1 171360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_310_30
timestamp 1624015447
transform 1 0 3864 0 -1 171360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_311_27
timestamp 1624015447
transform 1 0 3588 0 1 171360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_617
timestamp 1624015447
transform -1 0 5152 0 1 170272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_619
timestamp 1624015447
transform -1 0 5152 0 -1 171360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_621
timestamp 1624015447
transform -1 0 5152 0 1 171360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_309_39
timestamp 1624015447
transform 1 0 4692 0 1 170272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_310_38
timestamp 1624015447
transform 1 0 4600 0 -1 171360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_311_39
timestamp 1624015447
transform 1 0 4692 0 1 171360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1306
timestamp 1624015447
transform 1 0 84180 0 1 170272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1308
timestamp 1624015447
transform 1 0 84180 0 -1 171360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1310
timestamp 1624015447
transform 1 0 84180 0 1 171360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_309_906
timestamp 1624015447
transform 1 0 84456 0 1 170272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_310_906
timestamp 1624015447
transform 1 0 84456 0 -1 171360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_311_906
timestamp 1624015447
transform 1 0 84456 0 1 171360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_309_918
timestamp 1624015447
transform 1 0 85560 0 1 170272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_309_930
timestamp 1624015447
transform 1 0 86664 0 1 170272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_310_918
timestamp 1624015447
transform 1 0 85560 0 -1 171360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_310_930
timestamp 1624015447
transform 1 0 86664 0 -1 171360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_311_918
timestamp 1624015447
transform 1 0 85560 0 1 171360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_311_930
timestamp 1624015447
transform 1 0 86664 0 1 171360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1860
timestamp 1624015447
transform 1 0 86848 0 -1 171360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_309_942
timestamp 1624015447
transform 1 0 87768 0 1 170272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_310_933
timestamp 1624015447
transform 1 0 86940 0 -1 171360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_310_945
timestamp 1624015447
transform 1 0 88044 0 -1 171360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_311_942
timestamp 1624015447
transform 1 0 87768 0 1 171360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1859
timestamp 1624015447
transform 1 0 89424 0 1 170272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1861
timestamp 1624015447
transform 1 0 89424 0 1 171360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_309_954
timestamp 1624015447
transform 1 0 88872 0 1 170272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_309_961
timestamp 1624015447
transform 1 0 89516 0 1 170272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_310_957
timestamp 1624015447
transform 1 0 89148 0 -1 171360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_311_954
timestamp 1624015447
transform 1 0 88872 0 1 171360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_311_961
timestamp 1624015447
transform 1 0 89516 0 1 171360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1307
timestamp 1624015447
transform -1 0 90896 0 1 170272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1309
timestamp 1624015447
transform -1 0 90896 0 -1 171360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1311
timestamp 1624015447
transform -1 0 90896 0 1 171360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_310_969
timestamp 1624015447
transform 1 0 90252 0 -1 171360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_622
timestamp 1624015447
transform 1 0 1104 0 -1 172448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_624
timestamp 1624015447
transform 1 0 1104 0 1 172448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_626
timestamp 1624015447
transform 1 0 1104 0 -1 173536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_312_3
timestamp 1624015447
transform 1 0 1380 0 -1 172448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_312_15
timestamp 1624015447
transform 1 0 2484 0 -1 172448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_313_3
timestamp 1624015447
transform 1 0 1380 0 1 172448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_313_15
timestamp 1624015447
transform 1 0 2484 0 1 172448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_314_3
timestamp 1624015447
transform 1 0 1380 0 -1 173536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_314_15
timestamp 1624015447
transform 1 0 2484 0 -1 173536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1531
timestamp 1624015447
transform 1 0 3772 0 -1 172448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1532
timestamp 1624015447
transform 1 0 3772 0 -1 173536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_312_27
timestamp 1624015447
transform 1 0 3588 0 -1 172448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_312_30
timestamp 1624015447
transform 1 0 3864 0 -1 172448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_313_27
timestamp 1624015447
transform 1 0 3588 0 1 172448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_314_27
timestamp 1624015447
transform 1 0 3588 0 -1 173536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_314_30
timestamp 1624015447
transform 1 0 3864 0 -1 173536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_623
timestamp 1624015447
transform -1 0 5152 0 -1 172448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_625
timestamp 1624015447
transform -1 0 5152 0 1 172448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_627
timestamp 1624015447
transform -1 0 5152 0 -1 173536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_312_38
timestamp 1624015447
transform 1 0 4600 0 -1 172448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_313_39
timestamp 1624015447
transform 1 0 4692 0 1 172448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_314_38
timestamp 1624015447
transform 1 0 4600 0 -1 173536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1312
timestamp 1624015447
transform 1 0 84180 0 -1 172448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1314
timestamp 1624015447
transform 1 0 84180 0 1 172448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1316
timestamp 1624015447
transform 1 0 84180 0 -1 173536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_312_906
timestamp 1624015447
transform 1 0 84456 0 -1 172448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_313_906
timestamp 1624015447
transform 1 0 84456 0 1 172448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_314_906
timestamp 1624015447
transform 1 0 84456 0 -1 173536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_312_918
timestamp 1624015447
transform 1 0 85560 0 -1 172448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_312_930
timestamp 1624015447
transform 1 0 86664 0 -1 172448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_313_918
timestamp 1624015447
transform 1 0 85560 0 1 172448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_313_930
timestamp 1624015447
transform 1 0 86664 0 1 172448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_314_918
timestamp 1624015447
transform 1 0 85560 0 -1 173536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_314_930
timestamp 1624015447
transform 1 0 86664 0 -1 173536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1862
timestamp 1624015447
transform 1 0 86848 0 -1 172448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1864
timestamp 1624015447
transform 1 0 86848 0 -1 173536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_312_933
timestamp 1624015447
transform 1 0 86940 0 -1 172448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_312_945
timestamp 1624015447
transform 1 0 88044 0 -1 172448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_313_942
timestamp 1624015447
transform 1 0 87768 0 1 172448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_314_933
timestamp 1624015447
transform 1 0 86940 0 -1 173536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_314_945
timestamp 1624015447
transform 1 0 88044 0 -1 173536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1863
timestamp 1624015447
transform 1 0 89424 0 1 172448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_312_957
timestamp 1624015447
transform 1 0 89148 0 -1 172448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_313_954
timestamp 1624015447
transform 1 0 88872 0 1 172448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_313_961
timestamp 1624015447
transform 1 0 89516 0 1 172448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_314_957
timestamp 1624015447
transform 1 0 89148 0 -1 173536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1313
timestamp 1624015447
transform -1 0 90896 0 -1 172448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1315
timestamp 1624015447
transform -1 0 90896 0 1 172448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1317
timestamp 1624015447
transform -1 0 90896 0 -1 173536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_312_969
timestamp 1624015447
transform 1 0 90252 0 -1 172448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_314_969
timestamp 1624015447
transform 1 0 90252 0 -1 173536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_628
timestamp 1624015447
transform 1 0 1104 0 1 173536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_630
timestamp 1624015447
transform 1 0 1104 0 -1 174624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_632
timestamp 1624015447
transform 1 0 1104 0 1 174624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_315_3
timestamp 1624015447
transform 1 0 1380 0 1 173536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_315_15
timestamp 1624015447
transform 1 0 2484 0 1 173536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_316_3
timestamp 1624015447
transform 1 0 1380 0 -1 174624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_316_15
timestamp 1624015447
transform 1 0 2484 0 -1 174624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_317_3
timestamp 1624015447
transform 1 0 1380 0 1 174624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_317_15
timestamp 1624015447
transform 1 0 2484 0 1 174624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1533
timestamp 1624015447
transform 1 0 3772 0 -1 174624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_315_27
timestamp 1624015447
transform 1 0 3588 0 1 173536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_316_27
timestamp 1624015447
transform 1 0 3588 0 -1 174624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_316_30
timestamp 1624015447
transform 1 0 3864 0 -1 174624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_317_27
timestamp 1624015447
transform 1 0 3588 0 1 174624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_629
timestamp 1624015447
transform -1 0 5152 0 1 173536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_631
timestamp 1624015447
transform -1 0 5152 0 -1 174624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_633
timestamp 1624015447
transform -1 0 5152 0 1 174624
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_addr0[1]
timestamp 1624015447
transform -1 0 4876 0 -1 174624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_315_39
timestamp 1624015447
transform 1 0 4692 0 1 173536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_316_38
timestamp 1624015447
transform 1 0 4600 0 -1 174624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_317_39
timestamp 1624015447
transform 1 0 4692 0 1 174624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1318
timestamp 1624015447
transform 1 0 84180 0 1 173536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1320
timestamp 1624015447
transform 1 0 84180 0 -1 174624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1322
timestamp 1624015447
transform 1 0 84180 0 1 174624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_315_906
timestamp 1624015447
transform 1 0 84456 0 1 173536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_316_906
timestamp 1624015447
transform 1 0 84456 0 -1 174624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_317_906
timestamp 1624015447
transform 1 0 84456 0 1 174624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_315_918
timestamp 1624015447
transform 1 0 85560 0 1 173536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_315_930
timestamp 1624015447
transform 1 0 86664 0 1 173536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_316_918
timestamp 1624015447
transform 1 0 85560 0 -1 174624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_316_930
timestamp 1624015447
transform 1 0 86664 0 -1 174624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_317_918
timestamp 1624015447
transform 1 0 85560 0 1 174624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_317_930
timestamp 1624015447
transform 1 0 86664 0 1 174624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1866
timestamp 1624015447
transform 1 0 86848 0 -1 174624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_315_942
timestamp 1624015447
transform 1 0 87768 0 1 173536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_316_933
timestamp 1624015447
transform 1 0 86940 0 -1 174624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_316_945
timestamp 1624015447
transform 1 0 88044 0 -1 174624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_317_942
timestamp 1624015447
transform 1 0 87768 0 1 174624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1865
timestamp 1624015447
transform 1 0 89424 0 1 173536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1867
timestamp 1624015447
transform 1 0 89424 0 1 174624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_315_954
timestamp 1624015447
transform 1 0 88872 0 1 173536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_315_961
timestamp 1624015447
transform 1 0 89516 0 1 173536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_316_957
timestamp 1624015447
transform 1 0 89148 0 -1 174624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_317_954
timestamp 1624015447
transform 1 0 88872 0 1 174624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_317_961
timestamp 1624015447
transform 1 0 89516 0 1 174624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1319
timestamp 1624015447
transform -1 0 90896 0 1 173536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1321
timestamp 1624015447
transform -1 0 90896 0 -1 174624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1323
timestamp 1624015447
transform -1 0 90896 0 1 174624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_316_969
timestamp 1624015447
transform 1 0 90252 0 -1 174624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_634
timestamp 1624015447
transform 1 0 1104 0 -1 175712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_636
timestamp 1624015447
transform 1 0 1104 0 1 175712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_638
timestamp 1624015447
transform 1 0 1104 0 -1 176800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_318_3
timestamp 1624015447
transform 1 0 1380 0 -1 175712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_318_15
timestamp 1624015447
transform 1 0 2484 0 -1 175712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_319_3
timestamp 1624015447
transform 1 0 1380 0 1 175712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_319_15
timestamp 1624015447
transform 1 0 2484 0 1 175712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_320_3
timestamp 1624015447
transform 1 0 1380 0 -1 176800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_320_15
timestamp 1624015447
transform 1 0 2484 0 -1 176800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1534
timestamp 1624015447
transform 1 0 3772 0 -1 175712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1535
timestamp 1624015447
transform 1 0 3772 0 -1 176800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_318_27
timestamp 1624015447
transform 1 0 3588 0 -1 175712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_318_30
timestamp 1624015447
transform 1 0 3864 0 -1 175712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_319_27
timestamp 1624015447
transform 1 0 3588 0 1 175712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_320_27
timestamp 1624015447
transform 1 0 3588 0 -1 176800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_320_30
timestamp 1624015447
transform 1 0 3864 0 -1 176800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_635
timestamp 1624015447
transform -1 0 5152 0 -1 175712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_637
timestamp 1624015447
transform -1 0 5152 0 1 175712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_639
timestamp 1624015447
transform -1 0 5152 0 -1 176800
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_addr0[2]
timestamp 1624015447
transform -1 0 4876 0 1 175712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_318_38
timestamp 1624015447
transform 1 0 4600 0 -1 175712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_320_38
timestamp 1624015447
transform 1 0 4600 0 -1 176800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1324
timestamp 1624015447
transform 1 0 84180 0 -1 175712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1326
timestamp 1624015447
transform 1 0 84180 0 1 175712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1328
timestamp 1624015447
transform 1 0 84180 0 -1 176800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_318_906
timestamp 1624015447
transform 1 0 84456 0 -1 175712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_319_906
timestamp 1624015447
transform 1 0 84456 0 1 175712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_320_906
timestamp 1624015447
transform 1 0 84456 0 -1 176800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_318_918
timestamp 1624015447
transform 1 0 85560 0 -1 175712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_318_930
timestamp 1624015447
transform 1 0 86664 0 -1 175712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_319_918
timestamp 1624015447
transform 1 0 85560 0 1 175712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_319_930
timestamp 1624015447
transform 1 0 86664 0 1 175712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_320_918
timestamp 1624015447
transform 1 0 85560 0 -1 176800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_320_930
timestamp 1624015447
transform 1 0 86664 0 -1 176800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1868
timestamp 1624015447
transform 1 0 86848 0 -1 175712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1870
timestamp 1624015447
transform 1 0 86848 0 -1 176800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_318_933
timestamp 1624015447
transform 1 0 86940 0 -1 175712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_318_945
timestamp 1624015447
transform 1 0 88044 0 -1 175712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_319_942
timestamp 1624015447
transform 1 0 87768 0 1 175712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_320_933
timestamp 1624015447
transform 1 0 86940 0 -1 176800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_320_945
timestamp 1624015447
transform 1 0 88044 0 -1 176800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1869
timestamp 1624015447
transform 1 0 89424 0 1 175712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_318_957
timestamp 1624015447
transform 1 0 89148 0 -1 175712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_319_954
timestamp 1624015447
transform 1 0 88872 0 1 175712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_319_961
timestamp 1624015447
transform 1 0 89516 0 1 175712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_320_957
timestamp 1624015447
transform 1 0 89148 0 -1 176800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1325
timestamp 1624015447
transform -1 0 90896 0 -1 175712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1327
timestamp 1624015447
transform -1 0 90896 0 1 175712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1329
timestamp 1624015447
transform -1 0 90896 0 -1 176800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_318_969
timestamp 1624015447
transform 1 0 90252 0 -1 175712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_320_969
timestamp 1624015447
transform 1 0 90252 0 -1 176800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_640
timestamp 1624015447
transform 1 0 1104 0 1 176800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_642
timestamp 1624015447
transform 1 0 1104 0 -1 177888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_644
timestamp 1624015447
transform 1 0 1104 0 1 177888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_321_3
timestamp 1624015447
transform 1 0 1380 0 1 176800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_321_15
timestamp 1624015447
transform 1 0 2484 0 1 176800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_322_3
timestamp 1624015447
transform 1 0 1380 0 -1 177888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_322_15
timestamp 1624015447
transform 1 0 2484 0 -1 177888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_323_3
timestamp 1624015447
transform 1 0 1380 0 1 177888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_323_15
timestamp 1624015447
transform 1 0 2484 0 1 177888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1536
timestamp 1624015447
transform 1 0 3772 0 -1 177888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_321_27
timestamp 1624015447
transform 1 0 3588 0 1 176800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_322_27
timestamp 1624015447
transform 1 0 3588 0 -1 177888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_322_30
timestamp 1624015447
transform 1 0 3864 0 -1 177888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_323_27
timestamp 1624015447
transform 1 0 3588 0 1 177888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_641
timestamp 1624015447
transform -1 0 5152 0 1 176800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_643
timestamp 1624015447
transform -1 0 5152 0 -1 177888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_645
timestamp 1624015447
transform -1 0 5152 0 1 177888
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_addr0[3]
timestamp 1624015447
transform -1 0 4876 0 1 176800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_322_38
timestamp 1624015447
transform 1 0 4600 0 -1 177888
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_323_39
timestamp 1624015447
transform 1 0 4692 0 1 177888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1330
timestamp 1624015447
transform 1 0 84180 0 1 176800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1332
timestamp 1624015447
transform 1 0 84180 0 -1 177888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1334
timestamp 1624015447
transform 1 0 84180 0 1 177888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_321_906
timestamp 1624015447
transform 1 0 84456 0 1 176800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_322_906
timestamp 1624015447
transform 1 0 84456 0 -1 177888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_323_906
timestamp 1624015447
transform 1 0 84456 0 1 177888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_321_918
timestamp 1624015447
transform 1 0 85560 0 1 176800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_321_930
timestamp 1624015447
transform 1 0 86664 0 1 176800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_322_918
timestamp 1624015447
transform 1 0 85560 0 -1 177888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_322_930
timestamp 1624015447
transform 1 0 86664 0 -1 177888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_323_918
timestamp 1624015447
transform 1 0 85560 0 1 177888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_323_930
timestamp 1624015447
transform 1 0 86664 0 1 177888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1872
timestamp 1624015447
transform 1 0 86848 0 -1 177888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_321_942
timestamp 1624015447
transform 1 0 87768 0 1 176800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_322_933
timestamp 1624015447
transform 1 0 86940 0 -1 177888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_322_945
timestamp 1624015447
transform 1 0 88044 0 -1 177888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_323_942
timestamp 1624015447
transform 1 0 87768 0 1 177888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1871
timestamp 1624015447
transform 1 0 89424 0 1 176800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1873
timestamp 1624015447
transform 1 0 89424 0 1 177888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_321_954
timestamp 1624015447
transform 1 0 88872 0 1 176800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_321_961
timestamp 1624015447
transform 1 0 89516 0 1 176800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_322_957
timestamp 1624015447
transform 1 0 89148 0 -1 177888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_323_954
timestamp 1624015447
transform 1 0 88872 0 1 177888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_323_961
timestamp 1624015447
transform 1 0 89516 0 1 177888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1331
timestamp 1624015447
transform -1 0 90896 0 1 176800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1333
timestamp 1624015447
transform -1 0 90896 0 -1 177888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1335
timestamp 1624015447
transform -1 0 90896 0 1 177888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_322_969
timestamp 1624015447
transform 1 0 90252 0 -1 177888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_325_15
timestamp 1624015447
transform 1 0 2484 0 1 178976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_325_3
timestamp 1624015447
transform 1 0 1380 0 1 178976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_324_15
timestamp 1624015447
transform 1 0 2484 0 -1 178976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_324_3
timestamp 1624015447
transform 1 0 1380 0 -1 178976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_648
timestamp 1624015447
transform 1 0 1104 0 1 178976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_646
timestamp 1624015447
transform 1 0 1104 0 -1 178976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_326_15
timestamp 1624015447
transform 1 0 2484 0 -1 180064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_326_3
timestamp 1624015447
transform 1 0 1380 0 -1 180064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_650
timestamp 1624015447
transform 1 0 1104 0 -1 180064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_327_15
timestamp 1624015447
transform 1 0 2484 0 1 180064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_327_3
timestamp 1624015447
transform 1 0 1380 0 1 180064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_652
timestamp 1624015447
transform 1 0 1104 0 1 180064
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1537
timestamp 1624015447
transform 1 0 3772 0 -1 178976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1538
timestamp 1624015447
transform 1 0 3772 0 -1 180064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_324_27
timestamp 1624015447
transform 1 0 3588 0 -1 178976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_324_30
timestamp 1624015447
transform 1 0 3864 0 -1 178976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_325_27
timestamp 1624015447
transform 1 0 3588 0 1 178976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_326_27
timestamp 1624015447
transform 1 0 3588 0 -1 180064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_326_30
timestamp 1624015447
transform 1 0 3864 0 -1 180064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_327_27
timestamp 1624015447
transform 1 0 3588 0 1 180064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_647
timestamp 1624015447
transform -1 0 5152 0 -1 178976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_649
timestamp 1624015447
transform -1 0 5152 0 1 178976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_651
timestamp 1624015447
transform -1 0 5152 0 -1 180064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_653
timestamp 1624015447
transform -1 0 5152 0 1 180064
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_addr0[4]
timestamp 1624015447
transform -1 0 4876 0 1 178976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_addr0[5]
timestamp 1624015447
transform -1 0 4876 0 1 180064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_324_38
timestamp 1624015447
transform 1 0 4600 0 -1 178976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_326_38
timestamp 1624015447
transform 1 0 4600 0 -1 180064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _13_
timestamp 1624015447
transform -1 0 84732 0 -1 180064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1336
timestamp 1624015447
transform 1 0 84180 0 -1 178976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1338
timestamp 1624015447
transform 1 0 84180 0 1 178976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1340
timestamp 1624015447
transform 1 0 84180 0 -1 180064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1342
timestamp 1624015447
transform 1 0 84180 0 1 180064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_324_906
timestamp 1624015447
transform 1 0 84456 0 -1 178976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_325_906
timestamp 1624015447
transform 1 0 84456 0 1 178976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_326_909
timestamp 1624015447
transform 1 0 84732 0 -1 180064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_327_906
timestamp 1624015447
transform 1 0 84456 0 1 180064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_324_918
timestamp 1624015447
transform 1 0 85560 0 -1 178976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_324_930
timestamp 1624015447
transform 1 0 86664 0 -1 178976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_325_918
timestamp 1624015447
transform 1 0 85560 0 1 178976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_325_930
timestamp 1624015447
transform 1 0 86664 0 1 178976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_326_921
timestamp 1624015447
transform 1 0 85836 0 -1 180064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_326_929
timestamp 1624015447
transform 1 0 86572 0 -1 180064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_327_918
timestamp 1624015447
transform 1 0 85560 0 1 180064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_327_930
timestamp 1624015447
transform 1 0 86664 0 1 180064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1874
timestamp 1624015447
transform 1 0 86848 0 -1 178976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1876
timestamp 1624015447
transform 1 0 86848 0 -1 180064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_324_933
timestamp 1624015447
transform 1 0 86940 0 -1 178976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_324_945
timestamp 1624015447
transform 1 0 88044 0 -1 178976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_325_942
timestamp 1624015447
transform 1 0 87768 0 1 178976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_326_933
timestamp 1624015447
transform 1 0 86940 0 -1 180064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_326_945
timestamp 1624015447
transform 1 0 88044 0 -1 180064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_327_942
timestamp 1624015447
transform 1 0 87768 0 1 180064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1875
timestamp 1624015447
transform 1 0 89424 0 1 178976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1877
timestamp 1624015447
transform 1 0 89424 0 1 180064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_324_957
timestamp 1624015447
transform 1 0 89148 0 -1 178976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_325_954
timestamp 1624015447
transform 1 0 88872 0 1 178976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_325_961
timestamp 1624015447
transform 1 0 89516 0 1 178976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_326_957
timestamp 1624015447
transform 1 0 89148 0 -1 180064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_327_954
timestamp 1624015447
transform 1 0 88872 0 1 180064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_327_961
timestamp 1624015447
transform 1 0 89516 0 1 180064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1337
timestamp 1624015447
transform -1 0 90896 0 -1 178976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1339
timestamp 1624015447
transform -1 0 90896 0 1 178976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1341
timestamp 1624015447
transform -1 0 90896 0 -1 180064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1343
timestamp 1624015447
transform -1 0 90896 0 1 180064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_324_969
timestamp 1624015447
transform 1 0 90252 0 -1 178976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_326_969
timestamp 1624015447
transform 1 0 90252 0 -1 180064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_654
timestamp 1624015447
transform 1 0 1104 0 -1 181152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_656
timestamp 1624015447
transform 1 0 1104 0 1 181152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_658
timestamp 1624015447
transform 1 0 1104 0 -1 182240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_328_3
timestamp 1624015447
transform 1 0 1380 0 -1 181152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_328_15
timestamp 1624015447
transform 1 0 2484 0 -1 181152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_329_3
timestamp 1624015447
transform 1 0 1380 0 1 181152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_329_15
timestamp 1624015447
transform 1 0 2484 0 1 181152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_330_3
timestamp 1624015447
transform 1 0 1380 0 -1 182240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_330_15
timestamp 1624015447
transform 1 0 2484 0 -1 182240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1539
timestamp 1624015447
transform 1 0 3772 0 -1 181152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1540
timestamp 1624015447
transform 1 0 3772 0 -1 182240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_328_27
timestamp 1624015447
transform 1 0 3588 0 -1 181152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_328_30
timestamp 1624015447
transform 1 0 3864 0 -1 181152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_329_27
timestamp 1624015447
transform 1 0 3588 0 1 181152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_330_27
timestamp 1624015447
transform 1 0 3588 0 -1 182240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_330_30
timestamp 1624015447
transform 1 0 3864 0 -1 182240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_655
timestamp 1624015447
transform -1 0 5152 0 -1 181152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_657
timestamp 1624015447
transform -1 0 5152 0 1 181152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_659
timestamp 1624015447
transform -1 0 5152 0 -1 182240
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_addr0[6]
timestamp 1624015447
transform -1 0 4876 0 -1 182240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_328_38
timestamp 1624015447
transform 1 0 4600 0 -1 181152
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_329_39
timestamp 1624015447
transform 1 0 4692 0 1 181152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_330_38
timestamp 1624015447
transform 1 0 4600 0 -1 182240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1344
timestamp 1624015447
transform 1 0 84180 0 -1 181152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1346
timestamp 1624015447
transform 1 0 84180 0 1 181152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1348
timestamp 1624015447
transform 1 0 84180 0 -1 182240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_328_906
timestamp 1624015447
transform 1 0 84456 0 -1 181152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_329_906
timestamp 1624015447
transform 1 0 84456 0 1 181152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_330_906
timestamp 1624015447
transform 1 0 84456 0 -1 182240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_328_918
timestamp 1624015447
transform 1 0 85560 0 -1 181152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_328_930
timestamp 1624015447
transform 1 0 86664 0 -1 181152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_329_918
timestamp 1624015447
transform 1 0 85560 0 1 181152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_329_930
timestamp 1624015447
transform 1 0 86664 0 1 181152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_330_918
timestamp 1624015447
transform 1 0 85560 0 -1 182240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_330_930
timestamp 1624015447
transform 1 0 86664 0 -1 182240
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1878
timestamp 1624015447
transform 1 0 86848 0 -1 181152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1880
timestamp 1624015447
transform 1 0 86848 0 -1 182240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_328_933
timestamp 1624015447
transform 1 0 86940 0 -1 181152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_328_945
timestamp 1624015447
transform 1 0 88044 0 -1 181152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_329_942
timestamp 1624015447
transform 1 0 87768 0 1 181152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_330_933
timestamp 1624015447
transform 1 0 86940 0 -1 182240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_330_945
timestamp 1624015447
transform 1 0 88044 0 -1 182240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1879
timestamp 1624015447
transform 1 0 89424 0 1 181152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_328_957
timestamp 1624015447
transform 1 0 89148 0 -1 181152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_329_954
timestamp 1624015447
transform 1 0 88872 0 1 181152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_329_961
timestamp 1624015447
transform 1 0 89516 0 1 181152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_330_957
timestamp 1624015447
transform 1 0 89148 0 -1 182240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1345
timestamp 1624015447
transform -1 0 90896 0 -1 181152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1347
timestamp 1624015447
transform -1 0 90896 0 1 181152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1349
timestamp 1624015447
transform -1 0 90896 0 -1 182240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_328_969
timestamp 1624015447
transform 1 0 90252 0 -1 181152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_330_969
timestamp 1624015447
transform 1 0 90252 0 -1 182240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_660
timestamp 1624015447
transform 1 0 1104 0 1 182240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_662
timestamp 1624015447
transform 1 0 1104 0 -1 183328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_664
timestamp 1624015447
transform 1 0 1104 0 1 183328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_331_3
timestamp 1624015447
transform 1 0 1380 0 1 182240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_331_15
timestamp 1624015447
transform 1 0 2484 0 1 182240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_332_3
timestamp 1624015447
transform 1 0 1380 0 -1 183328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_332_15
timestamp 1624015447
transform 1 0 2484 0 -1 183328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_333_3
timestamp 1624015447
transform 1 0 1380 0 1 183328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_333_15
timestamp 1624015447
transform 1 0 2484 0 1 183328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1541
timestamp 1624015447
transform 1 0 3772 0 -1 183328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_331_27
timestamp 1624015447
transform 1 0 3588 0 1 182240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_332_27
timestamp 1624015447
transform 1 0 3588 0 -1 183328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_332_30
timestamp 1624015447
transform 1 0 3864 0 -1 183328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_333_27
timestamp 1624015447
transform 1 0 3588 0 1 183328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_661
timestamp 1624015447
transform -1 0 5152 0 1 182240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_663
timestamp 1624015447
transform -1 0 5152 0 -1 183328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_665
timestamp 1624015447
transform -1 0 5152 0 1 183328
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_addr0[7]
timestamp 1624015447
transform -1 0 4876 0 -1 183328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_331_39
timestamp 1624015447
transform 1 0 4692 0 1 182240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_332_38
timestamp 1624015447
transform 1 0 4600 0 -1 183328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_333_39
timestamp 1624015447
transform 1 0 4692 0 1 183328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1350
timestamp 1624015447
transform 1 0 84180 0 1 182240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1352
timestamp 1624015447
transform 1 0 84180 0 -1 183328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1354
timestamp 1624015447
transform 1 0 84180 0 1 183328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_331_906
timestamp 1624015447
transform 1 0 84456 0 1 182240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_332_906
timestamp 1624015447
transform 1 0 84456 0 -1 183328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_333_906
timestamp 1624015447
transform 1 0 84456 0 1 183328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_331_918
timestamp 1624015447
transform 1 0 85560 0 1 182240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_331_930
timestamp 1624015447
transform 1 0 86664 0 1 182240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_332_918
timestamp 1624015447
transform 1 0 85560 0 -1 183328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_332_930
timestamp 1624015447
transform 1 0 86664 0 -1 183328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_333_918
timestamp 1624015447
transform 1 0 85560 0 1 183328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_333_930
timestamp 1624015447
transform 1 0 86664 0 1 183328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1882
timestamp 1624015447
transform 1 0 86848 0 -1 183328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_331_942
timestamp 1624015447
transform 1 0 87768 0 1 182240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_332_933
timestamp 1624015447
transform 1 0 86940 0 -1 183328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_332_945
timestamp 1624015447
transform 1 0 88044 0 -1 183328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_333_942
timestamp 1624015447
transform 1 0 87768 0 1 183328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1881
timestamp 1624015447
transform 1 0 89424 0 1 182240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1883
timestamp 1624015447
transform 1 0 89424 0 1 183328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_331_954
timestamp 1624015447
transform 1 0 88872 0 1 182240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_331_961
timestamp 1624015447
transform 1 0 89516 0 1 182240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_332_957
timestamp 1624015447
transform 1 0 89148 0 -1 183328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_333_954
timestamp 1624015447
transform 1 0 88872 0 1 183328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_333_961
timestamp 1624015447
transform 1 0 89516 0 1 183328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1351
timestamp 1624015447
transform -1 0 90896 0 1 182240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1353
timestamp 1624015447
transform -1 0 90896 0 -1 183328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1355
timestamp 1624015447
transform -1 0 90896 0 1 183328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_332_969
timestamp 1624015447
transform 1 0 90252 0 -1 183328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_666
timestamp 1624015447
transform 1 0 1104 0 -1 184416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_668
timestamp 1624015447
transform 1 0 1104 0 1 184416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_334_3
timestamp 1624015447
transform 1 0 1380 0 -1 184416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_334_15
timestamp 1624015447
transform 1 0 2484 0 -1 184416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_335_3
timestamp 1624015447
transform 1 0 1380 0 1 184416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_335_15
timestamp 1624015447
transform 1 0 2484 0 1 184416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1542
timestamp 1624015447
transform 1 0 3772 0 -1 184416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_334_27
timestamp 1624015447
transform 1 0 3588 0 -1 184416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_334_30
timestamp 1624015447
transform 1 0 3864 0 -1 184416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_335_27
timestamp 1624015447
transform 1 0 3588 0 1 184416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_667
timestamp 1624015447
transform -1 0 5152 0 -1 184416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_669
timestamp 1624015447
transform -1 0 5152 0 1 184416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_334_38
timestamp 1624015447
transform 1 0 4600 0 -1 184416
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_335_39
timestamp 1624015447
transform 1 0 4692 0 1 184416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1356
timestamp 1624015447
transform 1 0 84180 0 -1 184416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1358
timestamp 1624015447
transform 1 0 84180 0 1 184416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_334_906
timestamp 1624015447
transform 1 0 84456 0 -1 184416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_335_906
timestamp 1624015447
transform 1 0 84456 0 1 184416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_334_918
timestamp 1624015447
transform 1 0 85560 0 -1 184416
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_334_930
timestamp 1624015447
transform 1 0 86664 0 -1 184416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_335_918
timestamp 1624015447
transform 1 0 85560 0 1 184416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_335_930
timestamp 1624015447
transform 1 0 86664 0 1 184416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1884
timestamp 1624015447
transform 1 0 86848 0 -1 184416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_334_933
timestamp 1624015447
transform 1 0 86940 0 -1 184416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_334_945
timestamp 1624015447
transform 1 0 88044 0 -1 184416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_335_942
timestamp 1624015447
transform 1 0 87768 0 1 184416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1885
timestamp 1624015447
transform 1 0 89424 0 1 184416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_334_957
timestamp 1624015447
transform 1 0 89148 0 -1 184416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_335_954
timestamp 1624015447
transform 1 0 88872 0 1 184416
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_335_961
timestamp 1624015447
transform 1 0 89516 0 1 184416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1357
timestamp 1624015447
transform -1 0 90896 0 -1 184416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1359
timestamp 1624015447
transform -1 0 90896 0 1 184416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_334_969
timestamp 1624015447
transform 1 0 90252 0 -1 184416
box -38 -48 406 592
use sram_1rw1r_32_256_8_sky130  SRAM_1
timestamp 1624446551
transform 1 0 6000 0 1 96408
box 0 0 77296 91247
use sky130_fd_sc_hd__decap_3  PHY_670
timestamp 1624015447
transform 1 0 1104 0 -1 185504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_672
timestamp 1624015447
transform 1 0 1104 0 1 185504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_336_3
timestamp 1624015447
transform 1 0 1380 0 -1 185504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_337_3
timestamp 1624015447
transform 1 0 1380 0 1 185504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_336_15
timestamp 1624015447
transform 1 0 2484 0 -1 185504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_337_15
timestamp 1624015447
transform 1 0 2484 0 1 185504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1543
timestamp 1624015447
transform 1 0 3772 0 -1 185504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_336_27
timestamp 1624015447
transform 1 0 3588 0 -1 185504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_336_30
timestamp 1624015447
transform 1 0 3864 0 -1 185504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_336_38
timestamp 1624015447
transform 1 0 4600 0 -1 185504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_337_27
timestamp 1624015447
transform 1 0 3588 0 1 185504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_671
timestamp 1624015447
transform -1 0 5152 0 -1 185504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_673
timestamp 1624015447
transform -1 0 5152 0 1 185504
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_337_39
timestamp 1624015447
transform 1 0 4692 0 1 185504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_674
timestamp 1624015447
transform 1 0 1104 0 -1 186592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_338_3
timestamp 1624015447
transform 1 0 1380 0 -1 186592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_338_15
timestamp 1624015447
transform 1 0 2484 0 -1 186592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1544
timestamp 1624015447
transform 1 0 3772 0 -1 186592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_338_27
timestamp 1624015447
transform 1 0 3588 0 -1 186592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_338_30
timestamp 1624015447
transform 1 0 3864 0 -1 186592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_338_38
timestamp 1624015447
transform 1 0 4600 0 -1 186592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_675
timestamp 1624015447
transform -1 0 5152 0 -1 186592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_676
timestamp 1624015447
transform 1 0 1104 0 1 186592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_678
timestamp 1624015447
transform 1 0 1104 0 -1 187680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_339_3
timestamp 1624015447
transform 1 0 1380 0 1 186592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_340_3
timestamp 1624015447
transform 1 0 1380 0 -1 187680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_339_15
timestamp 1624015447
transform 1 0 2484 0 1 186592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_340_15
timestamp 1624015447
transform 1 0 2484 0 -1 187680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1545
timestamp 1624015447
transform 1 0 3772 0 -1 187680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_339_27
timestamp 1624015447
transform 1 0 3588 0 1 186592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_340_27
timestamp 1624015447
transform 1 0 3588 0 -1 187680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_340_30
timestamp 1624015447
transform 1 0 3864 0 -1 187680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_340_38
timestamp 1624015447
transform 1 0 4600 0 -1 187680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_677
timestamp 1624015447
transform -1 0 5152 0 1 186592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_679
timestamp 1624015447
transform -1 0 5152 0 -1 187680
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_339_39
timestamp 1624015447
transform 1 0 4692 0 1 186592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_680
timestamp 1624015447
transform 1 0 1104 0 1 187680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_682
timestamp 1624015447
transform 1 0 1104 0 -1 188768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_341_3
timestamp 1624015447
transform 1 0 1380 0 1 187680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_342_3
timestamp 1624015447
transform 1 0 1380 0 -1 188768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_341_15
timestamp 1624015447
transform 1 0 2484 0 1 187680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_342_15
timestamp 1624015447
transform 1 0 2484 0 -1 188768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1546
timestamp 1624015447
transform 1 0 3772 0 -1 188768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_341_27
timestamp 1624015447
transform 1 0 3588 0 1 187680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_342_27
timestamp 1624015447
transform 1 0 3588 0 -1 188768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_342_30
timestamp 1624015447
transform 1 0 3864 0 -1 188768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_342_38
timestamp 1624015447
transform 1 0 4600 0 -1 188768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_681
timestamp 1624015447
transform -1 0 5152 0 1 187680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_683
timestamp 1624015447
transform -1 0 5152 0 -1 188768
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_341_39
timestamp 1624015447
transform 1 0 4692 0 1 187680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_684
timestamp 1624015447
transform 1 0 1104 0 1 188768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_343_3
timestamp 1624015447
transform 1 0 1380 0 1 188768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_343_15
timestamp 1624015447
transform 1 0 2484 0 1 188768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1547
timestamp 1624015447
transform 1 0 3772 0 1 188768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_343_27
timestamp 1624015447
transform 1 0 3588 0 1 188768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_343_30
timestamp 1624015447
transform 1 0 3864 0 1 188768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_343_38
timestamp 1624015447
transform 1 0 4600 0 1 188768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_685
timestamp 1624015447
transform -1 0 5152 0 1 188768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1360
timestamp 1624015447
transform 1 0 84180 0 -1 185504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1362
timestamp 1624015447
transform 1 0 84180 0 1 185504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1364
timestamp 1624015447
transform 1 0 84180 0 -1 186592
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_csb1
timestamp 1624015447
transform -1 0 84824 0 -1 186592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_336_906
timestamp 1624015447
transform 1 0 84456 0 -1 185504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_337_906
timestamp 1624015447
transform 1 0 84456 0 1 185504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_338_906
timestamp 1624015447
transform 1 0 84456 0 -1 186592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1366
timestamp 1624015447
transform 1 0 84180 0 1 186592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1368
timestamp 1624015447
transform 1 0 84180 0 -1 187680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1370
timestamp 1624015447
transform 1 0 84180 0 1 187680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1372
timestamp 1624015447
transform 1 0 84180 0 -1 188768
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_addr1[0]
timestamp 1624015447
transform -1 0 84824 0 -1 187680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_339_906
timestamp 1624015447
transform 1 0 84456 0 1 186592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_340_906
timestamp 1624015447
transform 1 0 84456 0 -1 187680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_341_906
timestamp 1624015447
transform 1 0 84456 0 1 187680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_342_906
timestamp 1624015447
transform 1 0 84456 0 -1 188768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1374
timestamp 1624015447
transform 1 0 84180 0 1 188768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_343_906
timestamp 1624015447
transform 1 0 84456 0 1 188768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_336_918
timestamp 1624015447
transform 1 0 85560 0 -1 185504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_337_918
timestamp 1624015447
transform 1 0 85560 0 1 185504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1886
timestamp 1624015447
transform 1 0 86848 0 -1 185504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_336_930
timestamp 1624015447
transform 1 0 86664 0 -1 185504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_336_933
timestamp 1624015447
transform 1 0 86940 0 -1 185504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_337_930
timestamp 1624015447
transform 1 0 86664 0 1 185504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_336_945
timestamp 1624015447
transform 1 0 88044 0 -1 185504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_337_942
timestamp 1624015447
transform 1 0 87768 0 1 185504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_336_957
timestamp 1624015447
transform 1 0 89148 0 -1 185504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_337_954
timestamp 1624015447
transform 1 0 88872 0 1 185504
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1887
timestamp 1624015447
transform 1 0 89424 0 1 185504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_336_969
timestamp 1624015447
transform 1 0 90252 0 -1 185504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_337_961
timestamp 1624015447
transform 1 0 89516 0 1 185504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1361
timestamp 1624015447
transform -1 0 90896 0 -1 185504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1363
timestamp 1624015447
transform -1 0 90896 0 1 185504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_338_910
timestamp 1624015447
transform 1 0 84824 0 -1 186592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1888
timestamp 1624015447
transform 1 0 86848 0 -1 186592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_338_922
timestamp 1624015447
transform 1 0 85928 0 -1 186592
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_338_930
timestamp 1624015447
transform 1 0 86664 0 -1 186592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_338_933
timestamp 1624015447
transform 1 0 86940 0 -1 186592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_338_945
timestamp 1624015447
transform 1 0 88044 0 -1 186592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_338_957
timestamp 1624015447
transform 1 0 89148 0 -1 186592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_338_969
timestamp 1624015447
transform 1 0 90252 0 -1 186592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1365
timestamp 1624015447
transform -1 0 90896 0 -1 186592
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_SRAM_1_clk1
timestamp 1624015447
transform -1 0 85192 0 -1 187680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_339_918
timestamp 1624015447
transform 1 0 85560 0 1 186592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_340_910
timestamp 1624015447
transform 1 0 84824 0 -1 187680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_340_914
timestamp 1624015447
transform 1 0 85192 0 -1 187680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1890
timestamp 1624015447
transform 1 0 86848 0 -1 187680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_339_930
timestamp 1624015447
transform 1 0 86664 0 1 186592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_340_926
timestamp 1624015447
transform 1 0 86296 0 -1 187680
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_340_933
timestamp 1624015447
transform 1 0 86940 0 -1 187680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_339_942
timestamp 1624015447
transform 1 0 87768 0 1 186592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_340_945
timestamp 1624015447
transform 1 0 88044 0 -1 187680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_339_954
timestamp 1624015447
transform 1 0 88872 0 1 186592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_340_957
timestamp 1624015447
transform 1 0 89148 0 -1 187680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1889
timestamp 1624015447
transform 1 0 89424 0 1 186592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_339_961
timestamp 1624015447
transform 1 0 89516 0 1 186592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_340_969
timestamp 1624015447
transform 1 0 90252 0 -1 187680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1367
timestamp 1624015447
transform -1 0 90896 0 1 186592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1369
timestamp 1624015447
transform -1 0 90896 0 -1 187680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_341_918
timestamp 1624015447
transform 1 0 85560 0 1 187680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_341_930
timestamp 1624015447
transform 1 0 86664 0 1 187680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_341_942
timestamp 1624015447
transform 1 0 87768 0 1 187680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_341_954
timestamp 1624015447
transform 1 0 88872 0 1 187680
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1891
timestamp 1624015447
transform 1 0 89424 0 1 187680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_341_961
timestamp 1624015447
transform 1 0 89516 0 1 187680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1371
timestamp 1624015447
transform -1 0 90896 0 1 187680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_342_918
timestamp 1624015447
transform 1 0 85560 0 -1 188768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_343_918
timestamp 1624015447
transform 1 0 85560 0 1 188768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1892
timestamp 1624015447
transform 1 0 86848 0 -1 188768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1893
timestamp 1624015447
transform 1 0 86848 0 1 188768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_342_930
timestamp 1624015447
transform 1 0 86664 0 -1 188768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_342_933
timestamp 1624015447
transform 1 0 86940 0 -1 188768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_343_930
timestamp 1624015447
transform 1 0 86664 0 1 188768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_343_933
timestamp 1624015447
transform 1 0 86940 0 1 188768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_342_945
timestamp 1624015447
transform 1 0 88044 0 -1 188768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_343_945
timestamp 1624015447
transform 1 0 88044 0 1 188768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_342_957
timestamp 1624015447
transform 1 0 89148 0 -1 188768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_343_957
timestamp 1624015447
transform 1 0 89148 0 1 188768
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1894
timestamp 1624015447
transform 1 0 89516 0 1 188768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_342_969
timestamp 1624015447
transform 1 0 90252 0 -1 188768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_343_962
timestamp 1624015447
transform 1 0 89608 0 1 188768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_343_970
timestamp 1624015447
transform 1 0 90344 0 1 188768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1373
timestamp 1624015447
transform -1 0 90896 0 -1 188768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1375
timestamp 1624015447
transform -1 0 90896 0 1 188768
box -38 -48 314 592
<< labels >>
rlabel metal3 s 91200 88000 92000 88120 6 mgmt_addr[0]
port 0 nsew signal input
rlabel metal3 s 91200 89224 92000 89344 6 mgmt_addr[1]
port 1 nsew signal input
rlabel metal3 s 91200 90448 92000 90568 6 mgmt_addr[2]
port 2 nsew signal input
rlabel metal3 s 91200 91672 92000 91792 6 mgmt_addr[3]
port 3 nsew signal input
rlabel metal3 s 91200 92896 92000 93016 6 mgmt_addr[4]
port 4 nsew signal input
rlabel metal3 s 91200 94120 92000 94240 6 mgmt_addr[5]
port 5 nsew signal input
rlabel metal3 s 91200 95344 92000 95464 6 mgmt_addr[6]
port 6 nsew signal input
rlabel metal3 s 91200 96568 92000 96688 6 mgmt_addr[7]
port 7 nsew signal input
rlabel metal3 s 91200 97656 92000 97776 6 mgmt_addr_ro[0]
port 8 nsew signal input
rlabel metal3 s 91200 98880 92000 99000 6 mgmt_addr_ro[1]
port 9 nsew signal input
rlabel metal3 s 91200 100104 92000 100224 6 mgmt_addr_ro[2]
port 10 nsew signal input
rlabel metal3 s 91200 101328 92000 101448 6 mgmt_addr_ro[3]
port 11 nsew signal input
rlabel metal3 s 91200 102552 92000 102672 6 mgmt_addr_ro[4]
port 12 nsew signal input
rlabel metal3 s 91200 103776 92000 103896 6 mgmt_addr_ro[5]
port 13 nsew signal input
rlabel metal3 s 91200 105000 92000 105120 6 mgmt_addr_ro[6]
port 14 nsew signal input
rlabel metal3 s 91200 106224 92000 106344 6 mgmt_addr_ro[7]
port 15 nsew signal input
rlabel metal3 s 91200 86776 92000 86896 6 mgmt_clk
port 16 nsew signal input
rlabel metal3 s 91200 552 92000 672 6 mgmt_ena[0]
port 17 nsew signal input
rlabel metal3 s 91200 146344 92000 146464 6 mgmt_ena[1]
port 18 nsew signal input
rlabel metal3 s 91200 1640 92000 1760 6 mgmt_ena_ro
port 19 nsew signal input
rlabel metal3 s 91200 8984 92000 9104 6 mgmt_rdata[0]
port 20 nsew signal tristate
rlabel metal3 s 91200 21088 92000 21208 6 mgmt_rdata[10]
port 21 nsew signal tristate
rlabel metal3 s 91200 22312 92000 22432 6 mgmt_rdata[11]
port 22 nsew signal tristate
rlabel metal3 s 91200 23536 92000 23656 6 mgmt_rdata[12]
port 23 nsew signal tristate
rlabel metal3 s 91200 24760 92000 24880 6 mgmt_rdata[13]
port 24 nsew signal tristate
rlabel metal3 s 91200 25984 92000 26104 6 mgmt_rdata[14]
port 25 nsew signal tristate
rlabel metal3 s 91200 27208 92000 27328 6 mgmt_rdata[15]
port 26 nsew signal tristate
rlabel metal3 s 91200 28432 92000 28552 6 mgmt_rdata[16]
port 27 nsew signal tristate
rlabel metal3 s 91200 29656 92000 29776 6 mgmt_rdata[17]
port 28 nsew signal tristate
rlabel metal3 s 91200 30880 92000 31000 6 mgmt_rdata[18]
port 29 nsew signal tristate
rlabel metal3 s 91200 32104 92000 32224 6 mgmt_rdata[19]
port 30 nsew signal tristate
rlabel metal3 s 91200 10208 92000 10328 6 mgmt_rdata[1]
port 31 nsew signal tristate
rlabel metal3 s 91200 33328 92000 33448 6 mgmt_rdata[20]
port 32 nsew signal tristate
rlabel metal3 s 91200 34552 92000 34672 6 mgmt_rdata[21]
port 33 nsew signal tristate
rlabel metal3 s 91200 35776 92000 35896 6 mgmt_rdata[22]
port 34 nsew signal tristate
rlabel metal3 s 91200 37000 92000 37120 6 mgmt_rdata[23]
port 35 nsew signal tristate
rlabel metal3 s 91200 38224 92000 38344 6 mgmt_rdata[24]
port 36 nsew signal tristate
rlabel metal3 s 91200 39312 92000 39432 6 mgmt_rdata[25]
port 37 nsew signal tristate
rlabel metal3 s 91200 40536 92000 40656 6 mgmt_rdata[26]
port 38 nsew signal tristate
rlabel metal3 s 91200 41760 92000 41880 6 mgmt_rdata[27]
port 39 nsew signal tristate
rlabel metal3 s 91200 42984 92000 43104 6 mgmt_rdata[28]
port 40 nsew signal tristate
rlabel metal3 s 91200 44208 92000 44328 6 mgmt_rdata[29]
port 41 nsew signal tristate
rlabel metal3 s 91200 11432 92000 11552 6 mgmt_rdata[2]
port 42 nsew signal tristate
rlabel metal3 s 91200 45432 92000 45552 6 mgmt_rdata[30]
port 43 nsew signal tristate
rlabel metal3 s 91200 46656 92000 46776 6 mgmt_rdata[31]
port 44 nsew signal tristate
rlabel metal3 s 91200 153688 92000 153808 6 mgmt_rdata[32]
port 45 nsew signal tristate
rlabel metal3 s 91200 154776 92000 154896 6 mgmt_rdata[33]
port 46 nsew signal tristate
rlabel metal3 s 91200 156000 92000 156120 6 mgmt_rdata[34]
port 47 nsew signal tristate
rlabel metal3 s 91200 157224 92000 157344 6 mgmt_rdata[35]
port 48 nsew signal tristate
rlabel metal3 s 91200 158448 92000 158568 6 mgmt_rdata[36]
port 49 nsew signal tristate
rlabel metal3 s 91200 159672 92000 159792 6 mgmt_rdata[37]
port 50 nsew signal tristate
rlabel metal3 s 91200 160896 92000 161016 6 mgmt_rdata[38]
port 51 nsew signal tristate
rlabel metal3 s 91200 162120 92000 162240 6 mgmt_rdata[39]
port 52 nsew signal tristate
rlabel metal3 s 91200 12656 92000 12776 6 mgmt_rdata[3]
port 53 nsew signal tristate
rlabel metal3 s 91200 163344 92000 163464 6 mgmt_rdata[40]
port 54 nsew signal tristate
rlabel metal3 s 91200 164568 92000 164688 6 mgmt_rdata[41]
port 55 nsew signal tristate
rlabel metal3 s 91200 165792 92000 165912 6 mgmt_rdata[42]
port 56 nsew signal tristate
rlabel metal3 s 91200 167016 92000 167136 6 mgmt_rdata[43]
port 57 nsew signal tristate
rlabel metal3 s 91200 168240 92000 168360 6 mgmt_rdata[44]
port 58 nsew signal tristate
rlabel metal3 s 91200 169464 92000 169584 6 mgmt_rdata[45]
port 59 nsew signal tristate
rlabel metal3 s 91200 170688 92000 170808 6 mgmt_rdata[46]
port 60 nsew signal tristate
rlabel metal3 s 91200 171912 92000 172032 6 mgmt_rdata[47]
port 61 nsew signal tristate
rlabel metal3 s 91200 173136 92000 173256 6 mgmt_rdata[48]
port 62 nsew signal tristate
rlabel metal3 s 91200 174224 92000 174344 6 mgmt_rdata[49]
port 63 nsew signal tristate
rlabel metal3 s 91200 13880 92000 14000 6 mgmt_rdata[4]
port 64 nsew signal tristate
rlabel metal3 s 91200 175448 92000 175568 6 mgmt_rdata[50]
port 65 nsew signal tristate
rlabel metal3 s 91200 176672 92000 176792 6 mgmt_rdata[51]
port 66 nsew signal tristate
rlabel metal3 s 91200 177896 92000 178016 6 mgmt_rdata[52]
port 67 nsew signal tristate
rlabel metal3 s 91200 179120 92000 179240 6 mgmt_rdata[53]
port 68 nsew signal tristate
rlabel metal3 s 91200 180344 92000 180464 6 mgmt_rdata[54]
port 69 nsew signal tristate
rlabel metal3 s 91200 181568 92000 181688 6 mgmt_rdata[55]
port 70 nsew signal tristate
rlabel metal3 s 91200 182792 92000 182912 6 mgmt_rdata[56]
port 71 nsew signal tristate
rlabel metal3 s 91200 184016 92000 184136 6 mgmt_rdata[57]
port 72 nsew signal tristate
rlabel metal3 s 91200 185240 92000 185360 6 mgmt_rdata[58]
port 73 nsew signal tristate
rlabel metal3 s 91200 186464 92000 186584 6 mgmt_rdata[59]
port 74 nsew signal tristate
rlabel metal3 s 91200 15104 92000 15224 6 mgmt_rdata[5]
port 75 nsew signal tristate
rlabel metal3 s 91200 187688 92000 187808 6 mgmt_rdata[60]
port 76 nsew signal tristate
rlabel metal3 s 91200 188912 92000 189032 6 mgmt_rdata[61]
port 77 nsew signal tristate
rlabel metal3 s 91200 190136 92000 190256 6 mgmt_rdata[62]
port 78 nsew signal tristate
rlabel metal3 s 91200 191360 92000 191480 6 mgmt_rdata[63]
port 79 nsew signal tristate
rlabel metal3 s 91200 16328 92000 16448 6 mgmt_rdata[6]
port 80 nsew signal tristate
rlabel metal3 s 91200 17552 92000 17672 6 mgmt_rdata[7]
port 81 nsew signal tristate
rlabel metal3 s 91200 18776 92000 18896 6 mgmt_rdata[8]
port 82 nsew signal tristate
rlabel metal3 s 91200 19864 92000 19984 6 mgmt_rdata[9]
port 83 nsew signal tristate
rlabel metal3 s 91200 47880 92000 48000 6 mgmt_rdata_ro[0]
port 84 nsew signal tristate
rlabel metal3 s 91200 59984 92000 60104 6 mgmt_rdata_ro[10]
port 85 nsew signal tristate
rlabel metal3 s 91200 61208 92000 61328 6 mgmt_rdata_ro[11]
port 86 nsew signal tristate
rlabel metal3 s 91200 62432 92000 62552 6 mgmt_rdata_ro[12]
port 87 nsew signal tristate
rlabel metal3 s 91200 63656 92000 63776 6 mgmt_rdata_ro[13]
port 88 nsew signal tristate
rlabel metal3 s 91200 64880 92000 65000 6 mgmt_rdata_ro[14]
port 89 nsew signal tristate
rlabel metal3 s 91200 66104 92000 66224 6 mgmt_rdata_ro[15]
port 90 nsew signal tristate
rlabel metal3 s 91200 67328 92000 67448 6 mgmt_rdata_ro[16]
port 91 nsew signal tristate
rlabel metal3 s 91200 68552 92000 68672 6 mgmt_rdata_ro[17]
port 92 nsew signal tristate
rlabel metal3 s 91200 69776 92000 69896 6 mgmt_rdata_ro[18]
port 93 nsew signal tristate
rlabel metal3 s 91200 71000 92000 71120 6 mgmt_rdata_ro[19]
port 94 nsew signal tristate
rlabel metal3 s 91200 49104 92000 49224 6 mgmt_rdata_ro[1]
port 95 nsew signal tristate
rlabel metal3 s 91200 72224 92000 72344 6 mgmt_rdata_ro[20]
port 96 nsew signal tristate
rlabel metal3 s 91200 73448 92000 73568 6 mgmt_rdata_ro[21]
port 97 nsew signal tristate
rlabel metal3 s 91200 74672 92000 74792 6 mgmt_rdata_ro[22]
port 98 nsew signal tristate
rlabel metal3 s 91200 75896 92000 76016 6 mgmt_rdata_ro[23]
port 99 nsew signal tristate
rlabel metal3 s 91200 77120 92000 77240 6 mgmt_rdata_ro[24]
port 100 nsew signal tristate
rlabel metal3 s 91200 78208 92000 78328 6 mgmt_rdata_ro[25]
port 101 nsew signal tristate
rlabel metal3 s 91200 79432 92000 79552 6 mgmt_rdata_ro[26]
port 102 nsew signal tristate
rlabel metal3 s 91200 80656 92000 80776 6 mgmt_rdata_ro[27]
port 103 nsew signal tristate
rlabel metal3 s 91200 81880 92000 82000 6 mgmt_rdata_ro[28]
port 104 nsew signal tristate
rlabel metal3 s 91200 83104 92000 83224 6 mgmt_rdata_ro[29]
port 105 nsew signal tristate
rlabel metal3 s 91200 50328 92000 50448 6 mgmt_rdata_ro[2]
port 106 nsew signal tristate
rlabel metal3 s 91200 84328 92000 84448 6 mgmt_rdata_ro[30]
port 107 nsew signal tristate
rlabel metal3 s 91200 85552 92000 85672 6 mgmt_rdata_ro[31]
port 108 nsew signal tristate
rlabel metal3 s 91200 51552 92000 51672 6 mgmt_rdata_ro[3]
port 109 nsew signal tristate
rlabel metal3 s 91200 52776 92000 52896 6 mgmt_rdata_ro[4]
port 110 nsew signal tristate
rlabel metal3 s 91200 54000 92000 54120 6 mgmt_rdata_ro[5]
port 111 nsew signal tristate
rlabel metal3 s 91200 55224 92000 55344 6 mgmt_rdata_ro[6]
port 112 nsew signal tristate
rlabel metal3 s 91200 56448 92000 56568 6 mgmt_rdata_ro[7]
port 113 nsew signal tristate
rlabel metal3 s 91200 57672 92000 57792 6 mgmt_rdata_ro[8]
port 114 nsew signal tristate
rlabel metal3 s 91200 58760 92000 58880 6 mgmt_rdata_ro[9]
port 115 nsew signal tristate
rlabel metal3 s 91200 107448 92000 107568 6 mgmt_wdata[0]
port 116 nsew signal input
rlabel metal3 s 91200 119552 92000 119672 6 mgmt_wdata[10]
port 117 nsew signal input
rlabel metal3 s 91200 120776 92000 120896 6 mgmt_wdata[11]
port 118 nsew signal input
rlabel metal3 s 91200 122000 92000 122120 6 mgmt_wdata[12]
port 119 nsew signal input
rlabel metal3 s 91200 123224 92000 123344 6 mgmt_wdata[13]
port 120 nsew signal input
rlabel metal3 s 91200 124448 92000 124568 6 mgmt_wdata[14]
port 121 nsew signal input
rlabel metal3 s 91200 125672 92000 125792 6 mgmt_wdata[15]
port 122 nsew signal input
rlabel metal3 s 91200 126896 92000 127016 6 mgmt_wdata[16]
port 123 nsew signal input
rlabel metal3 s 91200 128120 92000 128240 6 mgmt_wdata[17]
port 124 nsew signal input
rlabel metal3 s 91200 129344 92000 129464 6 mgmt_wdata[18]
port 125 nsew signal input
rlabel metal3 s 91200 130568 92000 130688 6 mgmt_wdata[19]
port 126 nsew signal input
rlabel metal3 s 91200 108672 92000 108792 6 mgmt_wdata[1]
port 127 nsew signal input
rlabel metal3 s 91200 131792 92000 131912 6 mgmt_wdata[20]
port 128 nsew signal input
rlabel metal3 s 91200 133016 92000 133136 6 mgmt_wdata[21]
port 129 nsew signal input
rlabel metal3 s 91200 134240 92000 134360 6 mgmt_wdata[22]
port 130 nsew signal input
rlabel metal3 s 91200 135328 92000 135448 6 mgmt_wdata[23]
port 131 nsew signal input
rlabel metal3 s 91200 136552 92000 136672 6 mgmt_wdata[24]
port 132 nsew signal input
rlabel metal3 s 91200 137776 92000 137896 6 mgmt_wdata[25]
port 133 nsew signal input
rlabel metal3 s 91200 139000 92000 139120 6 mgmt_wdata[26]
port 134 nsew signal input
rlabel metal3 s 91200 140224 92000 140344 6 mgmt_wdata[27]
port 135 nsew signal input
rlabel metal3 s 91200 141448 92000 141568 6 mgmt_wdata[28]
port 136 nsew signal input
rlabel metal3 s 91200 142672 92000 142792 6 mgmt_wdata[29]
port 137 nsew signal input
rlabel metal3 s 91200 109896 92000 110016 6 mgmt_wdata[2]
port 138 nsew signal input
rlabel metal3 s 91200 143896 92000 144016 6 mgmt_wdata[30]
port 139 nsew signal input
rlabel metal3 s 91200 145120 92000 145240 6 mgmt_wdata[31]
port 140 nsew signal input
rlabel metal3 s 91200 111120 92000 111240 6 mgmt_wdata[3]
port 141 nsew signal input
rlabel metal3 s 91200 112344 92000 112464 6 mgmt_wdata[4]
port 142 nsew signal input
rlabel metal3 s 91200 113568 92000 113688 6 mgmt_wdata[5]
port 143 nsew signal input
rlabel metal3 s 91200 114792 92000 114912 6 mgmt_wdata[6]
port 144 nsew signal input
rlabel metal3 s 91200 115880 92000 116000 6 mgmt_wdata[7]
port 145 nsew signal input
rlabel metal3 s 91200 117104 92000 117224 6 mgmt_wdata[8]
port 146 nsew signal input
rlabel metal3 s 91200 118328 92000 118448 6 mgmt_wdata[9]
port 147 nsew signal input
rlabel metal3 s 91200 2864 92000 2984 6 mgmt_wen[0]
port 148 nsew signal input
rlabel metal3 s 91200 147568 92000 147688 6 mgmt_wen[1]
port 149 nsew signal input
rlabel metal3 s 91200 4088 92000 4208 6 mgmt_wen_mask[0]
port 150 nsew signal input
rlabel metal3 s 91200 5312 92000 5432 6 mgmt_wen_mask[1]
port 151 nsew signal input
rlabel metal3 s 91200 6536 92000 6656 6 mgmt_wen_mask[2]
port 152 nsew signal input
rlabel metal3 s 91200 7760 92000 7880 6 mgmt_wen_mask[3]
port 153 nsew signal input
rlabel metal3 s 91200 148792 92000 148912 6 mgmt_wen_mask[4]
port 154 nsew signal input
rlabel metal3 s 91200 150016 92000 150136 6 mgmt_wen_mask[5]
port 155 nsew signal input
rlabel metal3 s 91200 151240 92000 151360 6 mgmt_wen_mask[6]
port 156 nsew signal input
rlabel metal3 s 91200 152464 92000 152584 6 mgmt_wen_mask[7]
port 157 nsew signal input
rlabel metal4 s 89944 2128 90264 189360 6 VPWR
port 158 nsew power bidirectional
rlabel metal4 s 85944 2128 86264 189360 6 VPWR
port 159 nsew power bidirectional
rlabel metal4 s 1944 2128 2264 189360 6 VPWR
port 160 nsew power bidirectional
rlabel metal5 s 1104 185298 90896 185618 6 VPWR
port 161 nsew power bidirectional
rlabel metal5 s 1104 175298 90896 175618 6 VPWR
port 162 nsew power bidirectional
rlabel metal5 s 1104 165298 90896 165618 6 VPWR
port 163 nsew power bidirectional
rlabel metal5 s 1104 155298 90896 155618 6 VPWR
port 164 nsew power bidirectional
rlabel metal5 s 1104 145298 90896 145618 6 VPWR
port 165 nsew power bidirectional
rlabel metal5 s 1104 135298 90896 135618 6 VPWR
port 166 nsew power bidirectional
rlabel metal5 s 1104 125298 90896 125618 6 VPWR
port 167 nsew power bidirectional
rlabel metal5 s 1104 115298 90896 115618 6 VPWR
port 168 nsew power bidirectional
rlabel metal5 s 1104 105298 90896 105618 6 VPWR
port 169 nsew power bidirectional
rlabel metal5 s 1104 95298 90896 95618 6 VPWR
port 170 nsew power bidirectional
rlabel metal5 s 1104 85298 90896 85618 6 VPWR
port 171 nsew power bidirectional
rlabel metal5 s 1104 75298 90896 75618 6 VPWR
port 172 nsew power bidirectional
rlabel metal5 s 1104 65298 90896 65618 6 VPWR
port 173 nsew power bidirectional
rlabel metal5 s 1104 55298 90896 55618 6 VPWR
port 174 nsew power bidirectional
rlabel metal5 s 1104 45298 90896 45618 6 VPWR
port 175 nsew power bidirectional
rlabel metal5 s 1104 35298 90896 35618 6 VPWR
port 176 nsew power bidirectional
rlabel metal5 s 1104 25298 90896 25618 6 VPWR
port 177 nsew power bidirectional
rlabel metal5 s 1104 15298 90896 15618 6 VPWR
port 178 nsew power bidirectional
rlabel metal5 s 1104 5298 90896 5618 6 VPWR
port 179 nsew power bidirectional
rlabel metal4 s 87944 2128 88264 189360 6 VGND
port 180 nsew ground bidirectional
rlabel metal4 s 3944 2128 4264 189360 6 VGND
port 181 nsew ground bidirectional
rlabel metal5 s 1104 180298 90896 180618 6 VGND
port 182 nsew ground bidirectional
rlabel metal5 s 1104 170298 90896 170618 6 VGND
port 183 nsew ground bidirectional
rlabel metal5 s 1104 160298 90896 160618 6 VGND
port 184 nsew ground bidirectional
rlabel metal5 s 1104 150298 90896 150618 6 VGND
port 185 nsew ground bidirectional
rlabel metal5 s 1104 140298 90896 140618 6 VGND
port 186 nsew ground bidirectional
rlabel metal5 s 1104 130298 90896 130618 6 VGND
port 187 nsew ground bidirectional
rlabel metal5 s 1104 120298 90896 120618 6 VGND
port 188 nsew ground bidirectional
rlabel metal5 s 1104 110298 90896 110618 6 VGND
port 189 nsew ground bidirectional
rlabel metal5 s 1104 100298 90896 100618 6 VGND
port 190 nsew ground bidirectional
rlabel metal5 s 1104 90298 90896 90618 6 VGND
port 191 nsew ground bidirectional
rlabel metal5 s 1104 80298 90896 80618 6 VGND
port 192 nsew ground bidirectional
rlabel metal5 s 1104 70298 90896 70618 6 VGND
port 193 nsew ground bidirectional
rlabel metal5 s 1104 60298 90896 60618 6 VGND
port 194 nsew ground bidirectional
rlabel metal5 s 1104 50298 90896 50618 6 VGND
port 195 nsew ground bidirectional
rlabel metal5 s 1104 40298 90896 40618 6 VGND
port 196 nsew ground bidirectional
rlabel metal5 s 1104 30298 90896 30618 6 VGND
port 197 nsew ground bidirectional
rlabel metal5 s 1104 20298 90896 20618 6 VGND
port 198 nsew ground bidirectional
rlabel metal5 s 1104 10298 90896 10618 6 VGND
port 199 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 92000 192000
<< end >>
