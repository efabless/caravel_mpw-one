magic
tech sky130A
magscale 1 2
timestamp 1624273664
<< obsli1 >>
rect 920 2159 9844 11441
<< obsm1 >>
rect 920 1028 14430 13252
<< obsm2 >>
rect 1172 167 14426 13705
<< metal3 >>
rect 14000 13608 34000 13728
rect 14000 13064 34000 13184
rect 14000 12520 34000 12640
rect 14000 12112 34000 12232
rect 14000 11568 34000 11688
rect 14000 11024 34000 11144
rect 14000 10616 34000 10736
rect 14000 10072 34000 10192
rect 14000 9528 34000 9648
rect 14000 9120 34000 9240
rect 14000 8576 34000 8696
rect 14000 8032 34000 8152
rect 14000 7624 34000 7744
rect 14000 7080 34000 7200
rect 14000 6536 34000 6656
rect 14000 6128 34000 6248
rect 14000 5584 34000 5704
rect 14000 5040 34000 5160
rect 14000 4632 34000 4752
rect 14000 4088 34000 4208
rect 14000 3544 34000 3664
rect 14000 3136 34000 3256
rect 14000 2592 34000 2712
rect 14000 2048 34000 2168
rect 14000 1640 34000 1760
rect 14000 1096 34000 1216
rect 14000 552 34000 672
rect 14000 144 34000 264
<< obsm3 >>
rect 1160 2143 9230 11457
<< metal4 >>
rect -1620 -364 -1300 13964
rect -960 296 -640 13304
rect -300 956 20 12644
rect 360 1616 680 11984
rect 1160 5632 1480 12644
rect 2060 5680 2380 13964
rect 2710 5632 3030 12644
rect 3610 5680 3930 13964
rect 1160 956 1480 2128
rect 2060 -364 2380 2080
rect 2710 956 3030 2128
rect 3610 -364 3930 2080
rect 4260 956 4580 12644
rect 5160 -364 5480 13964
rect 5810 956 6130 12644
rect 6710 -364 7030 13964
rect 7360 956 7680 12644
rect 8260 -364 8580 13964
rect 8910 956 9230 12644
rect 10084 1616 10404 11984
rect 10744 956 11064 12644
rect 11404 296 11724 13304
rect 12064 -364 12384 13964
<< obsm4 >>
rect 1478 2432 3314 5248
<< metal5 >>
rect -1620 13644 12384 13964
rect -960 12984 11724 13304
rect -300 12324 11064 12644
rect 360 11664 10404 11984
rect -300 10166 11064 10486
rect -1620 9516 12384 9836
rect -300 8616 11064 8936
rect -1620 7966 12384 8286
rect -300 7066 11064 7386
rect -1620 6416 12384 6736
rect -300 5516 11064 5836
rect -1620 4866 12384 5186
rect -300 3966 11064 4286
rect -1620 3316 12384 3636
rect -300 2416 11064 2736
rect 360 1616 10404 1936
rect -300 956 11064 1276
rect -960 296 11724 616
rect -1620 -364 12384 -44
<< labels >>
rlabel metal3 s 14000 1096 34000 1216 6 mgmt_gpio_in
port 1 nsew signal output
rlabel metal3 s 14000 1640 34000 1760 6 mgmt_gpio_oeb
port 2 nsew signal input
rlabel metal3 s 14000 2048 34000 2168 6 mgmt_gpio_out
port 3 nsew signal input
rlabel metal3 s 14000 552 34000 672 6 one
port 4 nsew signal output
rlabel metal3 s 14000 2592 34000 2712 6 pad_gpio_ana_en
port 5 nsew signal output
rlabel metal3 s 14000 3136 34000 3256 6 pad_gpio_ana_pol
port 6 nsew signal output
rlabel metal3 s 14000 3544 34000 3664 6 pad_gpio_ana_sel
port 7 nsew signal output
rlabel metal3 s 14000 4088 34000 4208 6 pad_gpio_dm[0]
port 8 nsew signal output
rlabel metal3 s 14000 4632 34000 4752 6 pad_gpio_dm[1]
port 9 nsew signal output
rlabel metal3 s 14000 5040 34000 5160 6 pad_gpio_dm[2]
port 10 nsew signal output
rlabel metal3 s 14000 5584 34000 5704 6 pad_gpio_holdover
port 11 nsew signal output
rlabel metal3 s 14000 6128 34000 6248 6 pad_gpio_ib_mode_sel
port 12 nsew signal output
rlabel metal3 s 14000 6536 34000 6656 6 pad_gpio_in
port 13 nsew signal input
rlabel metal3 s 14000 7080 34000 7200 6 pad_gpio_inenb
port 14 nsew signal output
rlabel metal3 s 14000 7624 34000 7744 6 pad_gpio_out
port 15 nsew signal output
rlabel metal3 s 14000 8032 34000 8152 6 pad_gpio_outenb
port 16 nsew signal output
rlabel metal3 s 14000 8576 34000 8696 6 pad_gpio_slow_sel
port 17 nsew signal output
rlabel metal3 s 14000 9120 34000 9240 6 pad_gpio_vtrip_sel
port 18 nsew signal output
rlabel metal3 s 14000 9528 34000 9648 6 resetn
port 19 nsew signal input
rlabel metal3 s 14000 10072 34000 10192 6 resetn_out
port 20 nsew signal output
rlabel metal3 s 14000 10616 34000 10736 6 serial_clock
port 21 nsew signal input
rlabel metal3 s 14000 11024 34000 11144 6 serial_clock_out
port 22 nsew signal output
rlabel metal3 s 14000 11568 34000 11688 6 serial_data_in
port 23 nsew signal input
rlabel metal3 s 14000 12112 34000 12232 6 serial_data_out
port 24 nsew signal output
rlabel metal3 s 14000 12520 34000 12640 6 user_gpio_in
port 25 nsew signal output
rlabel metal3 s 14000 13064 34000 13184 6 user_gpio_oeb
port 26 nsew signal input
rlabel metal3 s 14000 13608 34000 13728 6 user_gpio_out
port 27 nsew signal input
rlabel metal3 s 14000 144 34000 264 6 zero
port 28 nsew signal output
rlabel metal4 s 7360 956 7680 12644 6 vccd
port 29 nsew power bidirectional
rlabel metal4 s 4260 956 4580 12644 6 vccd
port 30 nsew power bidirectional
rlabel metal4 s 1160 5632 1480 12644 6 vccd
port 31 nsew power bidirectional
rlabel metal4 s 10084 1616 10404 11984 6 vccd
port 32 nsew power bidirectional
rlabel metal4 s 360 1616 680 11984 6 vccd
port 33 nsew power bidirectional
rlabel metal4 s 1160 956 1480 2128 6 vccd
port 34 nsew power bidirectional
rlabel metal5 s 360 11664 10404 11984 6 vccd
port 35 nsew power bidirectional
rlabel metal5 s -300 8616 11064 8936 6 vccd
port 36 nsew power bidirectional
rlabel metal5 s -300 5516 11064 5836 6 vccd
port 37 nsew power bidirectional
rlabel metal5 s -300 2416 11064 2736 6 vccd
port 38 nsew power bidirectional
rlabel metal5 s 360 1616 10404 1936 6 vccd
port 39 nsew power bidirectional
rlabel metal4 s 10744 956 11064 12644 6 vssd
port 40 nsew ground bidirectional
rlabel metal4 s 8910 956 9230 12644 6 vssd
port 41 nsew ground bidirectional
rlabel metal4 s 5810 956 6130 12644 6 vssd
port 42 nsew ground bidirectional
rlabel metal4 s 2710 5632 3030 12644 6 vssd
port 43 nsew ground bidirectional
rlabel metal4 s -300 956 20 12644 4 vssd
port 44 nsew ground bidirectional
rlabel metal4 s 2710 956 3030 2128 6 vssd
port 45 nsew ground bidirectional
rlabel metal5 s -300 12324 11064 12644 6 vssd
port 46 nsew ground bidirectional
rlabel metal5 s -300 10166 11064 10486 6 vssd
port 47 nsew ground bidirectional
rlabel metal5 s -300 7066 11064 7386 6 vssd
port 48 nsew ground bidirectional
rlabel metal5 s -300 3966 11064 4286 6 vssd
port 49 nsew ground bidirectional
rlabel metal5 s -300 956 11064 1276 6 vssd
port 50 nsew ground bidirectional
rlabel metal4 s 8260 -364 8580 13964 6 vccd1
port 51 nsew power bidirectional
rlabel metal4 s 5160 -364 5480 13964 6 vccd1
port 52 nsew power bidirectional
rlabel metal4 s 2060 5680 2380 13964 6 vccd1
port 53 nsew power bidirectional
rlabel metal4 s 11404 296 11724 13304 6 vccd1
port 54 nsew power bidirectional
rlabel metal4 s -960 296 -640 13304 4 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 2060 -364 2380 2080 6 vccd1
port 56 nsew power bidirectional
rlabel metal5 s -960 12984 11724 13304 6 vccd1
port 57 nsew power bidirectional
rlabel metal5 s -1620 9516 12384 9836 6 vccd1
port 58 nsew power bidirectional
rlabel metal5 s -1620 6416 12384 6736 6 vccd1
port 59 nsew power bidirectional
rlabel metal5 s -1620 3316 12384 3636 6 vccd1
port 60 nsew power bidirectional
rlabel metal5 s -960 296 11724 616 6 vccd1
port 61 nsew power bidirectional
rlabel metal4 s 12064 -364 12384 13964 6 vssd1
port 62 nsew ground bidirectional
rlabel metal4 s 6710 -364 7030 13964 6 vssd1
port 63 nsew ground bidirectional
rlabel metal4 s 3610 5680 3930 13964 6 vssd1
port 64 nsew ground bidirectional
rlabel metal4 s -1620 -364 -1300 13964 4 vssd1
port 65 nsew ground bidirectional
rlabel metal4 s 3610 -364 3930 2080 6 vssd1
port 66 nsew ground bidirectional
rlabel metal5 s -1620 13644 12384 13964 6 vssd1
port 67 nsew ground bidirectional
rlabel metal5 s -1620 7966 12384 8286 6 vssd1
port 68 nsew ground bidirectional
rlabel metal5 s -1620 4866 12384 5186 6 vssd1
port 69 nsew ground bidirectional
rlabel metal5 s -1620 -364 12384 -44 8 vssd1
port 70 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 34000 14000
string LEFview TRUE
string GDS_FILE ../gds/gpio_control_block.gds
string GDS_END 384068
string GDS_START 156762
<< end >>

